VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2866.790 89.660 2867.110 89.720 ;
        RECT 2898.990 89.660 2899.310 89.720 ;
        RECT 2866.790 89.520 2899.310 89.660 ;
        RECT 2866.790 89.460 2867.110 89.520 ;
        RECT 2898.990 89.460 2899.310 89.520 ;
      LAYER via ;
        RECT 2866.820 89.460 2867.080 89.720 ;
        RECT 2899.020 89.460 2899.280 89.720 ;
      LAYER met2 ;
        RECT 2866.810 159.275 2867.090 159.645 ;
        RECT 2866.880 89.750 2867.020 159.275 ;
        RECT 2866.820 89.430 2867.080 89.750 ;
        RECT 2899.020 89.430 2899.280 89.750 ;
        RECT 2899.080 88.245 2899.220 89.430 ;
        RECT 2899.010 87.875 2899.290 88.245 ;
      LAYER via2 ;
        RECT 2866.810 159.320 2867.090 159.600 ;
        RECT 2899.010 87.920 2899.290 88.200 ;
      LAYER met3 ;
        RECT 2841.000 159.610 2845.000 159.800 ;
        RECT 2866.785 159.610 2867.115 159.625 ;
        RECT 2841.000 159.310 2867.115 159.610 ;
        RECT 2841.000 159.200 2845.000 159.310 ;
        RECT 2866.785 159.295 2867.115 159.310 ;
        RECT 2898.985 88.210 2899.315 88.225 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2898.985 87.910 2924.800 88.210 ;
        RECT 2898.985 87.895 2899.315 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2839.725 3284.825 2839.895 3309.815 ;
        RECT 2839.725 3188.265 2839.895 3211.895 ;
        RECT 2839.725 3091.705 2839.895 3115.335 ;
        RECT 2839.725 2994.465 2839.895 3035.775 ;
        RECT 2839.725 2801.685 2839.895 2815.795 ;
        RECT 2839.725 2753.065 2839.895 2767.175 ;
        RECT 2840.185 2512.005 2840.355 2527.815 ;
        RECT 2840.185 2476.985 2840.355 2511.495 ;
      LAYER mcon ;
        RECT 2839.725 3309.645 2839.895 3309.815 ;
        RECT 2839.725 3211.725 2839.895 3211.895 ;
        RECT 2839.725 3115.165 2839.895 3115.335 ;
        RECT 2839.725 3035.605 2839.895 3035.775 ;
        RECT 2839.725 2815.625 2839.895 2815.795 ;
        RECT 2839.725 2767.005 2839.895 2767.175 ;
        RECT 2840.185 2527.645 2840.355 2527.815 ;
        RECT 2840.185 2511.325 2840.355 2511.495 ;
      LAYER met1 ;
        RECT 942.610 3431.180 942.930 3431.240 ;
        RECT 2839.190 3431.180 2839.510 3431.240 ;
        RECT 942.610 3431.040 2839.510 3431.180 ;
        RECT 942.610 3430.980 942.930 3431.040 ;
        RECT 2839.190 3430.980 2839.510 3431.040 ;
        RECT 2839.650 3309.800 2839.970 3309.860 ;
        RECT 2839.455 3309.660 2839.970 3309.800 ;
        RECT 2839.650 3309.600 2839.970 3309.660 ;
        RECT 2839.650 3284.980 2839.970 3285.040 ;
        RECT 2839.455 3284.840 2839.970 3284.980 ;
        RECT 2839.650 3284.780 2839.970 3284.840 ;
        RECT 2839.650 3211.880 2839.970 3211.940 ;
        RECT 2839.455 3211.740 2839.970 3211.880 ;
        RECT 2839.650 3211.680 2839.970 3211.740 ;
        RECT 2839.650 3188.420 2839.970 3188.480 ;
        RECT 2839.455 3188.280 2839.970 3188.420 ;
        RECT 2839.650 3188.220 2839.970 3188.280 ;
        RECT 2839.650 3115.320 2839.970 3115.380 ;
        RECT 2839.455 3115.180 2839.970 3115.320 ;
        RECT 2839.650 3115.120 2839.970 3115.180 ;
        RECT 2839.650 3091.860 2839.970 3091.920 ;
        RECT 2839.455 3091.720 2839.970 3091.860 ;
        RECT 2839.650 3091.660 2839.970 3091.720 ;
        RECT 2839.650 3035.760 2839.970 3035.820 ;
        RECT 2839.455 3035.620 2839.970 3035.760 ;
        RECT 2839.650 3035.560 2839.970 3035.620 ;
        RECT 2839.650 2994.620 2839.970 2994.680 ;
        RECT 2839.455 2994.480 2839.970 2994.620 ;
        RECT 2839.650 2994.420 2839.970 2994.480 ;
        RECT 2839.650 2863.520 2839.970 2863.780 ;
        RECT 2839.740 2863.100 2839.880 2863.520 ;
        RECT 2839.650 2862.840 2839.970 2863.100 ;
        RECT 2839.650 2815.780 2839.970 2815.840 ;
        RECT 2839.455 2815.640 2839.970 2815.780 ;
        RECT 2839.650 2815.580 2839.970 2815.640 ;
        RECT 2839.650 2801.840 2839.970 2801.900 ;
        RECT 2839.455 2801.700 2839.970 2801.840 ;
        RECT 2839.650 2801.640 2839.970 2801.700 ;
        RECT 2839.650 2767.160 2839.970 2767.220 ;
        RECT 2839.455 2767.020 2839.970 2767.160 ;
        RECT 2839.650 2766.960 2839.970 2767.020 ;
        RECT 2839.650 2753.220 2839.970 2753.280 ;
        RECT 2839.455 2753.080 2839.970 2753.220 ;
        RECT 2839.650 2753.020 2839.970 2753.080 ;
        RECT 2839.650 2670.400 2839.970 2670.660 ;
        RECT 2839.740 2669.980 2839.880 2670.400 ;
        RECT 2839.650 2669.720 2839.970 2669.980 ;
        RECT 2839.650 2574.040 2839.970 2574.100 ;
        RECT 2839.650 2573.900 2840.340 2574.040 ;
        RECT 2839.650 2573.840 2839.970 2573.900 ;
        RECT 2840.200 2573.420 2840.340 2573.900 ;
        RECT 2840.110 2573.160 2840.430 2573.420 ;
        RECT 2840.110 2527.800 2840.430 2527.860 ;
        RECT 2839.915 2527.660 2840.430 2527.800 ;
        RECT 2840.110 2527.600 2840.430 2527.660 ;
        RECT 2840.110 2512.160 2840.430 2512.220 ;
        RECT 2839.915 2512.020 2840.430 2512.160 ;
        RECT 2840.110 2511.960 2840.430 2512.020 ;
        RECT 2840.110 2511.480 2840.430 2511.540 ;
        RECT 2839.915 2511.340 2840.430 2511.480 ;
        RECT 2840.110 2511.280 2840.430 2511.340 ;
        RECT 2839.650 2477.140 2839.970 2477.200 ;
        RECT 2840.125 2477.140 2840.415 2477.185 ;
        RECT 2839.650 2477.000 2840.415 2477.140 ;
        RECT 2839.650 2476.940 2839.970 2477.000 ;
        RECT 2840.125 2476.955 2840.415 2477.000 ;
        RECT 2898.530 2435.660 2898.850 2435.720 ;
        RECT 2839.740 2435.520 2898.850 2435.660 ;
        RECT 2839.740 2435.380 2839.880 2435.520 ;
        RECT 2898.530 2435.460 2898.850 2435.520 ;
        RECT 2839.650 2435.120 2839.970 2435.380 ;
      LAYER via ;
        RECT 942.640 3430.980 942.900 3431.240 ;
        RECT 2839.220 3430.980 2839.480 3431.240 ;
        RECT 2839.680 3309.600 2839.940 3309.860 ;
        RECT 2839.680 3284.780 2839.940 3285.040 ;
        RECT 2839.680 3211.680 2839.940 3211.940 ;
        RECT 2839.680 3188.220 2839.940 3188.480 ;
        RECT 2839.680 3115.120 2839.940 3115.380 ;
        RECT 2839.680 3091.660 2839.940 3091.920 ;
        RECT 2839.680 3035.560 2839.940 3035.820 ;
        RECT 2839.680 2994.420 2839.940 2994.680 ;
        RECT 2839.680 2863.520 2839.940 2863.780 ;
        RECT 2839.680 2862.840 2839.940 2863.100 ;
        RECT 2839.680 2815.580 2839.940 2815.840 ;
        RECT 2839.680 2801.640 2839.940 2801.900 ;
        RECT 2839.680 2766.960 2839.940 2767.220 ;
        RECT 2839.680 2753.020 2839.940 2753.280 ;
        RECT 2839.680 2670.400 2839.940 2670.660 ;
        RECT 2839.680 2669.720 2839.940 2669.980 ;
        RECT 2839.680 2573.840 2839.940 2574.100 ;
        RECT 2840.140 2573.160 2840.400 2573.420 ;
        RECT 2840.140 2527.600 2840.400 2527.860 ;
        RECT 2840.140 2511.960 2840.400 2512.220 ;
        RECT 2840.140 2511.280 2840.400 2511.540 ;
        RECT 2839.680 2476.940 2839.940 2477.200 ;
        RECT 2898.560 2435.460 2898.820 2435.720 ;
        RECT 2839.680 2435.120 2839.940 2435.380 ;
      LAYER met2 ;
        RECT 942.640 3430.950 942.900 3431.270 ;
        RECT 2839.220 3430.950 2839.480 3431.270 ;
        RECT 940.970 3419.450 941.250 3420.000 ;
        RECT 942.700 3419.450 942.840 3430.950 ;
        RECT 940.970 3419.310 942.840 3419.450 ;
        RECT 940.970 3416.000 941.250 3419.310 ;
        RECT 2839.280 3347.370 2839.420 3430.950 ;
        RECT 2838.820 3347.230 2839.420 3347.370 ;
        RECT 2838.820 3309.970 2838.960 3347.230 ;
        RECT 2838.820 3309.890 2839.880 3309.970 ;
        RECT 2838.820 3309.830 2839.940 3309.890 ;
        RECT 2839.680 3309.570 2839.940 3309.830 ;
        RECT 2839.680 3284.980 2839.940 3285.070 ;
        RECT 2839.280 3284.840 2839.940 3284.980 ;
        RECT 2839.280 3250.810 2839.420 3284.840 ;
        RECT 2839.680 3284.750 2839.940 3284.840 ;
        RECT 2838.820 3250.670 2839.420 3250.810 ;
        RECT 2838.820 3212.050 2838.960 3250.670 ;
        RECT 2838.820 3211.970 2839.880 3212.050 ;
        RECT 2838.820 3211.910 2839.940 3211.970 ;
        RECT 2839.680 3211.650 2839.940 3211.910 ;
        RECT 2839.680 3188.250 2839.940 3188.510 ;
        RECT 2839.280 3188.190 2839.940 3188.250 ;
        RECT 2839.280 3188.110 2839.880 3188.190 ;
        RECT 2839.280 3152.890 2839.420 3188.110 ;
        RECT 2838.820 3152.750 2839.420 3152.890 ;
        RECT 2838.820 3115.490 2838.960 3152.750 ;
        RECT 2838.820 3115.410 2839.880 3115.490 ;
        RECT 2838.820 3115.350 2839.940 3115.410 ;
        RECT 2839.680 3115.090 2839.940 3115.350 ;
        RECT 2839.680 3091.690 2839.940 3091.950 ;
        RECT 2839.280 3091.630 2839.940 3091.690 ;
        RECT 2839.280 3091.550 2839.880 3091.630 ;
        RECT 2839.280 3067.210 2839.420 3091.550 ;
        RECT 2838.820 3067.070 2839.420 3067.210 ;
        RECT 2838.820 3035.930 2838.960 3067.070 ;
        RECT 2838.820 3035.850 2839.880 3035.930 ;
        RECT 2838.820 3035.790 2839.940 3035.850 ;
        RECT 2839.680 3035.530 2839.940 3035.790 ;
        RECT 2839.680 2994.620 2839.940 2994.710 ;
        RECT 2839.280 2994.480 2839.940 2994.620 ;
        RECT 2839.280 2873.410 2839.420 2994.480 ;
        RECT 2839.680 2994.390 2839.940 2994.480 ;
        RECT 2839.280 2873.270 2839.880 2873.410 ;
        RECT 2839.740 2863.810 2839.880 2873.270 ;
        RECT 2839.680 2863.490 2839.940 2863.810 ;
        RECT 2839.680 2862.810 2839.940 2863.130 ;
        RECT 2839.740 2849.610 2839.880 2862.810 ;
        RECT 2839.280 2849.470 2839.880 2849.610 ;
        RECT 2839.280 2816.290 2839.420 2849.470 ;
        RECT 2839.280 2816.150 2839.880 2816.290 ;
        RECT 2839.740 2815.870 2839.880 2816.150 ;
        RECT 2839.680 2815.550 2839.940 2815.870 ;
        RECT 2839.680 2801.610 2839.940 2801.930 ;
        RECT 2839.740 2767.250 2839.880 2801.610 ;
        RECT 2839.680 2766.930 2839.940 2767.250 ;
        RECT 2839.740 2753.310 2839.880 2753.465 ;
        RECT 2839.680 2753.050 2839.940 2753.310 ;
        RECT 2839.280 2752.990 2839.940 2753.050 ;
        RECT 2839.280 2752.910 2839.880 2752.990 ;
        RECT 2839.280 2680.970 2839.420 2752.910 ;
        RECT 2839.280 2680.830 2839.880 2680.970 ;
        RECT 2839.740 2670.690 2839.880 2680.830 ;
        RECT 2839.680 2670.370 2839.940 2670.690 ;
        RECT 2839.680 2669.690 2839.940 2670.010 ;
        RECT 2839.740 2656.490 2839.880 2669.690 ;
        RECT 2839.280 2656.350 2839.880 2656.490 ;
        RECT 2839.280 2574.210 2839.420 2656.350 ;
        RECT 2839.280 2574.130 2839.880 2574.210 ;
        RECT 2839.280 2574.070 2839.940 2574.130 ;
        RECT 2839.680 2573.810 2839.940 2574.070 ;
        RECT 2840.140 2573.130 2840.400 2573.450 ;
        RECT 2840.200 2527.890 2840.340 2573.130 ;
        RECT 2840.140 2527.570 2840.400 2527.890 ;
        RECT 2840.140 2511.930 2840.400 2512.250 ;
        RECT 2840.200 2511.570 2840.340 2511.930 ;
        RECT 2840.140 2511.250 2840.400 2511.570 ;
        RECT 2839.680 2476.910 2839.940 2477.230 ;
        RECT 2839.740 2463.370 2839.880 2476.910 ;
        RECT 2839.280 2463.230 2839.880 2463.370 ;
        RECT 2839.280 2435.490 2839.420 2463.230 ;
        RECT 2839.280 2435.410 2839.880 2435.490 ;
        RECT 2898.560 2435.430 2898.820 2435.750 ;
        RECT 2839.280 2435.350 2839.940 2435.410 ;
        RECT 2839.680 2435.090 2839.940 2435.350 ;
        RECT 2898.620 2434.245 2898.760 2435.430 ;
        RECT 2898.550 2433.875 2898.830 2434.245 ;
      LAYER via2 ;
        RECT 2898.550 2433.920 2898.830 2434.200 ;
      LAYER met3 ;
        RECT 2898.525 2434.210 2898.855 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2898.525 2433.910 2924.800 2434.210 ;
        RECT 2898.525 2433.895 2898.855 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2668.740 2924.800 2669.940 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2903.340 2924.800 2904.540 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3137.940 2924.800 3139.140 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3372.540 2924.800 3373.740 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 144.510 3501.560 144.830 3501.620 ;
        RECT 2798.250 3501.560 2798.570 3501.620 ;
        RECT 144.510 3501.420 2798.570 3501.560 ;
        RECT 144.510 3501.360 144.830 3501.420 ;
        RECT 2798.250 3501.360 2798.570 3501.420 ;
      LAYER via ;
        RECT 144.540 3501.360 144.800 3501.620 ;
        RECT 2798.280 3501.360 2798.540 3501.620 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3501.650 2798.480 3517.600 ;
        RECT 144.540 3501.330 144.800 3501.650 ;
        RECT 2798.280 3501.330 2798.540 3501.650 ;
        RECT 144.600 3420.810 144.740 3501.330 ;
        RECT 144.370 3420.670 144.740 3420.810 ;
        RECT 144.370 3420.000 144.510 3420.670 ;
        RECT 144.250 3416.000 144.530 3420.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 234.210 3501.900 234.530 3501.960 ;
        RECT 2473.950 3501.900 2474.270 3501.960 ;
        RECT 234.210 3501.760 2474.270 3501.900 ;
        RECT 234.210 3501.700 234.530 3501.760 ;
        RECT 2473.950 3501.700 2474.270 3501.760 ;
      LAYER via ;
        RECT 234.240 3501.700 234.500 3501.960 ;
        RECT 2473.980 3501.700 2474.240 3501.960 ;
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3501.990 2474.180 3517.600 ;
        RECT 234.240 3501.670 234.500 3501.990 ;
        RECT 2473.980 3501.670 2474.240 3501.990 ;
        RECT 232.570 3419.450 232.850 3420.000 ;
        RECT 234.300 3419.450 234.440 3501.670 ;
        RECT 232.570 3419.310 234.440 3419.450 ;
        RECT 232.570 3416.000 232.850 3419.310 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 323.910 3502.240 324.230 3502.300 ;
        RECT 2149.190 3502.240 2149.510 3502.300 ;
        RECT 323.910 3502.100 2149.510 3502.240 ;
        RECT 323.910 3502.040 324.230 3502.100 ;
        RECT 2149.190 3502.040 2149.510 3502.100 ;
      LAYER via ;
        RECT 323.940 3502.040 324.200 3502.300 ;
        RECT 2149.220 3502.040 2149.480 3502.300 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3502.330 2149.420 3517.600 ;
        RECT 323.940 3502.010 324.200 3502.330 ;
        RECT 2149.220 3502.010 2149.480 3502.330 ;
        RECT 320.890 3418.770 321.170 3420.000 ;
        RECT 324.000 3418.770 324.140 3502.010 ;
        RECT 320.890 3418.630 324.140 3418.770 ;
        RECT 320.890 3416.000 321.170 3418.630 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 413.610 3502.580 413.930 3502.640 ;
        RECT 1824.890 3502.580 1825.210 3502.640 ;
        RECT 413.610 3502.440 1825.210 3502.580 ;
        RECT 413.610 3502.380 413.930 3502.440 ;
        RECT 1824.890 3502.380 1825.210 3502.440 ;
        RECT 411.310 3435.940 411.630 3436.000 ;
        RECT 413.610 3435.940 413.930 3436.000 ;
        RECT 411.310 3435.800 413.930 3435.940 ;
        RECT 411.310 3435.740 411.630 3435.800 ;
        RECT 413.610 3435.740 413.930 3435.800 ;
      LAYER via ;
        RECT 413.640 3502.380 413.900 3502.640 ;
        RECT 1824.920 3502.380 1825.180 3502.640 ;
        RECT 411.340 3435.740 411.600 3436.000 ;
        RECT 413.640 3435.740 413.900 3436.000 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3502.670 1825.120 3517.600 ;
        RECT 413.640 3502.350 413.900 3502.670 ;
        RECT 1824.920 3502.350 1825.180 3502.670 ;
        RECT 413.700 3436.030 413.840 3502.350 ;
        RECT 411.340 3435.710 411.600 3436.030 ;
        RECT 413.640 3435.710 413.900 3436.030 ;
        RECT 409.670 3419.450 409.950 3420.000 ;
        RECT 411.400 3419.450 411.540 3435.710 ;
        RECT 409.670 3419.310 411.540 3419.450 ;
        RECT 409.670 3416.000 409.950 3419.310 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 503.310 3502.920 503.630 3502.980 ;
        RECT 1500.590 3502.920 1500.910 3502.980 ;
        RECT 503.310 3502.780 1500.910 3502.920 ;
        RECT 503.310 3502.720 503.630 3502.780 ;
        RECT 1500.590 3502.720 1500.910 3502.780 ;
        RECT 499.630 3434.240 499.950 3434.300 ;
        RECT 503.310 3434.240 503.630 3434.300 ;
        RECT 499.630 3434.100 503.630 3434.240 ;
        RECT 499.630 3434.040 499.950 3434.100 ;
        RECT 503.310 3434.040 503.630 3434.100 ;
      LAYER via ;
        RECT 503.340 3502.720 503.600 3502.980 ;
        RECT 1500.620 3502.720 1500.880 3502.980 ;
        RECT 499.660 3434.040 499.920 3434.300 ;
        RECT 503.340 3434.040 503.600 3434.300 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3503.010 1500.820 3517.600 ;
        RECT 503.340 3502.690 503.600 3503.010 ;
        RECT 1500.620 3502.690 1500.880 3503.010 ;
        RECT 503.400 3434.330 503.540 3502.690 ;
        RECT 499.660 3434.010 499.920 3434.330 ;
        RECT 503.340 3434.010 503.600 3434.330 ;
        RECT 497.990 3419.450 498.270 3420.000 ;
        RECT 499.720 3419.450 499.860 3434.010 ;
        RECT 497.990 3419.310 499.860 3419.450 ;
        RECT 497.990 3416.000 498.270 3419.310 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2887.030 317.800 2887.350 317.860 ;
        RECT 2900.830 317.800 2901.150 317.860 ;
        RECT 2887.030 317.660 2901.150 317.800 ;
        RECT 2887.030 317.600 2887.350 317.660 ;
        RECT 2900.830 317.600 2901.150 317.660 ;
        RECT 2856.210 276.660 2856.530 276.720 ;
        RECT 2887.030 276.660 2887.350 276.720 ;
        RECT 2856.210 276.520 2887.350 276.660 ;
        RECT 2856.210 276.460 2856.530 276.520 ;
        RECT 2887.030 276.460 2887.350 276.520 ;
      LAYER via ;
        RECT 2887.060 317.600 2887.320 317.860 ;
        RECT 2900.860 317.600 2901.120 317.860 ;
        RECT 2856.240 276.460 2856.500 276.720 ;
        RECT 2887.060 276.460 2887.320 276.720 ;
      LAYER met2 ;
        RECT 2900.850 322.475 2901.130 322.845 ;
        RECT 2900.920 317.890 2901.060 322.475 ;
        RECT 2887.060 317.570 2887.320 317.890 ;
        RECT 2900.860 317.570 2901.120 317.890 ;
        RECT 2887.120 276.750 2887.260 317.570 ;
        RECT 2856.240 276.605 2856.500 276.750 ;
        RECT 2856.230 276.235 2856.510 276.605 ;
        RECT 2887.060 276.430 2887.320 276.750 ;
      LAYER via2 ;
        RECT 2900.850 322.520 2901.130 322.800 ;
        RECT 2856.230 276.280 2856.510 276.560 ;
      LAYER met3 ;
        RECT 2900.825 322.810 2901.155 322.825 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2900.825 322.510 2924.800 322.810 ;
        RECT 2900.825 322.495 2901.155 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
        RECT 2841.000 277.520 2845.000 278.120 ;
        RECT 2843.110 276.570 2843.410 277.520 ;
        RECT 2856.205 276.570 2856.535 276.585 ;
        RECT 2843.110 276.270 2856.535 276.570 ;
        RECT 2856.205 276.255 2856.535 276.270 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 593.010 3503.260 593.330 3503.320 ;
        RECT 1175.830 3503.260 1176.150 3503.320 ;
        RECT 593.010 3503.120 1176.150 3503.260 ;
        RECT 593.010 3503.060 593.330 3503.120 ;
        RECT 1175.830 3503.060 1176.150 3503.120 ;
        RECT 588.410 3435.600 588.730 3435.660 ;
        RECT 593.010 3435.600 593.330 3435.660 ;
        RECT 588.410 3435.460 593.330 3435.600 ;
        RECT 588.410 3435.400 588.730 3435.460 ;
        RECT 593.010 3435.400 593.330 3435.460 ;
      LAYER via ;
        RECT 593.040 3503.060 593.300 3503.320 ;
        RECT 1175.860 3503.060 1176.120 3503.320 ;
        RECT 588.440 3435.400 588.700 3435.660 ;
        RECT 593.040 3435.400 593.300 3435.660 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3503.350 1176.060 3517.600 ;
        RECT 593.040 3503.030 593.300 3503.350 ;
        RECT 1175.860 3503.030 1176.120 3503.350 ;
        RECT 593.100 3435.690 593.240 3503.030 ;
        RECT 588.440 3435.370 588.700 3435.690 ;
        RECT 593.040 3435.370 593.300 3435.690 ;
        RECT 586.770 3419.450 587.050 3420.000 ;
        RECT 588.500 3419.450 588.640 3435.370 ;
        RECT 586.770 3419.310 588.640 3419.450 ;
        RECT 586.770 3416.000 587.050 3419.310 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 675.810 3503.600 676.130 3503.660 ;
        RECT 851.530 3503.600 851.850 3503.660 ;
        RECT 675.810 3503.460 851.850 3503.600 ;
        RECT 675.810 3503.400 676.130 3503.460 ;
        RECT 851.530 3503.400 851.850 3503.460 ;
      LAYER via ;
        RECT 675.840 3503.400 676.100 3503.660 ;
        RECT 851.560 3503.400 851.820 3503.660 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3503.690 851.760 3517.600 ;
        RECT 675.840 3503.370 676.100 3503.690 ;
        RECT 851.560 3503.370 851.820 3503.690 ;
        RECT 675.090 3419.450 675.370 3420.000 ;
        RECT 675.900 3419.450 676.040 3503.370 ;
        RECT 675.090 3419.310 676.040 3419.450 ;
        RECT 675.090 3416.000 675.370 3419.310 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 527.230 3503.260 527.550 3503.320 ;
        RECT 530.910 3503.260 531.230 3503.320 ;
        RECT 527.230 3503.120 531.230 3503.260 ;
        RECT 527.230 3503.060 527.550 3503.120 ;
        RECT 530.910 3503.060 531.230 3503.120 ;
        RECT 530.910 3433.560 531.230 3433.620 ;
        RECT 762.290 3433.560 762.610 3433.620 ;
        RECT 530.910 3433.420 762.610 3433.560 ;
        RECT 530.910 3433.360 531.230 3433.420 ;
        RECT 762.290 3433.360 762.610 3433.420 ;
      LAYER via ;
        RECT 527.260 3503.060 527.520 3503.320 ;
        RECT 530.940 3503.060 531.200 3503.320 ;
        RECT 530.940 3433.360 531.200 3433.620 ;
        RECT 762.320 3433.360 762.580 3433.620 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3503.350 527.460 3517.600 ;
        RECT 527.260 3503.030 527.520 3503.350 ;
        RECT 530.940 3503.030 531.200 3503.350 ;
        RECT 531.000 3433.650 531.140 3503.030 ;
        RECT 530.940 3433.330 531.200 3433.650 ;
        RECT 762.320 3433.330 762.580 3433.650 ;
        RECT 762.380 3419.450 762.520 3433.330 ;
        RECT 763.870 3419.450 764.150 3420.000 ;
        RECT 762.380 3419.310 764.150 3419.450 ;
        RECT 763.870 3416.000 764.150 3419.310 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 202.470 3502.240 202.790 3502.300 ;
        RECT 206.610 3502.240 206.930 3502.300 ;
        RECT 202.470 3502.100 206.930 3502.240 ;
        RECT 202.470 3502.040 202.790 3502.100 ;
        RECT 206.610 3502.040 206.930 3502.100 ;
        RECT 206.610 3433.220 206.930 3433.280 ;
        RECT 850.610 3433.220 850.930 3433.280 ;
        RECT 206.610 3433.080 850.930 3433.220 ;
        RECT 206.610 3433.020 206.930 3433.080 ;
        RECT 850.610 3433.020 850.930 3433.080 ;
      LAYER via ;
        RECT 202.500 3502.040 202.760 3502.300 ;
        RECT 206.640 3502.040 206.900 3502.300 ;
        RECT 206.640 3433.020 206.900 3433.280 ;
        RECT 850.640 3433.020 850.900 3433.280 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3502.330 202.700 3517.600 ;
        RECT 202.500 3502.010 202.760 3502.330 ;
        RECT 206.640 3502.010 206.900 3502.330 ;
        RECT 206.700 3433.310 206.840 3502.010 ;
        RECT 206.640 3432.990 206.900 3433.310 ;
        RECT 850.640 3432.990 850.900 3433.310 ;
        RECT 850.700 3419.450 850.840 3432.990 ;
        RECT 852.190 3419.450 852.470 3420.000 ;
        RECT 850.700 3419.310 852.470 3419.450 ;
        RECT 852.190 3416.000 852.470 3419.310 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3410.620 2.400 3411.820 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3123.660 2.400 3124.860 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2836.020 2.400 2837.220 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2549.060 2.400 2550.260 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2261.420 2.400 2262.620 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1974.460 2.400 1975.660 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2866.790 552.400 2867.110 552.460 ;
        RECT 2898.070 552.400 2898.390 552.460 ;
        RECT 2866.790 552.260 2898.390 552.400 ;
        RECT 2866.790 552.200 2867.110 552.260 ;
        RECT 2898.070 552.200 2898.390 552.260 ;
        RECT 2856.210 396.340 2856.530 396.400 ;
        RECT 2866.790 396.340 2867.110 396.400 ;
        RECT 2856.210 396.200 2867.110 396.340 ;
        RECT 2856.210 396.140 2856.530 396.200 ;
        RECT 2866.790 396.140 2867.110 396.200 ;
      LAYER via ;
        RECT 2866.820 552.200 2867.080 552.460 ;
        RECT 2898.100 552.200 2898.360 552.460 ;
        RECT 2856.240 396.140 2856.500 396.400 ;
        RECT 2866.820 396.140 2867.080 396.400 ;
      LAYER met2 ;
        RECT 2898.090 557.075 2898.370 557.445 ;
        RECT 2898.160 552.490 2898.300 557.075 ;
        RECT 2866.820 552.170 2867.080 552.490 ;
        RECT 2898.100 552.170 2898.360 552.490 ;
        RECT 2866.880 396.430 2867.020 552.170 ;
        RECT 2856.240 396.285 2856.500 396.430 ;
        RECT 2856.230 395.915 2856.510 396.285 ;
        RECT 2866.820 396.110 2867.080 396.430 ;
      LAYER via2 ;
        RECT 2898.090 557.120 2898.370 557.400 ;
        RECT 2856.230 395.960 2856.510 396.240 ;
      LAYER met3 ;
        RECT 2898.065 557.410 2898.395 557.425 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2898.065 557.110 2924.800 557.410 ;
        RECT 2898.065 557.095 2898.395 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
        RECT 2841.000 396.250 2845.000 396.440 ;
        RECT 2856.205 396.250 2856.535 396.265 ;
        RECT 2841.000 395.950 2856.535 396.250 ;
        RECT 2841.000 395.840 2845.000 395.950 ;
        RECT 2856.205 395.935 2856.535 395.950 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1686.820 2.400 1688.020 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1471.260 2.400 1472.460 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1255.700 2.400 1256.900 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1040.140 2.400 1041.340 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 824.580 2.400 825.780 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 609.700 2.400 610.900 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 394.140 2.400 395.340 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 178.580 2.400 179.780 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2873.690 787.000 2874.010 787.060 ;
        RECT 2898.070 787.000 2898.390 787.060 ;
        RECT 2873.690 786.860 2898.390 787.000 ;
        RECT 2873.690 786.800 2874.010 786.860 ;
        RECT 2898.070 786.800 2898.390 786.860 ;
        RECT 2856.210 515.340 2856.530 515.400 ;
        RECT 2873.690 515.340 2874.010 515.400 ;
        RECT 2856.210 515.200 2874.010 515.340 ;
        RECT 2856.210 515.140 2856.530 515.200 ;
        RECT 2873.690 515.140 2874.010 515.200 ;
      LAYER via ;
        RECT 2873.720 786.800 2873.980 787.060 ;
        RECT 2898.100 786.800 2898.360 787.060 ;
        RECT 2856.240 515.140 2856.500 515.400 ;
        RECT 2873.720 515.140 2873.980 515.400 ;
      LAYER met2 ;
        RECT 2898.090 791.675 2898.370 792.045 ;
        RECT 2898.160 787.090 2898.300 791.675 ;
        RECT 2873.720 786.770 2873.980 787.090 ;
        RECT 2898.100 786.770 2898.360 787.090 ;
        RECT 2873.780 515.430 2873.920 786.770 ;
        RECT 2856.240 515.285 2856.500 515.430 ;
        RECT 2856.230 514.915 2856.510 515.285 ;
        RECT 2873.720 515.110 2873.980 515.430 ;
      LAYER via2 ;
        RECT 2898.090 791.720 2898.370 792.000 ;
        RECT 2856.230 514.960 2856.510 515.240 ;
      LAYER met3 ;
        RECT 2898.065 792.010 2898.395 792.025 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2898.065 791.710 2924.800 792.010 ;
        RECT 2898.065 791.695 2898.395 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
        RECT 2841.000 515.250 2845.000 515.440 ;
        RECT 2856.205 515.250 2856.535 515.265 ;
        RECT 2841.000 514.950 2856.535 515.250 ;
        RECT 2841.000 514.840 2845.000 514.950 ;
        RECT 2856.205 514.935 2856.535 514.950 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2866.790 1021.600 2867.110 1021.660 ;
        RECT 2898.070 1021.600 2898.390 1021.660 ;
        RECT 2866.790 1021.460 2898.390 1021.600 ;
        RECT 2866.790 1021.400 2867.110 1021.460 ;
        RECT 2898.070 1021.400 2898.390 1021.460 ;
        RECT 2856.210 633.660 2856.530 633.720 ;
        RECT 2866.790 633.660 2867.110 633.720 ;
        RECT 2856.210 633.520 2867.110 633.660 ;
        RECT 2856.210 633.460 2856.530 633.520 ;
        RECT 2866.790 633.460 2867.110 633.520 ;
      LAYER via ;
        RECT 2866.820 1021.400 2867.080 1021.660 ;
        RECT 2898.100 1021.400 2898.360 1021.660 ;
        RECT 2856.240 633.460 2856.500 633.720 ;
        RECT 2866.820 633.460 2867.080 633.720 ;
      LAYER met2 ;
        RECT 2898.090 1026.275 2898.370 1026.645 ;
        RECT 2898.160 1021.690 2898.300 1026.275 ;
        RECT 2866.820 1021.370 2867.080 1021.690 ;
        RECT 2898.100 1021.370 2898.360 1021.690 ;
        RECT 2866.880 633.750 2867.020 1021.370 ;
        RECT 2856.240 633.605 2856.500 633.750 ;
        RECT 2856.230 633.235 2856.510 633.605 ;
        RECT 2866.820 633.430 2867.080 633.750 ;
      LAYER via2 ;
        RECT 2898.090 1026.320 2898.370 1026.600 ;
        RECT 2856.230 633.280 2856.510 633.560 ;
      LAYER met3 ;
        RECT 2898.065 1026.610 2898.395 1026.625 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2898.065 1026.310 2924.800 1026.610 ;
        RECT 2898.065 1026.295 2898.395 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
        RECT 2841.000 633.570 2845.000 633.760 ;
        RECT 2856.205 633.570 2856.535 633.585 ;
        RECT 2841.000 633.270 2856.535 633.570 ;
        RECT 2841.000 633.160 2845.000 633.270 ;
        RECT 2856.205 633.255 2856.535 633.270 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2880.590 1256.200 2880.910 1256.260 ;
        RECT 2898.070 1256.200 2898.390 1256.260 ;
        RECT 2880.590 1256.060 2898.390 1256.200 ;
        RECT 2880.590 1256.000 2880.910 1256.060 ;
        RECT 2898.070 1256.000 2898.390 1256.060 ;
        RECT 2856.210 751.980 2856.530 752.040 ;
        RECT 2880.590 751.980 2880.910 752.040 ;
        RECT 2856.210 751.840 2880.910 751.980 ;
        RECT 2856.210 751.780 2856.530 751.840 ;
        RECT 2880.590 751.780 2880.910 751.840 ;
      LAYER via ;
        RECT 2880.620 1256.000 2880.880 1256.260 ;
        RECT 2898.100 1256.000 2898.360 1256.260 ;
        RECT 2856.240 751.780 2856.500 752.040 ;
        RECT 2880.620 751.780 2880.880 752.040 ;
      LAYER met2 ;
        RECT 2898.090 1260.875 2898.370 1261.245 ;
        RECT 2898.160 1256.290 2898.300 1260.875 ;
        RECT 2880.620 1255.970 2880.880 1256.290 ;
        RECT 2898.100 1255.970 2898.360 1256.290 ;
        RECT 2880.680 752.070 2880.820 1255.970 ;
        RECT 2856.240 751.925 2856.500 752.070 ;
        RECT 2856.230 751.555 2856.510 751.925 ;
        RECT 2880.620 751.750 2880.880 752.070 ;
      LAYER via2 ;
        RECT 2898.090 1260.920 2898.370 1261.200 ;
        RECT 2856.230 751.600 2856.510 751.880 ;
      LAYER met3 ;
        RECT 2898.065 1261.210 2898.395 1261.225 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2898.065 1260.910 2924.800 1261.210 ;
        RECT 2898.065 1260.895 2898.395 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
        RECT 2841.000 751.890 2845.000 752.080 ;
        RECT 2856.205 751.890 2856.535 751.905 ;
        RECT 2841.000 751.590 2856.535 751.890 ;
        RECT 2841.000 751.480 2845.000 751.590 ;
        RECT 2856.205 751.575 2856.535 751.590 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2873.690 1490.800 2874.010 1490.860 ;
        RECT 2898.070 1490.800 2898.390 1490.860 ;
        RECT 2873.690 1490.660 2898.390 1490.800 ;
        RECT 2873.690 1490.600 2874.010 1490.660 ;
        RECT 2898.070 1490.600 2898.390 1490.660 ;
        RECT 2856.210 870.980 2856.530 871.040 ;
        RECT 2873.690 870.980 2874.010 871.040 ;
        RECT 2856.210 870.840 2874.010 870.980 ;
        RECT 2856.210 870.780 2856.530 870.840 ;
        RECT 2873.690 870.780 2874.010 870.840 ;
      LAYER via ;
        RECT 2873.720 1490.600 2873.980 1490.860 ;
        RECT 2898.100 1490.600 2898.360 1490.860 ;
        RECT 2856.240 870.780 2856.500 871.040 ;
        RECT 2873.720 870.780 2873.980 871.040 ;
      LAYER met2 ;
        RECT 2898.090 1495.475 2898.370 1495.845 ;
        RECT 2898.160 1490.890 2898.300 1495.475 ;
        RECT 2873.720 1490.570 2873.980 1490.890 ;
        RECT 2898.100 1490.570 2898.360 1490.890 ;
        RECT 2873.780 871.070 2873.920 1490.570 ;
        RECT 2856.240 870.925 2856.500 871.070 ;
        RECT 2856.230 870.555 2856.510 870.925 ;
        RECT 2873.720 870.750 2873.980 871.070 ;
      LAYER via2 ;
        RECT 2898.090 1495.520 2898.370 1495.800 ;
        RECT 2856.230 870.600 2856.510 870.880 ;
      LAYER met3 ;
        RECT 2898.065 1495.810 2898.395 1495.825 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2898.065 1495.510 2924.800 1495.810 ;
        RECT 2898.065 1495.495 2898.395 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
        RECT 2841.000 870.890 2845.000 871.080 ;
        RECT 2856.205 870.890 2856.535 870.905 ;
        RECT 2841.000 870.590 2856.535 870.890 ;
        RECT 2841.000 870.480 2845.000 870.590 ;
        RECT 2856.205 870.575 2856.535 870.590 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2887.490 1727.780 2887.810 1727.840 ;
        RECT 2898.070 1727.780 2898.390 1727.840 ;
        RECT 2887.490 1727.640 2898.390 1727.780 ;
        RECT 2887.490 1727.580 2887.810 1727.640 ;
        RECT 2898.070 1727.580 2898.390 1727.640 ;
        RECT 2856.210 987.260 2856.530 987.320 ;
        RECT 2887.490 987.260 2887.810 987.320 ;
        RECT 2856.210 987.120 2887.810 987.260 ;
        RECT 2856.210 987.060 2856.530 987.120 ;
        RECT 2887.490 987.060 2887.810 987.120 ;
      LAYER via ;
        RECT 2887.520 1727.580 2887.780 1727.840 ;
        RECT 2898.100 1727.580 2898.360 1727.840 ;
        RECT 2856.240 987.060 2856.500 987.320 ;
        RECT 2887.520 987.060 2887.780 987.320 ;
      LAYER met2 ;
        RECT 2898.090 1730.075 2898.370 1730.445 ;
        RECT 2898.160 1727.870 2898.300 1730.075 ;
        RECT 2887.520 1727.550 2887.780 1727.870 ;
        RECT 2898.100 1727.550 2898.360 1727.870 ;
        RECT 2856.230 987.515 2856.510 987.885 ;
        RECT 2856.300 987.350 2856.440 987.515 ;
        RECT 2887.580 987.350 2887.720 1727.550 ;
        RECT 2856.240 987.030 2856.500 987.350 ;
        RECT 2887.520 987.030 2887.780 987.350 ;
      LAYER via2 ;
        RECT 2898.090 1730.120 2898.370 1730.400 ;
        RECT 2856.230 987.560 2856.510 987.840 ;
      LAYER met3 ;
        RECT 2898.065 1730.410 2898.395 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2898.065 1730.110 2924.800 1730.410 ;
        RECT 2898.065 1730.095 2898.395 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
        RECT 2841.000 988.800 2845.000 989.400 ;
        RECT 2844.030 987.850 2844.330 988.800 ;
        RECT 2856.205 987.850 2856.535 987.865 ;
        RECT 2844.030 987.550 2856.535 987.850 ;
        RECT 2856.205 987.535 2856.535 987.550 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2866.790 1960.000 2867.110 1960.060 ;
        RECT 2898.070 1960.000 2898.390 1960.060 ;
        RECT 2866.790 1959.860 2898.390 1960.000 ;
        RECT 2866.790 1959.800 2867.110 1959.860 ;
        RECT 2898.070 1959.800 2898.390 1959.860 ;
        RECT 2856.210 1107.620 2856.530 1107.680 ;
        RECT 2866.790 1107.620 2867.110 1107.680 ;
        RECT 2856.210 1107.480 2867.110 1107.620 ;
        RECT 2856.210 1107.420 2856.530 1107.480 ;
        RECT 2866.790 1107.420 2867.110 1107.480 ;
      LAYER via ;
        RECT 2866.820 1959.800 2867.080 1960.060 ;
        RECT 2898.100 1959.800 2898.360 1960.060 ;
        RECT 2856.240 1107.420 2856.500 1107.680 ;
        RECT 2866.820 1107.420 2867.080 1107.680 ;
      LAYER met2 ;
        RECT 2898.090 1964.675 2898.370 1965.045 ;
        RECT 2898.160 1960.090 2898.300 1964.675 ;
        RECT 2866.820 1959.770 2867.080 1960.090 ;
        RECT 2898.100 1959.770 2898.360 1960.090 ;
        RECT 2866.880 1107.710 2867.020 1959.770 ;
        RECT 2856.240 1107.565 2856.500 1107.710 ;
        RECT 2856.230 1107.195 2856.510 1107.565 ;
        RECT 2866.820 1107.390 2867.080 1107.710 ;
      LAYER via2 ;
        RECT 2898.090 1964.720 2898.370 1965.000 ;
        RECT 2856.230 1107.240 2856.510 1107.520 ;
      LAYER met3 ;
        RECT 2898.065 1965.010 2898.395 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2898.065 1964.710 2924.800 1965.010 ;
        RECT 2898.065 1964.695 2898.395 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
        RECT 2841.000 1107.530 2845.000 1107.720 ;
        RECT 2856.205 1107.530 2856.535 1107.545 ;
        RECT 2841.000 1107.230 2856.535 1107.530 ;
        RECT 2841.000 1107.120 2845.000 1107.230 ;
        RECT 2856.205 1107.215 2856.535 1107.230 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2856.210 1221.860 2856.530 1221.920 ;
        RECT 2894.390 1221.860 2894.710 1221.920 ;
        RECT 2856.210 1221.720 2894.710 1221.860 ;
        RECT 2856.210 1221.660 2856.530 1221.720 ;
        RECT 2894.390 1221.660 2894.710 1221.720 ;
      LAYER via ;
        RECT 2856.240 1221.660 2856.500 1221.920 ;
        RECT 2894.420 1221.660 2894.680 1221.920 ;
      LAYER met2 ;
        RECT 2894.410 2199.275 2894.690 2199.645 ;
        RECT 2856.230 1223.475 2856.510 1223.845 ;
        RECT 2856.300 1221.950 2856.440 1223.475 ;
        RECT 2894.480 1221.950 2894.620 2199.275 ;
        RECT 2856.240 1221.630 2856.500 1221.950 ;
        RECT 2894.420 1221.630 2894.680 1221.950 ;
      LAYER via2 ;
        RECT 2894.410 2199.320 2894.690 2199.600 ;
        RECT 2856.230 1223.520 2856.510 1223.800 ;
      LAYER met3 ;
        RECT 2894.385 2199.610 2894.715 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2894.385 2199.310 2924.800 2199.610 ;
        RECT 2894.385 2199.295 2894.715 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
        RECT 2841.000 1226.120 2845.000 1226.720 ;
        RECT 2844.030 1223.810 2844.330 1226.120 ;
        RECT 2856.205 1223.810 2856.535 1223.825 ;
        RECT 2844.030 1223.510 2856.535 1223.810 ;
        RECT 2856.205 1223.495 2856.535 1223.510 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 204.420 2924.800 205.620 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2551.100 2924.800 2552.300 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2785.700 2924.800 2786.900 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3020.300 2924.800 3021.500 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3254.900 2924.800 3256.100 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3489.500 2924.800 3490.700 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 439.020 2924.800 440.220 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 3267.140 2.400 3268.340 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2979.500 2.400 2980.700 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2692.540 2.400 2693.740 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2404.900 2.400 2406.100 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2117.940 2.400 2119.140 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1830.300 2.400 1831.500 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 673.620 2924.800 674.820 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1543.340 2.400 1544.540 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1327.780 2.400 1328.980 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1112.220 2.400 1113.420 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 896.660 2.400 897.860 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 681.100 2.400 682.300 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 465.540 2.400 466.740 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 249.980 2.400 251.180 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 35.100 2.400 36.300 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 908.900 2924.800 910.100 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1143.500 2924.800 1144.700 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1378.100 2924.800 1379.300 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1612.700 2924.800 1613.900 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1847.300 2924.800 1848.500 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2081.900 2924.800 2083.100 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2316.500 2924.800 2317.700 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 145.940 2924.800 147.140 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2492.620 2924.800 2493.820 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 306.890 96.460 307.210 96.520 ;
        RECT 2902.670 96.460 2902.990 96.520 ;
        RECT 306.890 96.320 2902.990 96.460 ;
        RECT 306.890 96.260 307.210 96.320 ;
        RECT 2902.670 96.260 2902.990 96.320 ;
      LAYER via ;
        RECT 306.920 96.260 307.180 96.520 ;
        RECT 2902.700 96.260 2902.960 96.520 ;
      LAYER met2 ;
        RECT 2902.690 2727.635 2902.970 2728.005 ;
        RECT 305.250 100.370 305.530 104.000 ;
        RECT 305.250 100.230 307.120 100.370 ;
        RECT 305.250 100.000 305.530 100.230 ;
        RECT 306.980 96.550 307.120 100.230 ;
        RECT 2902.760 96.550 2902.900 2727.635 ;
        RECT 306.920 96.230 307.180 96.550 ;
        RECT 2902.700 96.230 2902.960 96.550 ;
      LAYER via2 ;
        RECT 2902.690 2727.680 2902.970 2727.960 ;
      LAYER met3 ;
        RECT 2902.665 2727.970 2902.995 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2902.665 2727.670 2924.800 2727.970 ;
        RECT 2902.665 2727.655 2902.995 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 351.050 96.120 351.370 96.180 ;
        RECT 2902.210 96.120 2902.530 96.180 ;
        RECT 351.050 95.980 2902.530 96.120 ;
        RECT 351.050 95.920 351.370 95.980 ;
        RECT 2902.210 95.920 2902.530 95.980 ;
      LAYER via ;
        RECT 351.080 95.920 351.340 96.180 ;
        RECT 2902.240 95.920 2902.500 96.180 ;
      LAYER met2 ;
        RECT 2902.230 2962.235 2902.510 2962.605 ;
        RECT 351.250 100.370 351.530 104.000 ;
        RECT 351.140 100.000 351.530 100.370 ;
        RECT 351.140 96.210 351.280 100.000 ;
        RECT 2902.300 96.210 2902.440 2962.235 ;
        RECT 351.080 95.890 351.340 96.210 ;
        RECT 2902.240 95.890 2902.500 96.210 ;
      LAYER via2 ;
        RECT 2902.230 2962.280 2902.510 2962.560 ;
      LAYER met3 ;
        RECT 2902.205 2962.570 2902.535 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2902.205 2962.270 2924.800 2962.570 ;
        RECT 2902.205 2962.255 2902.535 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 398.430 95.780 398.750 95.840 ;
        RECT 2901.750 95.780 2902.070 95.840 ;
        RECT 398.430 95.640 2902.070 95.780 ;
        RECT 398.430 95.580 398.750 95.640 ;
        RECT 2901.750 95.580 2902.070 95.640 ;
      LAYER via ;
        RECT 398.460 95.580 398.720 95.840 ;
        RECT 2901.780 95.580 2902.040 95.840 ;
      LAYER met2 ;
        RECT 2901.770 3196.835 2902.050 3197.205 ;
        RECT 396.790 100.370 397.070 104.000 ;
        RECT 396.790 100.230 398.660 100.370 ;
        RECT 396.790 100.000 397.070 100.230 ;
        RECT 398.520 95.870 398.660 100.230 ;
        RECT 2901.840 95.870 2901.980 3196.835 ;
        RECT 398.460 95.550 398.720 95.870 ;
        RECT 2901.780 95.550 2902.040 95.870 ;
      LAYER via2 ;
        RECT 2901.770 3196.880 2902.050 3197.160 ;
      LAYER met3 ;
        RECT 2901.745 3197.170 2902.075 3197.185 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2901.745 3196.870 2924.800 3197.170 ;
        RECT 2901.745 3196.855 2902.075 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 444.430 95.440 444.750 95.500 ;
        RECT 2901.290 95.440 2901.610 95.500 ;
        RECT 444.430 95.300 2901.610 95.440 ;
        RECT 444.430 95.240 444.750 95.300 ;
        RECT 2901.290 95.240 2901.610 95.300 ;
      LAYER via ;
        RECT 444.460 95.240 444.720 95.500 ;
        RECT 2901.320 95.240 2901.580 95.500 ;
      LAYER met2 ;
        RECT 2901.310 3431.435 2901.590 3431.805 ;
        RECT 442.790 100.370 443.070 104.000 ;
        RECT 442.790 100.230 444.660 100.370 ;
        RECT 442.790 100.000 443.070 100.230 ;
        RECT 444.520 95.530 444.660 100.230 ;
        RECT 2901.380 95.530 2901.520 3431.435 ;
        RECT 444.460 95.210 444.720 95.530 ;
        RECT 2901.320 95.210 2901.580 95.530 ;
      LAYER via2 ;
        RECT 2901.310 3431.480 2901.590 3431.760 ;
      LAYER met3 ;
        RECT 2901.285 3431.770 2901.615 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2901.285 3431.470 2924.800 3431.770 ;
        RECT 2901.285 3431.455 2901.615 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 380.540 2924.800 381.740 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3339.720 17.410 3339.780 ;
        RECT 99.890 3339.720 100.210 3339.780 ;
        RECT 17.090 3339.580 100.210 3339.720 ;
        RECT 17.090 3339.520 17.410 3339.580 ;
        RECT 99.890 3339.520 100.210 3339.580 ;
        RECT 99.890 103.260 100.210 103.320 ;
        RECT 121.050 103.260 121.370 103.320 ;
        RECT 99.890 103.120 121.370 103.260 ;
        RECT 99.890 103.060 100.210 103.120 ;
        RECT 121.050 103.060 121.370 103.120 ;
      LAYER via ;
        RECT 17.120 3339.520 17.380 3339.780 ;
        RECT 99.920 3339.520 100.180 3339.780 ;
        RECT 99.920 103.060 100.180 103.320 ;
        RECT 121.080 103.060 121.340 103.320 ;
      LAYER met2 ;
        RECT 17.110 3339.635 17.390 3340.005 ;
        RECT 17.120 3339.490 17.380 3339.635 ;
        RECT 99.920 3339.490 100.180 3339.810 ;
        RECT 99.980 103.350 100.120 3339.490 ;
        RECT 99.920 103.030 100.180 103.350 ;
        RECT 121.080 103.090 121.340 103.350 ;
        RECT 122.630 103.090 122.910 104.000 ;
        RECT 121.080 103.030 122.910 103.090 ;
        RECT 121.140 102.950 122.910 103.030 ;
        RECT 122.630 100.000 122.910 102.950 ;
      LAYER via2 ;
        RECT 17.110 3339.680 17.390 3339.960 ;
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 17.085 3339.970 17.415 3339.985 ;
        RECT -4.800 3339.670 17.415 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 17.085 3339.655 17.415 3339.670 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3050.040 17.410 3050.100 ;
        RECT 79.190 3050.040 79.510 3050.100 ;
        RECT 17.090 3049.900 79.510 3050.040 ;
        RECT 17.090 3049.840 17.410 3049.900 ;
        RECT 79.190 3049.840 79.510 3049.900 ;
        RECT 79.190 88.980 79.510 89.040 ;
        RECT 166.590 88.980 166.910 89.040 ;
        RECT 79.190 88.840 166.910 88.980 ;
        RECT 79.190 88.780 79.510 88.840 ;
        RECT 166.590 88.780 166.910 88.840 ;
      LAYER via ;
        RECT 17.120 3049.840 17.380 3050.100 ;
        RECT 79.220 3049.840 79.480 3050.100 ;
        RECT 79.220 88.780 79.480 89.040 ;
        RECT 166.620 88.780 166.880 89.040 ;
      LAYER met2 ;
        RECT 17.110 3051.995 17.390 3052.365 ;
        RECT 17.180 3050.130 17.320 3051.995 ;
        RECT 17.120 3049.810 17.380 3050.130 ;
        RECT 79.220 3049.810 79.480 3050.130 ;
        RECT 79.280 89.070 79.420 3049.810 ;
        RECT 168.170 100.370 168.450 104.000 ;
        RECT 166.680 100.230 168.450 100.370 ;
        RECT 166.680 89.070 166.820 100.230 ;
        RECT 168.170 100.000 168.450 100.230 ;
        RECT 79.220 88.750 79.480 89.070 ;
        RECT 166.620 88.750 166.880 89.070 ;
      LAYER via2 ;
        RECT 17.110 3052.040 17.390 3052.320 ;
      LAYER met3 ;
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 17.085 3052.330 17.415 3052.345 ;
        RECT -4.800 3052.030 17.415 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 17.085 3052.015 17.415 3052.030 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 2760.360 16.030 2760.420 ;
        RECT 92.990 2760.360 93.310 2760.420 ;
        RECT 15.710 2760.220 93.310 2760.360 ;
        RECT 15.710 2760.160 16.030 2760.220 ;
        RECT 92.990 2760.160 93.310 2760.220 ;
        RECT 92.990 89.320 93.310 89.380 ;
        RECT 212.130 89.320 212.450 89.380 ;
        RECT 92.990 89.180 212.450 89.320 ;
        RECT 92.990 89.120 93.310 89.180 ;
        RECT 212.130 89.120 212.450 89.180 ;
      LAYER via ;
        RECT 15.740 2760.160 16.000 2760.420 ;
        RECT 93.020 2760.160 93.280 2760.420 ;
        RECT 93.020 89.120 93.280 89.380 ;
        RECT 212.160 89.120 212.420 89.380 ;
      LAYER met2 ;
        RECT 15.730 2765.035 16.010 2765.405 ;
        RECT 15.800 2760.450 15.940 2765.035 ;
        RECT 15.740 2760.130 16.000 2760.450 ;
        RECT 93.020 2760.130 93.280 2760.450 ;
        RECT 93.080 89.410 93.220 2760.130 ;
        RECT 213.710 100.370 213.990 104.000 ;
        RECT 212.220 100.230 213.990 100.370 ;
        RECT 212.220 89.410 212.360 100.230 ;
        RECT 213.710 100.000 213.990 100.230 ;
        RECT 93.020 89.090 93.280 89.410 ;
        RECT 212.160 89.090 212.420 89.410 ;
      LAYER via2 ;
        RECT 15.730 2765.080 16.010 2765.360 ;
      LAYER met3 ;
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 15.705 2765.370 16.035 2765.385 ;
        RECT -4.800 2765.070 16.035 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 15.705 2765.055 16.035 2765.070 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 88.640 17.410 88.700 ;
        RECT 258.130 88.640 258.450 88.700 ;
        RECT 17.090 88.500 258.450 88.640 ;
        RECT 17.090 88.440 17.410 88.500 ;
        RECT 258.130 88.440 258.450 88.500 ;
      LAYER via ;
        RECT 17.120 88.440 17.380 88.700 ;
        RECT 258.160 88.440 258.420 88.700 ;
      LAYER met2 ;
        RECT 17.110 2477.395 17.390 2477.765 ;
        RECT 17.180 88.730 17.320 2477.395 ;
        RECT 259.710 100.370 259.990 104.000 ;
        RECT 258.220 100.230 259.990 100.370 ;
        RECT 258.220 88.730 258.360 100.230 ;
        RECT 259.710 100.000 259.990 100.230 ;
        RECT 17.120 88.410 17.380 88.730 ;
        RECT 258.160 88.410 258.420 88.730 ;
      LAYER via2 ;
        RECT 17.110 2477.440 17.390 2477.720 ;
      LAYER met3 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 17.085 2477.730 17.415 2477.745 ;
        RECT -4.800 2477.430 17.415 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 17.085 2477.415 17.415 2477.430 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 2187.460 17.870 2187.520 ;
        RECT 37.790 2187.460 38.110 2187.520 ;
        RECT 17.550 2187.320 38.110 2187.460 ;
        RECT 17.550 2187.260 17.870 2187.320 ;
        RECT 37.790 2187.260 38.110 2187.320 ;
        RECT 37.790 172.280 38.110 172.340 ;
        RECT 85.170 172.280 85.490 172.340 ;
        RECT 37.790 172.140 85.490 172.280 ;
        RECT 37.790 172.080 38.110 172.140 ;
        RECT 85.170 172.080 85.490 172.140 ;
      LAYER via ;
        RECT 17.580 2187.260 17.840 2187.520 ;
        RECT 37.820 2187.260 38.080 2187.520 ;
        RECT 37.820 172.080 38.080 172.340 ;
        RECT 85.200 172.080 85.460 172.340 ;
      LAYER met2 ;
        RECT 17.570 2189.755 17.850 2190.125 ;
        RECT 17.640 2187.550 17.780 2189.755 ;
        RECT 17.580 2187.230 17.840 2187.550 ;
        RECT 37.820 2187.230 38.080 2187.550 ;
        RECT 37.880 172.370 38.020 2187.230 ;
        RECT 37.820 172.050 38.080 172.370 ;
        RECT 85.200 172.050 85.460 172.370 ;
        RECT 85.260 166.445 85.400 172.050 ;
        RECT 85.190 166.075 85.470 166.445 ;
      LAYER via2 ;
        RECT 17.570 2189.800 17.850 2190.080 ;
        RECT 85.190 166.120 85.470 166.400 ;
      LAYER met3 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 17.545 2190.090 17.875 2190.105 ;
        RECT -4.800 2189.790 17.875 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 17.545 2189.775 17.875 2189.790 ;
        RECT 85.165 166.410 85.495 166.425 ;
        RECT 100.000 166.410 104.000 166.600 ;
        RECT 85.165 166.110 104.000 166.410 ;
        RECT 85.165 166.095 85.495 166.110 ;
        RECT 100.000 166.000 104.000 166.110 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 303.520 17.870 303.580 ;
        RECT 84.710 303.520 85.030 303.580 ;
        RECT 17.550 303.380 85.030 303.520 ;
        RECT 17.550 303.320 17.870 303.380 ;
        RECT 84.710 303.320 85.030 303.380 ;
      LAYER via ;
        RECT 17.580 303.320 17.840 303.580 ;
        RECT 84.740 303.320 85.000 303.580 ;
      LAYER met2 ;
        RECT 17.570 1902.795 17.850 1903.165 ;
        RECT 17.640 303.610 17.780 1902.795 ;
        RECT 17.580 303.290 17.840 303.610 ;
        RECT 84.740 303.290 85.000 303.610 ;
        RECT 84.800 299.045 84.940 303.290 ;
        RECT 84.730 298.675 85.010 299.045 ;
      LAYER via2 ;
        RECT 17.570 1902.840 17.850 1903.120 ;
        RECT 84.730 298.720 85.010 299.000 ;
      LAYER met3 ;
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 17.545 1903.130 17.875 1903.145 ;
        RECT -4.800 1902.830 17.875 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
        RECT 17.545 1902.815 17.875 1902.830 ;
        RECT 84.705 299.010 85.035 299.025 ;
        RECT 100.000 299.010 104.000 299.200 ;
        RECT 84.705 298.710 104.000 299.010 ;
        RECT 84.705 298.695 85.035 298.710 ;
        RECT 100.000 298.600 104.000 298.710 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 615.140 2924.800 616.340 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 1614.900 16.950 1614.960 ;
        RECT 51.590 1614.900 51.910 1614.960 ;
        RECT 16.630 1614.760 51.910 1614.900 ;
        RECT 16.630 1614.700 16.950 1614.760 ;
        RECT 51.590 1614.700 51.910 1614.760 ;
        RECT 51.590 433.060 51.910 433.120 ;
        RECT 85.170 433.060 85.490 433.120 ;
        RECT 51.590 432.920 85.490 433.060 ;
        RECT 51.590 432.860 51.910 432.920 ;
        RECT 85.170 432.860 85.490 432.920 ;
      LAYER via ;
        RECT 16.660 1614.700 16.920 1614.960 ;
        RECT 51.620 1614.700 51.880 1614.960 ;
        RECT 51.620 432.860 51.880 433.120 ;
        RECT 85.200 432.860 85.460 433.120 ;
      LAYER met2 ;
        RECT 16.650 1615.155 16.930 1615.525 ;
        RECT 16.720 1614.990 16.860 1615.155 ;
        RECT 16.660 1614.670 16.920 1614.990 ;
        RECT 51.620 1614.670 51.880 1614.990 ;
        RECT 51.680 433.150 51.820 1614.670 ;
        RECT 51.620 432.830 51.880 433.150 ;
        RECT 85.200 432.830 85.460 433.150 ;
        RECT 85.260 431.645 85.400 432.830 ;
        RECT 85.190 431.275 85.470 431.645 ;
      LAYER via2 ;
        RECT 16.650 1615.200 16.930 1615.480 ;
        RECT 85.190 431.320 85.470 431.600 ;
      LAYER met3 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 16.625 1615.490 16.955 1615.505 ;
        RECT -4.800 1615.190 16.955 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 16.625 1615.175 16.955 1615.190 ;
        RECT 85.165 431.610 85.495 431.625 ;
        RECT 100.000 431.610 104.000 431.800 ;
        RECT 85.165 431.310 104.000 431.610 ;
        RECT 85.165 431.295 85.495 431.310 ;
        RECT 100.000 431.200 104.000 431.310 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.010 565.660 18.330 565.720 ;
        RECT 85.170 565.660 85.490 565.720 ;
        RECT 18.010 565.520 85.490 565.660 ;
        RECT 18.010 565.460 18.330 565.520 ;
        RECT 85.170 565.460 85.490 565.520 ;
      LAYER via ;
        RECT 18.040 565.460 18.300 565.720 ;
        RECT 85.200 565.460 85.460 565.720 ;
      LAYER met2 ;
        RECT 18.030 1400.275 18.310 1400.645 ;
        RECT 18.100 565.750 18.240 1400.275 ;
        RECT 18.040 565.430 18.300 565.750 ;
        RECT 85.200 565.430 85.460 565.750 ;
        RECT 85.260 564.245 85.400 565.430 ;
        RECT 85.190 563.875 85.470 564.245 ;
      LAYER via2 ;
        RECT 18.030 1400.320 18.310 1400.600 ;
        RECT 85.190 563.920 85.470 564.200 ;
      LAYER met3 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 18.005 1400.610 18.335 1400.625 ;
        RECT -4.800 1400.310 18.335 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 18.005 1400.295 18.335 1400.310 ;
        RECT 85.165 564.210 85.495 564.225 ;
        RECT 100.000 564.210 104.000 564.400 ;
        RECT 85.165 563.910 104.000 564.210 ;
        RECT 85.165 563.895 85.495 563.910 ;
        RECT 100.000 563.800 104.000 563.910 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.470 703.700 18.790 703.760 ;
        RECT 83.790 703.700 84.110 703.760 ;
        RECT 18.470 703.560 84.110 703.700 ;
        RECT 18.470 703.500 18.790 703.560 ;
        RECT 83.790 703.500 84.110 703.560 ;
      LAYER via ;
        RECT 18.500 703.500 18.760 703.760 ;
        RECT 83.820 703.500 84.080 703.760 ;
      LAYER met2 ;
        RECT 18.490 1184.715 18.770 1185.085 ;
        RECT 18.560 703.790 18.700 1184.715 ;
        RECT 18.500 703.470 18.760 703.790 ;
        RECT 83.820 703.470 84.080 703.790 ;
        RECT 83.880 697.525 84.020 703.470 ;
        RECT 83.810 697.155 84.090 697.525 ;
      LAYER via2 ;
        RECT 18.490 1184.760 18.770 1185.040 ;
        RECT 83.810 697.200 84.090 697.480 ;
      LAYER met3 ;
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 18.465 1185.050 18.795 1185.065 ;
        RECT -4.800 1184.750 18.795 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 18.465 1184.735 18.795 1184.750 ;
        RECT 83.785 697.490 84.115 697.505 ;
        RECT 100.000 697.490 104.000 697.680 ;
        RECT 83.785 697.190 104.000 697.490 ;
        RECT 83.785 697.175 84.115 697.190 ;
        RECT 100.000 697.080 104.000 697.190 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.390 834.940 19.710 835.000 ;
        RECT 85.170 834.940 85.490 835.000 ;
        RECT 19.390 834.800 85.490 834.940 ;
        RECT 19.390 834.740 19.710 834.800 ;
        RECT 85.170 834.740 85.490 834.800 ;
      LAYER via ;
        RECT 19.420 834.740 19.680 835.000 ;
        RECT 85.200 834.740 85.460 835.000 ;
      LAYER met2 ;
        RECT 19.410 969.155 19.690 969.525 ;
        RECT 19.480 835.030 19.620 969.155 ;
        RECT 19.420 834.710 19.680 835.030 ;
        RECT 85.200 834.710 85.460 835.030 ;
        RECT 85.260 830.125 85.400 834.710 ;
        RECT 85.190 829.755 85.470 830.125 ;
      LAYER via2 ;
        RECT 19.410 969.200 19.690 969.480 ;
        RECT 85.190 829.800 85.470 830.080 ;
      LAYER met3 ;
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 19.385 969.490 19.715 969.505 ;
        RECT -4.800 969.190 19.715 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
        RECT 19.385 969.175 19.715 969.190 ;
        RECT 85.165 830.090 85.495 830.105 ;
        RECT 100.000 830.090 104.000 830.280 ;
        RECT 85.165 829.790 104.000 830.090 ;
        RECT 85.165 829.775 85.495 829.790 ;
        RECT 100.000 829.680 104.000 829.790 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.930 959.380 19.250 959.440 ;
        RECT 85.170 959.380 85.490 959.440 ;
        RECT 18.930 959.240 85.490 959.380 ;
        RECT 18.930 959.180 19.250 959.240 ;
        RECT 85.170 959.180 85.490 959.240 ;
      LAYER via ;
        RECT 18.960 959.180 19.220 959.440 ;
        RECT 85.200 959.180 85.460 959.440 ;
      LAYER met2 ;
        RECT 85.190 962.355 85.470 962.725 ;
        RECT 85.260 959.470 85.400 962.355 ;
        RECT 18.960 959.150 19.220 959.470 ;
        RECT 85.200 959.150 85.460 959.470 ;
        RECT 19.020 753.965 19.160 959.150 ;
        RECT 18.950 753.595 19.230 753.965 ;
      LAYER via2 ;
        RECT 85.190 962.400 85.470 962.680 ;
        RECT 18.950 753.640 19.230 753.920 ;
      LAYER met3 ;
        RECT 85.165 962.690 85.495 962.705 ;
        RECT 100.000 962.690 104.000 962.880 ;
        RECT 85.165 962.390 104.000 962.690 ;
        RECT 85.165 962.375 85.495 962.390 ;
        RECT 100.000 962.280 104.000 962.390 ;
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 18.925 753.930 19.255 753.945 ;
        RECT -4.800 753.630 19.255 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
        RECT 18.925 753.615 19.255 753.630 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 58.950 1090.280 59.270 1090.340 ;
        RECT 85.170 1090.280 85.490 1090.340 ;
        RECT 58.950 1090.140 85.490 1090.280 ;
        RECT 58.950 1090.080 59.270 1090.140 ;
        RECT 85.170 1090.080 85.490 1090.140 ;
        RECT 16.630 544.920 16.950 544.980 ;
        RECT 58.950 544.920 59.270 544.980 ;
        RECT 16.630 544.780 59.270 544.920 ;
        RECT 16.630 544.720 16.950 544.780 ;
        RECT 58.950 544.720 59.270 544.780 ;
      LAYER via ;
        RECT 58.980 1090.080 59.240 1090.340 ;
        RECT 85.200 1090.080 85.460 1090.340 ;
        RECT 16.660 544.720 16.920 544.980 ;
        RECT 58.980 544.720 59.240 544.980 ;
      LAYER met2 ;
        RECT 85.190 1094.955 85.470 1095.325 ;
        RECT 85.260 1090.370 85.400 1094.955 ;
        RECT 58.980 1090.050 59.240 1090.370 ;
        RECT 85.200 1090.050 85.460 1090.370 ;
        RECT 59.040 545.010 59.180 1090.050 ;
        RECT 16.660 544.690 16.920 545.010 ;
        RECT 58.980 544.690 59.240 545.010 ;
        RECT 16.720 538.405 16.860 544.690 ;
        RECT 16.650 538.035 16.930 538.405 ;
      LAYER via2 ;
        RECT 85.190 1095.000 85.470 1095.280 ;
        RECT 16.650 538.080 16.930 538.360 ;
      LAYER met3 ;
        RECT 85.165 1095.290 85.495 1095.305 ;
        RECT 100.000 1095.290 104.000 1095.480 ;
        RECT 85.165 1094.990 104.000 1095.290 ;
        RECT 85.165 1094.975 85.495 1094.990 ;
        RECT 100.000 1094.880 104.000 1094.990 ;
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 16.625 538.370 16.955 538.385 ;
        RECT -4.800 538.070 16.955 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
        RECT 16.625 538.055 16.955 538.070 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 72.750 1228.320 73.070 1228.380 ;
        RECT 85.170 1228.320 85.490 1228.380 ;
        RECT 72.750 1228.180 85.490 1228.320 ;
        RECT 72.750 1228.120 73.070 1228.180 ;
        RECT 85.170 1228.120 85.490 1228.180 ;
        RECT 16.630 324.260 16.950 324.320 ;
        RECT 72.750 324.260 73.070 324.320 ;
        RECT 16.630 324.120 73.070 324.260 ;
        RECT 16.630 324.060 16.950 324.120 ;
        RECT 72.750 324.060 73.070 324.120 ;
      LAYER via ;
        RECT 72.780 1228.120 73.040 1228.380 ;
        RECT 85.200 1228.120 85.460 1228.380 ;
        RECT 16.660 324.060 16.920 324.320 ;
        RECT 72.780 324.060 73.040 324.320 ;
      LAYER met2 ;
        RECT 72.780 1228.090 73.040 1228.410 ;
        RECT 85.190 1228.235 85.470 1228.605 ;
        RECT 85.200 1228.090 85.460 1228.235 ;
        RECT 72.840 324.350 72.980 1228.090 ;
        RECT 16.660 324.030 16.920 324.350 ;
        RECT 72.780 324.030 73.040 324.350 ;
        RECT 16.720 322.845 16.860 324.030 ;
        RECT 16.650 322.475 16.930 322.845 ;
      LAYER via2 ;
        RECT 85.190 1228.280 85.470 1228.560 ;
        RECT 16.650 322.520 16.930 322.800 ;
      LAYER met3 ;
        RECT 85.165 1228.570 85.495 1228.585 ;
        RECT 100.000 1228.570 104.000 1228.760 ;
        RECT 85.165 1228.270 104.000 1228.570 ;
        RECT 85.165 1228.255 85.495 1228.270 ;
        RECT 100.000 1228.160 104.000 1228.270 ;
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 16.625 322.810 16.955 322.825 ;
        RECT -4.800 322.510 16.955 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
        RECT 16.625 322.495 16.955 322.510 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 58.490 1359.560 58.810 1359.620 ;
        RECT 85.170 1359.560 85.490 1359.620 ;
        RECT 58.490 1359.420 85.490 1359.560 ;
        RECT 58.490 1359.360 58.810 1359.420 ;
        RECT 85.170 1359.360 85.490 1359.420 ;
        RECT 15.710 110.400 16.030 110.460 ;
        RECT 58.490 110.400 58.810 110.460 ;
        RECT 15.710 110.260 58.810 110.400 ;
        RECT 15.710 110.200 16.030 110.260 ;
        RECT 58.490 110.200 58.810 110.260 ;
      LAYER via ;
        RECT 58.520 1359.360 58.780 1359.620 ;
        RECT 85.200 1359.360 85.460 1359.620 ;
        RECT 15.740 110.200 16.000 110.460 ;
        RECT 58.520 110.200 58.780 110.460 ;
      LAYER met2 ;
        RECT 85.190 1360.835 85.470 1361.205 ;
        RECT 85.260 1359.650 85.400 1360.835 ;
        RECT 58.520 1359.330 58.780 1359.650 ;
        RECT 85.200 1359.330 85.460 1359.650 ;
        RECT 58.580 110.490 58.720 1359.330 ;
        RECT 15.740 110.170 16.000 110.490 ;
        RECT 58.520 110.170 58.780 110.490 ;
        RECT 15.800 107.285 15.940 110.170 ;
        RECT 15.730 106.915 16.010 107.285 ;
      LAYER via2 ;
        RECT 85.190 1360.880 85.470 1361.160 ;
        RECT 15.730 106.960 16.010 107.240 ;
      LAYER met3 ;
        RECT 85.165 1361.170 85.495 1361.185 ;
        RECT 100.000 1361.170 104.000 1361.360 ;
        RECT 85.165 1360.870 104.000 1361.170 ;
        RECT 85.165 1360.855 85.495 1360.870 ;
        RECT 100.000 1360.760 104.000 1360.870 ;
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 15.705 107.250 16.035 107.265 ;
        RECT -4.800 106.950 16.035 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
        RECT 15.705 106.935 16.035 106.950 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 849.740 2924.800 850.940 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1084.340 2924.800 1085.540 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1318.940 2924.800 1320.140 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1553.540 2924.800 1554.740 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1788.820 2924.800 1790.020 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2023.420 2924.800 2024.620 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2258.020 2924.800 2259.220 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 674.310 -4.800 674.870 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2.830 23.700 3.150 23.760 ;
        RECT 1945.870 23.700 1946.190 23.760 ;
        RECT 2.830 23.560 1946.190 23.700 ;
        RECT 2.830 23.500 3.150 23.560 ;
        RECT 1945.870 23.500 1946.190 23.560 ;
      LAYER via ;
        RECT 2.860 23.500 3.120 23.760 ;
        RECT 1945.900 23.500 1946.160 23.760 ;
      LAYER met2 ;
        RECT 1952.510 100.370 1952.790 104.000 ;
        RECT 1945.960 100.230 1952.790 100.370 ;
        RECT 1945.960 23.790 1946.100 100.230 ;
        RECT 1952.510 100.000 1952.790 100.230 ;
        RECT 2.860 23.470 3.120 23.790 ;
        RECT 1945.900 23.470 1946.160 23.790 ;
        RECT 2.920 2.400 3.060 23.470 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 8.350 27.440 8.670 27.500 ;
        RECT 1994.170 27.440 1994.490 27.500 ;
        RECT 8.350 27.300 1994.490 27.440 ;
        RECT 8.350 27.240 8.670 27.300 ;
        RECT 1994.170 27.240 1994.490 27.300 ;
      LAYER via ;
        RECT 8.380 27.240 8.640 27.500 ;
        RECT 1994.200 27.240 1994.460 27.500 ;
      LAYER met2 ;
        RECT 1998.050 100.370 1998.330 104.000 ;
        RECT 1994.260 100.230 1998.330 100.370 ;
        RECT 1994.260 27.530 1994.400 100.230 ;
        RECT 1998.050 100.000 1998.330 100.230 ;
        RECT 8.380 27.210 8.640 27.530 ;
        RECT 1994.200 27.210 1994.460 27.530 ;
        RECT 8.440 2.400 8.580 27.210 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 72.290 1490.800 72.610 1490.860 ;
        RECT 85.170 1490.800 85.490 1490.860 ;
        RECT 72.290 1490.660 85.490 1490.800 ;
        RECT 72.290 1490.600 72.610 1490.660 ;
        RECT 85.170 1490.600 85.490 1490.660 ;
        RECT 14.330 17.240 14.650 17.300 ;
        RECT 72.290 17.240 72.610 17.300 ;
        RECT 14.330 17.100 72.610 17.240 ;
        RECT 14.330 17.040 14.650 17.100 ;
        RECT 72.290 17.040 72.610 17.100 ;
      LAYER via ;
        RECT 72.320 1490.600 72.580 1490.860 ;
        RECT 85.200 1490.600 85.460 1490.860 ;
        RECT 14.360 17.040 14.620 17.300 ;
        RECT 72.320 17.040 72.580 17.300 ;
      LAYER met2 ;
        RECT 85.190 1493.435 85.470 1493.805 ;
        RECT 85.260 1490.890 85.400 1493.435 ;
        RECT 72.320 1490.570 72.580 1490.890 ;
        RECT 85.200 1490.570 85.460 1490.890 ;
        RECT 72.380 17.330 72.520 1490.570 ;
        RECT 14.360 17.010 14.620 17.330 ;
        RECT 72.320 17.010 72.580 17.330 ;
        RECT 14.420 2.400 14.560 17.010 ;
        RECT 14.210 -4.800 14.770 2.400 ;
      LAYER via2 ;
        RECT 85.190 1493.480 85.470 1493.760 ;
      LAYER met3 ;
        RECT 85.165 1493.770 85.495 1493.785 ;
        RECT 100.000 1493.770 104.000 1493.960 ;
        RECT 85.165 1493.470 104.000 1493.770 ;
        RECT 85.165 1493.455 85.495 1493.470 ;
        RECT 100.000 1493.360 104.000 1493.470 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 41.010 1621.700 41.330 1621.760 ;
        RECT 85.170 1621.700 85.490 1621.760 ;
        RECT 41.010 1621.560 85.490 1621.700 ;
        RECT 41.010 1621.500 41.330 1621.560 ;
        RECT 85.170 1621.500 85.490 1621.560 ;
        RECT 38.250 17.580 38.570 17.640 ;
        RECT 41.010 17.580 41.330 17.640 ;
        RECT 38.250 17.440 41.330 17.580 ;
        RECT 38.250 17.380 38.570 17.440 ;
        RECT 41.010 17.380 41.330 17.440 ;
      LAYER via ;
        RECT 41.040 1621.500 41.300 1621.760 ;
        RECT 85.200 1621.500 85.460 1621.760 ;
        RECT 38.280 17.380 38.540 17.640 ;
        RECT 41.040 17.380 41.300 17.640 ;
      LAYER met2 ;
        RECT 85.190 1626.715 85.470 1627.085 ;
        RECT 85.260 1621.790 85.400 1626.715 ;
        RECT 41.040 1621.470 41.300 1621.790 ;
        RECT 85.200 1621.470 85.460 1621.790 ;
        RECT 41.100 17.670 41.240 1621.470 ;
        RECT 38.280 17.350 38.540 17.670 ;
        RECT 41.040 17.350 41.300 17.670 ;
        RECT 38.340 2.400 38.480 17.350 ;
        RECT 38.130 -4.800 38.690 2.400 ;
      LAYER via2 ;
        RECT 85.190 1626.760 85.470 1627.040 ;
      LAYER met3 ;
        RECT 85.165 1627.050 85.495 1627.065 ;
        RECT 100.000 1627.050 104.000 1627.240 ;
        RECT 85.165 1626.750 104.000 1627.050 ;
        RECT 85.165 1626.735 85.495 1626.750 ;
        RECT 100.000 1626.640 104.000 1626.750 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 241.110 25.060 241.430 25.120 ;
        RECT 2861.730 25.060 2862.050 25.120 ;
        RECT 241.110 24.920 2862.050 25.060 ;
        RECT 241.110 24.860 241.430 24.920 ;
        RECT 2861.730 24.860 2862.050 24.920 ;
      LAYER via ;
        RECT 241.140 24.860 241.400 25.120 ;
        RECT 2861.760 24.860 2862.020 25.120 ;
      LAYER met2 ;
        RECT 2861.750 1700.155 2862.030 1700.525 ;
        RECT 2861.820 25.150 2861.960 1700.155 ;
        RECT 241.140 24.830 241.400 25.150 ;
        RECT 2861.760 24.830 2862.020 25.150 ;
        RECT 241.200 12.650 241.340 24.830 ;
        RECT 240.740 12.510 241.340 12.650 ;
        RECT 240.740 2.400 240.880 12.510 ;
        RECT 240.530 -4.800 241.090 2.400 ;
      LAYER via2 ;
        RECT 2861.750 1700.200 2862.030 1700.480 ;
      LAYER met3 ;
        RECT 2841.000 1700.490 2845.000 1700.680 ;
        RECT 2861.725 1700.490 2862.055 1700.505 ;
        RECT 2841.000 1700.190 2862.055 1700.490 ;
        RECT 2841.000 1700.080 2845.000 1700.190 ;
        RECT 2861.725 1700.175 2862.055 1700.190 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 258.130 22.000 258.450 22.060 ;
        RECT 2132.170 22.000 2132.490 22.060 ;
        RECT 258.130 21.860 2132.490 22.000 ;
        RECT 258.130 21.800 258.450 21.860 ;
        RECT 2132.170 21.800 2132.490 21.860 ;
      LAYER via ;
        RECT 258.160 21.800 258.420 22.060 ;
        RECT 2132.200 21.800 2132.460 22.060 ;
      LAYER met2 ;
        RECT 2135.130 100.370 2135.410 104.000 ;
        RECT 2132.260 100.230 2135.410 100.370 ;
        RECT 2132.260 22.090 2132.400 100.230 ;
        RECT 2135.130 100.000 2135.410 100.230 ;
        RECT 258.160 21.770 258.420 22.090 ;
        RECT 2132.200 21.770 2132.460 22.090 ;
        RECT 258.220 2.400 258.360 21.770 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 85.630 20.640 85.950 20.700 ;
        RECT 276.070 20.640 276.390 20.700 ;
        RECT 85.630 20.500 276.390 20.640 ;
        RECT 85.630 20.440 85.950 20.500 ;
        RECT 276.070 20.440 276.390 20.500 ;
      LAYER via ;
        RECT 85.660 20.440 85.920 20.700 ;
        RECT 276.100 20.440 276.360 20.700 ;
      LAYER met2 ;
        RECT 85.650 1891.915 85.930 1892.285 ;
        RECT 85.720 20.730 85.860 1891.915 ;
        RECT 85.660 20.410 85.920 20.730 ;
        RECT 276.100 20.410 276.360 20.730 ;
        RECT 276.160 2.400 276.300 20.410 ;
        RECT 275.950 -4.800 276.510 2.400 ;
      LAYER via2 ;
        RECT 85.650 1891.960 85.930 1892.240 ;
      LAYER met3 ;
        RECT 85.625 1892.250 85.955 1892.265 ;
        RECT 100.000 1892.250 104.000 1892.440 ;
        RECT 85.625 1891.950 104.000 1892.250 ;
        RECT 85.625 1891.935 85.955 1891.950 ;
        RECT 100.000 1891.840 104.000 1891.950 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 294.010 22.340 294.330 22.400 ;
        RECT 2180.470 22.340 2180.790 22.400 ;
        RECT 294.010 22.200 2180.790 22.340 ;
        RECT 294.010 22.140 294.330 22.200 ;
        RECT 2180.470 22.140 2180.790 22.200 ;
      LAYER via ;
        RECT 294.040 22.140 294.300 22.400 ;
        RECT 2180.500 22.140 2180.760 22.400 ;
      LAYER met2 ;
        RECT 2181.130 100.370 2181.410 104.000 ;
        RECT 2180.560 100.230 2181.410 100.370 ;
        RECT 2180.560 22.430 2180.700 100.230 ;
        RECT 2181.130 100.000 2181.410 100.230 ;
        RECT 294.040 22.110 294.300 22.430 ;
        RECT 2180.500 22.110 2180.760 22.430 ;
        RECT 294.100 2.400 294.240 22.110 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 311.950 23.020 312.270 23.080 ;
        RECT 2221.870 23.020 2222.190 23.080 ;
        RECT 311.950 22.880 2222.190 23.020 ;
        RECT 311.950 22.820 312.270 22.880 ;
        RECT 2221.870 22.820 2222.190 22.880 ;
      LAYER via ;
        RECT 311.980 22.820 312.240 23.080 ;
        RECT 2221.900 22.820 2222.160 23.080 ;
      LAYER met2 ;
        RECT 2226.670 100.370 2226.950 104.000 ;
        RECT 2221.960 100.230 2226.950 100.370 ;
        RECT 2221.960 23.110 2222.100 100.230 ;
        RECT 2226.670 100.000 2226.950 100.230 ;
        RECT 311.980 22.790 312.240 23.110 ;
        RECT 2221.900 22.790 2222.160 23.110 ;
        RECT 312.040 2.400 312.180 22.790 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 329.890 23.360 330.210 23.420 ;
        RECT 2270.170 23.360 2270.490 23.420 ;
        RECT 329.890 23.220 2270.490 23.360 ;
        RECT 329.890 23.160 330.210 23.220 ;
        RECT 2270.170 23.160 2270.490 23.220 ;
      LAYER via ;
        RECT 329.920 23.160 330.180 23.420 ;
        RECT 2270.200 23.160 2270.460 23.420 ;
      LAYER met2 ;
        RECT 2272.670 100.370 2272.950 104.000 ;
        RECT 2270.260 100.230 2272.950 100.370 ;
        RECT 2270.260 23.450 2270.400 100.230 ;
        RECT 2272.670 100.000 2272.950 100.230 ;
        RECT 329.920 23.130 330.180 23.450 ;
        RECT 2270.200 23.130 2270.460 23.450 ;
        RECT 329.980 2.400 330.120 23.130 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 347.370 25.400 347.690 25.460 ;
        RECT 2861.270 25.400 2861.590 25.460 ;
        RECT 347.370 25.260 2861.590 25.400 ;
        RECT 347.370 25.200 347.690 25.260 ;
        RECT 2861.270 25.200 2861.590 25.260 ;
      LAYER via ;
        RECT 347.400 25.200 347.660 25.460 ;
        RECT 2861.300 25.200 2861.560 25.460 ;
      LAYER met2 ;
        RECT 2861.290 1819.155 2861.570 1819.525 ;
        RECT 2861.360 25.490 2861.500 1819.155 ;
        RECT 347.400 25.170 347.660 25.490 ;
        RECT 2861.300 25.170 2861.560 25.490 ;
        RECT 347.460 2.400 347.600 25.170 ;
        RECT 347.250 -4.800 347.810 2.400 ;
      LAYER via2 ;
        RECT 2861.290 1819.200 2861.570 1819.480 ;
      LAYER met3 ;
        RECT 2841.000 1819.490 2845.000 1819.680 ;
        RECT 2861.265 1819.490 2861.595 1819.505 ;
        RECT 2841.000 1819.190 2861.595 1819.490 ;
        RECT 2841.000 1819.080 2845.000 1819.190 ;
        RECT 2861.265 1819.175 2861.595 1819.190 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1293.610 3430.075 1293.890 3430.445 ;
        RECT 1293.680 3419.450 1293.820 3430.075 ;
        RECT 1295.170 3419.450 1295.450 3420.000 ;
        RECT 1293.680 3419.310 1295.450 3419.450 ;
        RECT 1295.170 3416.000 1295.450 3419.310 ;
        RECT 364.870 17.835 365.150 18.205 ;
        RECT 364.940 16.050 365.080 17.835 ;
        RECT 364.940 15.910 365.540 16.050 ;
        RECT 365.400 2.400 365.540 15.910 ;
        RECT 365.190 -4.800 365.750 2.400 ;
      LAYER via2 ;
        RECT 1293.610 3430.120 1293.890 3430.400 ;
        RECT 364.870 17.880 365.150 18.160 ;
      LAYER met3 ;
        RECT 118.030 3430.410 118.410 3430.420 ;
        RECT 1293.585 3430.410 1293.915 3430.425 ;
        RECT 118.030 3430.110 1293.915 3430.410 ;
        RECT 118.030 3430.100 118.410 3430.110 ;
        RECT 1293.585 3430.095 1293.915 3430.110 ;
        RECT 118.030 18.170 118.410 18.180 ;
        RECT 364.845 18.170 365.175 18.185 ;
        RECT 118.030 17.870 365.175 18.170 ;
        RECT 118.030 17.860 118.410 17.870 ;
        RECT 364.845 17.855 365.175 17.870 ;
      LAYER via3 ;
        RECT 118.060 3430.100 118.380 3430.420 ;
        RECT 118.060 17.860 118.380 18.180 ;
      LAYER met4 ;
        RECT 118.055 3430.095 118.385 3430.425 ;
        RECT 118.070 18.185 118.370 3430.095 ;
        RECT 118.055 17.855 118.385 18.185 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 108.630 3432.540 108.950 3432.600 ;
        RECT 1381.910 3432.540 1382.230 3432.600 ;
        RECT 108.630 3432.400 1382.230 3432.540 ;
        RECT 108.630 3432.340 108.950 3432.400 ;
        RECT 1381.910 3432.340 1382.230 3432.400 ;
        RECT 108.630 20.300 108.950 20.360 ;
        RECT 383.250 20.300 383.570 20.360 ;
        RECT 108.630 20.160 383.570 20.300 ;
        RECT 108.630 20.100 108.950 20.160 ;
        RECT 383.250 20.100 383.570 20.160 ;
      LAYER via ;
        RECT 108.660 3432.340 108.920 3432.600 ;
        RECT 1381.940 3432.340 1382.200 3432.600 ;
        RECT 108.660 20.100 108.920 20.360 ;
        RECT 383.280 20.100 383.540 20.360 ;
      LAYER met2 ;
        RECT 108.660 3432.310 108.920 3432.630 ;
        RECT 1381.940 3432.310 1382.200 3432.630 ;
        RECT 108.720 20.390 108.860 3432.310 ;
        RECT 1382.000 3419.450 1382.140 3432.310 ;
        RECT 1383.490 3419.450 1383.770 3420.000 ;
        RECT 1382.000 3419.310 1383.770 3419.450 ;
        RECT 1383.490 3416.000 1383.770 3419.310 ;
        RECT 108.660 20.070 108.920 20.390 ;
        RECT 383.280 20.070 383.540 20.390 ;
        RECT 383.340 2.400 383.480 20.070 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 401.190 25.740 401.510 25.800 ;
        RECT 2860.810 25.740 2861.130 25.800 ;
        RECT 401.190 25.600 2861.130 25.740 ;
        RECT 401.190 25.540 401.510 25.600 ;
        RECT 2860.810 25.540 2861.130 25.600 ;
      LAYER via ;
        RECT 401.220 25.540 401.480 25.800 ;
        RECT 2860.840 25.540 2861.100 25.800 ;
      LAYER met2 ;
        RECT 2860.830 1937.475 2861.110 1937.845 ;
        RECT 2860.900 25.830 2861.040 1937.475 ;
        RECT 401.220 25.510 401.480 25.830 ;
        RECT 2860.840 25.510 2861.100 25.830 ;
        RECT 401.280 2.400 401.420 25.510 ;
        RECT 401.070 -4.800 401.630 2.400 ;
      LAYER via2 ;
        RECT 2860.830 1937.520 2861.110 1937.800 ;
      LAYER met3 ;
        RECT 2841.000 1937.810 2845.000 1938.000 ;
        RECT 2860.805 1937.810 2861.135 1937.825 ;
        RECT 2841.000 1937.510 2861.135 1937.810 ;
        RECT 2841.000 1937.400 2845.000 1937.510 ;
        RECT 2860.805 1937.495 2861.135 1937.510 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 68.150 1759.740 68.470 1759.800 ;
        RECT 85.170 1759.740 85.490 1759.800 ;
        RECT 68.150 1759.600 85.490 1759.740 ;
        RECT 68.150 1759.540 68.470 1759.600 ;
        RECT 85.170 1759.540 85.490 1759.600 ;
        RECT 62.170 17.920 62.490 17.980 ;
        RECT 68.150 17.920 68.470 17.980 ;
        RECT 62.170 17.780 68.470 17.920 ;
        RECT 62.170 17.720 62.490 17.780 ;
        RECT 68.150 17.720 68.470 17.780 ;
      LAYER via ;
        RECT 68.180 1759.540 68.440 1759.800 ;
        RECT 85.200 1759.540 85.460 1759.800 ;
        RECT 62.200 17.720 62.460 17.980 ;
        RECT 68.180 17.720 68.440 17.980 ;
      LAYER met2 ;
        RECT 68.180 1759.510 68.440 1759.830 ;
        RECT 85.200 1759.685 85.460 1759.830 ;
        RECT 68.240 18.010 68.380 1759.510 ;
        RECT 85.190 1759.315 85.470 1759.685 ;
        RECT 62.200 17.690 62.460 18.010 ;
        RECT 68.180 17.690 68.440 18.010 ;
        RECT 62.260 2.400 62.400 17.690 ;
        RECT 62.050 -4.800 62.610 2.400 ;
      LAYER via2 ;
        RECT 85.190 1759.360 85.470 1759.640 ;
      LAYER met3 ;
        RECT 85.165 1759.650 85.495 1759.665 ;
        RECT 100.000 1759.650 104.000 1759.840 ;
        RECT 85.165 1759.350 104.000 1759.650 ;
        RECT 85.165 1759.335 85.495 1759.350 ;
        RECT 100.000 1759.240 104.000 1759.350 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 419.130 22.680 419.450 22.740 ;
        RECT 2311.570 22.680 2311.890 22.740 ;
        RECT 419.130 22.540 2311.890 22.680 ;
        RECT 419.130 22.480 419.450 22.540 ;
        RECT 2311.570 22.480 2311.890 22.540 ;
      LAYER via ;
        RECT 419.160 22.480 419.420 22.740 ;
        RECT 2311.600 22.480 2311.860 22.740 ;
      LAYER met2 ;
        RECT 2318.210 100.370 2318.490 104.000 ;
        RECT 2311.660 100.230 2318.490 100.370 ;
        RECT 2311.660 22.770 2311.800 100.230 ;
        RECT 2318.210 100.000 2318.490 100.230 ;
        RECT 419.160 22.450 419.420 22.770 ;
        RECT 2311.600 22.450 2311.860 22.770 ;
        RECT 419.220 2.400 419.360 22.450 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 436.610 26.080 436.930 26.140 ;
        RECT 2860.350 26.080 2860.670 26.140 ;
        RECT 436.610 25.940 2860.670 26.080 ;
        RECT 436.610 25.880 436.930 25.940 ;
        RECT 2860.350 25.880 2860.670 25.940 ;
      LAYER via ;
        RECT 436.640 25.880 436.900 26.140 ;
        RECT 2860.380 25.880 2860.640 26.140 ;
      LAYER met2 ;
        RECT 2860.370 2055.795 2860.650 2056.165 ;
        RECT 2860.440 26.170 2860.580 2055.795 ;
        RECT 436.640 25.850 436.900 26.170 ;
        RECT 2860.380 25.850 2860.640 26.170 ;
        RECT 436.700 2.400 436.840 25.850 ;
        RECT 436.490 -4.800 437.050 2.400 ;
      LAYER via2 ;
        RECT 2860.370 2055.840 2860.650 2056.120 ;
      LAYER met3 ;
        RECT 2841.000 2056.130 2845.000 2056.320 ;
        RECT 2860.345 2056.130 2860.675 2056.145 ;
        RECT 2841.000 2055.830 2860.675 2056.130 ;
        RECT 2841.000 2055.720 2845.000 2055.830 ;
        RECT 2860.345 2055.815 2860.675 2055.830 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 86.090 26.420 86.410 26.480 ;
        RECT 454.550 26.420 454.870 26.480 ;
        RECT 86.090 26.280 454.870 26.420 ;
        RECT 86.090 26.220 86.410 26.280 ;
        RECT 454.550 26.220 454.870 26.280 ;
      LAYER via ;
        RECT 86.120 26.220 86.380 26.480 ;
        RECT 454.580 26.220 454.840 26.480 ;
      LAYER met2 ;
        RECT 86.110 2024.515 86.390 2024.885 ;
        RECT 86.180 26.510 86.320 2024.515 ;
        RECT 86.120 26.190 86.380 26.510 ;
        RECT 454.580 26.190 454.840 26.510 ;
        RECT 454.640 2.400 454.780 26.190 ;
        RECT 454.430 -4.800 454.990 2.400 ;
      LAYER via2 ;
        RECT 86.110 2024.560 86.390 2024.840 ;
      LAYER met3 ;
        RECT 86.085 2024.850 86.415 2024.865 ;
        RECT 100.000 2024.850 104.000 2025.040 ;
        RECT 86.085 2024.550 104.000 2024.850 ;
        RECT 86.085 2024.535 86.415 2024.550 ;
        RECT 100.000 2024.440 104.000 2024.550 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 111.850 96.460 112.170 96.520 ;
        RECT 120.590 96.460 120.910 96.520 ;
        RECT 111.850 96.320 120.910 96.460 ;
        RECT 111.850 96.260 112.170 96.320 ;
        RECT 120.590 96.260 120.910 96.320 ;
        RECT 120.590 24.720 120.910 24.780 ;
        RECT 124.270 24.720 124.590 24.780 ;
        RECT 120.590 24.580 124.590 24.720 ;
        RECT 120.590 24.520 120.910 24.580 ;
        RECT 124.270 24.520 124.590 24.580 ;
        RECT 124.270 14.860 124.590 14.920 ;
        RECT 472.490 14.860 472.810 14.920 ;
        RECT 124.270 14.720 472.810 14.860 ;
        RECT 124.270 14.660 124.590 14.720 ;
        RECT 472.490 14.660 472.810 14.720 ;
      LAYER via ;
        RECT 111.880 96.260 112.140 96.520 ;
        RECT 120.620 96.260 120.880 96.520 ;
        RECT 120.620 24.520 120.880 24.780 ;
        RECT 124.300 24.520 124.560 24.780 ;
        RECT 124.300 14.660 124.560 14.920 ;
        RECT 472.520 14.660 472.780 14.920 ;
      LAYER met2 ;
        RECT 1469.330 3418.770 1469.610 3418.885 ;
        RECT 1472.270 3418.770 1472.550 3420.000 ;
        RECT 1469.330 3418.630 1472.550 3418.770 ;
        RECT 1469.330 3418.515 1469.610 3418.630 ;
        RECT 1472.270 3416.000 1472.550 3418.630 ;
        RECT 111.870 3413.755 112.150 3414.125 ;
        RECT 111.940 96.550 112.080 3413.755 ;
        RECT 111.880 96.230 112.140 96.550 ;
        RECT 120.620 96.230 120.880 96.550 ;
        RECT 120.680 24.810 120.820 96.230 ;
        RECT 120.620 24.490 120.880 24.810 ;
        RECT 124.300 24.490 124.560 24.810 ;
        RECT 124.360 14.950 124.500 24.490 ;
        RECT 124.300 14.630 124.560 14.950 ;
        RECT 472.520 14.630 472.780 14.950 ;
        RECT 472.580 2.400 472.720 14.630 ;
        RECT 472.370 -4.800 472.930 2.400 ;
      LAYER via2 ;
        RECT 1469.330 3418.560 1469.610 3418.840 ;
        RECT 111.870 3413.800 112.150 3414.080 ;
      LAYER met3 ;
        RECT 1424.430 3418.850 1424.810 3418.860 ;
        RECT 1469.305 3418.850 1469.635 3418.865 ;
        RECT 1424.430 3418.550 1469.635 3418.850 ;
        RECT 1424.430 3418.540 1424.810 3418.550 ;
        RECT 1469.305 3418.535 1469.635 3418.550 ;
        RECT 111.845 3414.090 112.175 3414.105 ;
        RECT 1424.430 3414.090 1424.810 3414.100 ;
        RECT 111.845 3413.790 1424.810 3414.090 ;
        RECT 111.845 3413.775 112.175 3413.790 ;
        RECT 1424.430 3413.780 1424.810 3413.790 ;
      LAYER via3 ;
        RECT 1424.460 3418.540 1424.780 3418.860 ;
        RECT 1424.460 3413.780 1424.780 3414.100 ;
      LAYER met4 ;
        RECT 1424.455 3418.535 1424.785 3418.865 ;
        RECT 1424.470 3414.105 1424.770 3418.535 ;
        RECT 1424.455 3413.775 1424.785 3414.105 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 111.390 96.800 111.710 96.860 ;
        RECT 111.390 96.660 121.280 96.800 ;
        RECT 111.390 96.600 111.710 96.660 ;
        RECT 121.140 96.460 121.280 96.660 ;
        RECT 124.270 96.460 124.590 96.520 ;
        RECT 121.140 96.320 124.590 96.460 ;
        RECT 124.270 96.260 124.590 96.320 ;
        RECT 124.270 54.980 124.590 55.040 ;
        RECT 144.050 54.980 144.370 55.040 ;
        RECT 124.270 54.840 144.370 54.980 ;
        RECT 124.270 54.780 124.590 54.840 ;
        RECT 144.050 54.780 144.370 54.840 ;
        RECT 144.050 41.720 144.370 41.780 ;
        RECT 144.050 41.580 145.200 41.720 ;
        RECT 144.050 41.520 144.370 41.580 ;
        RECT 145.060 41.380 145.200 41.580 ;
        RECT 165.670 41.380 165.990 41.440 ;
        RECT 145.060 41.240 165.990 41.380 ;
        RECT 165.670 41.180 165.990 41.240 ;
        RECT 165.670 14.520 165.990 14.580 ;
        RECT 490.430 14.520 490.750 14.580 ;
        RECT 165.670 14.380 490.750 14.520 ;
        RECT 165.670 14.320 165.990 14.380 ;
        RECT 490.430 14.320 490.750 14.380 ;
      LAYER via ;
        RECT 111.420 96.600 111.680 96.860 ;
        RECT 124.300 96.260 124.560 96.520 ;
        RECT 124.300 54.780 124.560 55.040 ;
        RECT 144.080 54.780 144.340 55.040 ;
        RECT 144.080 41.520 144.340 41.780 ;
        RECT 165.700 41.180 165.960 41.440 ;
        RECT 165.700 14.320 165.960 14.580 ;
        RECT 490.460 14.320 490.720 14.580 ;
      LAYER met2 ;
        RECT 1559.030 3416.730 1559.310 3416.845 ;
        RECT 1560.590 3416.730 1560.870 3420.000 ;
        RECT 1559.030 3416.590 1560.870 3416.730 ;
        RECT 1559.030 3416.475 1559.310 3416.590 ;
        RECT 1560.590 3416.000 1560.870 3416.590 ;
        RECT 111.410 3413.075 111.690 3413.445 ;
        RECT 111.480 96.890 111.620 3413.075 ;
        RECT 111.420 96.570 111.680 96.890 ;
        RECT 124.300 96.230 124.560 96.550 ;
        RECT 124.360 55.070 124.500 96.230 ;
        RECT 124.300 54.750 124.560 55.070 ;
        RECT 144.080 54.750 144.340 55.070 ;
        RECT 144.140 41.810 144.280 54.750 ;
        RECT 144.080 41.490 144.340 41.810 ;
        RECT 165.700 41.150 165.960 41.470 ;
        RECT 165.760 14.610 165.900 41.150 ;
        RECT 165.700 14.290 165.960 14.610 ;
        RECT 490.460 14.290 490.720 14.610 ;
        RECT 490.520 2.400 490.660 14.290 ;
        RECT 490.310 -4.800 490.870 2.400 ;
      LAYER via2 ;
        RECT 1559.030 3416.520 1559.310 3416.800 ;
        RECT 111.410 3413.120 111.690 3413.400 ;
      LAYER met3 ;
        RECT 1559.005 3416.820 1559.335 3416.825 ;
        RECT 1558.750 3416.810 1559.335 3416.820 ;
        RECT 1558.550 3416.510 1559.335 3416.810 ;
        RECT 1558.750 3416.500 1559.335 3416.510 ;
        RECT 1559.005 3416.495 1559.335 3416.500 ;
        RECT 111.385 3413.410 111.715 3413.425 ;
        RECT 1558.750 3413.410 1559.130 3413.420 ;
        RECT 111.385 3413.110 1559.130 3413.410 ;
        RECT 111.385 3413.095 111.715 3413.110 ;
        RECT 1558.750 3413.100 1559.130 3413.110 ;
      LAYER via3 ;
        RECT 1558.780 3416.500 1559.100 3416.820 ;
        RECT 1558.780 3413.100 1559.100 3413.420 ;
      LAYER met4 ;
        RECT 1558.775 3416.495 1559.105 3416.825 ;
        RECT 1558.790 3413.425 1559.090 3416.495 ;
        RECT 1558.775 3413.095 1559.105 3413.425 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 507.910 26.420 508.230 26.480 ;
        RECT 2859.890 26.420 2860.210 26.480 ;
        RECT 507.910 26.280 2860.210 26.420 ;
        RECT 507.910 26.220 508.230 26.280 ;
        RECT 2859.890 26.220 2860.210 26.280 ;
      LAYER via ;
        RECT 507.940 26.220 508.200 26.480 ;
        RECT 2859.920 26.220 2860.180 26.480 ;
      LAYER met2 ;
        RECT 2859.910 2174.795 2860.190 2175.165 ;
        RECT 2859.980 26.510 2860.120 2174.795 ;
        RECT 507.940 26.190 508.200 26.510 ;
        RECT 2859.920 26.190 2860.180 26.510 ;
        RECT 508.000 2.400 508.140 26.190 ;
        RECT 507.790 -4.800 508.350 2.400 ;
      LAYER via2 ;
        RECT 2859.910 2174.840 2860.190 2175.120 ;
      LAYER met3 ;
        RECT 2841.000 2175.130 2845.000 2175.320 ;
        RECT 2859.885 2175.130 2860.215 2175.145 ;
        RECT 2841.000 2174.830 2860.215 2175.130 ;
        RECT 2841.000 2174.720 2845.000 2174.830 ;
        RECT 2859.885 2174.815 2860.215 2174.830 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 112.770 48.180 113.090 48.240 ;
        RECT 124.270 48.180 124.590 48.240 ;
        RECT 112.770 48.040 124.590 48.180 ;
        RECT 112.770 47.980 113.090 48.040 ;
        RECT 124.270 47.980 124.590 48.040 ;
        RECT 124.270 25.400 124.590 25.460 ;
        RECT 248.010 25.400 248.330 25.460 ;
        RECT 124.270 25.260 248.330 25.400 ;
        RECT 124.270 25.200 124.590 25.260 ;
        RECT 248.010 25.200 248.330 25.260 ;
        RECT 525.850 14.180 526.170 14.240 ;
        RECT 255.920 14.040 526.170 14.180 ;
        RECT 248.010 13.840 248.330 13.900 ;
        RECT 255.920 13.840 256.060 14.040 ;
        RECT 525.850 13.980 526.170 14.040 ;
        RECT 248.010 13.700 256.060 13.840 ;
        RECT 248.010 13.640 248.330 13.700 ;
      LAYER via ;
        RECT 112.800 47.980 113.060 48.240 ;
        RECT 124.300 47.980 124.560 48.240 ;
        RECT 124.300 25.200 124.560 25.460 ;
        RECT 248.040 25.200 248.300 25.460 ;
        RECT 248.040 13.640 248.300 13.900 ;
        RECT 525.880 13.980 526.140 14.240 ;
      LAYER met2 ;
        RECT 1648.730 3417.410 1649.010 3417.525 ;
        RECT 1649.370 3417.410 1649.650 3420.000 ;
        RECT 1648.730 3417.270 1649.650 3417.410 ;
        RECT 1648.730 3417.155 1649.010 3417.270 ;
        RECT 1649.370 3416.000 1649.650 3417.270 ;
        RECT 112.790 3412.395 113.070 3412.765 ;
        RECT 112.860 48.270 113.000 3412.395 ;
        RECT 112.800 47.950 113.060 48.270 ;
        RECT 124.300 47.950 124.560 48.270 ;
        RECT 124.360 25.490 124.500 47.950 ;
        RECT 124.300 25.170 124.560 25.490 ;
        RECT 248.040 25.170 248.300 25.490 ;
        RECT 248.100 13.930 248.240 25.170 ;
        RECT 525.880 13.950 526.140 14.270 ;
        RECT 248.040 13.610 248.300 13.930 ;
        RECT 525.940 2.400 526.080 13.950 ;
        RECT 525.730 -4.800 526.290 2.400 ;
      LAYER via2 ;
        RECT 1648.730 3417.200 1649.010 3417.480 ;
        RECT 112.790 3412.440 113.070 3412.720 ;
      LAYER met3 ;
        RECT 1615.790 3417.490 1616.170 3417.500 ;
        RECT 1648.705 3417.490 1649.035 3417.505 ;
        RECT 1615.790 3417.190 1649.035 3417.490 ;
        RECT 1615.790 3417.180 1616.170 3417.190 ;
        RECT 1648.705 3417.175 1649.035 3417.190 ;
        RECT 112.765 3412.730 113.095 3412.745 ;
        RECT 1615.790 3412.730 1616.170 3412.740 ;
        RECT 112.765 3412.430 1616.170 3412.730 ;
        RECT 112.765 3412.415 113.095 3412.430 ;
        RECT 1615.790 3412.420 1616.170 3412.430 ;
      LAYER via3 ;
        RECT 1615.820 3417.180 1616.140 3417.500 ;
        RECT 1615.820 3412.420 1616.140 3412.740 ;
      LAYER met4 ;
        RECT 1615.815 3417.175 1616.145 3417.505 ;
        RECT 1615.830 3412.745 1616.130 3417.175 ;
        RECT 1615.815 3412.415 1616.145 3412.745 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 543.790 26.760 544.110 26.820 ;
        RECT 2859.430 26.760 2859.750 26.820 ;
        RECT 543.790 26.620 2859.750 26.760 ;
        RECT 543.790 26.560 544.110 26.620 ;
        RECT 2859.430 26.560 2859.750 26.620 ;
      LAYER via ;
        RECT 543.820 26.560 544.080 26.820 ;
        RECT 2859.460 26.560 2859.720 26.820 ;
      LAYER met2 ;
        RECT 2859.450 2293.115 2859.730 2293.485 ;
        RECT 2859.520 26.850 2859.660 2293.115 ;
        RECT 543.820 26.530 544.080 26.850 ;
        RECT 2859.460 26.530 2859.720 26.850 ;
        RECT 543.880 2.400 544.020 26.530 ;
        RECT 543.670 -4.800 544.230 2.400 ;
      LAYER via2 ;
        RECT 2859.450 2293.160 2859.730 2293.440 ;
      LAYER met3 ;
        RECT 2841.000 2293.450 2845.000 2293.640 ;
        RECT 2859.425 2293.450 2859.755 2293.465 ;
        RECT 2841.000 2293.150 2859.755 2293.450 ;
        RECT 2841.000 2293.040 2845.000 2293.150 ;
        RECT 2859.425 2293.135 2859.755 2293.150 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 561.730 21.660 562.050 21.720 ;
        RECT 2359.870 21.660 2360.190 21.720 ;
        RECT 561.730 21.520 2360.190 21.660 ;
        RECT 561.730 21.460 562.050 21.520 ;
        RECT 2359.870 21.460 2360.190 21.520 ;
      LAYER via ;
        RECT 561.760 21.460 562.020 21.720 ;
        RECT 2359.900 21.460 2360.160 21.720 ;
      LAYER met2 ;
        RECT 2364.210 100.370 2364.490 104.000 ;
        RECT 2359.960 100.230 2364.490 100.370 ;
        RECT 2359.960 21.750 2360.100 100.230 ;
        RECT 2364.210 100.000 2364.490 100.230 ;
        RECT 561.760 21.430 562.020 21.750 ;
        RECT 2359.900 21.430 2360.160 21.750 ;
        RECT 561.820 2.400 561.960 21.430 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 580.130 27.100 580.450 27.160 ;
        RECT 2858.970 27.100 2859.290 27.160 ;
        RECT 580.130 26.960 2859.290 27.100 ;
        RECT 580.130 26.900 580.450 26.960 ;
        RECT 2858.970 26.900 2859.290 26.960 ;
      LAYER via ;
        RECT 580.160 26.900 580.420 27.160 ;
        RECT 2859.000 26.900 2859.260 27.160 ;
      LAYER met2 ;
        RECT 2858.990 2411.435 2859.270 2411.805 ;
        RECT 2859.060 27.190 2859.200 2411.435 ;
        RECT 580.160 26.870 580.420 27.190 ;
        RECT 2859.000 26.870 2859.260 27.190 ;
        RECT 580.220 14.010 580.360 26.870 ;
        RECT 579.760 13.870 580.360 14.010 ;
        RECT 579.760 2.400 579.900 13.870 ;
        RECT 579.550 -4.800 580.110 2.400 ;
      LAYER via2 ;
        RECT 2858.990 2411.480 2859.270 2411.760 ;
      LAYER met3 ;
        RECT 2841.000 2411.770 2845.000 2411.960 ;
        RECT 2858.965 2411.770 2859.295 2411.785 ;
        RECT 2841.000 2411.470 2859.295 2411.770 ;
        RECT 2841.000 2411.360 2845.000 2411.470 ;
        RECT 2858.965 2411.455 2859.295 2411.470 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 86.090 24.040 86.410 24.100 ;
        RECT 2863.110 24.040 2863.430 24.100 ;
        RECT 86.090 23.900 2863.430 24.040 ;
        RECT 86.090 23.840 86.410 23.900 ;
        RECT 2863.110 23.840 2863.430 23.900 ;
      LAYER via ;
        RECT 86.120 23.840 86.380 24.100 ;
        RECT 2863.140 23.840 2863.400 24.100 ;
      LAYER met2 ;
        RECT 2863.130 1344.515 2863.410 1344.885 ;
        RECT 2863.200 24.130 2863.340 1344.515 ;
        RECT 86.120 23.810 86.380 24.130 ;
        RECT 2863.140 23.810 2863.400 24.130 ;
        RECT 86.180 2.400 86.320 23.810 ;
        RECT 85.970 -4.800 86.530 2.400 ;
      LAYER via2 ;
        RECT 2863.130 1344.560 2863.410 1344.840 ;
      LAYER met3 ;
        RECT 2841.000 1344.850 2845.000 1345.040 ;
        RECT 2863.105 1344.850 2863.435 1344.865 ;
        RECT 2841.000 1344.550 2863.435 1344.850 ;
        RECT 2841.000 1344.440 2845.000 1344.550 ;
        RECT 2863.105 1344.535 2863.435 1344.550 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 112.310 90.000 112.630 90.060 ;
        RECT 112.310 89.860 117.600 90.000 ;
        RECT 112.310 89.800 112.630 89.860 ;
        RECT 117.460 89.660 117.600 89.860 ;
        RECT 130.710 89.660 131.030 89.720 ;
        RECT 117.460 89.520 131.030 89.660 ;
        RECT 130.710 89.460 131.030 89.520 ;
        RECT 131.170 54.640 131.490 54.700 ;
        RECT 138.530 54.640 138.850 54.700 ;
        RECT 131.170 54.500 138.850 54.640 ;
        RECT 131.170 54.440 131.490 54.500 ;
        RECT 138.530 54.440 138.850 54.500 ;
        RECT 138.530 41.040 138.850 41.100 ;
        RECT 145.430 41.040 145.750 41.100 ;
        RECT 138.530 40.900 145.750 41.040 ;
        RECT 138.530 40.840 138.850 40.900 ;
        RECT 145.430 40.840 145.750 40.900 ;
        RECT 145.430 21.320 145.750 21.380 ;
        RECT 597.150 21.320 597.470 21.380 ;
        RECT 145.430 21.180 597.470 21.320 ;
        RECT 145.430 21.120 145.750 21.180 ;
        RECT 597.150 21.120 597.470 21.180 ;
      LAYER via ;
        RECT 112.340 89.800 112.600 90.060 ;
        RECT 130.740 89.460 131.000 89.720 ;
        RECT 131.200 54.440 131.460 54.700 ;
        RECT 138.560 54.440 138.820 54.700 ;
        RECT 138.560 40.840 138.820 41.100 ;
        RECT 145.460 40.840 145.720 41.100 ;
        RECT 145.460 21.120 145.720 21.380 ;
        RECT 597.180 21.120 597.440 21.380 ;
      LAYER met2 ;
        RECT 1736.130 3430.075 1736.410 3430.445 ;
        RECT 1736.200 3419.450 1736.340 3430.075 ;
        RECT 1737.690 3419.450 1737.970 3420.000 ;
        RECT 1736.200 3419.310 1737.970 3419.450 ;
        RECT 1737.690 3416.000 1737.970 3419.310 ;
        RECT 112.330 3411.715 112.610 3412.085 ;
        RECT 112.400 90.090 112.540 3411.715 ;
        RECT 112.340 89.770 112.600 90.090 ;
        RECT 130.740 89.430 131.000 89.750 ;
        RECT 130.800 75.890 130.940 89.430 ;
        RECT 130.800 75.750 131.400 75.890 ;
        RECT 131.260 54.730 131.400 75.750 ;
        RECT 131.200 54.410 131.460 54.730 ;
        RECT 138.560 54.410 138.820 54.730 ;
        RECT 138.620 41.130 138.760 54.410 ;
        RECT 138.560 40.810 138.820 41.130 ;
        RECT 145.460 40.810 145.720 41.130 ;
        RECT 145.520 21.410 145.660 40.810 ;
        RECT 145.460 21.090 145.720 21.410 ;
        RECT 597.180 21.090 597.440 21.410 ;
        RECT 597.240 2.400 597.380 21.090 ;
        RECT 597.030 -4.800 597.590 2.400 ;
      LAYER via2 ;
        RECT 1736.130 3430.120 1736.410 3430.400 ;
        RECT 112.330 3411.760 112.610 3412.040 ;
      LAYER met3 ;
        RECT 1686.630 3430.410 1687.010 3430.420 ;
        RECT 1736.105 3430.410 1736.435 3430.425 ;
        RECT 1686.630 3430.110 1736.435 3430.410 ;
        RECT 1686.630 3430.100 1687.010 3430.110 ;
        RECT 1736.105 3430.095 1736.435 3430.110 ;
        RECT 112.305 3412.050 112.635 3412.065 ;
        RECT 1686.630 3412.050 1687.010 3412.060 ;
        RECT 112.305 3411.750 1687.010 3412.050 ;
        RECT 112.305 3411.735 112.635 3411.750 ;
        RECT 1686.630 3411.740 1687.010 3411.750 ;
      LAYER via3 ;
        RECT 1686.660 3430.100 1686.980 3430.420 ;
        RECT 1686.660 3411.740 1686.980 3412.060 ;
      LAYER met4 ;
        RECT 1686.655 3430.095 1686.985 3430.425 ;
        RECT 1686.670 3412.065 1686.970 3430.095 ;
        RECT 1686.655 3411.735 1686.985 3412.065 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 615.090 31.860 615.410 31.920 ;
        RECT 2858.510 31.860 2858.830 31.920 ;
        RECT 615.090 31.720 2858.830 31.860 ;
        RECT 615.090 31.660 615.410 31.720 ;
        RECT 2858.510 31.660 2858.830 31.720 ;
      LAYER via ;
        RECT 615.120 31.660 615.380 31.920 ;
        RECT 2858.540 31.660 2858.800 31.920 ;
      LAYER met2 ;
        RECT 2858.530 2530.435 2858.810 2530.805 ;
        RECT 2858.600 31.950 2858.740 2530.435 ;
        RECT 615.120 31.630 615.380 31.950 ;
        RECT 2858.540 31.630 2858.800 31.950 ;
        RECT 615.180 2.400 615.320 31.630 ;
        RECT 614.970 -4.800 615.530 2.400 ;
      LAYER via2 ;
        RECT 2858.530 2530.480 2858.810 2530.760 ;
      LAYER met3 ;
        RECT 2841.000 2530.770 2845.000 2530.960 ;
        RECT 2858.505 2530.770 2858.835 2530.785 ;
        RECT 2841.000 2530.470 2858.835 2530.770 ;
        RECT 2841.000 2530.360 2845.000 2530.470 ;
        RECT 2858.505 2530.455 2858.835 2530.470 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 109.550 24.380 109.870 24.440 ;
        RECT 2862.650 24.380 2862.970 24.440 ;
        RECT 109.550 24.240 2862.970 24.380 ;
        RECT 109.550 24.180 109.870 24.240 ;
        RECT 2862.650 24.180 2862.970 24.240 ;
      LAYER via ;
        RECT 109.580 24.180 109.840 24.440 ;
        RECT 2862.680 24.180 2862.940 24.440 ;
      LAYER met2 ;
        RECT 2862.670 1462.835 2862.950 1463.205 ;
        RECT 2862.740 24.470 2862.880 1462.835 ;
        RECT 109.580 24.150 109.840 24.470 ;
        RECT 2862.680 24.150 2862.940 24.470 ;
        RECT 109.640 2.400 109.780 24.150 ;
        RECT 109.430 -4.800 109.990 2.400 ;
      LAYER via2 ;
        RECT 2862.670 1462.880 2862.950 1463.160 ;
      LAYER met3 ;
        RECT 2841.000 1463.170 2845.000 1463.360 ;
        RECT 2862.645 1463.170 2862.975 1463.185 ;
        RECT 2841.000 1462.870 2862.975 1463.170 ;
        RECT 2841.000 1462.760 2845.000 1462.870 ;
        RECT 2862.645 1462.855 2862.975 1462.870 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 133.470 24.720 133.790 24.780 ;
        RECT 2862.190 24.720 2862.510 24.780 ;
        RECT 133.470 24.580 2862.510 24.720 ;
        RECT 133.470 24.520 133.790 24.580 ;
        RECT 2862.190 24.520 2862.510 24.580 ;
      LAYER via ;
        RECT 133.500 24.520 133.760 24.780 ;
        RECT 2862.220 24.520 2862.480 24.780 ;
      LAYER met2 ;
        RECT 2862.210 1581.835 2862.490 1582.205 ;
        RECT 2862.280 24.810 2862.420 1581.835 ;
        RECT 133.500 24.490 133.760 24.810 ;
        RECT 2862.220 24.490 2862.480 24.810 ;
        RECT 133.560 2.400 133.700 24.490 ;
        RECT 133.350 -4.800 133.910 2.400 ;
      LAYER via2 ;
        RECT 2862.210 1581.880 2862.490 1582.160 ;
      LAYER met3 ;
        RECT 2841.000 1582.170 2845.000 1582.360 ;
        RECT 2862.185 1582.170 2862.515 1582.185 ;
        RECT 2841.000 1581.870 2862.515 1582.170 ;
        RECT 2841.000 1581.760 2845.000 1581.870 ;
        RECT 2862.185 1581.855 2862.515 1581.870 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 107.710 3432.880 108.030 3432.940 ;
        RECT 1028.170 3432.880 1028.490 3432.940 ;
        RECT 107.710 3432.740 1028.490 3432.880 ;
        RECT 107.710 3432.680 108.030 3432.740 ;
        RECT 1028.170 3432.680 1028.490 3432.740 ;
        RECT 107.710 18.260 108.030 18.320 ;
        RECT 107.710 18.120 124.500 18.260 ;
        RECT 107.710 18.060 108.030 18.120 ;
        RECT 124.360 17.920 124.500 18.120 ;
        RECT 151.410 17.920 151.730 17.980 ;
        RECT 124.360 17.780 151.730 17.920 ;
        RECT 151.410 17.720 151.730 17.780 ;
      LAYER via ;
        RECT 107.740 3432.680 108.000 3432.940 ;
        RECT 1028.200 3432.680 1028.460 3432.940 ;
        RECT 107.740 18.060 108.000 18.320 ;
        RECT 151.440 17.720 151.700 17.980 ;
      LAYER met2 ;
        RECT 107.740 3432.650 108.000 3432.970 ;
        RECT 1028.200 3432.650 1028.460 3432.970 ;
        RECT 107.800 18.350 107.940 3432.650 ;
        RECT 1028.260 3419.450 1028.400 3432.650 ;
        RECT 1029.290 3419.450 1029.570 3420.000 ;
        RECT 1028.260 3419.310 1029.570 3419.450 ;
        RECT 1029.290 3416.000 1029.570 3419.310 ;
        RECT 107.740 18.030 108.000 18.350 ;
        RECT 151.440 17.690 151.700 18.010 ;
        RECT 151.500 2.400 151.640 17.690 ;
        RECT 151.290 -4.800 151.850 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 172.110 87.280 172.430 87.340 ;
        RECT 2042.470 87.280 2042.790 87.340 ;
        RECT 172.110 87.140 2042.790 87.280 ;
        RECT 172.110 87.080 172.430 87.140 ;
        RECT 2042.470 87.080 2042.790 87.140 ;
        RECT 169.350 17.920 169.670 17.980 ;
        RECT 172.110 17.920 172.430 17.980 ;
        RECT 169.350 17.780 172.430 17.920 ;
        RECT 169.350 17.720 169.670 17.780 ;
        RECT 172.110 17.720 172.430 17.780 ;
      LAYER via ;
        RECT 172.140 87.080 172.400 87.340 ;
        RECT 2042.500 87.080 2042.760 87.340 ;
        RECT 169.380 17.720 169.640 17.980 ;
        RECT 172.140 17.720 172.400 17.980 ;
      LAYER met2 ;
        RECT 2043.590 100.370 2043.870 104.000 ;
        RECT 2042.560 100.230 2043.870 100.370 ;
        RECT 2042.560 87.370 2042.700 100.230 ;
        RECT 2043.590 100.000 2043.870 100.230 ;
        RECT 172.140 87.050 172.400 87.370 ;
        RECT 2042.500 87.050 2042.760 87.370 ;
        RECT 172.200 18.010 172.340 87.050 ;
        RECT 169.380 17.690 169.640 18.010 ;
        RECT 172.140 17.690 172.400 18.010 ;
        RECT 169.440 2.400 169.580 17.690 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1117.890 3431.435 1118.170 3431.805 ;
        RECT 1117.960 3420.000 1118.100 3431.435 ;
        RECT 1117.960 3419.310 1118.350 3420.000 ;
        RECT 1118.070 3416.000 1118.350 3419.310 ;
        RECT 186.850 16.475 187.130 16.845 ;
        RECT 186.920 2.400 187.060 16.475 ;
        RECT 186.710 -4.800 187.270 2.400 ;
      LAYER via2 ;
        RECT 1117.890 3431.480 1118.170 3431.760 ;
        RECT 186.850 16.520 187.130 16.800 ;
      LAYER met3 ;
        RECT 116.190 3431.770 116.570 3431.780 ;
        RECT 1117.865 3431.770 1118.195 3431.785 ;
        RECT 116.190 3431.470 1118.195 3431.770 ;
        RECT 116.190 3431.460 116.570 3431.470 ;
        RECT 1117.865 3431.455 1118.195 3431.470 ;
        RECT 116.190 16.810 116.570 16.820 ;
        RECT 186.825 16.810 187.155 16.825 ;
        RECT 116.190 16.510 187.155 16.810 ;
        RECT 116.190 16.500 116.570 16.510 ;
        RECT 186.825 16.495 187.155 16.510 ;
      LAYER via3 ;
        RECT 116.220 3431.460 116.540 3431.780 ;
        RECT 116.220 16.500 116.540 16.820 ;
      LAYER met4 ;
        RECT 116.215 3431.455 116.545 3431.785 ;
        RECT 116.230 16.825 116.530 3431.455 ;
        RECT 116.215 16.495 116.545 16.825 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 206.610 86.940 206.930 87.000 ;
        RECT 2088.010 86.940 2088.330 87.000 ;
        RECT 206.610 86.800 2088.330 86.940 ;
        RECT 206.610 86.740 206.930 86.800 ;
        RECT 2088.010 86.740 2088.330 86.800 ;
      LAYER via ;
        RECT 206.640 86.740 206.900 87.000 ;
        RECT 2088.040 86.740 2088.300 87.000 ;
      LAYER met2 ;
        RECT 2089.590 100.370 2089.870 104.000 ;
        RECT 2088.100 100.230 2089.870 100.370 ;
        RECT 2088.100 87.030 2088.240 100.230 ;
        RECT 2089.590 100.000 2089.870 100.230 ;
        RECT 206.640 86.710 206.900 87.030 ;
        RECT 2088.040 86.710 2088.300 87.030 ;
        RECT 206.700 17.410 206.840 86.710 ;
        RECT 204.860 17.270 206.840 17.410 ;
        RECT 204.860 2.400 205.000 17.270 ;
        RECT 204.650 -4.800 205.210 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1204.830 3430.755 1205.110 3431.125 ;
        RECT 1204.900 3419.450 1205.040 3430.755 ;
        RECT 1206.390 3419.450 1206.670 3420.000 ;
        RECT 1204.900 3419.310 1206.670 3419.450 ;
        RECT 1206.390 3416.000 1206.670 3419.310 ;
        RECT 222.730 19.195 223.010 19.565 ;
        RECT 222.800 2.400 222.940 19.195 ;
        RECT 222.590 -4.800 223.150 2.400 ;
      LAYER via2 ;
        RECT 1204.830 3430.800 1205.110 3431.080 ;
        RECT 222.730 19.240 223.010 19.520 ;
      LAYER met3 ;
        RECT 115.270 3431.090 115.650 3431.100 ;
        RECT 1204.805 3431.090 1205.135 3431.105 ;
        RECT 115.270 3430.790 1205.135 3431.090 ;
        RECT 115.270 3430.780 115.650 3430.790 ;
        RECT 1204.805 3430.775 1205.135 3430.790 ;
        RECT 115.270 19.530 115.650 19.540 ;
        RECT 222.705 19.530 223.035 19.545 ;
        RECT 115.270 19.230 223.035 19.530 ;
        RECT 115.270 19.220 115.650 19.230 ;
        RECT 222.705 19.215 223.035 19.230 ;
      LAYER via3 ;
        RECT 115.300 3430.780 115.620 3431.100 ;
        RECT 115.300 19.220 115.620 19.540 ;
      LAYER met4 ;
        RECT 115.295 3430.775 115.625 3431.105 ;
        RECT 115.310 19.545 115.610 3430.775 ;
        RECT 115.295 19.215 115.625 19.545 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 20.310 30.840 20.630 30.900 ;
        RECT 2858.050 30.840 2858.370 30.900 ;
        RECT 20.310 30.700 2858.370 30.840 ;
        RECT 20.310 30.640 20.630 30.700 ;
        RECT 2858.050 30.640 2858.370 30.700 ;
      LAYER via ;
        RECT 20.340 30.640 20.600 30.900 ;
        RECT 2858.080 30.640 2858.340 30.900 ;
      LAYER met2 ;
        RECT 2858.070 2648.755 2858.350 2649.125 ;
        RECT 2858.140 30.930 2858.280 2648.755 ;
        RECT 20.340 30.610 20.600 30.930 ;
        RECT 2858.080 30.610 2858.340 30.930 ;
        RECT 20.400 2.400 20.540 30.610 ;
        RECT 20.190 -4.800 20.750 2.400 ;
      LAYER via2 ;
        RECT 2858.070 2648.800 2858.350 2649.080 ;
      LAYER met3 ;
        RECT 2841.000 2649.090 2845.000 2649.280 ;
        RECT 2858.045 2649.090 2858.375 2649.105 ;
        RECT 2841.000 2648.790 2858.375 2649.090 ;
        RECT 2841.000 2648.680 2845.000 2648.790 ;
        RECT 2858.045 2648.775 2858.375 2648.790 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 47.910 3432.200 48.230 3432.260 ;
        RECT 1824.890 3432.200 1825.210 3432.260 ;
        RECT 47.910 3432.060 1825.210 3432.200 ;
        RECT 47.910 3432.000 48.230 3432.060 ;
        RECT 1824.890 3432.000 1825.210 3432.060 ;
        RECT 44.230 17.580 44.550 17.640 ;
        RECT 47.910 17.580 48.230 17.640 ;
        RECT 44.230 17.440 48.230 17.580 ;
        RECT 44.230 17.380 44.550 17.440 ;
        RECT 47.910 17.380 48.230 17.440 ;
      LAYER via ;
        RECT 47.940 3432.000 48.200 3432.260 ;
        RECT 1824.920 3432.000 1825.180 3432.260 ;
        RECT 44.260 17.380 44.520 17.640 ;
        RECT 47.940 17.380 48.200 17.640 ;
      LAYER met2 ;
        RECT 47.940 3431.970 48.200 3432.290 ;
        RECT 1824.920 3431.970 1825.180 3432.290 ;
        RECT 48.000 17.670 48.140 3431.970 ;
        RECT 1824.980 3419.450 1825.120 3431.970 ;
        RECT 1826.470 3419.450 1826.750 3420.000 ;
        RECT 1824.980 3419.310 1826.750 3419.450 ;
        RECT 1826.470 3416.000 1826.750 3419.310 ;
        RECT 44.260 17.350 44.520 17.670 ;
        RECT 47.940 17.350 48.200 17.670 ;
        RECT 44.320 2.400 44.460 17.350 ;
        RECT 44.110 -4.800 44.670 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 107.250 3430.840 107.570 3430.900 ;
        RECT 2090.770 3430.840 2091.090 3430.900 ;
        RECT 107.250 3430.700 2091.090 3430.840 ;
        RECT 107.250 3430.640 107.570 3430.700 ;
        RECT 2090.770 3430.640 2091.090 3430.700 ;
        RECT 107.250 14.180 107.570 14.240 ;
        RECT 246.630 14.180 246.950 14.240 ;
        RECT 107.250 14.040 246.950 14.180 ;
        RECT 107.250 13.980 107.570 14.040 ;
        RECT 246.630 13.980 246.950 14.040 ;
      LAYER via ;
        RECT 107.280 3430.640 107.540 3430.900 ;
        RECT 2090.800 3430.640 2091.060 3430.900 ;
        RECT 107.280 13.980 107.540 14.240 ;
        RECT 246.660 13.980 246.920 14.240 ;
      LAYER met2 ;
        RECT 107.280 3430.610 107.540 3430.930 ;
        RECT 2090.800 3430.610 2091.060 3430.930 ;
        RECT 107.340 14.270 107.480 3430.610 ;
        RECT 2090.860 3419.450 2091.000 3430.610 ;
        RECT 2091.890 3419.450 2092.170 3420.000 ;
        RECT 2090.860 3419.310 2092.170 3419.450 ;
        RECT 2091.890 3416.000 2092.170 3419.310 ;
        RECT 107.280 13.950 107.540 14.270 ;
        RECT 246.660 13.950 246.920 14.270 ;
        RECT 246.720 2.400 246.860 13.950 ;
        RECT 246.510 -4.800 247.070 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 109.550 3430.500 109.870 3430.560 ;
        RECT 2180.470 3430.500 2180.790 3430.560 ;
        RECT 109.550 3430.360 2180.790 3430.500 ;
        RECT 109.550 3430.300 109.870 3430.360 ;
        RECT 2180.470 3430.300 2180.790 3430.360 ;
        RECT 110.010 16.220 110.330 16.280 ;
        RECT 264.110 16.220 264.430 16.280 ;
        RECT 110.010 16.080 264.430 16.220 ;
        RECT 110.010 16.020 110.330 16.080 ;
        RECT 264.110 16.020 264.430 16.080 ;
      LAYER via ;
        RECT 109.580 3430.300 109.840 3430.560 ;
        RECT 2180.500 3430.300 2180.760 3430.560 ;
        RECT 110.040 16.020 110.300 16.280 ;
        RECT 264.140 16.020 264.400 16.280 ;
      LAYER met2 ;
        RECT 109.580 3430.270 109.840 3430.590 ;
        RECT 2180.500 3430.270 2180.760 3430.590 ;
        RECT 109.640 25.570 109.780 3430.270 ;
        RECT 2180.560 3420.000 2180.700 3430.270 ;
        RECT 2180.560 3419.310 2180.950 3420.000 ;
        RECT 2180.670 3416.000 2180.950 3419.310 ;
        RECT 109.640 25.430 110.240 25.570 ;
        RECT 110.100 16.310 110.240 25.430 ;
        RECT 110.040 15.990 110.300 16.310 ;
        RECT 264.140 15.990 264.400 16.310 ;
        RECT 264.200 2.400 264.340 15.990 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 128.025 15.725 128.195 16.575 ;
      LAYER mcon ;
        RECT 128.025 16.405 128.195 16.575 ;
      LAYER met1 ;
        RECT 127.965 16.560 128.255 16.605 ;
        RECT 282.050 16.560 282.370 16.620 ;
        RECT 127.965 16.420 282.370 16.560 ;
        RECT 127.965 16.375 128.255 16.420 ;
        RECT 282.050 16.360 282.370 16.420 ;
        RECT 96.210 15.880 96.530 15.940 ;
        RECT 127.965 15.880 128.255 15.925 ;
        RECT 96.210 15.740 128.255 15.880 ;
        RECT 96.210 15.680 96.530 15.740 ;
        RECT 127.965 15.695 128.255 15.740 ;
      LAYER via ;
        RECT 282.080 16.360 282.340 16.620 ;
        RECT 96.240 15.680 96.500 15.940 ;
      LAYER met2 ;
        RECT 96.230 2290.395 96.510 2290.765 ;
        RECT 96.300 15.970 96.440 2290.395 ;
        RECT 282.080 16.330 282.340 16.650 ;
        RECT 96.240 15.650 96.500 15.970 ;
        RECT 282.140 2.400 282.280 16.330 ;
        RECT 281.930 -4.800 282.490 2.400 ;
      LAYER via2 ;
        RECT 96.230 2290.440 96.510 2290.720 ;
      LAYER met3 ;
        RECT 96.205 2290.730 96.535 2290.745 ;
        RECT 100.000 2290.730 104.000 2290.920 ;
        RECT 96.205 2290.430 104.000 2290.730 ;
        RECT 96.205 2290.415 96.535 2290.430 ;
        RECT 100.000 2290.320 104.000 2290.430 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 106.330 3430.160 106.650 3430.220 ;
        RECT 2267.410 3430.160 2267.730 3430.220 ;
        RECT 106.330 3430.020 2267.730 3430.160 ;
        RECT 106.330 3429.960 106.650 3430.020 ;
        RECT 2267.410 3429.960 2267.730 3430.020 ;
        RECT 106.330 16.900 106.650 16.960 ;
        RECT 299.990 16.900 300.310 16.960 ;
        RECT 106.330 16.760 300.310 16.900 ;
        RECT 106.330 16.700 106.650 16.760 ;
        RECT 299.990 16.700 300.310 16.760 ;
      LAYER via ;
        RECT 106.360 3429.960 106.620 3430.220 ;
        RECT 2267.440 3429.960 2267.700 3430.220 ;
        RECT 106.360 16.700 106.620 16.960 ;
        RECT 300.020 16.700 300.280 16.960 ;
      LAYER met2 ;
        RECT 106.360 3429.930 106.620 3430.250 ;
        RECT 2267.440 3429.930 2267.700 3430.250 ;
        RECT 106.420 16.990 106.560 3429.930 ;
        RECT 2267.500 3419.450 2267.640 3429.930 ;
        RECT 2268.990 3419.450 2269.270 3420.000 ;
        RECT 2267.500 3419.310 2269.270 3419.450 ;
        RECT 2268.990 3416.000 2269.270 3419.310 ;
        RECT 106.360 16.670 106.620 16.990 ;
        RECT 300.020 16.670 300.280 16.990 ;
        RECT 300.080 2.400 300.220 16.670 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 317.930 20.640 318.250 20.700 ;
        RECT 323.910 20.640 324.230 20.700 ;
        RECT 317.930 20.500 324.230 20.640 ;
        RECT 317.930 20.440 318.250 20.500 ;
        RECT 323.910 20.440 324.230 20.500 ;
      LAYER via ;
        RECT 317.960 20.440 318.220 20.700 ;
        RECT 323.940 20.440 324.200 20.700 ;
      LAYER met2 ;
        RECT 2638.370 100.370 2638.650 104.000 ;
        RECT 2636.880 100.230 2638.650 100.370 ;
        RECT 2636.880 87.565 2637.020 100.230 ;
        RECT 2638.370 100.000 2638.650 100.230 ;
        RECT 323.930 87.195 324.210 87.565 ;
        RECT 2636.810 87.195 2637.090 87.565 ;
        RECT 324.000 20.730 324.140 87.195 ;
        RECT 317.960 20.410 318.220 20.730 ;
        RECT 323.940 20.410 324.200 20.730 ;
        RECT 318.020 2.400 318.160 20.410 ;
        RECT 317.810 -4.800 318.370 2.400 ;
      LAYER via2 ;
        RECT 323.930 87.240 324.210 87.520 ;
        RECT 2636.810 87.240 2637.090 87.520 ;
      LAYER met3 ;
        RECT 323.905 87.530 324.235 87.545 ;
        RECT 2636.785 87.530 2637.115 87.545 ;
        RECT 323.905 87.230 2637.115 87.530 ;
        RECT 323.905 87.215 324.235 87.230 ;
        RECT 2636.785 87.215 2637.115 87.230 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 335.870 31.180 336.190 31.240 ;
        RECT 2857.130 31.180 2857.450 31.240 ;
        RECT 335.870 31.040 2857.450 31.180 ;
        RECT 335.870 30.980 336.190 31.040 ;
        RECT 2857.130 30.980 2857.450 31.040 ;
      LAYER via ;
        RECT 335.900 30.980 336.160 31.240 ;
        RECT 2857.160 30.980 2857.420 31.240 ;
      LAYER met2 ;
        RECT 2857.150 2886.075 2857.430 2886.445 ;
        RECT 2857.220 31.270 2857.360 2886.075 ;
        RECT 335.900 30.950 336.160 31.270 ;
        RECT 2857.160 30.950 2857.420 31.270 ;
        RECT 335.960 2.400 336.100 30.950 ;
        RECT 335.750 -4.800 336.310 2.400 ;
      LAYER via2 ;
        RECT 2857.150 2886.120 2857.430 2886.400 ;
      LAYER met3 ;
        RECT 2841.000 2886.410 2845.000 2886.600 ;
        RECT 2857.125 2886.410 2857.455 2886.425 ;
        RECT 2841.000 2886.110 2857.455 2886.410 ;
        RECT 2841.000 2886.000 2845.000 2886.110 ;
        RECT 2857.125 2886.095 2857.455 2886.110 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2356.210 3429.395 2356.490 3429.765 ;
        RECT 2356.280 3419.450 2356.420 3429.395 ;
        RECT 2357.770 3419.450 2358.050 3420.000 ;
        RECT 2356.280 3419.310 2358.050 3419.450 ;
        RECT 2357.770 3416.000 2358.050 3419.310 ;
        RECT 353.370 18.515 353.650 18.885 ;
        RECT 353.440 2.400 353.580 18.515 ;
        RECT 353.230 -4.800 353.790 2.400 ;
      LAYER via2 ;
        RECT 2356.210 3429.440 2356.490 3429.720 ;
        RECT 353.370 18.560 353.650 18.840 ;
      LAYER met3 ;
        RECT 114.350 3429.730 114.730 3429.740 ;
        RECT 2356.185 3429.730 2356.515 3429.745 ;
        RECT 114.350 3429.430 2356.515 3429.730 ;
        RECT 114.350 3429.420 114.730 3429.430 ;
        RECT 2356.185 3429.415 2356.515 3429.430 ;
        RECT 114.350 18.850 114.730 18.860 ;
        RECT 353.345 18.850 353.675 18.865 ;
        RECT 114.350 18.550 353.675 18.850 ;
        RECT 114.350 18.540 114.730 18.550 ;
        RECT 353.345 18.535 353.675 18.550 ;
      LAYER via3 ;
        RECT 114.380 3429.420 114.700 3429.740 ;
        RECT 114.380 18.540 114.700 18.860 ;
      LAYER met4 ;
        RECT 114.375 3429.415 114.705 3429.745 ;
        RECT 114.390 18.865 114.690 3429.415 ;
        RECT 114.375 18.535 114.705 18.865 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 108.170 3429.820 108.490 3429.880 ;
        RECT 2444.510 3429.820 2444.830 3429.880 ;
        RECT 108.170 3429.680 2444.830 3429.820 ;
        RECT 108.170 3429.620 108.490 3429.680 ;
        RECT 2444.510 3429.620 2444.830 3429.680 ;
      LAYER via ;
        RECT 108.200 3429.620 108.460 3429.880 ;
        RECT 2444.540 3429.620 2444.800 3429.880 ;
      LAYER met2 ;
        RECT 108.200 3429.590 108.460 3429.910 ;
        RECT 2444.540 3429.590 2444.800 3429.910 ;
        RECT 108.260 17.525 108.400 3429.590 ;
        RECT 2444.600 3419.450 2444.740 3429.590 ;
        RECT 2446.090 3419.450 2446.370 3420.000 ;
        RECT 2444.600 3419.310 2446.370 3419.450 ;
        RECT 2446.090 3416.000 2446.370 3419.310 ;
        RECT 108.190 17.155 108.470 17.525 ;
        RECT 371.310 17.155 371.590 17.525 ;
        RECT 371.380 2.400 371.520 17.155 ;
        RECT 371.170 -4.800 371.730 2.400 ;
      LAYER via2 ;
        RECT 108.190 17.200 108.470 17.480 ;
        RECT 371.310 17.200 371.590 17.480 ;
      LAYER met3 ;
        RECT 108.165 17.490 108.495 17.505 ;
        RECT 371.285 17.490 371.615 17.505 ;
        RECT 108.165 17.190 371.615 17.490 ;
        RECT 108.165 17.175 108.495 17.190 ;
        RECT 371.285 17.175 371.615 17.190 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 389.230 31.520 389.550 31.580 ;
        RECT 2856.670 31.520 2856.990 31.580 ;
        RECT 389.230 31.380 2856.990 31.520 ;
        RECT 389.230 31.320 389.550 31.380 ;
        RECT 2856.670 31.320 2856.990 31.380 ;
      LAYER via ;
        RECT 389.260 31.320 389.520 31.580 ;
        RECT 2856.700 31.320 2856.960 31.580 ;
      LAYER met2 ;
        RECT 2856.690 3004.395 2856.970 3004.765 ;
        RECT 2856.760 31.610 2856.900 3004.395 ;
        RECT 389.260 31.290 389.520 31.610 ;
        RECT 2856.700 31.290 2856.960 31.610 ;
        RECT 389.320 2.400 389.460 31.290 ;
        RECT 389.110 -4.800 389.670 2.400 ;
      LAYER via2 ;
        RECT 2856.690 3004.440 2856.970 3004.720 ;
      LAYER met3 ;
        RECT 2841.000 3004.730 2845.000 3004.920 ;
        RECT 2856.665 3004.730 2856.995 3004.745 ;
        RECT 2841.000 3004.430 2856.995 3004.730 ;
        RECT 2841.000 3004.320 2845.000 3004.430 ;
        RECT 2856.665 3004.415 2856.995 3004.430 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 407.190 17.155 407.470 17.525 ;
        RECT 407.260 2.400 407.400 17.155 ;
        RECT 407.050 -4.800 407.610 2.400 ;
      LAYER via2 ;
        RECT 407.190 17.200 407.470 17.480 ;
      LAYER met3 ;
        RECT 2841.000 3123.050 2845.000 3123.240 ;
        RECT 2858.710 3123.050 2859.090 3123.060 ;
        RECT 2841.000 3122.750 2859.090 3123.050 ;
        RECT 2841.000 3122.640 2845.000 3122.750 ;
        RECT 2858.710 3122.740 2859.090 3122.750 ;
        RECT 407.165 17.490 407.495 17.505 ;
        RECT 2858.710 17.490 2859.090 17.500 ;
        RECT 407.165 17.190 2859.090 17.490 ;
        RECT 407.165 17.175 407.495 17.190 ;
        RECT 2858.710 17.180 2859.090 17.190 ;
      LAYER via3 ;
        RECT 2858.740 3122.740 2859.060 3123.060 ;
        RECT 2858.740 17.180 2859.060 17.500 ;
      LAYER met4 ;
        RECT 2858.735 3122.735 2859.065 3123.065 ;
        RECT 2858.750 17.505 2859.050 3122.735 ;
        RECT 2858.735 17.175 2859.065 17.505 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 68.610 3431.860 68.930 3431.920 ;
        RECT 1913.210 3431.860 1913.530 3431.920 ;
        RECT 68.610 3431.720 1913.530 3431.860 ;
        RECT 68.610 3431.660 68.930 3431.720 ;
        RECT 1913.210 3431.660 1913.530 3431.720 ;
      LAYER via ;
        RECT 68.640 3431.660 68.900 3431.920 ;
        RECT 1913.240 3431.660 1913.500 3431.920 ;
      LAYER met2 ;
        RECT 68.640 3431.630 68.900 3431.950 ;
        RECT 1913.240 3431.630 1913.500 3431.950 ;
        RECT 68.700 17.410 68.840 3431.630 ;
        RECT 1913.300 3419.450 1913.440 3431.630 ;
        RECT 1914.790 3419.450 1915.070 3420.000 ;
        RECT 1913.300 3419.310 1915.070 3419.450 ;
        RECT 1914.790 3416.000 1915.070 3419.310 ;
        RECT 68.240 17.270 68.840 17.410 ;
        RECT 68.240 2.400 68.380 17.270 ;
        RECT 68.030 -4.800 68.590 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 424.650 20.300 424.970 20.360 ;
        RECT 394.840 20.160 424.970 20.300 ;
        RECT 87.010 19.960 87.330 20.020 ;
        RECT 394.840 19.960 394.980 20.160 ;
        RECT 424.650 20.100 424.970 20.160 ;
        RECT 87.010 19.820 394.980 19.960 ;
        RECT 87.010 19.760 87.330 19.820 ;
      LAYER via ;
        RECT 87.040 19.760 87.300 20.020 ;
        RECT 424.680 20.100 424.940 20.360 ;
      LAYER met2 ;
        RECT 87.030 2422.995 87.310 2423.365 ;
        RECT 87.100 20.050 87.240 2422.995 ;
        RECT 424.680 20.070 424.940 20.390 ;
        RECT 87.040 19.730 87.300 20.050 ;
        RECT 424.740 2.400 424.880 20.070 ;
        RECT 424.530 -4.800 425.090 2.400 ;
      LAYER via2 ;
        RECT 87.030 2423.040 87.310 2423.320 ;
      LAYER met3 ;
        RECT 87.005 2423.330 87.335 2423.345 ;
        RECT 100.000 2423.330 104.000 2423.520 ;
        RECT 87.005 2423.030 104.000 2423.330 ;
        RECT 87.005 2423.015 87.335 2423.030 ;
        RECT 100.000 2422.920 104.000 2423.030 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 87.470 19.620 87.790 19.680 ;
        RECT 442.590 19.620 442.910 19.680 ;
        RECT 87.470 19.480 442.910 19.620 ;
        RECT 87.470 19.420 87.790 19.480 ;
        RECT 442.590 19.420 442.910 19.480 ;
      LAYER via ;
        RECT 87.500 19.420 87.760 19.680 ;
        RECT 442.620 19.420 442.880 19.680 ;
      LAYER met2 ;
        RECT 87.490 2556.275 87.770 2556.645 ;
        RECT 87.560 19.710 87.700 2556.275 ;
        RECT 87.500 19.390 87.760 19.710 ;
        RECT 442.620 19.390 442.880 19.710 ;
        RECT 442.680 2.400 442.820 19.390 ;
        RECT 442.470 -4.800 443.030 2.400 ;
      LAYER via2 ;
        RECT 87.490 2556.320 87.770 2556.600 ;
      LAYER met3 ;
        RECT 87.465 2556.610 87.795 2556.625 ;
        RECT 100.000 2556.610 104.000 2556.800 ;
        RECT 87.465 2556.310 104.000 2556.610 ;
        RECT 87.465 2556.295 87.795 2556.310 ;
        RECT 100.000 2556.200 104.000 2556.310 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 430.245 19.125 430.415 20.315 ;
      LAYER mcon ;
        RECT 430.245 20.145 430.415 20.315 ;
      LAYER met1 ;
        RECT 430.185 20.300 430.475 20.345 ;
        RECT 460.530 20.300 460.850 20.360 ;
        RECT 430.185 20.160 460.850 20.300 ;
        RECT 430.185 20.115 430.475 20.160 ;
        RECT 460.530 20.100 460.850 20.160 ;
        RECT 87.930 19.280 88.250 19.340 ;
        RECT 430.185 19.280 430.475 19.325 ;
        RECT 87.930 19.140 430.475 19.280 ;
        RECT 87.930 19.080 88.250 19.140 ;
        RECT 430.185 19.095 430.475 19.140 ;
      LAYER via ;
        RECT 460.560 20.100 460.820 20.360 ;
        RECT 87.960 19.080 88.220 19.340 ;
      LAYER met2 ;
        RECT 87.950 2688.875 88.230 2689.245 ;
        RECT 88.020 19.370 88.160 2688.875 ;
        RECT 460.560 20.070 460.820 20.390 ;
        RECT 87.960 19.050 88.220 19.370 ;
        RECT 460.620 2.400 460.760 20.070 ;
        RECT 460.410 -4.800 460.970 2.400 ;
      LAYER via2 ;
        RECT 87.950 2688.920 88.230 2689.200 ;
      LAYER met3 ;
        RECT 87.925 2689.210 88.255 2689.225 ;
        RECT 100.000 2689.210 104.000 2689.400 ;
        RECT 87.925 2688.910 104.000 2689.210 ;
        RECT 87.925 2688.895 88.255 2688.910 ;
        RECT 100.000 2688.800 104.000 2688.910 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 478.490 17.835 478.770 18.205 ;
        RECT 478.560 2.400 478.700 17.835 ;
        RECT 478.350 -4.800 478.910 2.400 ;
      LAYER via2 ;
        RECT 478.490 17.880 478.770 18.160 ;
      LAYER met3 ;
        RECT 2841.000 3242.050 2845.000 3242.240 ;
        RECT 2857.790 3242.050 2858.170 3242.060 ;
        RECT 2841.000 3241.750 2858.170 3242.050 ;
        RECT 2841.000 3241.640 2845.000 3241.750 ;
        RECT 2857.790 3241.740 2858.170 3241.750 ;
        RECT 478.465 18.170 478.795 18.185 ;
        RECT 2857.790 18.170 2858.170 18.180 ;
        RECT 478.465 17.870 2858.170 18.170 ;
        RECT 478.465 17.855 478.795 17.870 ;
        RECT 2857.790 17.860 2858.170 17.870 ;
      LAYER via3 ;
        RECT 2857.820 3241.740 2858.140 3242.060 ;
        RECT 2857.820 17.860 2858.140 18.180 ;
      LAYER met4 ;
        RECT 2857.815 3241.735 2858.145 3242.065 ;
        RECT 2857.830 18.185 2858.130 3241.735 ;
        RECT 2857.815 17.855 2858.145 18.185 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2536.530 3429.395 2536.810 3429.765 ;
        RECT 2534.870 3419.450 2535.150 3420.000 ;
        RECT 2536.600 3419.450 2536.740 3429.395 ;
        RECT 2534.870 3419.310 2536.740 3419.450 ;
        RECT 2534.870 3416.000 2535.150 3419.310 ;
        RECT 496.430 18.515 496.710 18.885 ;
        RECT 496.500 2.400 496.640 18.515 ;
        RECT 496.290 -4.800 496.850 2.400 ;
      LAYER via2 ;
        RECT 2536.530 3429.440 2536.810 3429.720 ;
        RECT 496.430 18.560 496.710 18.840 ;
      LAYER met3 ;
        RECT 2536.505 3429.730 2536.835 3429.745 ;
        RECT 2815.470 3429.730 2815.850 3429.740 ;
        RECT 2536.505 3429.430 2815.850 3429.730 ;
        RECT 2536.505 3429.415 2536.835 3429.430 ;
        RECT 2815.470 3429.420 2815.850 3429.430 ;
        RECT 496.405 18.850 496.735 18.865 ;
        RECT 2815.470 18.850 2815.850 18.860 ;
        RECT 496.405 18.550 2815.850 18.850 ;
        RECT 496.405 18.535 496.735 18.550 ;
        RECT 2815.470 18.540 2815.850 18.550 ;
      LAYER via3 ;
        RECT 2815.500 3429.420 2815.820 3429.740 ;
        RECT 2815.500 18.540 2815.820 18.860 ;
      LAYER met4 ;
        RECT 2815.495 3429.415 2815.825 3429.745 ;
        RECT 2815.510 18.865 2815.810 3429.415 ;
        RECT 2815.495 18.535 2815.825 18.865 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 88.390 18.940 88.710 19.000 ;
        RECT 513.890 18.940 514.210 19.000 ;
        RECT 88.390 18.800 514.210 18.940 ;
        RECT 88.390 18.740 88.710 18.800 ;
        RECT 513.890 18.740 514.210 18.800 ;
      LAYER via ;
        RECT 88.420 18.740 88.680 19.000 ;
        RECT 513.920 18.740 514.180 19.000 ;
      LAYER met2 ;
        RECT 88.410 2821.475 88.690 2821.845 ;
        RECT 88.480 19.030 88.620 2821.475 ;
        RECT 88.420 18.710 88.680 19.030 ;
        RECT 513.920 18.710 514.180 19.030 ;
        RECT 513.980 2.400 514.120 18.710 ;
        RECT 513.770 -4.800 514.330 2.400 ;
      LAYER via2 ;
        RECT 88.410 2821.520 88.690 2821.800 ;
      LAYER met3 ;
        RECT 88.385 2821.810 88.715 2821.825 ;
        RECT 100.000 2821.810 104.000 2822.000 ;
        RECT 88.385 2821.510 104.000 2821.810 ;
        RECT 88.385 2821.495 88.715 2821.510 ;
        RECT 100.000 2821.400 104.000 2821.510 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2624.850 3430.075 2625.130 3430.445 ;
        RECT 2623.190 3419.450 2623.470 3420.000 ;
        RECT 2624.920 3419.450 2625.060 3430.075 ;
        RECT 2623.190 3419.310 2625.060 3419.450 ;
        RECT 2623.190 3416.000 2623.470 3419.310 ;
        RECT 531.850 19.875 532.130 20.245 ;
        RECT 531.920 2.400 532.060 19.875 ;
        RECT 531.710 -4.800 532.270 2.400 ;
      LAYER via2 ;
        RECT 2624.850 3430.120 2625.130 3430.400 ;
        RECT 531.850 19.920 532.130 20.200 ;
      LAYER met3 ;
        RECT 2624.825 3430.410 2625.155 3430.425 ;
        RECT 2816.390 3430.410 2816.770 3430.420 ;
        RECT 2624.825 3430.110 2816.770 3430.410 ;
        RECT 2624.825 3430.095 2625.155 3430.110 ;
        RECT 2816.390 3430.100 2816.770 3430.110 ;
        RECT 531.825 20.210 532.155 20.225 ;
        RECT 2816.390 20.210 2816.770 20.220 ;
        RECT 531.825 19.910 2816.770 20.210 ;
        RECT 531.825 19.895 532.155 19.910 ;
        RECT 2816.390 19.900 2816.770 19.910 ;
      LAYER via3 ;
        RECT 2816.420 3430.100 2816.740 3430.420 ;
        RECT 2816.420 19.900 2816.740 20.220 ;
      LAYER met4 ;
        RECT 2816.415 3430.095 2816.745 3430.425 ;
        RECT 2816.430 20.225 2816.730 3430.095 ;
        RECT 2816.415 19.895 2816.745 20.225 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 549.790 19.195 550.070 19.565 ;
        RECT 549.860 2.400 550.000 19.195 ;
        RECT 549.650 -4.800 550.210 2.400 ;
      LAYER via2 ;
        RECT 549.790 19.240 550.070 19.520 ;
      LAYER met3 ;
        RECT 2841.000 3360.370 2845.000 3360.560 ;
        RECT 2856.870 3360.370 2857.250 3360.380 ;
        RECT 2841.000 3360.070 2857.250 3360.370 ;
        RECT 2841.000 3359.960 2845.000 3360.070 ;
        RECT 2856.870 3360.060 2857.250 3360.070 ;
        RECT 549.765 19.530 550.095 19.545 ;
        RECT 2856.870 19.530 2857.250 19.540 ;
        RECT 549.765 19.230 2857.250 19.530 ;
        RECT 549.765 19.215 550.095 19.230 ;
        RECT 2856.870 19.220 2857.250 19.230 ;
      LAYER via3 ;
        RECT 2856.900 3360.060 2857.220 3360.380 ;
        RECT 2856.900 19.220 2857.220 19.540 ;
      LAYER met4 ;
        RECT 2856.895 3360.055 2857.225 3360.385 ;
        RECT 2856.910 19.545 2857.210 3360.055 ;
        RECT 2856.895 19.215 2857.225 19.545 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 567.710 18.600 568.030 18.660 ;
        RECT 572.310 18.600 572.630 18.660 ;
        RECT 567.710 18.460 572.630 18.600 ;
        RECT 567.710 18.400 568.030 18.460 ;
        RECT 572.310 18.400 572.630 18.460 ;
      LAYER via ;
        RECT 567.740 18.400 568.000 18.660 ;
        RECT 572.340 18.400 572.600 18.660 ;
      LAYER met2 ;
        RECT 2713.630 3430.755 2713.910 3431.125 ;
        RECT 2711.970 3419.450 2712.250 3420.000 ;
        RECT 2713.700 3419.450 2713.840 3430.755 ;
        RECT 2711.970 3419.310 2713.840 3419.450 ;
        RECT 2711.970 3416.000 2712.250 3419.310 ;
        RECT 572.330 99.435 572.610 99.805 ;
        RECT 572.400 18.690 572.540 99.435 ;
        RECT 567.740 18.370 568.000 18.690 ;
        RECT 572.340 18.370 572.600 18.690 ;
        RECT 567.800 2.400 567.940 18.370 ;
        RECT 567.590 -4.800 568.150 2.400 ;
      LAYER via2 ;
        RECT 2713.630 3430.800 2713.910 3431.080 ;
        RECT 572.330 99.480 572.610 99.760 ;
      LAYER met3 ;
        RECT 2713.605 3431.090 2713.935 3431.105 ;
        RECT 2808.110 3431.090 2808.490 3431.100 ;
        RECT 2713.605 3430.790 2808.490 3431.090 ;
        RECT 2713.605 3430.775 2713.935 3430.790 ;
        RECT 2808.110 3430.780 2808.490 3430.790 ;
        RECT 572.305 99.770 572.635 99.785 ;
        RECT 2808.110 99.770 2808.490 99.780 ;
        RECT 572.305 99.470 2808.490 99.770 ;
        RECT 572.305 99.455 572.635 99.470 ;
        RECT 2808.110 99.460 2808.490 99.470 ;
      LAYER via3 ;
        RECT 2808.140 3430.780 2808.460 3431.100 ;
        RECT 2808.140 99.460 2808.460 99.780 ;
      LAYER met4 ;
        RECT 2808.135 3430.775 2808.465 3431.105 ;
        RECT 2808.150 99.785 2808.450 3430.775 ;
        RECT 2808.135 99.455 2808.465 99.785 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 585.650 86.600 585.970 86.660 ;
        RECT 2684.170 86.600 2684.490 86.660 ;
        RECT 585.650 86.460 2684.490 86.600 ;
        RECT 585.650 86.400 585.970 86.460 ;
        RECT 2684.170 86.400 2684.490 86.460 ;
      LAYER via ;
        RECT 585.680 86.400 585.940 86.660 ;
        RECT 2684.200 86.400 2684.460 86.660 ;
      LAYER met2 ;
        RECT 2684.370 100.370 2684.650 104.000 ;
        RECT 2684.260 100.000 2684.650 100.370 ;
        RECT 2684.260 86.690 2684.400 100.000 ;
        RECT 585.680 86.370 585.940 86.690 ;
        RECT 2684.200 86.370 2684.460 86.690 ;
        RECT 585.740 2.400 585.880 86.370 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 91.610 17.920 91.930 17.980 ;
        RECT 95.750 17.920 96.070 17.980 ;
        RECT 91.610 17.780 96.070 17.920 ;
        RECT 91.610 17.720 91.930 17.780 ;
        RECT 95.750 17.720 96.070 17.780 ;
      LAYER via ;
        RECT 91.640 17.720 91.900 17.980 ;
        RECT 95.780 17.720 96.040 17.980 ;
      LAYER met2 ;
        RECT 2409.750 100.370 2410.030 104.000 ;
        RECT 2408.260 100.230 2410.030 100.370 ;
        RECT 2408.260 86.885 2408.400 100.230 ;
        RECT 2409.750 100.000 2410.030 100.230 ;
        RECT 95.770 86.515 96.050 86.885 ;
        RECT 2408.190 86.515 2408.470 86.885 ;
        RECT 95.840 18.010 95.980 86.515 ;
        RECT 91.640 17.690 91.900 18.010 ;
        RECT 95.780 17.690 96.040 18.010 ;
        RECT 91.700 2.400 91.840 17.690 ;
        RECT 91.490 -4.800 92.050 2.400 ;
      LAYER via2 ;
        RECT 95.770 86.560 96.050 86.840 ;
        RECT 2408.190 86.560 2408.470 86.840 ;
      LAYER met3 ;
        RECT 95.745 86.850 96.075 86.865 ;
        RECT 2408.165 86.850 2408.495 86.865 ;
        RECT 95.745 86.550 2408.495 86.850 ;
        RECT 95.745 86.535 96.075 86.550 ;
        RECT 2408.165 86.535 2408.495 86.550 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 88.850 15.200 89.170 15.260 ;
        RECT 603.130 15.200 603.450 15.260 ;
        RECT 88.850 15.060 603.450 15.200 ;
        RECT 88.850 15.000 89.170 15.060 ;
        RECT 603.130 15.000 603.450 15.060 ;
      LAYER via ;
        RECT 88.880 15.000 89.140 15.260 ;
        RECT 603.160 15.000 603.420 15.260 ;
      LAYER met2 ;
        RECT 88.870 2954.075 89.150 2954.445 ;
        RECT 88.940 15.290 89.080 2954.075 ;
        RECT 88.880 14.970 89.140 15.290 ;
        RECT 603.160 14.970 603.420 15.290 ;
        RECT 603.220 2.400 603.360 14.970 ;
        RECT 603.010 -4.800 603.570 2.400 ;
      LAYER via2 ;
        RECT 88.870 2954.120 89.150 2954.400 ;
      LAYER met3 ;
        RECT 88.845 2954.410 89.175 2954.425 ;
        RECT 100.000 2954.410 104.000 2954.600 ;
        RECT 88.845 2954.110 104.000 2954.410 ;
        RECT 88.845 2954.095 89.175 2954.110 ;
        RECT 100.000 2954.000 104.000 2954.110 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 627.050 86.260 627.370 86.320 ;
        RECT 2728.330 86.260 2728.650 86.320 ;
        RECT 627.050 86.120 2728.650 86.260 ;
        RECT 627.050 86.060 627.370 86.120 ;
        RECT 2728.330 86.060 2728.650 86.120 ;
        RECT 621.070 18.600 621.390 18.660 ;
        RECT 627.050 18.600 627.370 18.660 ;
        RECT 621.070 18.460 627.370 18.600 ;
        RECT 621.070 18.400 621.390 18.460 ;
        RECT 627.050 18.400 627.370 18.460 ;
      LAYER via ;
        RECT 627.080 86.060 627.340 86.320 ;
        RECT 2728.360 86.060 2728.620 86.320 ;
        RECT 621.100 18.400 621.360 18.660 ;
        RECT 627.080 18.400 627.340 18.660 ;
      LAYER met2 ;
        RECT 2729.910 100.370 2730.190 104.000 ;
        RECT 2728.420 100.230 2730.190 100.370 ;
        RECT 2728.420 86.350 2728.560 100.230 ;
        RECT 2729.910 100.000 2730.190 100.230 ;
        RECT 627.080 86.030 627.340 86.350 ;
        RECT 2728.360 86.030 2728.620 86.350 ;
        RECT 627.140 18.690 627.280 86.030 ;
        RECT 621.100 18.370 621.360 18.690 ;
        RECT 627.080 18.370 627.340 18.690 ;
        RECT 621.160 2.400 621.300 18.370 ;
        RECT 620.950 -4.800 621.510 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 86.550 14.860 86.870 14.920 ;
        RECT 115.530 14.860 115.850 14.920 ;
        RECT 86.550 14.720 115.850 14.860 ;
        RECT 86.550 14.660 86.870 14.720 ;
        RECT 115.530 14.660 115.850 14.720 ;
      LAYER via ;
        RECT 86.580 14.660 86.840 14.920 ;
        RECT 115.560 14.660 115.820 14.920 ;
      LAYER met2 ;
        RECT 86.570 2157.795 86.850 2158.165 ;
        RECT 86.640 14.950 86.780 2157.795 ;
        RECT 86.580 14.630 86.840 14.950 ;
        RECT 115.560 14.630 115.820 14.950 ;
        RECT 115.620 2.400 115.760 14.630 ;
        RECT 115.410 -4.800 115.970 2.400 ;
      LAYER via2 ;
        RECT 86.570 2157.840 86.850 2158.120 ;
      LAYER met3 ;
        RECT 86.545 2158.130 86.875 2158.145 ;
        RECT 100.000 2158.130 104.000 2158.320 ;
        RECT 86.545 2157.830 104.000 2158.130 ;
        RECT 86.545 2157.815 86.875 2157.830 ;
        RECT 100.000 2157.720 104.000 2157.830 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 106.790 3431.520 107.110 3431.580 ;
        RECT 2001.990 3431.520 2002.310 3431.580 ;
        RECT 106.790 3431.380 2002.310 3431.520 ;
        RECT 106.790 3431.320 107.110 3431.380 ;
        RECT 2001.990 3431.320 2002.310 3431.380 ;
        RECT 106.790 102.920 107.110 102.980 ;
        RECT 138.070 102.920 138.390 102.980 ;
        RECT 106.790 102.780 138.390 102.920 ;
        RECT 106.790 102.720 107.110 102.780 ;
        RECT 138.070 102.720 138.390 102.780 ;
      LAYER via ;
        RECT 106.820 3431.320 107.080 3431.580 ;
        RECT 2002.020 3431.320 2002.280 3431.580 ;
        RECT 106.820 102.720 107.080 102.980 ;
        RECT 138.100 102.720 138.360 102.980 ;
      LAYER met2 ;
        RECT 106.820 3431.290 107.080 3431.610 ;
        RECT 2002.020 3431.290 2002.280 3431.610 ;
        RECT 106.880 103.010 107.020 3431.290 ;
        RECT 2002.080 3419.450 2002.220 3431.290 ;
        RECT 2003.570 3419.450 2003.850 3420.000 ;
        RECT 2002.080 3419.310 2003.850 3419.450 ;
        RECT 2003.570 3416.000 2003.850 3419.310 ;
        RECT 106.820 102.690 107.080 103.010 ;
        RECT 138.100 102.690 138.360 103.010 ;
        RECT 138.160 16.730 138.300 102.690 ;
        RECT 138.160 16.590 139.680 16.730 ;
        RECT 139.540 2.400 139.680 16.590 ;
        RECT 139.330 -4.800 139.890 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2455.290 100.370 2455.570 104.000 ;
        RECT 2453.800 100.230 2455.570 100.370 ;
        RECT 2453.800 88.245 2453.940 100.230 ;
        RECT 2455.290 100.000 2455.570 100.230 ;
        RECT 158.330 87.875 158.610 88.245 ;
        RECT 2453.730 87.875 2454.010 88.245 ;
        RECT 158.400 16.730 158.540 87.875 ;
        RECT 157.480 16.590 158.540 16.730 ;
        RECT 157.480 2.400 157.620 16.590 ;
        RECT 157.270 -4.800 157.830 2.400 ;
      LAYER via2 ;
        RECT 158.330 87.920 158.610 88.200 ;
        RECT 2453.730 87.920 2454.010 88.200 ;
      LAYER met3 ;
        RECT 158.305 88.210 158.635 88.225 ;
        RECT 2453.705 88.210 2454.035 88.225 ;
        RECT 158.305 87.910 2454.035 88.210 ;
        RECT 158.305 87.895 158.635 87.910 ;
        RECT 2453.705 87.895 2454.035 87.910 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 174.870 18.260 175.190 18.320 ;
        RECT 2497.870 18.260 2498.190 18.320 ;
        RECT 174.870 18.120 2498.190 18.260 ;
        RECT 174.870 18.060 175.190 18.120 ;
        RECT 2497.870 18.060 2498.190 18.120 ;
      LAYER via ;
        RECT 174.900 18.060 175.160 18.320 ;
        RECT 2497.900 18.060 2498.160 18.320 ;
      LAYER met2 ;
        RECT 2501.290 100.370 2501.570 104.000 ;
        RECT 2497.960 100.230 2501.570 100.370 ;
        RECT 2497.960 18.350 2498.100 100.230 ;
        RECT 2501.290 100.000 2501.570 100.230 ;
        RECT 174.900 18.030 175.160 18.350 ;
        RECT 2497.900 18.030 2498.160 18.350 ;
        RECT 174.960 2.400 175.100 18.030 ;
        RECT 174.750 -4.800 175.310 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2857.610 2767.075 2857.890 2767.445 ;
        RECT 2857.680 16.845 2857.820 2767.075 ;
        RECT 192.830 16.475 193.110 16.845 ;
        RECT 2857.610 16.475 2857.890 16.845 ;
        RECT 192.900 2.400 193.040 16.475 ;
        RECT 192.690 -4.800 193.250 2.400 ;
      LAYER via2 ;
        RECT 2857.610 2767.120 2857.890 2767.400 ;
        RECT 192.830 16.520 193.110 16.800 ;
        RECT 2857.610 16.520 2857.890 16.800 ;
      LAYER met3 ;
        RECT 2841.000 2767.410 2845.000 2767.600 ;
        RECT 2857.585 2767.410 2857.915 2767.425 ;
        RECT 2841.000 2767.110 2857.915 2767.410 ;
        RECT 2841.000 2767.000 2845.000 2767.110 ;
        RECT 2857.585 2767.095 2857.915 2767.110 ;
        RECT 192.805 16.810 193.135 16.825 ;
        RECT 2857.585 16.810 2857.915 16.825 ;
        RECT 192.805 16.510 2857.915 16.810 ;
        RECT 192.805 16.495 193.135 16.510 ;
        RECT 2857.585 16.495 2857.915 16.510 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 210.750 17.920 211.070 17.980 ;
        RECT 213.510 17.920 213.830 17.980 ;
        RECT 210.750 17.780 213.830 17.920 ;
        RECT 210.750 17.720 211.070 17.780 ;
        RECT 213.510 17.720 213.830 17.780 ;
      LAYER via ;
        RECT 210.780 17.720 211.040 17.980 ;
        RECT 213.540 17.720 213.800 17.980 ;
      LAYER met2 ;
        RECT 2546.830 100.370 2547.110 104.000 ;
        RECT 2546.260 100.230 2547.110 100.370 ;
        RECT 2546.260 86.205 2546.400 100.230 ;
        RECT 2546.830 100.000 2547.110 100.230 ;
        RECT 213.530 85.835 213.810 86.205 ;
        RECT 2546.190 85.835 2546.470 86.205 ;
        RECT 213.600 18.010 213.740 85.835 ;
        RECT 210.780 17.690 211.040 18.010 ;
        RECT 213.540 17.690 213.800 18.010 ;
        RECT 210.840 2.400 210.980 17.690 ;
        RECT 210.630 -4.800 211.190 2.400 ;
      LAYER via2 ;
        RECT 213.530 85.880 213.810 86.160 ;
        RECT 2546.190 85.880 2546.470 86.160 ;
      LAYER met3 ;
        RECT 213.505 86.170 213.835 86.185 ;
        RECT 2546.165 86.170 2546.495 86.185 ;
        RECT 213.505 85.870 2546.495 86.170 ;
        RECT 213.505 85.855 213.835 85.870 ;
        RECT 2546.165 85.855 2546.495 85.870 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 255.445 14.025 255.615 17.935 ;
      LAYER mcon ;
        RECT 255.445 17.765 255.615 17.935 ;
      LAYER met1 ;
        RECT 255.385 17.920 255.675 17.965 ;
        RECT 2587.570 17.920 2587.890 17.980 ;
        RECT 255.385 17.780 2587.890 17.920 ;
        RECT 255.385 17.735 255.675 17.780 ;
        RECT 2587.570 17.720 2587.890 17.780 ;
        RECT 255.385 14.180 255.675 14.225 ;
        RECT 247.180 14.040 255.675 14.180 ;
        RECT 228.690 13.840 229.010 13.900 ;
        RECT 247.180 13.840 247.320 14.040 ;
        RECT 255.385 13.995 255.675 14.040 ;
        RECT 228.690 13.700 247.320 13.840 ;
        RECT 228.690 13.640 229.010 13.700 ;
      LAYER via ;
        RECT 2587.600 17.720 2587.860 17.980 ;
        RECT 228.720 13.640 228.980 13.900 ;
      LAYER met2 ;
        RECT 2592.830 100.370 2593.110 104.000 ;
        RECT 2587.660 100.230 2593.110 100.370 ;
        RECT 2587.660 18.010 2587.800 100.230 ;
        RECT 2592.830 100.000 2593.110 100.230 ;
        RECT 2587.600 17.690 2587.860 18.010 ;
        RECT 228.720 13.610 228.980 13.930 ;
        RECT 228.780 2.400 228.920 13.610 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 54.810 87.620 55.130 87.680 ;
        RECT 486.750 87.620 487.070 87.680 ;
        RECT 54.810 87.480 487.070 87.620 ;
        RECT 54.810 87.420 55.130 87.480 ;
        RECT 486.750 87.420 487.070 87.480 ;
        RECT 50.210 17.580 50.530 17.640 ;
        RECT 54.810 17.580 55.130 17.640 ;
        RECT 50.210 17.440 55.130 17.580 ;
        RECT 50.210 17.380 50.530 17.440 ;
        RECT 54.810 17.380 55.130 17.440 ;
      LAYER via ;
        RECT 54.840 87.420 55.100 87.680 ;
        RECT 486.780 87.420 487.040 87.680 ;
        RECT 50.240 17.380 50.500 17.640 ;
        RECT 54.840 17.380 55.100 17.640 ;
      LAYER met2 ;
        RECT 488.330 100.370 488.610 104.000 ;
        RECT 486.840 100.230 488.610 100.370 ;
        RECT 486.840 87.710 486.980 100.230 ;
        RECT 488.330 100.000 488.610 100.230 ;
        RECT 54.840 87.390 55.100 87.710 ;
        RECT 486.780 87.390 487.040 87.710 ;
        RECT 54.900 17.670 55.040 87.390 ;
        RECT 50.240 17.350 50.500 17.670 ;
        RECT 54.840 17.350 55.100 17.670 ;
        RECT 50.300 2.400 50.440 17.350 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 254.910 84.560 255.230 84.620 ;
        RECT 945.370 84.560 945.690 84.620 ;
        RECT 254.910 84.420 945.690 84.560 ;
        RECT 254.910 84.360 255.230 84.420 ;
        RECT 945.370 84.360 945.690 84.420 ;
        RECT 252.610 17.920 252.930 17.980 ;
        RECT 254.910 17.920 255.230 17.980 ;
        RECT 252.610 17.780 255.230 17.920 ;
        RECT 252.610 17.720 252.930 17.780 ;
        RECT 254.910 17.720 255.230 17.780 ;
      LAYER via ;
        RECT 254.940 84.360 255.200 84.620 ;
        RECT 945.400 84.360 945.660 84.620 ;
        RECT 252.640 17.720 252.900 17.980 ;
        RECT 254.940 17.720 255.200 17.980 ;
      LAYER met2 ;
        RECT 946.030 100.370 946.310 104.000 ;
        RECT 945.460 100.230 946.310 100.370 ;
        RECT 945.460 84.650 945.600 100.230 ;
        RECT 946.030 100.000 946.310 100.230 ;
        RECT 254.940 84.330 255.200 84.650 ;
        RECT 945.400 84.330 945.660 84.650 ;
        RECT 255.000 18.010 255.140 84.330 ;
        RECT 252.640 17.690 252.900 18.010 ;
        RECT 254.940 17.690 255.200 18.010 ;
        RECT 252.700 2.400 252.840 17.690 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 270.090 16.220 270.410 16.280 ;
        RECT 986.770 16.220 987.090 16.280 ;
        RECT 270.090 16.080 987.090 16.220 ;
        RECT 270.090 16.020 270.410 16.080 ;
        RECT 986.770 16.020 987.090 16.080 ;
      LAYER via ;
        RECT 270.120 16.020 270.380 16.280 ;
        RECT 986.800 16.020 987.060 16.280 ;
      LAYER met2 ;
        RECT 991.570 100.370 991.850 104.000 ;
        RECT 986.860 100.230 991.850 100.370 ;
        RECT 986.860 16.310 987.000 100.230 ;
        RECT 991.570 100.000 991.850 100.230 ;
        RECT 270.120 15.990 270.380 16.310 ;
        RECT 986.800 15.990 987.060 16.310 ;
        RECT 270.180 2.400 270.320 15.990 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 289.410 84.900 289.730 84.960 ;
        RECT 1035.990 84.900 1036.310 84.960 ;
        RECT 289.410 84.760 1036.310 84.900 ;
        RECT 289.410 84.700 289.730 84.760 ;
        RECT 1035.990 84.700 1036.310 84.760 ;
      LAYER via ;
        RECT 289.440 84.700 289.700 84.960 ;
        RECT 1036.020 84.700 1036.280 84.960 ;
      LAYER met2 ;
        RECT 1037.570 100.370 1037.850 104.000 ;
        RECT 1036.080 100.230 1037.850 100.370 ;
        RECT 1036.080 84.990 1036.220 100.230 ;
        RECT 1037.570 100.000 1037.850 100.230 ;
        RECT 289.440 84.670 289.700 84.990 ;
        RECT 1036.020 84.670 1036.280 84.990 ;
        RECT 289.500 17.410 289.640 84.670 ;
        RECT 288.120 17.270 289.640 17.410 ;
        RECT 288.120 2.400 288.260 17.270 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 305.970 16.560 306.290 16.620 ;
        RECT 1076.470 16.560 1076.790 16.620 ;
        RECT 305.970 16.420 1076.790 16.560 ;
        RECT 305.970 16.360 306.290 16.420 ;
        RECT 1076.470 16.360 1076.790 16.420 ;
      LAYER via ;
        RECT 306.000 16.360 306.260 16.620 ;
        RECT 1076.500 16.360 1076.760 16.620 ;
      LAYER met2 ;
        RECT 1083.110 100.370 1083.390 104.000 ;
        RECT 1076.560 100.230 1083.390 100.370 ;
        RECT 1076.560 16.650 1076.700 100.230 ;
        RECT 1083.110 100.000 1083.390 100.230 ;
        RECT 306.000 16.330 306.260 16.650 ;
        RECT 1076.500 16.330 1076.760 16.650 ;
        RECT 306.060 2.400 306.200 16.330 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 323.450 85.240 323.770 85.300 ;
        RECT 1127.070 85.240 1127.390 85.300 ;
        RECT 323.450 85.100 1127.390 85.240 ;
        RECT 323.450 85.040 323.770 85.100 ;
        RECT 1127.070 85.040 1127.390 85.100 ;
      LAYER via ;
        RECT 323.480 85.040 323.740 85.300 ;
        RECT 1127.100 85.040 1127.360 85.300 ;
      LAYER met2 ;
        RECT 1128.650 100.370 1128.930 104.000 ;
        RECT 1127.160 100.230 1128.930 100.370 ;
        RECT 1127.160 85.330 1127.300 100.230 ;
        RECT 1128.650 100.000 1128.930 100.230 ;
        RECT 323.480 85.010 323.740 85.330 ;
        RECT 1127.100 85.010 1127.360 85.330 ;
        RECT 323.540 17.410 323.680 85.010 ;
        RECT 323.540 17.270 324.140 17.410 ;
        RECT 324.000 2.400 324.140 17.270 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 365.845 16.745 366.015 20.655 ;
      LAYER mcon ;
        RECT 365.845 20.485 366.015 20.655 ;
      LAYER met1 ;
        RECT 341.390 20.640 341.710 20.700 ;
        RECT 365.785 20.640 366.075 20.685 ;
        RECT 341.390 20.500 366.075 20.640 ;
        RECT 341.390 20.440 341.710 20.500 ;
        RECT 365.785 20.455 366.075 20.500 ;
        RECT 365.785 16.900 366.075 16.945 ;
        RECT 1173.070 16.900 1173.390 16.960 ;
        RECT 365.785 16.760 1173.390 16.900 ;
        RECT 365.785 16.715 366.075 16.760 ;
        RECT 1173.070 16.700 1173.390 16.760 ;
      LAYER via ;
        RECT 341.420 20.440 341.680 20.700 ;
        RECT 1173.100 16.700 1173.360 16.960 ;
      LAYER met2 ;
        RECT 1174.650 100.370 1174.930 104.000 ;
        RECT 1173.160 100.230 1174.930 100.370 ;
        RECT 341.420 20.410 341.680 20.730 ;
        RECT 341.480 2.400 341.620 20.410 ;
        RECT 1173.160 16.990 1173.300 100.230 ;
        RECT 1174.650 100.000 1174.930 100.230 ;
        RECT 1173.100 16.670 1173.360 16.990 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 365.310 85.580 365.630 85.640 ;
        RECT 1218.610 85.580 1218.930 85.640 ;
        RECT 365.310 85.440 1218.930 85.580 ;
        RECT 365.310 85.380 365.630 85.440 ;
        RECT 1218.610 85.380 1218.930 85.440 ;
        RECT 359.330 16.900 359.650 16.960 ;
        RECT 365.310 16.900 365.630 16.960 ;
        RECT 359.330 16.760 365.630 16.900 ;
        RECT 359.330 16.700 359.650 16.760 ;
        RECT 365.310 16.700 365.630 16.760 ;
      LAYER via ;
        RECT 365.340 85.380 365.600 85.640 ;
        RECT 1218.640 85.380 1218.900 85.640 ;
        RECT 359.360 16.700 359.620 16.960 ;
        RECT 365.340 16.700 365.600 16.960 ;
      LAYER met2 ;
        RECT 1220.190 100.370 1220.470 104.000 ;
        RECT 1218.700 100.230 1220.470 100.370 ;
        RECT 1218.700 85.670 1218.840 100.230 ;
        RECT 1220.190 100.000 1220.470 100.230 ;
        RECT 365.340 85.350 365.600 85.670 ;
        RECT 1218.640 85.350 1218.900 85.670 ;
        RECT 365.400 16.990 365.540 85.350 ;
        RECT 359.360 16.670 359.620 16.990 ;
        RECT 365.340 16.670 365.600 16.990 ;
        RECT 359.420 2.400 359.560 16.670 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 377.270 20.640 377.590 20.700 ;
        RECT 1262.770 20.640 1263.090 20.700 ;
        RECT 377.270 20.500 1263.090 20.640 ;
        RECT 377.270 20.440 377.590 20.500 ;
        RECT 1262.770 20.440 1263.090 20.500 ;
      LAYER via ;
        RECT 377.300 20.440 377.560 20.700 ;
        RECT 1262.800 20.440 1263.060 20.700 ;
      LAYER met2 ;
        RECT 1266.190 100.370 1266.470 104.000 ;
        RECT 1262.860 100.230 1266.470 100.370 ;
        RECT 1262.860 20.730 1263.000 100.230 ;
        RECT 1266.190 100.000 1266.470 100.230 ;
        RECT 377.300 20.410 377.560 20.730 ;
        RECT 1262.800 20.410 1263.060 20.730 ;
        RECT 377.360 2.400 377.500 20.410 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 399.810 85.920 400.130 85.980 ;
        RECT 1311.070 85.920 1311.390 85.980 ;
        RECT 399.810 85.780 1311.390 85.920 ;
        RECT 399.810 85.720 400.130 85.780 ;
        RECT 1311.070 85.720 1311.390 85.780 ;
        RECT 395.210 19.960 395.530 20.020 ;
        RECT 399.810 19.960 400.130 20.020 ;
        RECT 395.210 19.820 400.130 19.960 ;
        RECT 395.210 19.760 395.530 19.820 ;
        RECT 399.810 19.760 400.130 19.820 ;
      LAYER via ;
        RECT 399.840 85.720 400.100 85.980 ;
        RECT 1311.100 85.720 1311.360 85.980 ;
        RECT 395.240 19.760 395.500 20.020 ;
        RECT 399.840 19.760 400.100 20.020 ;
      LAYER met2 ;
        RECT 1311.730 100.370 1312.010 104.000 ;
        RECT 1311.160 100.230 1312.010 100.370 ;
        RECT 1311.160 86.010 1311.300 100.230 ;
        RECT 1311.730 100.000 1312.010 100.230 ;
        RECT 399.840 85.690 400.100 86.010 ;
        RECT 1311.100 85.690 1311.360 86.010 ;
        RECT 399.900 20.050 400.040 85.690 ;
        RECT 395.240 19.730 395.500 20.050 ;
        RECT 399.840 19.730 400.100 20.050 ;
        RECT 395.300 2.400 395.440 19.730 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 421.045 19.805 421.215 20.995 ;
        RECT 434.845 19.125 435.015 20.995 ;
        RECT 461.065 19.125 461.235 20.315 ;
      LAYER mcon ;
        RECT 421.045 20.825 421.215 20.995 ;
        RECT 434.845 20.825 435.015 20.995 ;
        RECT 461.065 20.145 461.235 20.315 ;
      LAYER met1 ;
        RECT 420.985 20.980 421.275 21.025 ;
        RECT 434.785 20.980 435.075 21.025 ;
        RECT 420.985 20.840 435.075 20.980 ;
        RECT 420.985 20.795 421.275 20.840 ;
        RECT 434.785 20.795 435.075 20.840 ;
        RECT 461.005 20.300 461.295 20.345 ;
        RECT 1352.470 20.300 1352.790 20.360 ;
        RECT 461.005 20.160 1352.790 20.300 ;
        RECT 461.005 20.115 461.295 20.160 ;
        RECT 1352.470 20.100 1352.790 20.160 ;
        RECT 413.150 19.960 413.470 20.020 ;
        RECT 420.985 19.960 421.275 20.005 ;
        RECT 413.150 19.820 421.275 19.960 ;
        RECT 413.150 19.760 413.470 19.820 ;
        RECT 420.985 19.775 421.275 19.820 ;
        RECT 434.785 19.280 435.075 19.325 ;
        RECT 461.005 19.280 461.295 19.325 ;
        RECT 434.785 19.140 461.295 19.280 ;
        RECT 434.785 19.095 435.075 19.140 ;
        RECT 461.005 19.095 461.295 19.140 ;
      LAYER via ;
        RECT 1352.500 20.100 1352.760 20.360 ;
        RECT 413.180 19.760 413.440 20.020 ;
      LAYER met2 ;
        RECT 1357.730 100.370 1358.010 104.000 ;
        RECT 1352.560 100.230 1358.010 100.370 ;
        RECT 1352.560 20.390 1352.700 100.230 ;
        RECT 1357.730 100.000 1358.010 100.230 ;
        RECT 1352.500 20.070 1352.760 20.390 ;
        RECT 413.180 19.730 413.440 20.050 ;
        RECT 413.240 2.400 413.380 19.730 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 75.510 86.600 75.830 86.660 ;
        RECT 532.750 86.600 533.070 86.660 ;
        RECT 75.510 86.460 533.070 86.600 ;
        RECT 75.510 86.400 75.830 86.460 ;
        RECT 532.750 86.400 533.070 86.460 ;
      LAYER via ;
        RECT 75.540 86.400 75.800 86.660 ;
        RECT 532.780 86.400 533.040 86.660 ;
      LAYER met2 ;
        RECT 534.330 100.370 534.610 104.000 ;
        RECT 532.840 100.230 534.610 100.370 ;
        RECT 532.840 86.690 532.980 100.230 ;
        RECT 534.330 100.000 534.610 100.230 ;
        RECT 75.540 86.370 75.800 86.690 ;
        RECT 532.780 86.370 533.040 86.690 ;
        RECT 75.600 17.410 75.740 86.370 ;
        RECT 74.220 17.270 75.740 17.410 ;
        RECT 74.220 2.400 74.360 17.270 ;
        RECT 74.010 -4.800 74.570 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 434.310 89.660 434.630 89.720 ;
        RECT 1401.690 89.660 1402.010 89.720 ;
        RECT 434.310 89.520 1402.010 89.660 ;
        RECT 434.310 89.460 434.630 89.520 ;
        RECT 1401.690 89.460 1402.010 89.520 ;
        RECT 430.630 19.280 430.950 19.340 ;
        RECT 434.310 19.280 434.630 19.340 ;
        RECT 430.630 19.140 434.630 19.280 ;
        RECT 430.630 19.080 430.950 19.140 ;
        RECT 434.310 19.080 434.630 19.140 ;
      LAYER via ;
        RECT 434.340 89.460 434.600 89.720 ;
        RECT 1401.720 89.460 1401.980 89.720 ;
        RECT 430.660 19.080 430.920 19.340 ;
        RECT 434.340 19.080 434.600 19.340 ;
      LAYER met2 ;
        RECT 1403.270 100.370 1403.550 104.000 ;
        RECT 1401.780 100.230 1403.550 100.370 ;
        RECT 1401.780 89.750 1401.920 100.230 ;
        RECT 1403.270 100.000 1403.550 100.230 ;
        RECT 434.340 89.430 434.600 89.750 ;
        RECT 1401.720 89.430 1401.980 89.750 ;
        RECT 434.400 19.370 434.540 89.430 ;
        RECT 430.660 19.050 430.920 19.370 ;
        RECT 434.340 19.050 434.600 19.370 ;
        RECT 430.720 2.400 430.860 19.050 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1449.070 19.960 1449.390 20.020 ;
        RECT 489.140 19.820 1449.390 19.960 ;
        RECT 448.570 19.620 448.890 19.680 ;
        RECT 489.140 19.620 489.280 19.820 ;
        RECT 1449.070 19.760 1449.390 19.820 ;
        RECT 448.570 19.480 489.280 19.620 ;
        RECT 448.570 19.420 448.890 19.480 ;
      LAYER via ;
        RECT 448.600 19.420 448.860 19.680 ;
        RECT 1449.100 19.760 1449.360 20.020 ;
      LAYER met2 ;
        RECT 1449.270 100.370 1449.550 104.000 ;
        RECT 1449.160 100.000 1449.550 100.370 ;
        RECT 1449.160 20.050 1449.300 100.000 ;
        RECT 1449.100 19.730 1449.360 20.050 ;
        RECT 448.600 19.390 448.860 19.710 ;
        RECT 448.660 2.400 448.800 19.390 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 468.810 89.320 469.130 89.380 ;
        RECT 1493.230 89.320 1493.550 89.380 ;
        RECT 468.810 89.180 1493.550 89.320 ;
        RECT 468.810 89.120 469.130 89.180 ;
        RECT 1493.230 89.120 1493.550 89.180 ;
        RECT 466.510 19.280 466.830 19.340 ;
        RECT 468.810 19.280 469.130 19.340 ;
        RECT 466.510 19.140 469.130 19.280 ;
        RECT 466.510 19.080 466.830 19.140 ;
        RECT 468.810 19.080 469.130 19.140 ;
      LAYER via ;
        RECT 468.840 89.120 469.100 89.380 ;
        RECT 1493.260 89.120 1493.520 89.380 ;
        RECT 466.540 19.080 466.800 19.340 ;
        RECT 468.840 19.080 469.100 19.340 ;
      LAYER met2 ;
        RECT 1494.810 100.370 1495.090 104.000 ;
        RECT 1493.320 100.230 1495.090 100.370 ;
        RECT 1493.320 89.410 1493.460 100.230 ;
        RECT 1494.810 100.000 1495.090 100.230 ;
        RECT 468.840 89.090 469.100 89.410 ;
        RECT 1493.260 89.090 1493.520 89.410 ;
        RECT 468.900 19.370 469.040 89.090 ;
        RECT 466.540 19.050 466.800 19.370 ;
        RECT 468.840 19.050 469.100 19.370 ;
        RECT 466.600 2.400 466.740 19.050 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 489.510 19.620 489.830 19.680 ;
        RECT 1538.770 19.620 1539.090 19.680 ;
        RECT 489.510 19.480 1539.090 19.620 ;
        RECT 489.510 19.420 489.830 19.480 ;
        RECT 1538.770 19.420 1539.090 19.480 ;
        RECT 484.450 14.860 484.770 14.920 ;
        RECT 489.510 14.860 489.830 14.920 ;
        RECT 484.450 14.720 489.830 14.860 ;
        RECT 484.450 14.660 484.770 14.720 ;
        RECT 489.510 14.660 489.830 14.720 ;
      LAYER via ;
        RECT 489.540 19.420 489.800 19.680 ;
        RECT 1538.800 19.420 1539.060 19.680 ;
        RECT 484.480 14.660 484.740 14.920 ;
        RECT 489.540 14.660 489.800 14.920 ;
      LAYER met2 ;
        RECT 1540.350 100.370 1540.630 104.000 ;
        RECT 1538.860 100.230 1540.630 100.370 ;
        RECT 1538.860 19.710 1539.000 100.230 ;
        RECT 1540.350 100.000 1540.630 100.230 ;
        RECT 489.540 19.390 489.800 19.710 ;
        RECT 1538.800 19.390 1539.060 19.710 ;
        RECT 489.600 14.950 489.740 19.390 ;
        RECT 484.480 14.630 484.740 14.950 ;
        RECT 489.540 14.630 489.800 14.950 ;
        RECT 484.540 2.400 484.680 14.630 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 503.310 88.980 503.630 89.040 ;
        RECT 1584.770 88.980 1585.090 89.040 ;
        RECT 503.310 88.840 1585.090 88.980 ;
        RECT 503.310 88.780 503.630 88.840 ;
        RECT 1584.770 88.780 1585.090 88.840 ;
      LAYER via ;
        RECT 503.340 88.780 503.600 89.040 ;
        RECT 1584.800 88.780 1585.060 89.040 ;
      LAYER met2 ;
        RECT 1586.350 100.370 1586.630 104.000 ;
        RECT 1584.860 100.230 1586.630 100.370 ;
        RECT 1584.860 89.070 1585.000 100.230 ;
        RECT 1586.350 100.000 1586.630 100.230 ;
        RECT 503.340 88.750 503.600 89.070 ;
        RECT 1584.800 88.750 1585.060 89.070 ;
        RECT 503.400 17.410 503.540 88.750 ;
        RECT 502.480 17.270 503.540 17.410 ;
        RECT 502.480 2.400 502.620 17.270 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 519.870 19.280 520.190 19.340 ;
        RECT 1628.470 19.280 1628.790 19.340 ;
        RECT 519.870 19.140 1628.790 19.280 ;
        RECT 519.870 19.080 520.190 19.140 ;
        RECT 1628.470 19.080 1628.790 19.140 ;
      LAYER via ;
        RECT 519.900 19.080 520.160 19.340 ;
        RECT 1628.500 19.080 1628.760 19.340 ;
      LAYER met2 ;
        RECT 1631.890 100.370 1632.170 104.000 ;
        RECT 1628.560 100.230 1632.170 100.370 ;
        RECT 1628.560 19.370 1628.700 100.230 ;
        RECT 1631.890 100.000 1632.170 100.230 ;
        RECT 519.900 19.050 520.160 19.370 ;
        RECT 1628.500 19.050 1628.760 19.370 ;
        RECT 519.960 2.400 520.100 19.050 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 537.810 88.640 538.130 88.700 ;
        RECT 1677.230 88.640 1677.550 88.700 ;
        RECT 537.810 88.500 1677.550 88.640 ;
        RECT 537.810 88.440 538.130 88.500 ;
        RECT 1677.230 88.440 1677.550 88.500 ;
      LAYER via ;
        RECT 537.840 88.440 538.100 88.700 ;
        RECT 1677.260 88.440 1677.520 88.700 ;
      LAYER met2 ;
        RECT 1677.890 100.370 1678.170 104.000 ;
        RECT 1677.320 100.230 1678.170 100.370 ;
        RECT 1677.320 88.730 1677.460 100.230 ;
        RECT 1677.890 100.000 1678.170 100.230 ;
        RECT 537.840 88.410 538.100 88.730 ;
        RECT 1677.260 88.410 1677.520 88.730 ;
        RECT 537.900 2.400 538.040 88.410 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 583.885 14.705 584.055 18.955 ;
      LAYER mcon ;
        RECT 583.885 18.785 584.055 18.955 ;
      LAYER met1 ;
        RECT 583.825 18.940 584.115 18.985 ;
        RECT 1718.170 18.940 1718.490 19.000 ;
        RECT 583.825 18.800 1718.490 18.940 ;
        RECT 583.825 18.755 584.115 18.800 ;
        RECT 1718.170 18.740 1718.490 18.800 ;
        RECT 555.750 14.860 556.070 14.920 ;
        RECT 583.825 14.860 584.115 14.905 ;
        RECT 555.750 14.720 584.115 14.860 ;
        RECT 555.750 14.660 556.070 14.720 ;
        RECT 583.825 14.675 584.115 14.720 ;
      LAYER via ;
        RECT 1718.200 18.740 1718.460 19.000 ;
        RECT 555.780 14.660 556.040 14.920 ;
      LAYER met2 ;
        RECT 1723.430 100.370 1723.710 104.000 ;
        RECT 1718.260 100.230 1723.710 100.370 ;
        RECT 1718.260 19.030 1718.400 100.230 ;
        RECT 1723.430 100.000 1723.710 100.230 ;
        RECT 1718.200 18.710 1718.460 19.030 ;
        RECT 555.780 14.630 556.040 14.950 ;
        RECT 555.840 2.400 555.980 14.630 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 579.210 88.300 579.530 88.360 ;
        RECT 1767.850 88.300 1768.170 88.360 ;
        RECT 579.210 88.160 1768.170 88.300 ;
        RECT 579.210 88.100 579.530 88.160 ;
        RECT 1767.850 88.100 1768.170 88.160 ;
        RECT 573.690 18.600 574.010 18.660 ;
        RECT 579.210 18.600 579.530 18.660 ;
        RECT 573.690 18.460 579.530 18.600 ;
        RECT 573.690 18.400 574.010 18.460 ;
        RECT 579.210 18.400 579.530 18.460 ;
      LAYER via ;
        RECT 579.240 88.100 579.500 88.360 ;
        RECT 1767.880 88.100 1768.140 88.360 ;
        RECT 573.720 18.400 573.980 18.660 ;
        RECT 579.240 18.400 579.500 18.660 ;
      LAYER met2 ;
        RECT 1769.430 100.370 1769.710 104.000 ;
        RECT 1767.940 100.230 1769.710 100.370 ;
        RECT 1767.940 88.390 1768.080 100.230 ;
        RECT 1769.430 100.000 1769.710 100.230 ;
        RECT 579.240 88.070 579.500 88.390 ;
        RECT 1767.880 88.070 1768.140 88.390 ;
        RECT 579.300 18.690 579.440 88.070 ;
        RECT 573.720 18.370 573.980 18.690 ;
        RECT 579.240 18.370 579.500 18.690 ;
        RECT 573.780 2.400 573.920 18.370 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 638.165 14.705 638.335 18.615 ;
      LAYER mcon ;
        RECT 638.165 18.445 638.335 18.615 ;
      LAYER met1 ;
        RECT 638.105 18.600 638.395 18.645 ;
        RECT 1814.770 18.600 1815.090 18.660 ;
        RECT 638.105 18.460 1815.090 18.600 ;
        RECT 638.105 18.415 638.395 18.460 ;
        RECT 1814.770 18.400 1815.090 18.460 ;
        RECT 591.170 14.860 591.490 14.920 ;
        RECT 638.105 14.860 638.395 14.905 ;
        RECT 591.170 14.720 638.395 14.860 ;
        RECT 591.170 14.660 591.490 14.720 ;
        RECT 638.105 14.675 638.395 14.720 ;
      LAYER via ;
        RECT 1814.800 18.400 1815.060 18.660 ;
        RECT 591.200 14.660 591.460 14.920 ;
      LAYER met2 ;
        RECT 1814.970 100.370 1815.250 104.000 ;
        RECT 1814.860 100.000 1815.250 100.370 ;
        RECT 1814.860 18.690 1815.000 100.000 ;
        RECT 1814.800 18.370 1815.060 18.690 ;
        RECT 591.200 14.630 591.460 14.950 ;
        RECT 591.260 2.400 591.400 14.630 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 565.945 14.365 566.115 18.615 ;
      LAYER mcon ;
        RECT 565.945 18.445 566.115 18.615 ;
      LAYER met1 ;
        RECT 97.590 18.600 97.910 18.660 ;
        RECT 565.885 18.600 566.175 18.645 ;
        RECT 97.590 18.460 566.175 18.600 ;
        RECT 97.590 18.400 97.910 18.460 ;
        RECT 565.885 18.415 566.175 18.460 ;
        RECT 565.885 14.520 566.175 14.565 ;
        RECT 579.670 14.520 579.990 14.580 ;
        RECT 565.885 14.380 579.990 14.520 ;
        RECT 565.885 14.335 566.175 14.380 ;
        RECT 579.670 14.320 579.990 14.380 ;
      LAYER via ;
        RECT 97.620 18.400 97.880 18.660 ;
        RECT 579.700 14.320 579.960 14.580 ;
      LAYER met2 ;
        RECT 579.870 100.370 580.150 104.000 ;
        RECT 579.760 100.000 580.150 100.370 ;
        RECT 97.620 18.370 97.880 18.690 ;
        RECT 97.680 2.400 97.820 18.370 ;
        RECT 579.760 14.610 579.900 100.000 ;
        RECT 579.700 14.290 579.960 14.610 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 613.710 87.960 614.030 88.020 ;
        RECT 1859.390 87.960 1859.710 88.020 ;
        RECT 613.710 87.820 1859.710 87.960 ;
        RECT 613.710 87.760 614.030 87.820 ;
        RECT 1859.390 87.760 1859.710 87.820 ;
        RECT 609.110 18.600 609.430 18.660 ;
        RECT 613.710 18.600 614.030 18.660 ;
        RECT 609.110 18.460 614.030 18.600 ;
        RECT 609.110 18.400 609.430 18.460 ;
        RECT 613.710 18.400 614.030 18.460 ;
      LAYER via ;
        RECT 613.740 87.760 614.000 88.020 ;
        RECT 1859.420 87.760 1859.680 88.020 ;
        RECT 609.140 18.400 609.400 18.660 ;
        RECT 613.740 18.400 614.000 18.660 ;
      LAYER met2 ;
        RECT 1860.970 100.370 1861.250 104.000 ;
        RECT 1859.480 100.230 1861.250 100.370 ;
        RECT 1859.480 88.050 1859.620 100.230 ;
        RECT 1860.970 100.000 1861.250 100.230 ;
        RECT 613.740 87.730 614.000 88.050 ;
        RECT 1859.420 87.730 1859.680 88.050 ;
        RECT 613.800 18.690 613.940 87.730 ;
        RECT 609.140 18.370 609.400 18.690 ;
        RECT 613.740 18.370 614.000 18.690 ;
        RECT 609.200 2.400 609.340 18.370 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 627.510 87.620 627.830 87.680 ;
        RECT 1904.930 87.620 1905.250 87.680 ;
        RECT 627.510 87.480 1905.250 87.620 ;
        RECT 627.510 87.420 627.830 87.480 ;
        RECT 1904.930 87.420 1905.250 87.480 ;
      LAYER via ;
        RECT 627.540 87.420 627.800 87.680 ;
        RECT 1904.960 87.420 1905.220 87.680 ;
      LAYER met2 ;
        RECT 1906.510 100.370 1906.790 104.000 ;
        RECT 1905.020 100.230 1906.790 100.370 ;
        RECT 1905.020 87.710 1905.160 100.230 ;
        RECT 1906.510 100.000 1906.790 100.230 ;
        RECT 627.540 87.390 627.800 87.710 ;
        RECT 1904.960 87.390 1905.220 87.710 ;
        RECT 627.600 17.410 627.740 87.390 ;
        RECT 627.140 17.270 627.740 17.410 ;
        RECT 627.140 2.400 627.280 17.270 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 123.810 86.260 124.130 86.320 ;
        RECT 623.830 86.260 624.150 86.320 ;
        RECT 123.810 86.120 624.150 86.260 ;
        RECT 123.810 86.060 124.130 86.120 ;
        RECT 623.830 86.060 624.150 86.120 ;
        RECT 121.510 17.920 121.830 17.980 ;
        RECT 123.810 17.920 124.130 17.980 ;
        RECT 121.510 17.780 124.130 17.920 ;
        RECT 121.510 17.720 121.830 17.780 ;
        RECT 123.810 17.720 124.130 17.780 ;
      LAYER via ;
        RECT 123.840 86.060 124.100 86.320 ;
        RECT 623.860 86.060 624.120 86.320 ;
        RECT 121.540 17.720 121.800 17.980 ;
        RECT 123.840 17.720 124.100 17.980 ;
      LAYER met2 ;
        RECT 625.410 100.370 625.690 104.000 ;
        RECT 623.920 100.230 625.690 100.370 ;
        RECT 623.920 86.350 624.060 100.230 ;
        RECT 625.410 100.000 625.690 100.230 ;
        RECT 123.840 86.030 124.100 86.350 ;
        RECT 623.860 86.030 624.120 86.350 ;
        RECT 123.900 18.010 124.040 86.030 ;
        RECT 121.540 17.690 121.800 18.010 ;
        RECT 123.840 17.690 124.100 18.010 ;
        RECT 121.600 2.400 121.740 17.690 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 145.430 15.540 145.750 15.600 ;
        RECT 669.370 15.540 669.690 15.600 ;
        RECT 145.430 15.400 669.690 15.540 ;
        RECT 145.430 15.340 145.750 15.400 ;
        RECT 669.370 15.340 669.690 15.400 ;
      LAYER via ;
        RECT 145.460 15.340 145.720 15.600 ;
        RECT 669.400 15.340 669.660 15.600 ;
      LAYER met2 ;
        RECT 671.410 100.370 671.690 104.000 ;
        RECT 669.460 100.230 671.690 100.370 ;
        RECT 669.460 15.630 669.600 100.230 ;
        RECT 671.410 100.000 671.690 100.230 ;
        RECT 145.460 15.310 145.720 15.630 ;
        RECT 669.400 15.310 669.660 15.630 ;
        RECT 145.520 2.400 145.660 15.310 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 165.210 83.200 165.530 83.260 ;
        RECT 715.370 83.200 715.690 83.260 ;
        RECT 165.210 83.060 715.690 83.200 ;
        RECT 165.210 83.000 165.530 83.060 ;
        RECT 715.370 83.000 715.690 83.060 ;
      LAYER via ;
        RECT 165.240 83.000 165.500 83.260 ;
        RECT 715.400 83.000 715.660 83.260 ;
      LAYER met2 ;
        RECT 716.950 100.370 717.230 104.000 ;
        RECT 715.460 100.230 717.230 100.370 ;
        RECT 715.460 83.290 715.600 100.230 ;
        RECT 716.950 100.000 717.230 100.230 ;
        RECT 165.240 82.970 165.500 83.290 ;
        RECT 715.400 82.970 715.660 83.290 ;
        RECT 165.300 16.730 165.440 82.970 ;
        RECT 163.460 16.590 165.440 16.730 ;
        RECT 163.460 2.400 163.600 16.590 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 180.850 15.880 181.170 15.940 ;
        RECT 759.070 15.880 759.390 15.940 ;
        RECT 180.850 15.740 759.390 15.880 ;
        RECT 180.850 15.680 181.170 15.740 ;
        RECT 759.070 15.680 759.390 15.740 ;
      LAYER via ;
        RECT 180.880 15.680 181.140 15.940 ;
        RECT 759.100 15.680 759.360 15.940 ;
      LAYER met2 ;
        RECT 762.950 100.370 763.230 104.000 ;
        RECT 759.160 100.230 763.230 100.370 ;
        RECT 759.160 15.970 759.300 100.230 ;
        RECT 762.950 100.000 763.230 100.230 ;
        RECT 180.880 15.650 181.140 15.970 ;
        RECT 759.100 15.650 759.360 15.970 ;
        RECT 180.940 2.400 181.080 15.650 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 199.710 83.540 200.030 83.600 ;
        RECT 807.830 83.540 808.150 83.600 ;
        RECT 199.710 83.400 808.150 83.540 ;
        RECT 199.710 83.340 200.030 83.400 ;
        RECT 807.830 83.340 808.150 83.400 ;
      LAYER via ;
        RECT 199.740 83.340 200.000 83.600 ;
        RECT 807.860 83.340 808.120 83.600 ;
      LAYER met2 ;
        RECT 808.490 100.370 808.770 104.000 ;
        RECT 807.920 100.230 808.770 100.370 ;
        RECT 807.920 83.630 808.060 100.230 ;
        RECT 808.490 100.000 808.770 100.230 ;
        RECT 199.740 83.310 200.000 83.630 ;
        RECT 807.860 83.310 808.120 83.630 ;
        RECT 199.800 17.410 199.940 83.310 ;
        RECT 198.880 17.270 199.940 17.410 ;
        RECT 198.880 2.400 199.020 17.270 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 220.410 83.880 220.730 83.940 ;
        RECT 852.910 83.880 853.230 83.940 ;
        RECT 220.410 83.740 853.230 83.880 ;
        RECT 220.410 83.680 220.730 83.740 ;
        RECT 852.910 83.680 853.230 83.740 ;
        RECT 216.730 17.920 217.050 17.980 ;
        RECT 220.410 17.920 220.730 17.980 ;
        RECT 216.730 17.780 220.730 17.920 ;
        RECT 216.730 17.720 217.050 17.780 ;
        RECT 220.410 17.720 220.730 17.780 ;
      LAYER via ;
        RECT 220.440 83.680 220.700 83.940 ;
        RECT 852.940 83.680 853.200 83.940 ;
        RECT 216.760 17.720 217.020 17.980 ;
        RECT 220.440 17.720 220.700 17.980 ;
      LAYER met2 ;
        RECT 854.490 100.370 854.770 104.000 ;
        RECT 853.000 100.230 854.770 100.370 ;
        RECT 853.000 83.970 853.140 100.230 ;
        RECT 854.490 100.000 854.770 100.230 ;
        RECT 220.440 83.650 220.700 83.970 ;
        RECT 852.940 83.650 853.200 83.970 ;
        RECT 220.500 18.010 220.640 83.650 ;
        RECT 216.760 17.690 217.020 18.010 ;
        RECT 220.440 17.690 220.700 18.010 ;
        RECT 216.820 2.400 216.960 17.690 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 240.650 84.220 240.970 84.280 ;
        RECT 898.450 84.220 898.770 84.280 ;
        RECT 240.650 84.080 898.770 84.220 ;
        RECT 240.650 84.020 240.970 84.080 ;
        RECT 898.450 84.020 898.770 84.080 ;
        RECT 234.670 17.920 234.990 17.980 ;
        RECT 240.650 17.920 240.970 17.980 ;
        RECT 234.670 17.780 240.970 17.920 ;
        RECT 234.670 17.720 234.990 17.780 ;
        RECT 240.650 17.720 240.970 17.780 ;
      LAYER via ;
        RECT 240.680 84.020 240.940 84.280 ;
        RECT 898.480 84.020 898.740 84.280 ;
        RECT 234.700 17.720 234.960 17.980 ;
        RECT 240.680 17.720 240.940 17.980 ;
      LAYER met2 ;
        RECT 900.030 100.370 900.310 104.000 ;
        RECT 898.540 100.230 900.310 100.370 ;
        RECT 898.540 84.310 898.680 100.230 ;
        RECT 900.030 100.000 900.310 100.230 ;
        RECT 240.680 83.990 240.940 84.310 ;
        RECT 898.480 83.990 898.740 84.310 ;
        RECT 240.740 18.010 240.880 83.990 ;
        RECT 234.700 17.690 234.960 18.010 ;
        RECT 240.680 17.690 240.940 18.010 ;
        RECT 234.760 2.400 234.900 17.690 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 56.190 17.580 56.510 17.640 ;
        RECT 2773.870 17.580 2774.190 17.640 ;
        RECT 56.190 17.440 2774.190 17.580 ;
        RECT 56.190 17.380 56.510 17.440 ;
        RECT 2773.870 17.380 2774.190 17.440 ;
      LAYER via ;
        RECT 56.220 17.380 56.480 17.640 ;
        RECT 2773.900 17.380 2774.160 17.640 ;
      LAYER met2 ;
        RECT 2775.910 100.370 2776.190 104.000 ;
        RECT 2773.960 100.230 2776.190 100.370 ;
        RECT 2773.960 17.670 2774.100 100.230 ;
        RECT 2775.910 100.000 2776.190 100.230 ;
        RECT 56.220 17.350 56.480 17.670 ;
        RECT 2773.900 17.350 2774.160 17.670 ;
        RECT 56.280 2.400 56.420 17.350 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 80.110 17.240 80.430 17.300 ;
        RECT 2815.270 17.240 2815.590 17.300 ;
        RECT 80.110 17.100 2815.590 17.240 ;
        RECT 80.110 17.040 80.430 17.100 ;
        RECT 2815.270 17.040 2815.590 17.100 ;
      LAYER via ;
        RECT 80.140 17.040 80.400 17.300 ;
        RECT 2815.300 17.040 2815.560 17.300 ;
      LAYER met2 ;
        RECT 2821.450 100.370 2821.730 104.000 ;
        RECT 2815.360 100.230 2821.730 100.370 ;
        RECT 2815.360 17.330 2815.500 100.230 ;
        RECT 2821.450 100.000 2821.730 100.230 ;
        RECT 80.140 17.010 80.400 17.330 ;
        RECT 2815.300 17.010 2815.560 17.330 ;
        RECT 80.200 2.400 80.340 17.010 ;
        RECT 79.990 -4.800 80.550 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 109.090 3433.900 109.410 3433.960 ;
        RECT 2798.710 3433.900 2799.030 3433.960 ;
        RECT 109.090 3433.760 2799.030 3433.900 ;
        RECT 109.090 3433.700 109.410 3433.760 ;
        RECT 2798.710 3433.700 2799.030 3433.760 ;
        RECT 103.570 17.920 103.890 17.980 ;
        RECT 109.090 17.920 109.410 17.980 ;
        RECT 103.570 17.780 109.410 17.920 ;
        RECT 103.570 17.720 103.890 17.780 ;
        RECT 109.090 17.720 109.410 17.780 ;
      LAYER via ;
        RECT 109.120 3433.700 109.380 3433.960 ;
        RECT 2798.740 3433.700 2799.000 3433.960 ;
        RECT 103.600 17.720 103.860 17.980 ;
        RECT 109.120 17.720 109.380 17.980 ;
      LAYER met2 ;
        RECT 109.120 3433.670 109.380 3433.990 ;
        RECT 2798.740 3433.670 2799.000 3433.990 ;
        RECT 109.180 18.010 109.320 3433.670 ;
        RECT 2798.800 3419.450 2798.940 3433.670 ;
        RECT 2800.290 3419.450 2800.570 3420.000 ;
        RECT 2798.800 3419.310 2800.570 3419.450 ;
        RECT 2800.290 3416.000 2800.570 3419.310 ;
        RECT 103.600 17.690 103.860 18.010 ;
        RECT 109.120 17.690 109.380 18.010 ;
        RECT 103.660 2.400 103.800 17.690 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 89.310 16.560 89.630 16.620 ;
        RECT 127.490 16.560 127.810 16.620 ;
        RECT 89.310 16.420 127.810 16.560 ;
        RECT 89.310 16.360 89.630 16.420 ;
        RECT 127.490 16.360 127.810 16.420 ;
      LAYER via ;
        RECT 89.340 16.360 89.600 16.620 ;
        RECT 127.520 16.360 127.780 16.620 ;
      LAYER met2 ;
        RECT 89.330 3087.355 89.610 3087.725 ;
        RECT 89.400 16.650 89.540 3087.355 ;
        RECT 89.340 16.330 89.600 16.650 ;
        RECT 127.520 16.330 127.780 16.650 ;
        RECT 127.580 2.400 127.720 16.330 ;
        RECT 127.370 -4.800 127.930 2.400 ;
      LAYER via2 ;
        RECT 89.330 3087.400 89.610 3087.680 ;
      LAYER met3 ;
        RECT 89.305 3087.690 89.635 3087.705 ;
        RECT 100.000 3087.690 104.000 3087.880 ;
        RECT 89.305 3087.390 104.000 3087.690 ;
        RECT 89.305 3087.375 89.635 3087.390 ;
        RECT 100.000 3087.280 104.000 3087.390 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 27.210 3215.620 27.530 3215.680 ;
        RECT 89.310 3215.620 89.630 3215.680 ;
        RECT 27.210 3215.480 89.630 3215.620 ;
        RECT 27.210 3215.420 27.530 3215.480 ;
        RECT 89.310 3215.420 89.630 3215.480 ;
        RECT 26.290 2.960 26.610 3.020 ;
        RECT 27.210 2.960 27.530 3.020 ;
        RECT 26.290 2.820 27.530 2.960 ;
        RECT 26.290 2.760 26.610 2.820 ;
        RECT 27.210 2.760 27.530 2.820 ;
      LAYER via ;
        RECT 27.240 3215.420 27.500 3215.680 ;
        RECT 89.340 3215.420 89.600 3215.680 ;
        RECT 26.320 2.760 26.580 3.020 ;
        RECT 27.240 2.760 27.500 3.020 ;
      LAYER met2 ;
        RECT 89.330 3219.955 89.610 3220.325 ;
        RECT 89.400 3215.710 89.540 3219.955 ;
        RECT 27.240 3215.390 27.500 3215.710 ;
        RECT 89.340 3215.390 89.600 3215.710 ;
        RECT 27.300 3.050 27.440 3215.390 ;
        RECT 26.320 2.730 26.580 3.050 ;
        RECT 27.240 2.730 27.500 3.050 ;
        RECT 26.380 2.400 26.520 2.730 ;
        RECT 26.170 -4.800 26.730 2.400 ;
      LAYER via2 ;
        RECT 89.330 3220.000 89.610 3220.280 ;
      LAYER met3 ;
        RECT 89.305 3220.290 89.635 3220.305 ;
        RECT 100.000 3220.290 104.000 3220.480 ;
        RECT 89.305 3219.990 104.000 3220.290 ;
        RECT 89.305 3219.975 89.635 3219.990 ;
        RECT 100.000 3219.880 104.000 3219.990 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 34.110 3346.860 34.430 3346.920 ;
        RECT 89.310 3346.860 89.630 3346.920 ;
        RECT 34.110 3346.720 89.630 3346.860 ;
        RECT 34.110 3346.660 34.430 3346.720 ;
        RECT 89.310 3346.660 89.630 3346.720 ;
      LAYER via ;
        RECT 34.140 3346.660 34.400 3346.920 ;
        RECT 89.340 3346.660 89.600 3346.920 ;
      LAYER met2 ;
        RECT 89.330 3352.555 89.610 3352.925 ;
        RECT 89.400 3346.950 89.540 3352.555 ;
        RECT 34.140 3346.630 34.400 3346.950 ;
        RECT 89.340 3346.630 89.600 3346.950 ;
        RECT 34.200 3.130 34.340 3346.630 ;
        RECT 32.360 2.990 34.340 3.130 ;
        RECT 32.360 2.400 32.500 2.990 ;
        RECT 32.150 -4.800 32.710 2.400 ;
      LAYER via2 ;
        RECT 89.330 3352.600 89.610 3352.880 ;
      LAYER met3 ;
        RECT 89.305 3352.890 89.635 3352.905 ;
        RECT 100.000 3352.890 104.000 3353.080 ;
        RECT 89.305 3352.590 104.000 3352.890 ;
        RECT 89.305 3352.575 89.635 3352.590 ;
        RECT 100.000 3352.480 104.000 3352.590 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 185.360 -9.320 188.360 3529.000 ;
        RECT 924.070 -9.320 927.070 3529.000 ;
        RECT 1662.780 -9.320 1665.780 3529.000 ;
        RECT 2401.490 -9.320 2404.490 3529.000 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 186.270 3523.010 187.450 3524.190 ;
        RECT 186.270 3521.410 187.450 3522.590 ;
        RECT 186.270 3431.090 187.450 3432.270 ;
        RECT 186.270 3429.490 187.450 3430.670 ;
        RECT 186.270 11.090 187.450 12.270 ;
        RECT 186.270 9.490 187.450 10.670 ;
        RECT 186.270 -2.910 187.450 -1.730 ;
        RECT 186.270 -4.510 187.450 -3.330 ;
        RECT 924.980 3523.010 926.160 3524.190 ;
        RECT 924.980 3521.410 926.160 3522.590 ;
        RECT 924.980 3431.090 926.160 3432.270 ;
        RECT 924.980 3429.490 926.160 3430.670 ;
        RECT 924.980 11.090 926.160 12.270 ;
        RECT 924.980 9.490 926.160 10.670 ;
        RECT 924.980 -2.910 926.160 -1.730 ;
        RECT 924.980 -4.510 926.160 -3.330 ;
        RECT 1663.690 3523.010 1664.870 3524.190 ;
        RECT 1663.690 3521.410 1664.870 3522.590 ;
        RECT 1663.690 3431.090 1664.870 3432.270 ;
        RECT 1663.690 3429.490 1664.870 3430.670 ;
        RECT 1663.690 11.090 1664.870 12.270 ;
        RECT 1663.690 9.490 1664.870 10.670 ;
        RECT 1663.690 -2.910 1664.870 -1.730 ;
        RECT 1663.690 -4.510 1664.870 -3.330 ;
        RECT 2402.400 3523.010 2403.580 3524.190 ;
        RECT 2402.400 3521.410 2403.580 3522.590 ;
        RECT 2402.400 3431.090 2403.580 3432.270 ;
        RECT 2402.400 3429.490 2403.580 3430.670 ;
        RECT 2402.400 11.090 2403.580 12.270 ;
        RECT 2402.400 9.490 2403.580 10.670 ;
        RECT 2402.400 -2.910 2403.580 -1.730 ;
        RECT 2402.400 -4.510 2403.580 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 185.360 3524.300 188.360 3524.310 ;
        RECT 924.070 3524.300 927.070 3524.310 ;
        RECT 1662.780 3524.300 1665.780 3524.310 ;
        RECT 2401.490 3524.300 2404.490 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 185.360 3521.290 188.360 3521.300 ;
        RECT 924.070 3521.290 927.070 3521.300 ;
        RECT 1662.780 3521.290 1665.780 3521.300 ;
        RECT 2401.490 3521.290 2404.490 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 185.360 3432.380 188.360 3432.390 ;
        RECT 924.070 3432.380 927.070 3432.390 ;
        RECT 1662.780 3432.380 1665.780 3432.390 ;
        RECT 2401.490 3432.380 2404.490 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.680 3429.380 2934.300 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 185.360 3429.370 188.360 3429.380 ;
        RECT 924.070 3429.370 927.070 3429.380 ;
        RECT 1662.780 3429.370 1665.780 3429.380 ;
        RECT 2401.490 3429.370 2404.490 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.680 3249.380 100.000 3252.380 ;
        RECT 2845.000 3249.380 2934.300 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.680 3069.380 100.000 3072.380 ;
        RECT 2845.000 3069.380 2934.300 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.680 2889.380 100.000 2892.380 ;
        RECT 2845.000 2889.380 2934.300 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.680 2709.380 100.000 2712.380 ;
        RECT 2845.000 2709.380 2934.300 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.680 2529.380 100.000 2532.380 ;
        RECT 2845.000 2529.380 2934.300 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.680 2349.380 100.000 2352.380 ;
        RECT 2845.000 2349.380 2934.300 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.680 2169.380 100.000 2172.380 ;
        RECT 2845.000 2169.380 2934.300 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.680 1989.380 100.000 1992.380 ;
        RECT 2845.000 1989.380 2934.300 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.680 1809.380 100.000 1812.380 ;
        RECT 2845.000 1809.380 2934.300 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.680 1629.380 100.000 1632.380 ;
        RECT 2845.000 1629.380 2934.300 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.680 1449.380 100.000 1452.380 ;
        RECT 2845.000 1449.380 2934.300 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.680 1269.380 100.000 1272.380 ;
        RECT 2845.000 1269.380 2934.300 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.680 1089.380 100.000 1092.380 ;
        RECT 2845.000 1089.380 2934.300 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.680 909.380 100.000 912.380 ;
        RECT 2845.000 909.380 2934.300 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.680 729.380 100.000 732.380 ;
        RECT 2845.000 729.380 2934.300 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.680 549.380 100.000 552.380 ;
        RECT 2845.000 549.380 2934.300 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.680 369.380 100.000 372.380 ;
        RECT 2845.000 369.380 2934.300 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.680 189.380 100.000 192.380 ;
        RECT 2845.000 189.380 2934.300 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 185.360 12.380 188.360 12.390 ;
        RECT 924.070 12.380 927.070 12.390 ;
        RECT 1662.780 12.380 1665.780 12.390 ;
        RECT 2401.490 12.380 2404.490 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.680 9.380 2934.300 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 185.360 9.370 188.360 9.380 ;
        RECT 924.070 9.370 927.070 9.380 ;
        RECT 1662.780 9.370 1665.780 9.380 ;
        RECT 2401.490 9.370 2404.490 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 185.360 -1.620 188.360 -1.610 ;
        RECT 924.070 -1.620 927.070 -1.610 ;
        RECT 1662.780 -1.620 1665.780 -1.610 ;
        RECT 2401.490 -1.620 2404.490 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 185.360 -4.630 188.360 -4.620 ;
        RECT 924.070 -4.630 927.070 -4.620 ;
        RECT 1662.780 -4.630 1665.780 -4.620 ;
        RECT 2401.490 -4.630 2404.490 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -14.680 -9.320 -11.680 3529.000 ;
        RECT 554.715 -9.320 557.715 3529.000 ;
        RECT 1293.425 -9.320 1296.425 3529.000 ;
        RECT 2032.135 -9.320 2035.135 3529.000 ;
        RECT 2770.845 -9.320 2773.845 3529.000 ;
        RECT 2931.300 -9.320 2934.300 3529.000 ;
      LAYER via4 ;
        RECT -13.770 3527.710 -12.590 3528.890 ;
        RECT -13.770 3526.110 -12.590 3527.290 ;
        RECT -13.770 3341.090 -12.590 3342.270 ;
        RECT -13.770 3339.490 -12.590 3340.670 ;
        RECT -13.770 3161.090 -12.590 3162.270 ;
        RECT -13.770 3159.490 -12.590 3160.670 ;
        RECT -13.770 2981.090 -12.590 2982.270 ;
        RECT -13.770 2979.490 -12.590 2980.670 ;
        RECT -13.770 2801.090 -12.590 2802.270 ;
        RECT -13.770 2799.490 -12.590 2800.670 ;
        RECT -13.770 2621.090 -12.590 2622.270 ;
        RECT -13.770 2619.490 -12.590 2620.670 ;
        RECT -13.770 2441.090 -12.590 2442.270 ;
        RECT -13.770 2439.490 -12.590 2440.670 ;
        RECT -13.770 2261.090 -12.590 2262.270 ;
        RECT -13.770 2259.490 -12.590 2260.670 ;
        RECT -13.770 2081.090 -12.590 2082.270 ;
        RECT -13.770 2079.490 -12.590 2080.670 ;
        RECT -13.770 1901.090 -12.590 1902.270 ;
        RECT -13.770 1899.490 -12.590 1900.670 ;
        RECT -13.770 1721.090 -12.590 1722.270 ;
        RECT -13.770 1719.490 -12.590 1720.670 ;
        RECT -13.770 1541.090 -12.590 1542.270 ;
        RECT -13.770 1539.490 -12.590 1540.670 ;
        RECT -13.770 1361.090 -12.590 1362.270 ;
        RECT -13.770 1359.490 -12.590 1360.670 ;
        RECT -13.770 1181.090 -12.590 1182.270 ;
        RECT -13.770 1179.490 -12.590 1180.670 ;
        RECT -13.770 1001.090 -12.590 1002.270 ;
        RECT -13.770 999.490 -12.590 1000.670 ;
        RECT -13.770 821.090 -12.590 822.270 ;
        RECT -13.770 819.490 -12.590 820.670 ;
        RECT -13.770 641.090 -12.590 642.270 ;
        RECT -13.770 639.490 -12.590 640.670 ;
        RECT -13.770 461.090 -12.590 462.270 ;
        RECT -13.770 459.490 -12.590 460.670 ;
        RECT -13.770 281.090 -12.590 282.270 ;
        RECT -13.770 279.490 -12.590 280.670 ;
        RECT -13.770 101.090 -12.590 102.270 ;
        RECT -13.770 99.490 -12.590 100.670 ;
        RECT -13.770 -7.610 -12.590 -6.430 ;
        RECT -13.770 -9.210 -12.590 -8.030 ;
        RECT 555.625 3527.710 556.805 3528.890 ;
        RECT 555.625 3526.110 556.805 3527.290 ;
        RECT 555.625 -7.610 556.805 -6.430 ;
        RECT 555.625 -9.210 556.805 -8.030 ;
        RECT 1294.335 3527.710 1295.515 3528.890 ;
        RECT 1294.335 3526.110 1295.515 3527.290 ;
        RECT 1294.335 -7.610 1295.515 -6.430 ;
        RECT 1294.335 -9.210 1295.515 -8.030 ;
        RECT 2033.045 3527.710 2034.225 3528.890 ;
        RECT 2033.045 3526.110 2034.225 3527.290 ;
        RECT 2033.045 -7.610 2034.225 -6.430 ;
        RECT 2033.045 -9.210 2034.225 -8.030 ;
        RECT 2771.755 3527.710 2772.935 3528.890 ;
        RECT 2771.755 3526.110 2772.935 3527.290 ;
        RECT 2771.755 -7.610 2772.935 -6.430 ;
        RECT 2771.755 -9.210 2772.935 -8.030 ;
        RECT 2932.210 3527.710 2933.390 3528.890 ;
        RECT 2932.210 3526.110 2933.390 3527.290 ;
        RECT 2932.210 3341.090 2933.390 3342.270 ;
        RECT 2932.210 3339.490 2933.390 3340.670 ;
        RECT 2932.210 3161.090 2933.390 3162.270 ;
        RECT 2932.210 3159.490 2933.390 3160.670 ;
        RECT 2932.210 2981.090 2933.390 2982.270 ;
        RECT 2932.210 2979.490 2933.390 2980.670 ;
        RECT 2932.210 2801.090 2933.390 2802.270 ;
        RECT 2932.210 2799.490 2933.390 2800.670 ;
        RECT 2932.210 2621.090 2933.390 2622.270 ;
        RECT 2932.210 2619.490 2933.390 2620.670 ;
        RECT 2932.210 2441.090 2933.390 2442.270 ;
        RECT 2932.210 2439.490 2933.390 2440.670 ;
        RECT 2932.210 2261.090 2933.390 2262.270 ;
        RECT 2932.210 2259.490 2933.390 2260.670 ;
        RECT 2932.210 2081.090 2933.390 2082.270 ;
        RECT 2932.210 2079.490 2933.390 2080.670 ;
        RECT 2932.210 1901.090 2933.390 1902.270 ;
        RECT 2932.210 1899.490 2933.390 1900.670 ;
        RECT 2932.210 1721.090 2933.390 1722.270 ;
        RECT 2932.210 1719.490 2933.390 1720.670 ;
        RECT 2932.210 1541.090 2933.390 1542.270 ;
        RECT 2932.210 1539.490 2933.390 1540.670 ;
        RECT 2932.210 1361.090 2933.390 1362.270 ;
        RECT 2932.210 1359.490 2933.390 1360.670 ;
        RECT 2932.210 1181.090 2933.390 1182.270 ;
        RECT 2932.210 1179.490 2933.390 1180.670 ;
        RECT 2932.210 1001.090 2933.390 1002.270 ;
        RECT 2932.210 999.490 2933.390 1000.670 ;
        RECT 2932.210 821.090 2933.390 822.270 ;
        RECT 2932.210 819.490 2933.390 820.670 ;
        RECT 2932.210 641.090 2933.390 642.270 ;
        RECT 2932.210 639.490 2933.390 640.670 ;
        RECT 2932.210 461.090 2933.390 462.270 ;
        RECT 2932.210 459.490 2933.390 460.670 ;
        RECT 2932.210 281.090 2933.390 282.270 ;
        RECT 2932.210 279.490 2933.390 280.670 ;
        RECT 2932.210 101.090 2933.390 102.270 ;
        RECT 2932.210 99.490 2933.390 100.670 ;
        RECT 2932.210 -7.610 2933.390 -6.430 ;
        RECT 2932.210 -9.210 2933.390 -8.030 ;
      LAYER met5 ;
        RECT -14.680 3529.000 -11.680 3529.010 ;
        RECT 554.715 3529.000 557.715 3529.010 ;
        RECT 1293.425 3529.000 1296.425 3529.010 ;
        RECT 2032.135 3529.000 2035.135 3529.010 ;
        RECT 2770.845 3529.000 2773.845 3529.010 ;
        RECT 2931.300 3529.000 2934.300 3529.010 ;
        RECT -14.680 3526.000 2934.300 3529.000 ;
        RECT -14.680 3525.990 -11.680 3526.000 ;
        RECT 554.715 3525.990 557.715 3526.000 ;
        RECT 1293.425 3525.990 1296.425 3526.000 ;
        RECT 2032.135 3525.990 2035.135 3526.000 ;
        RECT 2770.845 3525.990 2773.845 3526.000 ;
        RECT 2931.300 3525.990 2934.300 3526.000 ;
        RECT -14.680 3342.380 -11.680 3342.390 ;
        RECT 2931.300 3342.380 2934.300 3342.390 ;
        RECT -14.680 3339.380 100.000 3342.380 ;
        RECT 2845.000 3339.380 2934.300 3342.380 ;
        RECT -14.680 3339.370 -11.680 3339.380 ;
        RECT 2931.300 3339.370 2934.300 3339.380 ;
        RECT -14.680 3162.380 -11.680 3162.390 ;
        RECT 2931.300 3162.380 2934.300 3162.390 ;
        RECT -14.680 3159.380 100.000 3162.380 ;
        RECT 2845.000 3159.380 2934.300 3162.380 ;
        RECT -14.680 3159.370 -11.680 3159.380 ;
        RECT 2931.300 3159.370 2934.300 3159.380 ;
        RECT -14.680 2982.380 -11.680 2982.390 ;
        RECT 2931.300 2982.380 2934.300 2982.390 ;
        RECT -14.680 2979.380 100.000 2982.380 ;
        RECT 2845.000 2979.380 2934.300 2982.380 ;
        RECT -14.680 2979.370 -11.680 2979.380 ;
        RECT 2931.300 2979.370 2934.300 2979.380 ;
        RECT -14.680 2802.380 -11.680 2802.390 ;
        RECT 2931.300 2802.380 2934.300 2802.390 ;
        RECT -14.680 2799.380 100.000 2802.380 ;
        RECT 2845.000 2799.380 2934.300 2802.380 ;
        RECT -14.680 2799.370 -11.680 2799.380 ;
        RECT 2931.300 2799.370 2934.300 2799.380 ;
        RECT -14.680 2622.380 -11.680 2622.390 ;
        RECT 2931.300 2622.380 2934.300 2622.390 ;
        RECT -14.680 2619.380 100.000 2622.380 ;
        RECT 2845.000 2619.380 2934.300 2622.380 ;
        RECT -14.680 2619.370 -11.680 2619.380 ;
        RECT 2931.300 2619.370 2934.300 2619.380 ;
        RECT -14.680 2442.380 -11.680 2442.390 ;
        RECT 2931.300 2442.380 2934.300 2442.390 ;
        RECT -14.680 2439.380 100.000 2442.380 ;
        RECT 2845.000 2439.380 2934.300 2442.380 ;
        RECT -14.680 2439.370 -11.680 2439.380 ;
        RECT 2931.300 2439.370 2934.300 2439.380 ;
        RECT -14.680 2262.380 -11.680 2262.390 ;
        RECT 2931.300 2262.380 2934.300 2262.390 ;
        RECT -14.680 2259.380 100.000 2262.380 ;
        RECT 2845.000 2259.380 2934.300 2262.380 ;
        RECT -14.680 2259.370 -11.680 2259.380 ;
        RECT 2931.300 2259.370 2934.300 2259.380 ;
        RECT -14.680 2082.380 -11.680 2082.390 ;
        RECT 2931.300 2082.380 2934.300 2082.390 ;
        RECT -14.680 2079.380 100.000 2082.380 ;
        RECT 2845.000 2079.380 2934.300 2082.380 ;
        RECT -14.680 2079.370 -11.680 2079.380 ;
        RECT 2931.300 2079.370 2934.300 2079.380 ;
        RECT -14.680 1902.380 -11.680 1902.390 ;
        RECT 2931.300 1902.380 2934.300 1902.390 ;
        RECT -14.680 1899.380 100.000 1902.380 ;
        RECT 2845.000 1899.380 2934.300 1902.380 ;
        RECT -14.680 1899.370 -11.680 1899.380 ;
        RECT 2931.300 1899.370 2934.300 1899.380 ;
        RECT -14.680 1722.380 -11.680 1722.390 ;
        RECT 2931.300 1722.380 2934.300 1722.390 ;
        RECT -14.680 1719.380 100.000 1722.380 ;
        RECT 2845.000 1719.380 2934.300 1722.380 ;
        RECT -14.680 1719.370 -11.680 1719.380 ;
        RECT 2931.300 1719.370 2934.300 1719.380 ;
        RECT -14.680 1542.380 -11.680 1542.390 ;
        RECT 2931.300 1542.380 2934.300 1542.390 ;
        RECT -14.680 1539.380 100.000 1542.380 ;
        RECT 2845.000 1539.380 2934.300 1542.380 ;
        RECT -14.680 1539.370 -11.680 1539.380 ;
        RECT 2931.300 1539.370 2934.300 1539.380 ;
        RECT -14.680 1362.380 -11.680 1362.390 ;
        RECT 2931.300 1362.380 2934.300 1362.390 ;
        RECT -14.680 1359.380 100.000 1362.380 ;
        RECT 2845.000 1359.380 2934.300 1362.380 ;
        RECT -14.680 1359.370 -11.680 1359.380 ;
        RECT 2931.300 1359.370 2934.300 1359.380 ;
        RECT -14.680 1182.380 -11.680 1182.390 ;
        RECT 2931.300 1182.380 2934.300 1182.390 ;
        RECT -14.680 1179.380 100.000 1182.380 ;
        RECT 2845.000 1179.380 2934.300 1182.380 ;
        RECT -14.680 1179.370 -11.680 1179.380 ;
        RECT 2931.300 1179.370 2934.300 1179.380 ;
        RECT -14.680 1002.380 -11.680 1002.390 ;
        RECT 2931.300 1002.380 2934.300 1002.390 ;
        RECT -14.680 999.380 100.000 1002.380 ;
        RECT 2845.000 999.380 2934.300 1002.380 ;
        RECT -14.680 999.370 -11.680 999.380 ;
        RECT 2931.300 999.370 2934.300 999.380 ;
        RECT -14.680 822.380 -11.680 822.390 ;
        RECT 2931.300 822.380 2934.300 822.390 ;
        RECT -14.680 819.380 100.000 822.380 ;
        RECT 2845.000 819.380 2934.300 822.380 ;
        RECT -14.680 819.370 -11.680 819.380 ;
        RECT 2931.300 819.370 2934.300 819.380 ;
        RECT -14.680 642.380 -11.680 642.390 ;
        RECT 2931.300 642.380 2934.300 642.390 ;
        RECT -14.680 639.380 100.000 642.380 ;
        RECT 2845.000 639.380 2934.300 642.380 ;
        RECT -14.680 639.370 -11.680 639.380 ;
        RECT 2931.300 639.370 2934.300 639.380 ;
        RECT -14.680 462.380 -11.680 462.390 ;
        RECT 2931.300 462.380 2934.300 462.390 ;
        RECT -14.680 459.380 100.000 462.380 ;
        RECT 2845.000 459.380 2934.300 462.380 ;
        RECT -14.680 459.370 -11.680 459.380 ;
        RECT 2931.300 459.370 2934.300 459.380 ;
        RECT -14.680 282.380 -11.680 282.390 ;
        RECT 2931.300 282.380 2934.300 282.390 ;
        RECT -14.680 279.380 100.000 282.380 ;
        RECT 2845.000 279.380 2934.300 282.380 ;
        RECT -14.680 279.370 -11.680 279.380 ;
        RECT 2931.300 279.370 2934.300 279.380 ;
        RECT -14.680 102.380 -11.680 102.390 ;
        RECT 2931.300 102.380 2934.300 102.390 ;
        RECT -14.680 99.380 100.000 102.380 ;
        RECT 2845.000 99.380 2934.300 102.380 ;
        RECT -14.680 99.370 -11.680 99.380 ;
        RECT 2931.300 99.370 2934.300 99.380 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 554.715 -6.320 557.715 -6.310 ;
        RECT 1293.425 -6.320 1296.425 -6.310 ;
        RECT 2032.135 -6.320 2035.135 -6.310 ;
        RECT 2770.845 -6.320 2773.845 -6.310 ;
        RECT 2931.300 -6.320 2934.300 -6.310 ;
        RECT -14.680 -9.320 2934.300 -6.320 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 554.715 -9.330 557.715 -9.320 ;
        RECT 1293.425 -9.330 1296.425 -9.320 ;
        RECT 2032.135 -9.330 2035.135 -9.320 ;
        RECT 2770.845 -9.330 2773.845 -9.320 ;
        RECT 2931.300 -9.330 2934.300 -9.320 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 105.520 110.795 2839.300 3407.605 ;
      LAYER met1 ;
        RECT 105.520 110.640 2839.300 3415.640 ;
      LAYER met2 ;
        RECT 113.440 3415.720 143.970 3416.000 ;
        RECT 144.810 3415.720 232.290 3416.000 ;
        RECT 233.130 3415.720 320.610 3416.000 ;
        RECT 321.450 3415.720 409.390 3416.000 ;
        RECT 410.230 3415.720 497.710 3416.000 ;
        RECT 498.550 3415.720 586.490 3416.000 ;
        RECT 587.330 3415.720 674.810 3416.000 ;
        RECT 675.650 3415.720 763.590 3416.000 ;
        RECT 764.430 3415.720 851.910 3416.000 ;
        RECT 852.750 3415.720 940.690 3416.000 ;
        RECT 941.530 3415.720 1029.010 3416.000 ;
        RECT 1029.850 3415.720 1117.790 3416.000 ;
        RECT 1118.630 3415.720 1206.110 3416.000 ;
        RECT 1206.950 3415.720 1294.890 3416.000 ;
        RECT 1295.730 3415.720 1383.210 3416.000 ;
        RECT 1384.050 3415.720 1471.990 3416.000 ;
        RECT 1472.830 3415.720 1560.310 3416.000 ;
        RECT 1561.150 3415.720 1649.090 3416.000 ;
        RECT 1649.930 3415.720 1737.410 3416.000 ;
        RECT 1738.250 3415.720 1826.190 3416.000 ;
        RECT 1827.030 3415.720 1914.510 3416.000 ;
        RECT 1915.350 3415.720 2003.290 3416.000 ;
        RECT 2004.130 3415.720 2091.610 3416.000 ;
        RECT 2092.450 3415.720 2180.390 3416.000 ;
        RECT 2181.230 3415.720 2268.710 3416.000 ;
        RECT 2269.550 3415.720 2357.490 3416.000 ;
        RECT 2358.330 3415.720 2445.810 3416.000 ;
        RECT 2446.650 3415.720 2534.590 3416.000 ;
        RECT 2535.430 3415.720 2622.910 3416.000 ;
        RECT 2623.750 3415.720 2711.690 3416.000 ;
        RECT 2712.530 3415.720 2800.010 3416.000 ;
        RECT 2800.850 3415.720 2825.410 3416.000 ;
        RECT 113.440 104.280 2825.410 3415.720 ;
        RECT 113.440 104.000 122.350 104.280 ;
        RECT 123.190 104.000 167.890 104.280 ;
        RECT 168.730 104.000 213.430 104.280 ;
        RECT 214.270 104.000 259.430 104.280 ;
        RECT 260.270 104.000 304.970 104.280 ;
        RECT 305.810 104.000 350.970 104.280 ;
        RECT 351.810 104.000 396.510 104.280 ;
        RECT 397.350 104.000 442.510 104.280 ;
        RECT 443.350 104.000 488.050 104.280 ;
        RECT 488.890 104.000 534.050 104.280 ;
        RECT 534.890 104.000 579.590 104.280 ;
        RECT 580.430 104.000 625.130 104.280 ;
        RECT 625.970 104.000 671.130 104.280 ;
        RECT 671.970 104.000 716.670 104.280 ;
        RECT 717.510 104.000 762.670 104.280 ;
        RECT 763.510 104.000 808.210 104.280 ;
        RECT 809.050 104.000 854.210 104.280 ;
        RECT 855.050 104.000 899.750 104.280 ;
        RECT 900.590 104.000 945.750 104.280 ;
        RECT 946.590 104.000 991.290 104.280 ;
        RECT 992.130 104.000 1037.290 104.280 ;
        RECT 1038.130 104.000 1082.830 104.280 ;
        RECT 1083.670 104.000 1128.370 104.280 ;
        RECT 1129.210 104.000 1174.370 104.280 ;
        RECT 1175.210 104.000 1219.910 104.280 ;
        RECT 1220.750 104.000 1265.910 104.280 ;
        RECT 1266.750 104.000 1311.450 104.280 ;
        RECT 1312.290 104.000 1357.450 104.280 ;
        RECT 1358.290 104.000 1402.990 104.280 ;
        RECT 1403.830 104.000 1448.990 104.280 ;
        RECT 1449.830 104.000 1494.530 104.280 ;
        RECT 1495.370 104.000 1540.070 104.280 ;
        RECT 1540.910 104.000 1586.070 104.280 ;
        RECT 1586.910 104.000 1631.610 104.280 ;
        RECT 1632.450 104.000 1677.610 104.280 ;
        RECT 1678.450 104.000 1723.150 104.280 ;
        RECT 1723.990 104.000 1769.150 104.280 ;
        RECT 1769.990 104.000 1814.690 104.280 ;
        RECT 1815.530 104.000 1860.690 104.280 ;
        RECT 1861.530 104.000 1906.230 104.280 ;
        RECT 1907.070 104.000 1952.230 104.280 ;
        RECT 1953.070 104.000 1997.770 104.280 ;
        RECT 1998.610 104.000 2043.310 104.280 ;
        RECT 2044.150 104.000 2089.310 104.280 ;
        RECT 2090.150 104.000 2134.850 104.280 ;
        RECT 2135.690 104.000 2180.850 104.280 ;
        RECT 2181.690 104.000 2226.390 104.280 ;
        RECT 2227.230 104.000 2272.390 104.280 ;
        RECT 2273.230 104.000 2317.930 104.280 ;
        RECT 2318.770 104.000 2363.930 104.280 ;
        RECT 2364.770 104.000 2409.470 104.280 ;
        RECT 2410.310 104.000 2455.010 104.280 ;
        RECT 2455.850 104.000 2501.010 104.280 ;
        RECT 2501.850 104.000 2546.550 104.280 ;
        RECT 2547.390 104.000 2592.550 104.280 ;
        RECT 2593.390 104.000 2638.090 104.280 ;
        RECT 2638.930 104.000 2684.090 104.280 ;
        RECT 2684.930 104.000 2729.630 104.280 ;
        RECT 2730.470 104.000 2775.630 104.280 ;
        RECT 2776.470 104.000 2821.170 104.280 ;
        RECT 2822.010 104.000 2825.410 104.280 ;
      LAYER met3 ;
        RECT 104.000 3360.960 2841.000 3407.685 ;
        RECT 104.000 3359.560 2840.600 3360.960 ;
        RECT 104.000 3353.480 2841.000 3359.560 ;
        RECT 104.400 3352.080 2841.000 3353.480 ;
        RECT 104.000 3242.640 2841.000 3352.080 ;
        RECT 104.000 3241.240 2840.600 3242.640 ;
        RECT 104.000 3220.880 2841.000 3241.240 ;
        RECT 104.400 3219.480 2841.000 3220.880 ;
        RECT 104.000 3123.640 2841.000 3219.480 ;
        RECT 104.000 3122.240 2840.600 3123.640 ;
        RECT 104.000 3088.280 2841.000 3122.240 ;
        RECT 104.400 3086.880 2841.000 3088.280 ;
        RECT 104.000 3005.320 2841.000 3086.880 ;
        RECT 104.000 3003.920 2840.600 3005.320 ;
        RECT 104.000 2955.000 2841.000 3003.920 ;
        RECT 104.400 2953.600 2841.000 2955.000 ;
        RECT 104.000 2887.000 2841.000 2953.600 ;
        RECT 104.000 2885.600 2840.600 2887.000 ;
        RECT 104.000 2822.400 2841.000 2885.600 ;
        RECT 104.400 2821.000 2841.000 2822.400 ;
        RECT 104.000 2768.000 2841.000 2821.000 ;
        RECT 104.000 2766.600 2840.600 2768.000 ;
        RECT 104.000 2689.800 2841.000 2766.600 ;
        RECT 104.400 2688.400 2841.000 2689.800 ;
        RECT 104.000 2649.680 2841.000 2688.400 ;
        RECT 104.000 2648.280 2840.600 2649.680 ;
        RECT 104.000 2557.200 2841.000 2648.280 ;
        RECT 104.400 2555.800 2841.000 2557.200 ;
        RECT 104.000 2531.360 2841.000 2555.800 ;
        RECT 104.000 2529.960 2840.600 2531.360 ;
        RECT 104.000 2423.920 2841.000 2529.960 ;
        RECT 104.400 2422.520 2841.000 2423.920 ;
        RECT 104.000 2412.360 2841.000 2422.520 ;
        RECT 104.000 2410.960 2840.600 2412.360 ;
        RECT 104.000 2294.040 2841.000 2410.960 ;
        RECT 104.000 2292.640 2840.600 2294.040 ;
        RECT 104.000 2291.320 2841.000 2292.640 ;
        RECT 104.400 2289.920 2841.000 2291.320 ;
        RECT 104.000 2175.720 2841.000 2289.920 ;
        RECT 104.000 2174.320 2840.600 2175.720 ;
        RECT 104.000 2158.720 2841.000 2174.320 ;
        RECT 104.400 2157.320 2841.000 2158.720 ;
        RECT 104.000 2056.720 2841.000 2157.320 ;
        RECT 104.000 2055.320 2840.600 2056.720 ;
        RECT 104.000 2025.440 2841.000 2055.320 ;
        RECT 104.400 2024.040 2841.000 2025.440 ;
        RECT 104.000 1938.400 2841.000 2024.040 ;
        RECT 104.000 1937.000 2840.600 1938.400 ;
        RECT 104.000 1892.840 2841.000 1937.000 ;
        RECT 104.400 1891.440 2841.000 1892.840 ;
        RECT 104.000 1820.080 2841.000 1891.440 ;
        RECT 104.000 1818.680 2840.600 1820.080 ;
        RECT 104.000 1760.240 2841.000 1818.680 ;
        RECT 104.400 1758.840 2841.000 1760.240 ;
        RECT 104.000 1701.080 2841.000 1758.840 ;
        RECT 104.000 1699.680 2840.600 1701.080 ;
        RECT 104.000 1627.640 2841.000 1699.680 ;
        RECT 104.400 1626.240 2841.000 1627.640 ;
        RECT 104.000 1582.760 2841.000 1626.240 ;
        RECT 104.000 1581.360 2840.600 1582.760 ;
        RECT 104.000 1494.360 2841.000 1581.360 ;
        RECT 104.400 1492.960 2841.000 1494.360 ;
        RECT 104.000 1463.760 2841.000 1492.960 ;
        RECT 104.000 1462.360 2840.600 1463.760 ;
        RECT 104.000 1361.760 2841.000 1462.360 ;
        RECT 104.400 1360.360 2841.000 1361.760 ;
        RECT 104.000 1345.440 2841.000 1360.360 ;
        RECT 104.000 1344.040 2840.600 1345.440 ;
        RECT 104.000 1229.160 2841.000 1344.040 ;
        RECT 104.400 1227.760 2841.000 1229.160 ;
        RECT 104.000 1227.120 2841.000 1227.760 ;
        RECT 104.000 1225.720 2840.600 1227.120 ;
        RECT 104.000 1108.120 2841.000 1225.720 ;
        RECT 104.000 1106.720 2840.600 1108.120 ;
        RECT 104.000 1095.880 2841.000 1106.720 ;
        RECT 104.400 1094.480 2841.000 1095.880 ;
        RECT 104.000 989.800 2841.000 1094.480 ;
        RECT 104.000 988.400 2840.600 989.800 ;
        RECT 104.000 963.280 2841.000 988.400 ;
        RECT 104.400 961.880 2841.000 963.280 ;
        RECT 104.000 871.480 2841.000 961.880 ;
        RECT 104.000 870.080 2840.600 871.480 ;
        RECT 104.000 830.680 2841.000 870.080 ;
        RECT 104.400 829.280 2841.000 830.680 ;
        RECT 104.000 752.480 2841.000 829.280 ;
        RECT 104.000 751.080 2840.600 752.480 ;
        RECT 104.000 698.080 2841.000 751.080 ;
        RECT 104.400 696.680 2841.000 698.080 ;
        RECT 104.000 634.160 2841.000 696.680 ;
        RECT 104.000 632.760 2840.600 634.160 ;
        RECT 104.000 564.800 2841.000 632.760 ;
        RECT 104.400 563.400 2841.000 564.800 ;
        RECT 104.000 515.840 2841.000 563.400 ;
        RECT 104.000 514.440 2840.600 515.840 ;
        RECT 104.000 432.200 2841.000 514.440 ;
        RECT 104.400 430.800 2841.000 432.200 ;
        RECT 104.000 396.840 2841.000 430.800 ;
        RECT 104.000 395.440 2840.600 396.840 ;
        RECT 104.000 299.600 2841.000 395.440 ;
        RECT 104.400 298.200 2841.000 299.600 ;
        RECT 104.000 278.520 2841.000 298.200 ;
        RECT 104.000 277.120 2840.600 278.520 ;
        RECT 104.000 167.000 2841.000 277.120 ;
        RECT 104.400 165.600 2841.000 167.000 ;
        RECT 104.000 160.200 2841.000 165.600 ;
        RECT 104.000 158.800 2840.600 160.200 ;
        RECT 104.000 104.255 2841.000 158.800 ;
      LAYER met4 ;
        RECT 118.905 110.640 185.360 3407.760 ;
        RECT 188.360 110.640 554.715 3407.760 ;
        RECT 557.715 110.640 924.070 3407.760 ;
        RECT 927.070 110.640 1293.425 3407.760 ;
        RECT 1296.425 110.640 1662.780 3407.760 ;
        RECT 1665.780 110.640 2032.135 3407.760 ;
        RECT 2035.135 110.640 2401.490 3407.760 ;
        RECT 2404.490 110.640 2770.845 3407.760 ;
        RECT 2773.845 110.640 2806.705 3407.760 ;
      LAYER met5 ;
        RECT 105.520 192.700 2839.300 3383.165 ;
      LAYER met5 ;
        RECT 105.520 164.785 2839.300 166.385 ;
        RECT 105.520 126.490 2839.300 128.090 ;
  END
END user_project_wrapper
END LIBRARY


magic
tech sky130A
magscale 1 2
timestamp 1608322654
<< locali >>
rect 567945 656999 567979 661929
rect 567945 637687 567979 642345
rect 567945 618375 567979 623033
rect 567945 598927 567979 607121
rect 567945 560371 567979 563125
rect 567945 550647 567979 553401
rect 568037 502435 568071 505529
rect 568037 495431 568071 502265
rect 25605 3179 25639 3281
rect 51089 2839 51123 3553
rect 73169 3383 73203 4097
rect 84209 3995 84243 4165
rect 86049 3859 86083 4029
rect 86969 3859 87003 4165
rect 92213 3859 92247 4029
rect 113189 2907 113223 3689
rect 116777 2975 116811 3757
rect 127633 2975 127667 3689
<< viali >>
rect 567945 661929 567979 661963
rect 567945 656965 567979 656999
rect 567945 642345 567979 642379
rect 567945 637653 567979 637687
rect 567945 623033 567979 623067
rect 567945 618341 567979 618375
rect 567945 607121 567979 607155
rect 567945 598893 567979 598927
rect 567945 563125 567979 563159
rect 567945 560337 567979 560371
rect 567945 553401 567979 553435
rect 567945 550613 567979 550647
rect 568037 505529 568071 505563
rect 568037 502401 568071 502435
rect 568037 502265 568071 502299
rect 568037 495397 568071 495431
rect 84209 4165 84243 4199
rect 73169 4097 73203 4131
rect 51089 3553 51123 3587
rect 25605 3281 25639 3315
rect 25605 3145 25639 3179
rect 86969 4165 87003 4199
rect 84209 3961 84243 3995
rect 86049 4029 86083 4063
rect 86049 3825 86083 3859
rect 86969 3825 87003 3859
rect 92213 4029 92247 4063
rect 92213 3825 92247 3859
rect 116777 3757 116811 3791
rect 73169 3349 73203 3383
rect 113189 3689 113223 3723
rect 116777 2941 116811 2975
rect 127633 3689 127667 3723
rect 127633 2941 127667 2975
rect 113189 2873 113223 2907
rect 51089 2805 51123 2839
<< metal1 >>
rect 135162 700680 135168 700732
rect 135220 700720 135226 700732
rect 170306 700720 170312 700732
rect 135220 700692 170312 700720
rect 135220 700680 135226 700692
rect 170306 700680 170312 700692
rect 170364 700680 170370 700732
rect 105446 700612 105452 700664
rect 105504 700652 105510 700664
rect 106182 700652 106188 700664
rect 105504 700624 106188 700652
rect 105504 700612 105510 700624
rect 106182 700612 106188 700624
rect 106240 700612 106246 700664
rect 118602 700612 118608 700664
rect 118660 700652 118666 700664
rect 235166 700652 235172 700664
rect 118660 700624 235172 700652
rect 118660 700612 118666 700624
rect 235166 700612 235172 700624
rect 235224 700612 235230 700664
rect 100662 700544 100668 700596
rect 100720 700584 100726 700596
rect 300118 700584 300124 700596
rect 100720 700556 300124 700584
rect 100720 700544 100726 700556
rect 300118 700544 300124 700556
rect 300176 700544 300182 700596
rect 82722 700476 82728 700528
rect 82780 700516 82786 700528
rect 364978 700516 364984 700528
rect 82780 700488 364984 700516
rect 82780 700476 82786 700488
rect 364978 700476 364984 700488
rect 365036 700476 365042 700528
rect 40494 700408 40500 700460
rect 40552 700448 40558 700460
rect 41322 700448 41328 700460
rect 40552 700420 41328 700448
rect 40552 700408 40558 700420
rect 41322 700408 41328 700420
rect 41380 700408 41386 700460
rect 64782 700408 64788 700460
rect 64840 700448 64846 700460
rect 429838 700448 429844 700460
rect 64840 700420 429844 700448
rect 64840 700408 64846 700420
rect 429838 700408 429844 700420
rect 429896 700408 429902 700460
rect 46842 700340 46848 700392
rect 46900 700380 46906 700392
rect 494790 700380 494796 700392
rect 46900 700352 494796 700380
rect 46900 700340 46906 700352
rect 494790 700340 494796 700352
rect 494848 700340 494854 700392
rect 28902 700272 28908 700324
rect 28960 700312 28966 700324
rect 559650 700312 559656 700324
rect 28960 700284 559656 700312
rect 28960 700272 28966 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 82262 687148 82268 687200
rect 82320 687188 82326 687200
rect 82722 687188 82728 687200
rect 82320 687160 82728 687188
rect 82320 687148 82326 687160
rect 82722 687148 82728 687160
rect 82780 687148 82786 687200
rect 117682 687080 117688 687132
rect 117740 687120 117746 687132
rect 118602 687120 118608 687132
rect 117740 687092 118608 687120
rect 117740 687080 117746 687092
rect 118602 687080 118608 687092
rect 118660 687080 118666 687132
rect 99926 686808 99932 686860
rect 99984 686848 99990 686860
rect 100662 686848 100668 686860
rect 99984 686820 100668 686848
rect 99984 686808 99990 686820
rect 100662 686808 100668 686820
rect 100720 686808 100726 686860
rect 21818 686740 21824 686792
rect 21876 686780 21882 686792
rect 559742 686780 559748 686792
rect 21876 686752 559748 686780
rect 21876 686740 21882 686752
rect 559742 686740 559748 686752
rect 559800 686740 559806 686792
rect 106182 686672 106188 686724
rect 106240 686712 106246 686724
rect 152458 686712 152464 686724
rect 106240 686684 152464 686712
rect 106240 686672 106246 686684
rect 152458 686672 152464 686684
rect 152516 686672 152522 686724
rect 41322 686604 41328 686656
rect 41380 686644 41386 686656
rect 170122 686644 170128 686656
rect 41380 686616 170128 686644
rect 41380 686604 41386 686616
rect 170122 686604 170128 686616
rect 170180 686604 170186 686656
rect 21542 686536 21548 686588
rect 21600 686576 21606 686588
rect 205634 686576 205640 686588
rect 21600 686548 205640 686576
rect 21600 686536 21606 686548
rect 205634 686536 205640 686548
rect 205692 686536 205698 686588
rect 21726 686468 21732 686520
rect 21784 686508 21790 686520
rect 276382 686508 276388 686520
rect 21784 686480 276388 686508
rect 21784 686468 21790 686480
rect 276382 686468 276388 686480
rect 276440 686468 276446 686520
rect 9582 686400 9588 686452
rect 9640 686440 9646 686452
rect 364978 686440 364984 686452
rect 9640 686412 364984 686440
rect 9640 686400 9646 686412
rect 364978 686400 364984 686412
rect 365036 686400 365042 686452
rect 13722 686332 13728 686384
rect 13780 686372 13786 686384
rect 382642 686372 382648 686384
rect 13780 686344 382648 686372
rect 13780 686332 13786 686344
rect 382642 686332 382648 686344
rect 382700 686332 382706 686384
rect 21358 686264 21364 686316
rect 21416 686304 21422 686316
rect 400398 686304 400404 686316
rect 21416 686276 400404 686304
rect 21416 686264 21422 686276
rect 400398 686264 400404 686276
rect 400456 686264 400462 686316
rect 188522 686196 188528 686248
rect 188580 686236 188586 686248
rect 567838 686236 567844 686248
rect 188580 686208 567844 686236
rect 188580 686196 188586 686208
rect 567838 686196 567844 686208
rect 567896 686196 567902 686248
rect 21450 686128 21456 686180
rect 21508 686168 21514 686180
rect 418154 686168 418160 686180
rect 21508 686140 418160 686168
rect 21508 686128 21514 686140
rect 418154 686128 418160 686140
rect 418212 686128 418218 686180
rect 21910 686060 21916 686112
rect 21968 686100 21974 686112
rect 436094 686100 436100 686112
rect 21968 686072 436100 686100
rect 21968 686060 21974 686072
rect 436094 686060 436100 686072
rect 436152 686060 436158 686112
rect 21266 685992 21272 686044
rect 21324 686032 21330 686044
rect 453482 686032 453488 686044
rect 21324 686004 453488 686032
rect 21324 685992 21330 686004
rect 453482 685992 453488 686004
rect 453540 685992 453546 686044
rect 21634 685924 21640 685976
rect 21692 685964 21698 685976
rect 488902 685964 488908 685976
rect 21692 685936 488908 685964
rect 21692 685924 21698 685936
rect 488902 685924 488908 685936
rect 488960 685924 488966 685976
rect 6822 669332 6828 669384
rect 6880 669372 6886 669384
rect 17862 669372 17868 669384
rect 6880 669344 17868 669372
rect 6880 669332 6886 669344
rect 17862 669332 17868 669344
rect 17920 669332 17926 669384
rect 3418 667904 3424 667956
rect 3476 667944 3482 667956
rect 19978 667944 19984 667956
rect 3476 667916 19984 667944
rect 3476 667904 3482 667916
rect 19978 667904 19984 667916
rect 20036 667904 20042 667956
rect 567930 661960 567936 661972
rect 567891 661932 567936 661960
rect 567930 661920 567936 661932
rect 567988 661920 567994 661972
rect 567930 656996 567936 657008
rect 567891 656968 567936 656996
rect 567930 656956 567936 656968
rect 567988 656956 567994 657008
rect 5442 643084 5448 643136
rect 5500 643124 5506 643136
rect 17862 643124 17868 643136
rect 5500 643096 17868 643124
rect 5500 643084 5506 643096
rect 17862 643084 17868 643096
rect 17920 643084 17926 643136
rect 567930 642376 567936 642388
rect 567891 642348 567936 642376
rect 567930 642336 567936 642348
rect 567988 642336 567994 642388
rect 567930 637684 567936 637696
rect 567891 637656 567936 637684
rect 567930 637644 567936 637656
rect 567988 637644 567994 637696
rect 567930 623064 567936 623076
rect 567891 623036 567936 623064
rect 567930 623024 567936 623036
rect 567988 623024 567994 623076
rect 567930 618372 567936 618384
rect 567891 618344 567936 618372
rect 567930 618332 567936 618344
rect 567988 618332 567994 618384
rect 3418 609968 3424 610020
rect 3476 610008 3482 610020
rect 15838 610008 15844 610020
rect 3476 609980 15844 610008
rect 3476 609968 3482 609980
rect 15838 609968 15844 609980
rect 15896 609968 15902 610020
rect 567930 607152 567936 607164
rect 567891 607124 567936 607152
rect 567930 607112 567936 607124
rect 567988 607112 567994 607164
rect 567930 598924 567936 598936
rect 567891 598896 567936 598924
rect 567930 598884 567936 598896
rect 567988 598884 567994 598936
rect 567930 572704 567936 572756
rect 567988 572704 567994 572756
rect 567948 572620 567976 572704
rect 567930 572568 567936 572620
rect 567988 572568 567994 572620
rect 567930 563156 567936 563168
rect 567891 563128 567936 563156
rect 567930 563116 567936 563128
rect 567988 563116 567994 563168
rect 567930 560368 567936 560380
rect 567891 560340 567936 560368
rect 567930 560328 567936 560340
rect 567988 560328 567994 560380
rect 567930 553432 567936 553444
rect 567891 553404 567936 553432
rect 567930 553392 567936 553404
rect 567988 553392 567994 553444
rect 3142 552032 3148 552084
rect 3200 552072 3206 552084
rect 18598 552072 18604 552084
rect 3200 552044 18604 552072
rect 3200 552032 3206 552044
rect 18598 552032 18604 552044
rect 18656 552032 18662 552084
rect 567930 550644 567936 550656
rect 567891 550616 567936 550644
rect 567930 550604 567936 550616
rect 567988 550604 567994 550656
rect 567930 534080 567936 534132
rect 567988 534080 567994 534132
rect 567948 533996 567976 534080
rect 567930 533944 567936 533996
rect 567988 533944 567994 533996
rect 567930 514768 567936 514820
rect 567988 514808 567994 514820
rect 567988 514780 568068 514808
rect 567988 514768 567994 514780
rect 568040 514684 568068 514780
rect 568022 514632 568028 514684
rect 568080 514632 568086 514684
rect 568022 505560 568028 505572
rect 567983 505532 568028 505560
rect 568022 505520 568028 505532
rect 568080 505520 568086 505572
rect 568022 502432 568028 502444
rect 567983 502404 568028 502432
rect 568022 502392 568028 502404
rect 568080 502392 568086 502444
rect 568022 502296 568028 502308
rect 567983 502268 568028 502296
rect 568022 502256 568028 502268
rect 568080 502256 568086 502308
rect 567930 495388 567936 495440
rect 567988 495428 567994 495440
rect 568025 495431 568083 495437
rect 568025 495428 568037 495431
rect 567988 495400 568037 495428
rect 567988 495388 567994 495400
rect 568025 495397 568037 495400
rect 568071 495397 568083 495431
rect 568025 495391 568083 495397
rect 579706 487132 579712 487144
rect 567948 487104 579712 487132
rect 567948 487076 567976 487104
rect 579706 487092 579712 487104
rect 579764 487092 579770 487144
rect 567930 487024 567936 487076
rect 567988 487024 567994 487076
rect 3510 437452 3516 437504
rect 3568 437492 3574 437504
rect 7558 437492 7564 437504
rect 3568 437464 7564 437492
rect 3568 437452 3574 437464
rect 7558 437452 7564 437464
rect 7616 437452 7622 437504
rect 573358 391960 573364 392012
rect 573416 392000 573422 392012
rect 579614 392000 579620 392012
rect 573416 391972 579620 392000
rect 573416 391960 573422 391972
rect 579614 391960 579620 391972
rect 579672 391960 579678 392012
rect 13630 351908 13636 351960
rect 13688 351948 13694 351960
rect 17034 351948 17040 351960
rect 13688 351920 17040 351948
rect 13688 351908 13694 351920
rect 17034 351908 17040 351920
rect 17092 351908 17098 351960
rect 577498 345516 577504 345568
rect 577556 345556 577562 345568
rect 579614 345556 579620 345568
rect 577556 345528 579620 345556
rect 577556 345516 577562 345528
rect 579614 345516 579620 345528
rect 579672 345516 579678 345568
rect 8202 324300 8208 324352
rect 8260 324340 8266 324352
rect 17034 324340 17040 324352
rect 8260 324312 17040 324340
rect 8260 324300 8266 324312
rect 17034 324300 17040 324312
rect 17092 324300 17098 324352
rect 3326 322940 3332 322992
rect 3384 322980 3390 322992
rect 10318 322980 10324 322992
rect 3384 322952 10324 322980
rect 3384 322940 3390 322952
rect 10318 322940 10324 322952
rect 10376 322940 10382 322992
rect 14458 298120 14464 298172
rect 14516 298160 14522 298172
rect 17034 298160 17040 298172
rect 14516 298132 17040 298160
rect 14516 298120 14522 298132
rect 17034 298120 17040 298132
rect 17092 298120 17098 298172
rect 574738 298120 574744 298172
rect 574796 298160 574802 298172
rect 579614 298160 579620 298172
rect 574796 298132 579620 298160
rect 574796 298120 574802 298132
rect 579614 298120 579620 298132
rect 579672 298120 579678 298172
rect 11698 271872 11704 271924
rect 11756 271912 11762 271924
rect 17034 271912 17040 271924
rect 11756 271884 17040 271912
rect 11756 271872 11762 271884
rect 17034 271872 17040 271884
rect 17092 271872 17098 271924
rect 576118 251200 576124 251252
rect 576176 251240 576182 251252
rect 579614 251240 579620 251252
rect 576176 251212 579620 251240
rect 576176 251200 576182 251212
rect 579614 251200 579620 251212
rect 579672 251200 579678 251252
rect 14550 245624 14556 245676
rect 14608 245664 14614 245676
rect 17034 245664 17040 245676
rect 14608 245636 17040 245664
rect 14608 245624 14614 245636
rect 17034 245624 17040 245636
rect 17092 245624 17098 245676
rect 571242 244332 571248 244384
rect 571300 244372 571306 244384
rect 578878 244372 578884 244384
rect 571300 244344 578884 244372
rect 571300 244332 571306 244344
rect 578878 244332 578884 244344
rect 578936 244332 578942 244384
rect 571242 221484 571248 221536
rect 571300 221524 571306 221536
rect 573358 221524 573364 221536
rect 571300 221496 573364 221524
rect 571300 221484 571306 221496
rect 573358 221484 573364 221496
rect 573416 221484 573422 221536
rect 11790 218016 11796 218068
rect 11848 218056 11854 218068
rect 17034 218056 17040 218068
rect 11848 218028 17040 218056
rect 11848 218016 11854 218028
rect 17034 218016 17040 218028
rect 17092 218016 17098 218068
rect 573358 204280 573364 204332
rect 573416 204320 573422 204332
rect 579614 204320 579620 204332
rect 573416 204292 579620 204320
rect 573416 204280 573422 204292
rect 579614 204280 579620 204292
rect 579672 204280 579678 204332
rect 571242 197412 571248 197464
rect 571300 197452 571306 197464
rect 577498 197452 577504 197464
rect 571300 197424 577504 197452
rect 571300 197412 571306 197424
rect 577498 197412 577504 197424
rect 577556 197412 577562 197464
rect 3786 191836 3792 191888
rect 3844 191876 3850 191888
rect 17034 191876 17040 191888
rect 3844 191848 17040 191876
rect 3844 191836 3850 191848
rect 17034 191836 17040 191848
rect 17092 191836 17098 191888
rect 571242 174156 571248 174208
rect 571300 174196 571306 174208
rect 574738 174196 574744 174208
rect 571300 174168 574744 174196
rect 571300 174156 571306 174168
rect 574738 174156 574744 174168
rect 574796 174156 574802 174208
rect 3878 166948 3884 167000
rect 3936 166988 3942 167000
rect 17034 166988 17040 167000
rect 3936 166960 17040 166988
rect 3936 166948 3942 166960
rect 17034 166948 17040 166960
rect 17092 166948 17098 167000
rect 574738 157360 574744 157412
rect 574796 157400 574802 157412
rect 579614 157400 579620 157412
rect 574796 157372 579620 157400
rect 574796 157360 574802 157372
rect 579614 157360 579620 157372
rect 579672 157360 579678 157412
rect 571242 150356 571248 150408
rect 571300 150396 571306 150408
rect 576118 150396 576124 150408
rect 571300 150368 576124 150396
rect 571300 150356 571306 150368
rect 576118 150356 576124 150368
rect 576176 150356 576182 150408
rect 3694 140700 3700 140752
rect 3752 140740 3758 140752
rect 16758 140740 16764 140752
rect 3752 140712 16764 140740
rect 3752 140700 3758 140712
rect 16758 140700 16764 140712
rect 16816 140700 16822 140752
rect 571242 126692 571248 126744
rect 571300 126732 571306 126744
rect 573358 126732 573364 126744
rect 571300 126704 573364 126732
rect 571300 126692 571306 126704
rect 573358 126692 573364 126704
rect 573416 126692 573422 126744
rect 3602 113092 3608 113144
rect 3660 113132 3666 113144
rect 17034 113132 17040 113144
rect 3660 113104 17040 113132
rect 3660 113092 3666 113104
rect 17034 113092 17040 113104
rect 17092 113092 17098 113144
rect 573358 110440 573364 110492
rect 573416 110480 573422 110492
rect 579614 110480 579620 110492
rect 573416 110452 579620 110480
rect 573416 110440 573422 110452
rect 579614 110440 579620 110452
rect 579672 110440 579678 110492
rect 3326 108944 3332 108996
rect 3384 108984 3390 108996
rect 11790 108984 11796 108996
rect 3384 108956 11796 108984
rect 3384 108944 3390 108956
rect 11790 108944 11796 108956
rect 11848 108944 11854 108996
rect 571242 103028 571248 103080
rect 571300 103068 571306 103080
rect 574738 103068 574744 103080
rect 571300 103040 574744 103068
rect 571300 103028 571306 103040
rect 574738 103028 574744 103040
rect 574796 103028 574802 103080
rect 10318 86572 10324 86624
rect 10376 86612 10382 86624
rect 17034 86612 17040 86624
rect 10376 86584 17040 86612
rect 10376 86572 10382 86584
rect 17034 86572 17040 86584
rect 17092 86572 17098 86624
rect 571242 79228 571248 79280
rect 571300 79268 571306 79280
rect 573358 79268 573364 79280
rect 571300 79240 573364 79268
rect 571300 79228 571306 79240
rect 573358 79228 573364 79240
rect 573416 79228 573422 79280
rect 3326 64812 3332 64864
rect 3384 64852 3390 64864
rect 14550 64852 14556 64864
rect 3384 64824 14556 64852
rect 3384 64812 3390 64824
rect 14550 64812 14556 64824
rect 14608 64812 14614 64864
rect 577406 63520 577412 63572
rect 577464 63560 577470 63572
rect 580166 63560 580172 63572
rect 577464 63532 580172 63560
rect 577464 63520 577470 63532
rect 580166 63520 580172 63532
rect 580224 63520 580230 63572
rect 3510 60664 3516 60716
rect 3568 60704 3574 60716
rect 16942 60704 16948 60716
rect 3568 60676 16948 60704
rect 3568 60664 3574 60676
rect 16942 60664 16948 60676
rect 17000 60664 17006 60716
rect 571242 55292 571248 55344
rect 571300 55332 571306 55344
rect 577406 55332 577412 55344
rect 571300 55304 577412 55332
rect 571300 55292 571306 55304
rect 577406 55292 577412 55304
rect 577464 55292 577470 55344
rect 7558 34416 7564 34468
rect 7616 34456 7622 34468
rect 17034 34456 17040 34468
rect 7616 34428 17040 34456
rect 7616 34416 7622 34428
rect 17034 34416 17040 34428
rect 17092 34416 17098 34468
rect 3142 22040 3148 22092
rect 3200 22080 3206 22092
rect 11698 22080 11704 22092
rect 3200 22052 11704 22080
rect 3200 22040 3206 22052
rect 11698 22040 11704 22052
rect 11756 22040 11762 22092
rect 19978 20612 19984 20664
rect 20036 20652 20042 20664
rect 24210 20652 24216 20664
rect 20036 20624 24216 20652
rect 20036 20612 20042 20624
rect 24210 20612 24216 20624
rect 24268 20612 24274 20664
rect 21358 20544 21364 20596
rect 21416 20584 21422 20596
rect 27614 20584 27620 20596
rect 21416 20556 27620 20584
rect 21416 20544 21422 20556
rect 27614 20544 27620 20556
rect 27672 20544 27678 20596
rect 22278 19320 22284 19372
rect 22336 19360 22342 19372
rect 22336 19332 24256 19360
rect 22336 19320 22342 19332
rect 22370 19252 22376 19304
rect 22428 19292 22434 19304
rect 24118 19292 24124 19304
rect 22428 19264 24124 19292
rect 22428 19252 22434 19264
rect 24118 19252 24124 19264
rect 24176 19252 24182 19304
rect 24228 19292 24256 19332
rect 24854 19292 24860 19304
rect 24228 19264 24860 19292
rect 24854 19252 24860 19264
rect 24912 19252 24918 19304
rect 61378 19252 61384 19304
rect 61436 19292 61442 19304
rect 580534 19292 580540 19304
rect 61436 19264 580540 19292
rect 61436 19252 61442 19264
rect 580534 19252 580540 19264
rect 580592 19252 580598 19304
rect 70210 19184 70216 19236
rect 70268 19224 70274 19236
rect 580442 19224 580448 19236
rect 70268 19196 580448 19224
rect 70268 19184 70274 19196
rect 580442 19184 580448 19196
rect 580500 19184 580506 19236
rect 79686 19116 79692 19168
rect 79744 19156 79750 19168
rect 580350 19156 580356 19168
rect 79744 19128 580356 19156
rect 79744 19116 79750 19128
rect 580350 19116 580356 19128
rect 580408 19116 580414 19168
rect 88886 19048 88892 19100
rect 88944 19088 88950 19100
rect 580258 19088 580264 19100
rect 88944 19060 580264 19088
rect 88944 19048 88950 19060
rect 580258 19048 580264 19060
rect 580316 19048 580322 19100
rect 22462 17960 22468 18012
rect 22520 18000 22526 18012
rect 22520 17972 23520 18000
rect 22520 17960 22526 17972
rect 23492 17932 23520 17972
rect 26142 17932 26148 17944
rect 23492 17904 26148 17932
rect 26142 17892 26148 17904
rect 26200 17892 26206 17944
rect 86862 17892 86868 17944
rect 86920 17932 86926 17944
rect 280338 17932 280344 17944
rect 86920 17904 280344 17932
rect 86920 17892 86926 17904
rect 280338 17892 280344 17904
rect 280396 17892 280402 17944
rect 573358 17892 573364 17944
rect 573416 17932 573422 17944
rect 579798 17932 579804 17944
rect 573416 17904 579804 17932
rect 573416 17892 573422 17904
rect 579798 17892 579804 17904
rect 579856 17892 579862 17944
rect 18598 17824 18604 17876
rect 18656 17864 18662 17876
rect 42426 17864 42432 17876
rect 18656 17836 42432 17864
rect 18656 17824 18662 17836
rect 42426 17824 42432 17836
rect 42484 17824 42490 17876
rect 93762 17824 93768 17876
rect 93820 17864 93826 17876
rect 298646 17864 298652 17876
rect 93820 17836 298652 17864
rect 93820 17824 93826 17836
rect 298646 17824 298652 17836
rect 298704 17824 298710 17876
rect 15838 17756 15844 17808
rect 15896 17796 15902 17808
rect 33318 17796 33324 17808
rect 15896 17768 33324 17796
rect 15896 17756 15902 17768
rect 33318 17756 33324 17768
rect 33376 17756 33382 17808
rect 100662 17756 100668 17808
rect 100720 17796 100726 17808
rect 316954 17796 316960 17808
rect 100720 17768 316960 17796
rect 100720 17756 100726 17768
rect 316954 17756 316960 17768
rect 317012 17756 317018 17808
rect 3418 17688 3424 17740
rect 3476 17728 3482 17740
rect 51626 17728 51632 17740
rect 3476 17700 51632 17728
rect 3476 17688 3482 17700
rect 51626 17688 51632 17700
rect 51684 17688 51690 17740
rect 107562 17688 107568 17740
rect 107620 17728 107626 17740
rect 335446 17728 335452 17740
rect 107620 17700 335452 17728
rect 107620 17688 107626 17700
rect 335446 17688 335452 17700
rect 335504 17688 335510 17740
rect 115842 17620 115848 17672
rect 115900 17660 115906 17672
rect 353570 17660 353576 17672
rect 115900 17632 353576 17660
rect 115900 17620 115906 17632
rect 353570 17620 353576 17632
rect 353628 17620 353634 17672
rect 122742 17552 122748 17604
rect 122800 17592 122806 17604
rect 371878 17592 371884 17604
rect 122800 17564 371884 17592
rect 122800 17552 122806 17564
rect 371878 17552 371884 17564
rect 371936 17552 371942 17604
rect 10962 17484 10968 17536
rect 11020 17524 11026 17536
rect 97350 17524 97356 17536
rect 11020 17496 97356 17524
rect 11020 17484 11026 17496
rect 97350 17484 97356 17496
rect 97408 17484 97414 17536
rect 125502 17484 125508 17536
rect 125560 17524 125566 17536
rect 380986 17524 380992 17536
rect 125560 17496 380992 17524
rect 125560 17484 125566 17496
rect 380986 17484 380992 17496
rect 381044 17484 381050 17536
rect 34422 17416 34428 17468
rect 34480 17456 34486 17468
rect 408494 17456 408500 17468
rect 34480 17428 408500 17456
rect 34480 17416 34486 17428
rect 408494 17416 408500 17428
rect 408552 17416 408558 17468
rect 41322 17348 41328 17400
rect 41380 17388 41386 17400
rect 417602 17388 417608 17400
rect 41380 17360 417608 17388
rect 41380 17348 41386 17360
rect 417602 17348 417608 17360
rect 417660 17348 417666 17400
rect 15102 17280 15108 17332
rect 15160 17320 15166 17332
rect 106550 17320 106556 17332
rect 15160 17292 106556 17320
rect 15160 17280 15166 17292
rect 106550 17280 106556 17292
rect 106608 17280 106614 17332
rect 117130 17280 117136 17332
rect 117188 17320 117194 17332
rect 536834 17320 536840 17332
rect 117188 17292 536840 17320
rect 117188 17280 117194 17292
rect 536834 17280 536840 17292
rect 536892 17280 536898 17332
rect 24762 17212 24768 17264
rect 24820 17252 24826 17264
rect 124766 17252 124772 17264
rect 24820 17224 124772 17252
rect 24820 17212 24826 17224
rect 124766 17212 124772 17224
rect 124824 17212 124830 17264
rect 125410 17212 125416 17264
rect 125468 17252 125474 17264
rect 545666 17252 545672 17264
rect 125468 17224 545672 17252
rect 125468 17212 125474 17224
rect 545666 17212 545672 17224
rect 545724 17212 545730 17264
rect 79962 17144 79968 17196
rect 80020 17184 80026 17196
rect 262214 17184 262220 17196
rect 80020 17156 262220 17184
rect 80020 17144 80026 17156
rect 262214 17144 262220 17156
rect 262272 17144 262278 17196
rect 73062 17076 73068 17128
rect 73120 17116 73126 17128
rect 243722 17116 243728 17128
rect 73120 17088 243728 17116
rect 73120 17076 73126 17088
rect 243722 17076 243728 17088
rect 243780 17076 243786 17128
rect 64690 17008 64696 17060
rect 64748 17048 64754 17060
rect 225414 17048 225420 17060
rect 64748 17020 225420 17048
rect 64748 17008 64754 17020
rect 225414 17008 225420 17020
rect 225472 17008 225478 17060
rect 57882 16940 57888 16992
rect 57940 16980 57946 16992
rect 207198 16980 207204 16992
rect 57940 16952 207204 16980
rect 57940 16940 57946 16952
rect 207198 16940 207204 16952
rect 207256 16940 207262 16992
rect 50982 16872 50988 16924
rect 51040 16912 51046 16924
rect 189074 16912 189080 16924
rect 51040 16884 189080 16912
rect 51040 16872 51046 16884
rect 189074 16872 189080 16884
rect 189132 16872 189138 16924
rect 48130 16804 48136 16856
rect 48188 16844 48194 16856
rect 179690 16844 179696 16856
rect 48188 16816 179696 16844
rect 48188 16804 48194 16816
rect 179690 16804 179696 16816
rect 179748 16804 179754 16856
rect 44082 16736 44088 16788
rect 44140 16776 44146 16788
rect 170582 16776 170588 16788
rect 44140 16748 170588 16776
rect 44140 16736 44146 16748
rect 170582 16736 170588 16748
rect 170640 16736 170646 16788
rect 39942 16668 39948 16720
rect 40000 16708 40006 16720
rect 161566 16708 161572 16720
rect 40000 16680 161572 16708
rect 40000 16668 40006 16680
rect 161566 16668 161572 16680
rect 161624 16668 161630 16720
rect 33042 16600 33048 16652
rect 33100 16640 33106 16652
rect 143074 16640 143080 16652
rect 33100 16612 143080 16640
rect 33100 16600 33106 16612
rect 143074 16600 143080 16612
rect 143132 16600 143138 16652
rect 24854 10956 24860 11008
rect 24912 10996 24918 11008
rect 28810 10996 28816 11008
rect 24912 10968 28816 10996
rect 24912 10956 24918 10968
rect 28810 10956 28816 10968
rect 28868 10956 28874 11008
rect 26234 10888 26240 10940
rect 26292 10928 26298 10940
rect 27706 10928 27712 10940
rect 26292 10900 27712 10928
rect 26292 10888 26298 10900
rect 27706 10888 27712 10900
rect 27764 10888 27770 10940
rect 22554 9596 22560 9648
rect 22612 9636 22618 9648
rect 24854 9636 24860 9648
rect 22612 9608 24860 9636
rect 22612 9596 22618 9608
rect 24854 9596 24860 9608
rect 24912 9596 24918 9648
rect 28810 8304 28816 8356
rect 28868 8344 28874 8356
rect 28868 8316 29040 8344
rect 28868 8304 28874 8316
rect 29012 8276 29040 8316
rect 33134 8276 33140 8288
rect 29012 8248 33140 8276
rect 33134 8236 33140 8248
rect 33192 8236 33198 8288
rect 27706 8168 27712 8220
rect 27764 8208 27770 8220
rect 29086 8208 29092 8220
rect 27764 8180 29092 8208
rect 27764 8168 27770 8180
rect 29086 8168 29092 8180
rect 29144 8168 29150 8220
rect 123018 6332 123024 6384
rect 123076 6372 123082 6384
rect 571702 6372 571708 6384
rect 123076 6344 571708 6372
rect 123076 6332 123082 6344
rect 571702 6332 571708 6344
rect 571760 6332 571766 6384
rect 77846 6264 77852 6316
rect 77904 6304 77910 6316
rect 571334 6304 571340 6316
rect 77904 6276 571340 6304
rect 77904 6264 77910 6276
rect 571334 6264 571340 6276
rect 571392 6264 571398 6316
rect 67174 6196 67180 6248
rect 67232 6236 67238 6248
rect 571426 6236 571432 6248
rect 67232 6208 571432 6236
rect 67232 6196 67238 6208
rect 571426 6196 571432 6208
rect 571484 6196 571490 6248
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 571610 6168 571616 6180
rect 4120 6140 571616 6168
rect 4120 6128 4126 6140
rect 571610 6128 571616 6140
rect 571668 6128 571674 6180
rect 1670 5448 1676 5500
rect 1728 5488 1734 5500
rect 398834 5488 398840 5500
rect 1728 5460 398840 5488
rect 1728 5448 1734 5460
rect 398834 5448 398840 5460
rect 398892 5448 398898 5500
rect 116026 5380 116032 5432
rect 116084 5420 116090 5432
rect 571794 5420 571800 5432
rect 116084 5392 571800 5420
rect 116084 5380 116090 5392
rect 571794 5380 571800 5392
rect 571852 5380 571858 5432
rect 108758 5312 108764 5364
rect 108816 5352 108822 5364
rect 571886 5352 571892 5364
rect 108816 5324 571892 5352
rect 108816 5312 108822 5324
rect 571886 5312 571892 5324
rect 571944 5312 571950 5364
rect 17218 5244 17224 5296
rect 17276 5284 17282 5296
rect 90910 5284 90916 5296
rect 17276 5256 90916 5284
rect 17276 5244 17282 5256
rect 90910 5244 90916 5256
rect 90968 5244 90974 5296
rect 101582 5244 101588 5296
rect 101640 5284 101646 5296
rect 571978 5284 571984 5296
rect 101640 5256 571984 5284
rect 101640 5244 101646 5256
rect 571978 5244 571984 5256
rect 572036 5244 572042 5296
rect 87322 5176 87328 5228
rect 87380 5216 87386 5228
rect 572070 5216 572076 5228
rect 87380 5188 572076 5216
rect 87380 5176 87386 5188
rect 572070 5176 572076 5188
rect 572128 5176 572134 5228
rect 80238 5108 80244 5160
rect 80296 5148 80302 5160
rect 572162 5148 572168 5160
rect 80296 5120 572168 5148
rect 80296 5108 80302 5120
rect 572162 5108 572168 5120
rect 572220 5108 572226 5160
rect 24854 5040 24860 5092
rect 24912 5080 24918 5092
rect 49602 5080 49608 5092
rect 24912 5052 49608 5080
rect 24912 5040 24918 5052
rect 49602 5040 49608 5052
rect 49660 5040 49666 5092
rect 69474 5040 69480 5092
rect 69532 5080 69538 5092
rect 572254 5080 572260 5092
rect 69532 5052 572260 5080
rect 69532 5040 69538 5052
rect 572254 5040 572260 5052
rect 572312 5040 572318 5092
rect 48222 4972 48228 5024
rect 48280 5012 48286 5024
rect 572346 5012 572352 5024
rect 48280 4984 572352 5012
rect 48280 4972 48286 4984
rect 572346 4972 572352 4984
rect 572404 4972 572410 5024
rect 24118 4904 24124 4956
rect 24176 4944 24182 4956
rect 24854 4944 24860 4956
rect 24176 4916 24860 4944
rect 24176 4904 24182 4916
rect 24854 4904 24860 4916
rect 24912 4904 24918 4956
rect 26694 4904 26700 4956
rect 26752 4944 26758 4956
rect 572438 4944 572444 4956
rect 26752 4916 572444 4944
rect 26752 4904 26758 4916
rect 572438 4904 572444 4916
rect 572496 4904 572502 4956
rect 21910 4836 21916 4888
rect 21968 4876 21974 4888
rect 572530 4876 572536 4888
rect 21968 4848 572536 4876
rect 21968 4836 21974 4848
rect 572530 4836 572536 4848
rect 572588 4836 572594 4888
rect 17218 4768 17224 4820
rect 17276 4808 17282 4820
rect 572622 4808 572628 4820
rect 17276 4780 572628 4808
rect 17276 4768 17282 4780
rect 572622 4768 572628 4780
rect 572680 4768 572686 4820
rect 566 4700 572 4752
rect 624 4740 630 4752
rect 389174 4740 389180 4752
rect 624 4712 389180 4740
rect 624 4700 630 4712
rect 389174 4700 389180 4712
rect 389232 4700 389238 4752
rect 65978 4632 65984 4684
rect 66036 4672 66042 4684
rect 454034 4672 454040 4684
rect 66036 4644 454040 4672
rect 66036 4632 66042 4644
rect 454034 4632 454040 4644
rect 454092 4632 454098 4684
rect 62390 4564 62396 4616
rect 62448 4604 62454 4616
rect 444374 4604 444380 4616
rect 62448 4576 444380 4604
rect 62448 4564 62454 4576
rect 444374 4564 444380 4576
rect 444432 4564 444438 4616
rect 83826 4496 83832 4548
rect 83884 4536 83890 4548
rect 462314 4536 462320 4548
rect 83884 4508 462320 4536
rect 83884 4496 83890 4508
rect 462314 4496 462320 4508
rect 462372 4496 462378 4548
rect 58802 4428 58808 4480
rect 58860 4468 58866 4480
rect 436094 4468 436100 4480
rect 58860 4440 436100 4468
rect 58860 4428 58866 4440
rect 436094 4428 436100 4440
rect 436152 4428 436158 4480
rect 51626 4360 51632 4412
rect 51684 4400 51690 4412
rect 426434 4400 426440 4412
rect 51684 4372 426440 4400
rect 51684 4360 51690 4372
rect 426434 4360 426440 4372
rect 426492 4360 426498 4412
rect 112346 4292 112352 4344
rect 112404 4332 112410 4344
rect 471974 4332 471980 4344
rect 112404 4304 471980 4332
rect 112404 4292 112410 4304
rect 471974 4292 471980 4304
rect 472032 4292 472038 4344
rect 29086 4224 29092 4276
rect 29144 4264 29150 4276
rect 119430 4264 119436 4276
rect 29144 4236 119436 4264
rect 29144 4224 29150 4236
rect 119430 4224 119436 4236
rect 119488 4224 119494 4276
rect 84197 4199 84255 4205
rect 84197 4165 84209 4199
rect 84243 4196 84255 4199
rect 86957 4199 87015 4205
rect 86957 4196 86969 4199
rect 84243 4168 86969 4196
rect 84243 4165 84255 4168
rect 84197 4159 84255 4165
rect 86957 4165 86969 4168
rect 87003 4165 87015 4199
rect 86957 4159 87015 4165
rect 17126 4088 17132 4140
rect 17184 4128 17190 4140
rect 55214 4128 55220 4140
rect 17184 4100 55220 4128
rect 17184 4088 17190 4100
rect 55214 4088 55220 4100
rect 55272 4088 55278 4140
rect 63586 4088 63592 4140
rect 63644 4128 63650 4140
rect 64782 4128 64788 4140
rect 63644 4100 64788 4128
rect 63644 4088 63650 4100
rect 64782 4088 64788 4100
rect 64840 4088 64846 4140
rect 68278 4088 68284 4140
rect 68336 4128 68342 4140
rect 73157 4131 73215 4137
rect 73157 4128 73169 4131
rect 68336 4100 73169 4128
rect 68336 4088 68342 4100
rect 73157 4097 73169 4100
rect 73203 4097 73215 4131
rect 73157 4091 73215 4097
rect 75454 4088 75460 4140
rect 75512 4128 75518 4140
rect 252554 4128 252560 4140
rect 75512 4100 252560 4128
rect 75512 4088 75518 4100
rect 252554 4088 252560 4100
rect 252612 4088 252618 4140
rect 21726 4020 21732 4072
rect 21784 4060 21790 4072
rect 76650 4060 76656 4072
rect 21784 4032 76656 4060
rect 21784 4020 21790 4032
rect 76650 4020 76656 4032
rect 76708 4020 76714 4072
rect 84930 4060 84936 4072
rect 78968 4032 84936 4060
rect 17402 3952 17408 4004
rect 17460 3992 17466 4004
rect 78968 3992 78996 4032
rect 84930 4020 84936 4032
rect 84988 4020 84994 4072
rect 86037 4063 86095 4069
rect 86037 4029 86049 4063
rect 86083 4060 86095 4063
rect 92106 4060 92112 4072
rect 86083 4032 92112 4060
rect 86083 4029 86095 4032
rect 86037 4023 86095 4029
rect 92106 4020 92112 4032
rect 92164 4020 92170 4072
rect 92201 4063 92259 4069
rect 92201 4029 92213 4063
rect 92247 4060 92259 4063
rect 270494 4060 270500 4072
rect 92247 4032 270500 4060
rect 92247 4029 92259 4032
rect 92201 4023 92259 4029
rect 270494 4020 270500 4032
rect 270552 4020 270558 4072
rect 17460 3964 78996 3992
rect 17460 3952 17466 3964
rect 79042 3952 79048 4004
rect 79100 3992 79106 4004
rect 79962 3992 79968 4004
rect 79100 3964 79968 3992
rect 79100 3952 79106 3964
rect 79962 3952 79968 3964
rect 80020 3952 80026 4004
rect 82630 3952 82636 4004
rect 82688 3992 82694 4004
rect 84197 3995 84255 4001
rect 84197 3992 84209 3995
rect 82688 3964 84209 3992
rect 82688 3952 82694 3964
rect 84197 3961 84209 3964
rect 84243 3961 84255 3995
rect 289814 3992 289820 4004
rect 84197 3955 84255 3961
rect 97828 3964 289820 3992
rect 17494 3884 17500 3936
rect 17552 3924 17558 3936
rect 88518 3924 88524 3936
rect 17552 3896 88524 3924
rect 17552 3884 17558 3896
rect 88518 3884 88524 3896
rect 88576 3884 88582 3936
rect 89714 3884 89720 3936
rect 89772 3924 89778 3936
rect 97828 3924 97856 3964
rect 289814 3952 289820 3964
rect 289872 3952 289878 4004
rect 89772 3896 97856 3924
rect 89772 3884 89778 3896
rect 97902 3884 97908 3936
rect 97960 3924 97966 3936
rect 307754 3924 307760 3936
rect 97960 3896 307760 3924
rect 97960 3884 97966 3896
rect 307754 3884 307760 3896
rect 307812 3884 307818 3936
rect 17586 3816 17592 3868
rect 17644 3856 17650 3868
rect 86037 3859 86095 3865
rect 86037 3856 86049 3859
rect 17644 3828 86049 3856
rect 17644 3816 17650 3828
rect 86037 3825 86049 3828
rect 86083 3825 86095 3859
rect 86037 3819 86095 3825
rect 86126 3816 86132 3868
rect 86184 3856 86190 3868
rect 86862 3856 86868 3868
rect 86184 3828 86868 3856
rect 86184 3816 86190 3828
rect 86862 3816 86868 3828
rect 86920 3816 86926 3868
rect 86957 3859 87015 3865
rect 86957 3825 86969 3859
rect 87003 3856 87015 3859
rect 92201 3859 92259 3865
rect 92201 3856 92213 3859
rect 87003 3828 92213 3856
rect 87003 3825 87015 3828
rect 86957 3819 87015 3825
rect 92201 3825 92213 3828
rect 92247 3825 92259 3859
rect 92201 3819 92259 3825
rect 93302 3816 93308 3868
rect 93360 3856 93366 3868
rect 93762 3856 93768 3868
rect 93360 3828 93768 3856
rect 93360 3816 93366 3828
rect 93762 3816 93768 3828
rect 93820 3816 93826 3868
rect 103974 3816 103980 3868
rect 104032 3856 104038 3868
rect 325694 3856 325700 3868
rect 104032 3828 325700 3856
rect 104032 3816 104038 3828
rect 325694 3816 325700 3828
rect 325752 3816 325758 3868
rect 17678 3748 17684 3800
rect 17736 3788 17742 3800
rect 102778 3788 102784 3800
rect 17736 3760 102784 3788
rect 17736 3748 17742 3760
rect 102778 3748 102784 3760
rect 102836 3748 102842 3800
rect 116765 3791 116823 3797
rect 116765 3757 116777 3791
rect 116811 3788 116823 3791
rect 343634 3788 343640 3800
rect 116811 3760 343640 3788
rect 116811 3757 116823 3760
rect 116765 3751 116823 3757
rect 343634 3748 343640 3760
rect 343692 3748 343698 3800
rect 19518 3680 19524 3732
rect 19576 3720 19582 3732
rect 113177 3723 113235 3729
rect 113177 3720 113189 3723
rect 19576 3692 113189 3720
rect 19576 3680 19582 3692
rect 113177 3689 113189 3692
rect 113223 3689 113235 3723
rect 113177 3683 113235 3689
rect 113542 3680 113548 3732
rect 113600 3720 113606 3732
rect 114462 3720 114468 3732
rect 113600 3692 114468 3720
rect 113600 3680 113606 3692
rect 114462 3680 114468 3692
rect 114520 3680 114526 3732
rect 114738 3680 114744 3732
rect 114796 3720 114802 3732
rect 115842 3720 115848 3732
rect 114796 3692 115848 3720
rect 114796 3680 114802 3692
rect 115842 3680 115848 3692
rect 115900 3680 115906 3732
rect 121822 3680 121828 3732
rect 121880 3720 121886 3732
rect 122742 3720 122748 3732
rect 121880 3692 122748 3720
rect 121880 3680 121886 3692
rect 122742 3680 122748 3692
rect 122800 3680 122806 3732
rect 124214 3680 124220 3732
rect 124272 3720 124278 3732
rect 125410 3720 125416 3732
rect 124272 3692 125416 3720
rect 124272 3680 124278 3692
rect 125410 3680 125416 3692
rect 125468 3680 125474 3732
rect 127621 3723 127679 3729
rect 127621 3689 127633 3723
rect 127667 3720 127679 3723
rect 362954 3720 362960 3732
rect 127667 3692 362960 3720
rect 127667 3689 127679 3692
rect 127621 3683 127679 3689
rect 362954 3680 362960 3692
rect 363012 3680 363018 3732
rect 21542 3612 21548 3664
rect 21600 3652 21606 3664
rect 21600 3624 24900 3652
rect 21600 3612 21606 3624
rect 12434 3544 12440 3596
rect 12492 3584 12498 3596
rect 13630 3584 13636 3596
rect 12492 3556 13636 3584
rect 12492 3544 12498 3556
rect 13630 3544 13636 3556
rect 13688 3544 13694 3596
rect 18322 3544 18328 3596
rect 18380 3584 18386 3596
rect 19150 3584 19156 3596
rect 18380 3556 19156 3584
rect 18380 3544 18386 3556
rect 19150 3544 19156 3556
rect 19208 3544 19214 3596
rect 20714 3544 20720 3596
rect 20772 3584 20778 3596
rect 21818 3584 21824 3596
rect 20772 3556 21824 3584
rect 20772 3544 20778 3556
rect 21818 3544 21824 3556
rect 21876 3544 21882 3596
rect 24302 3544 24308 3596
rect 24360 3584 24366 3596
rect 24762 3584 24768 3596
rect 24360 3556 24768 3584
rect 24360 3544 24366 3556
rect 24762 3544 24768 3556
rect 24820 3544 24826 3596
rect 24872 3584 24900 3624
rect 34974 3612 34980 3664
rect 35032 3652 35038 3664
rect 499574 3652 499580 3664
rect 35032 3624 499580 3652
rect 35032 3612 35038 3624
rect 499574 3612 499580 3624
rect 499632 3612 499638 3664
rect 30282 3584 30288 3596
rect 24872 3556 30288 3584
rect 30282 3544 30288 3556
rect 30340 3544 30346 3596
rect 33870 3544 33876 3596
rect 33928 3584 33934 3596
rect 34422 3584 34428 3596
rect 33928 3556 34428 3584
rect 33928 3544 33934 3556
rect 34422 3544 34428 3556
rect 34480 3544 34486 3596
rect 42150 3544 42156 3596
rect 42208 3584 42214 3596
rect 42702 3584 42708 3596
rect 42208 3556 42708 3584
rect 42208 3544 42214 3556
rect 42702 3544 42708 3556
rect 42760 3544 42766 3596
rect 43346 3544 43352 3596
rect 43404 3584 43410 3596
rect 44082 3584 44088 3596
rect 43404 3556 44088 3584
rect 43404 3544 43410 3556
rect 44082 3544 44088 3556
rect 44140 3544 44146 3596
rect 46934 3544 46940 3596
rect 46992 3584 46998 3596
rect 48130 3584 48136 3596
rect 46992 3556 48136 3584
rect 46992 3544 46998 3556
rect 48130 3544 48136 3556
rect 48188 3544 48194 3596
rect 50522 3544 50528 3596
rect 50580 3584 50586 3596
rect 50982 3584 50988 3596
rect 50580 3556 50988 3584
rect 50580 3544 50586 3556
rect 50982 3544 50988 3556
rect 51040 3544 51046 3596
rect 51077 3587 51135 3593
rect 51077 3553 51089 3587
rect 51123 3584 51135 3587
rect 517514 3584 517520 3596
rect 51123 3556 517520 3584
rect 51123 3553 51135 3556
rect 51077 3547 51135 3553
rect 517514 3544 517520 3556
rect 517572 3544 517578 3596
rect 7650 3476 7656 3528
rect 7708 3516 7714 3528
rect 8202 3516 8208 3528
rect 7708 3488 8208 3516
rect 7708 3476 7714 3488
rect 8202 3476 8208 3488
rect 8260 3476 8266 3528
rect 8846 3476 8852 3528
rect 8904 3516 8910 3528
rect 9582 3516 9588 3528
rect 8904 3488 9588 3516
rect 8904 3476 8910 3488
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 10042 3476 10048 3528
rect 10100 3516 10106 3528
rect 10962 3516 10968 3528
rect 10100 3488 10968 3516
rect 10100 3476 10106 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 11238 3476 11244 3528
rect 11296 3516 11302 3528
rect 554774 3516 554780 3528
rect 11296 3488 554780 3516
rect 11296 3476 11302 3488
rect 554774 3476 554780 3488
rect 554832 3476 554838 3528
rect 2866 3408 2872 3460
rect 2924 3448 2930 3460
rect 14458 3448 14464 3460
rect 2924 3420 14464 3448
rect 2924 3408 2930 3420
rect 14458 3408 14464 3420
rect 14516 3408 14522 3460
rect 16022 3408 16028 3460
rect 16080 3448 16086 3460
rect 563054 3448 563060 3460
rect 16080 3420 563060 3448
rect 16080 3408 16086 3420
rect 563054 3408 563060 3420
rect 563112 3408 563118 3460
rect 21266 3340 21272 3392
rect 21324 3380 21330 3392
rect 59998 3380 60004 3392
rect 21324 3352 60004 3380
rect 21324 3340 21330 3352
rect 59998 3340 60004 3352
rect 60056 3340 60062 3392
rect 71866 3340 71872 3392
rect 71924 3380 71930 3392
rect 73062 3380 73068 3392
rect 71924 3352 73068 3380
rect 71924 3340 71930 3352
rect 73062 3340 73068 3352
rect 73120 3340 73126 3392
rect 73157 3383 73215 3389
rect 73157 3349 73169 3383
rect 73203 3380 73215 3383
rect 234614 3380 234620 3392
rect 73203 3352 234620 3380
rect 73203 3349 73215 3352
rect 73157 3343 73215 3349
rect 234614 3340 234620 3352
rect 234672 3340 234678 3392
rect 17862 3272 17868 3324
rect 17920 3312 17926 3324
rect 25498 3312 25504 3324
rect 17920 3284 25504 3312
rect 17920 3272 17926 3284
rect 25498 3272 25504 3284
rect 25556 3272 25562 3324
rect 25593 3315 25651 3321
rect 25593 3281 25605 3315
rect 25639 3312 25651 3315
rect 56410 3312 56416 3324
rect 25639 3284 56416 3312
rect 25639 3281 25651 3284
rect 25593 3275 25651 3281
rect 56410 3272 56416 3284
rect 56468 3272 56474 3324
rect 61194 3272 61200 3324
rect 61252 3312 61258 3324
rect 215294 3312 215300 3324
rect 61252 3284 215300 3312
rect 61252 3272 61258 3284
rect 215294 3272 215300 3284
rect 215352 3272 215358 3324
rect 22002 3204 22008 3256
rect 22060 3244 22066 3256
rect 52822 3244 52828 3256
rect 22060 3216 52828 3244
rect 22060 3204 22066 3216
rect 52822 3204 52828 3216
rect 52880 3204 52886 3256
rect 54018 3204 54024 3256
rect 54076 3244 54082 3256
rect 197354 3244 197360 3256
rect 54076 3216 197360 3244
rect 54076 3204 54082 3216
rect 197354 3204 197360 3216
rect 197412 3204 197418 3256
rect 19242 3136 19248 3188
rect 19300 3176 19306 3188
rect 25593 3179 25651 3185
rect 25593 3176 25605 3179
rect 19300 3148 25605 3176
rect 19300 3136 19306 3148
rect 25593 3145 25605 3148
rect 25639 3145 25651 3179
rect 25593 3139 25651 3145
rect 36170 3136 36176 3188
rect 36228 3176 36234 3188
rect 151814 3176 151820 3188
rect 36228 3148 151820 3176
rect 36228 3136 36234 3148
rect 151814 3136 151820 3148
rect 151872 3136 151878 3188
rect 29086 3068 29092 3120
rect 29144 3108 29150 3120
rect 133874 3108 133880 3120
rect 29144 3080 133880 3108
rect 29144 3068 29150 3080
rect 133874 3068 133880 3080
rect 133932 3068 133938 3120
rect 17770 3000 17776 3052
rect 17828 3040 17834 3052
rect 120626 3040 120632 3052
rect 17828 3012 120632 3040
rect 17828 3000 17834 3012
rect 120626 3000 120632 3012
rect 120684 3000 120690 3052
rect 17310 2932 17316 2984
rect 17368 2972 17374 2984
rect 23106 2972 23112 2984
rect 17368 2944 23112 2972
rect 17368 2932 17374 2944
rect 23106 2932 23112 2944
rect 23164 2932 23170 2984
rect 24854 2932 24860 2984
rect 24912 2972 24918 2984
rect 94498 2972 94504 2984
rect 24912 2944 94504 2972
rect 24912 2932 24918 2944
rect 94498 2932 94504 2944
rect 94556 2932 94562 2984
rect 96890 2932 96896 2984
rect 96948 2972 96954 2984
rect 97902 2972 97908 2984
rect 96948 2944 97908 2972
rect 96948 2932 96954 2944
rect 97902 2932 97908 2944
rect 97960 2932 97966 2984
rect 111150 2932 111156 2984
rect 111208 2972 111214 2984
rect 116765 2975 116823 2981
rect 116765 2972 116777 2975
rect 111208 2944 116777 2972
rect 111208 2932 111214 2944
rect 116765 2941 116777 2944
rect 116811 2941 116823 2975
rect 116765 2935 116823 2941
rect 118234 2932 118240 2984
rect 118292 2972 118298 2984
rect 127621 2975 127679 2981
rect 127621 2972 127633 2975
rect 118292 2944 127633 2972
rect 118292 2932 118298 2944
rect 127621 2941 127633 2944
rect 127667 2941 127679 2975
rect 127621 2935 127679 2941
rect 33134 2864 33140 2916
rect 33192 2904 33198 2916
rect 98086 2904 98092 2916
rect 33192 2876 98092 2904
rect 33192 2864 33198 2876
rect 98086 2864 98092 2876
rect 98144 2864 98150 2916
rect 113177 2907 113235 2913
rect 113177 2873 113189 2907
rect 113223 2904 113235 2907
rect 115934 2904 115940 2916
rect 113223 2876 115940 2904
rect 113223 2873 113235 2876
rect 113177 2867 113235 2873
rect 115934 2864 115940 2876
rect 115992 2864 115998 2916
rect 21450 2796 21456 2848
rect 21508 2836 21514 2848
rect 49326 2836 49332 2848
rect 21508 2808 49332 2836
rect 21508 2796 21514 2808
rect 49326 2796 49332 2808
rect 49384 2796 49390 2848
rect 51077 2839 51135 2845
rect 51077 2836 51089 2839
rect 49436 2808 51089 2836
rect 45738 2728 45744 2780
rect 45796 2768 45802 2780
rect 49436 2768 49464 2808
rect 51077 2805 51089 2808
rect 51123 2805 51135 2839
rect 105170 2836 105176 2848
rect 51077 2799 51135 2805
rect 51184 2808 105176 2836
rect 45796 2740 49464 2768
rect 45796 2728 45802 2740
rect 49602 2728 49608 2780
rect 49660 2768 49666 2780
rect 51184 2768 51212 2808
rect 105170 2796 105176 2808
rect 105228 2796 105234 2848
rect 49660 2740 51212 2768
rect 49660 2728 49666 2740
rect 5258 552 5264 604
rect 5316 592 5322 604
rect 5442 592 5448 604
rect 5316 564 5448 592
rect 5316 552 5322 564
rect 5442 552 5448 564
rect 5500 552 5506 604
<< via1 >>
rect 135168 700680 135220 700732
rect 170312 700680 170364 700732
rect 105452 700612 105504 700664
rect 106188 700612 106240 700664
rect 118608 700612 118660 700664
rect 235172 700612 235224 700664
rect 100668 700544 100720 700596
rect 300124 700544 300176 700596
rect 82728 700476 82780 700528
rect 364984 700476 365036 700528
rect 40500 700408 40552 700460
rect 41328 700408 41380 700460
rect 64788 700408 64840 700460
rect 429844 700408 429896 700460
rect 46848 700340 46900 700392
rect 494796 700340 494848 700392
rect 28908 700272 28960 700324
rect 559656 700272 559708 700324
rect 82268 687148 82320 687200
rect 82728 687148 82780 687200
rect 117688 687080 117740 687132
rect 118608 687080 118660 687132
rect 99932 686808 99984 686860
rect 100668 686808 100720 686860
rect 21824 686740 21876 686792
rect 559748 686740 559800 686792
rect 106188 686672 106240 686724
rect 152464 686672 152516 686724
rect 41328 686604 41380 686656
rect 170128 686604 170180 686656
rect 21548 686536 21600 686588
rect 205640 686536 205692 686588
rect 21732 686468 21784 686520
rect 276388 686468 276440 686520
rect 9588 686400 9640 686452
rect 364984 686400 365036 686452
rect 13728 686332 13780 686384
rect 382648 686332 382700 686384
rect 21364 686264 21416 686316
rect 400404 686264 400456 686316
rect 188528 686196 188580 686248
rect 567844 686196 567896 686248
rect 21456 686128 21508 686180
rect 418160 686128 418212 686180
rect 21916 686060 21968 686112
rect 436100 686060 436152 686112
rect 21272 685992 21324 686044
rect 453488 685992 453540 686044
rect 21640 685924 21692 685976
rect 488908 685924 488960 685976
rect 6828 669332 6880 669384
rect 17868 669332 17920 669384
rect 3424 667904 3476 667956
rect 19984 667904 20036 667956
rect 567936 661963 567988 661972
rect 567936 661929 567945 661963
rect 567945 661929 567979 661963
rect 567979 661929 567988 661963
rect 567936 661920 567988 661929
rect 567936 656999 567988 657008
rect 567936 656965 567945 656999
rect 567945 656965 567979 656999
rect 567979 656965 567988 656999
rect 567936 656956 567988 656965
rect 5448 643084 5500 643136
rect 17868 643084 17920 643136
rect 567936 642379 567988 642388
rect 567936 642345 567945 642379
rect 567945 642345 567979 642379
rect 567979 642345 567988 642379
rect 567936 642336 567988 642345
rect 567936 637687 567988 637696
rect 567936 637653 567945 637687
rect 567945 637653 567979 637687
rect 567979 637653 567988 637687
rect 567936 637644 567988 637653
rect 567936 623067 567988 623076
rect 567936 623033 567945 623067
rect 567945 623033 567979 623067
rect 567979 623033 567988 623067
rect 567936 623024 567988 623033
rect 567936 618375 567988 618384
rect 567936 618341 567945 618375
rect 567945 618341 567979 618375
rect 567979 618341 567988 618375
rect 567936 618332 567988 618341
rect 3424 609968 3476 610020
rect 15844 609968 15896 610020
rect 567936 607155 567988 607164
rect 567936 607121 567945 607155
rect 567945 607121 567979 607155
rect 567979 607121 567988 607155
rect 567936 607112 567988 607121
rect 567936 598927 567988 598936
rect 567936 598893 567945 598927
rect 567945 598893 567979 598927
rect 567979 598893 567988 598927
rect 567936 598884 567988 598893
rect 567936 572704 567988 572756
rect 567936 572568 567988 572620
rect 567936 563159 567988 563168
rect 567936 563125 567945 563159
rect 567945 563125 567979 563159
rect 567979 563125 567988 563159
rect 567936 563116 567988 563125
rect 567936 560371 567988 560380
rect 567936 560337 567945 560371
rect 567945 560337 567979 560371
rect 567979 560337 567988 560371
rect 567936 560328 567988 560337
rect 567936 553435 567988 553444
rect 567936 553401 567945 553435
rect 567945 553401 567979 553435
rect 567979 553401 567988 553435
rect 567936 553392 567988 553401
rect 3148 552032 3200 552084
rect 18604 552032 18656 552084
rect 567936 550647 567988 550656
rect 567936 550613 567945 550647
rect 567945 550613 567979 550647
rect 567979 550613 567988 550647
rect 567936 550604 567988 550613
rect 567936 534080 567988 534132
rect 567936 533944 567988 533996
rect 567936 514768 567988 514820
rect 568028 514632 568080 514684
rect 568028 505563 568080 505572
rect 568028 505529 568037 505563
rect 568037 505529 568071 505563
rect 568071 505529 568080 505563
rect 568028 505520 568080 505529
rect 568028 502435 568080 502444
rect 568028 502401 568037 502435
rect 568037 502401 568071 502435
rect 568071 502401 568080 502435
rect 568028 502392 568080 502401
rect 568028 502299 568080 502308
rect 568028 502265 568037 502299
rect 568037 502265 568071 502299
rect 568071 502265 568080 502299
rect 568028 502256 568080 502265
rect 567936 495388 567988 495440
rect 579712 487092 579764 487144
rect 567936 487024 567988 487076
rect 3516 437452 3568 437504
rect 7564 437452 7616 437504
rect 573364 391960 573416 392012
rect 579620 391960 579672 392012
rect 13636 351908 13688 351960
rect 17040 351908 17092 351960
rect 577504 345516 577556 345568
rect 579620 345516 579672 345568
rect 8208 324300 8260 324352
rect 17040 324300 17092 324352
rect 3332 322940 3384 322992
rect 10324 322940 10376 322992
rect 14464 298120 14516 298172
rect 17040 298120 17092 298172
rect 574744 298120 574796 298172
rect 579620 298120 579672 298172
rect 11704 271872 11756 271924
rect 17040 271872 17092 271924
rect 576124 251200 576176 251252
rect 579620 251200 579672 251252
rect 14556 245624 14608 245676
rect 17040 245624 17092 245676
rect 571248 244332 571300 244384
rect 578884 244332 578936 244384
rect 571248 221484 571300 221536
rect 573364 221484 573416 221536
rect 11796 218016 11848 218068
rect 17040 218016 17092 218068
rect 573364 204280 573416 204332
rect 579620 204280 579672 204332
rect 571248 197412 571300 197464
rect 577504 197412 577556 197464
rect 3792 191836 3844 191888
rect 17040 191836 17092 191888
rect 571248 174156 571300 174208
rect 574744 174156 574796 174208
rect 3884 166948 3936 167000
rect 17040 166948 17092 167000
rect 574744 157360 574796 157412
rect 579620 157360 579672 157412
rect 571248 150356 571300 150408
rect 576124 150356 576176 150408
rect 3700 140700 3752 140752
rect 16764 140700 16816 140752
rect 571248 126692 571300 126744
rect 573364 126692 573416 126744
rect 3608 113092 3660 113144
rect 17040 113092 17092 113144
rect 573364 110440 573416 110492
rect 579620 110440 579672 110492
rect 3332 108944 3384 108996
rect 11796 108944 11848 108996
rect 571248 103028 571300 103080
rect 574744 103028 574796 103080
rect 10324 86572 10376 86624
rect 17040 86572 17092 86624
rect 571248 79228 571300 79280
rect 573364 79228 573416 79280
rect 3332 64812 3384 64864
rect 14556 64812 14608 64864
rect 577412 63520 577464 63572
rect 580172 63520 580224 63572
rect 3516 60664 3568 60716
rect 16948 60664 17000 60716
rect 571248 55292 571300 55344
rect 577412 55292 577464 55344
rect 7564 34416 7616 34468
rect 17040 34416 17092 34468
rect 3148 22040 3200 22092
rect 11704 22040 11756 22092
rect 19984 20612 20036 20664
rect 24216 20612 24268 20664
rect 21364 20544 21416 20596
rect 27620 20544 27672 20596
rect 22284 19320 22336 19372
rect 22376 19252 22428 19304
rect 24124 19252 24176 19304
rect 24860 19252 24912 19304
rect 61384 19252 61436 19304
rect 580540 19252 580592 19304
rect 70216 19184 70268 19236
rect 580448 19184 580500 19236
rect 79692 19116 79744 19168
rect 580356 19116 580408 19168
rect 88892 19048 88944 19100
rect 580264 19048 580316 19100
rect 22468 17960 22520 18012
rect 26148 17892 26200 17944
rect 86868 17892 86920 17944
rect 280344 17892 280396 17944
rect 573364 17892 573416 17944
rect 579804 17892 579856 17944
rect 18604 17824 18656 17876
rect 42432 17824 42484 17876
rect 93768 17824 93820 17876
rect 298652 17824 298704 17876
rect 15844 17756 15896 17808
rect 33324 17756 33376 17808
rect 100668 17756 100720 17808
rect 316960 17756 317012 17808
rect 3424 17688 3476 17740
rect 51632 17688 51684 17740
rect 107568 17688 107620 17740
rect 335452 17688 335504 17740
rect 115848 17620 115900 17672
rect 353576 17620 353628 17672
rect 122748 17552 122800 17604
rect 371884 17552 371936 17604
rect 10968 17484 11020 17536
rect 97356 17484 97408 17536
rect 125508 17484 125560 17536
rect 380992 17484 381044 17536
rect 34428 17416 34480 17468
rect 408500 17416 408552 17468
rect 41328 17348 41380 17400
rect 417608 17348 417660 17400
rect 15108 17280 15160 17332
rect 106556 17280 106608 17332
rect 117136 17280 117188 17332
rect 536840 17280 536892 17332
rect 24768 17212 24820 17264
rect 124772 17212 124824 17264
rect 125416 17212 125468 17264
rect 545672 17212 545724 17264
rect 79968 17144 80020 17196
rect 262220 17144 262272 17196
rect 73068 17076 73120 17128
rect 243728 17076 243780 17128
rect 64696 17008 64748 17060
rect 225420 17008 225472 17060
rect 57888 16940 57940 16992
rect 207204 16940 207256 16992
rect 50988 16872 51040 16924
rect 189080 16872 189132 16924
rect 48136 16804 48188 16856
rect 179696 16804 179748 16856
rect 44088 16736 44140 16788
rect 170588 16736 170640 16788
rect 39948 16668 40000 16720
rect 161572 16668 161624 16720
rect 33048 16600 33100 16652
rect 143080 16600 143132 16652
rect 24860 10956 24912 11008
rect 28816 10956 28868 11008
rect 26240 10888 26292 10940
rect 27712 10888 27764 10940
rect 22560 9596 22612 9648
rect 24860 9596 24912 9648
rect 28816 8304 28868 8356
rect 33140 8236 33192 8288
rect 27712 8168 27764 8220
rect 29092 8168 29144 8220
rect 123024 6332 123076 6384
rect 571708 6332 571760 6384
rect 77852 6264 77904 6316
rect 571340 6264 571392 6316
rect 67180 6196 67232 6248
rect 571432 6196 571484 6248
rect 4068 6128 4120 6180
rect 571616 6128 571668 6180
rect 1676 5448 1728 5500
rect 398840 5448 398892 5500
rect 116032 5380 116084 5432
rect 571800 5380 571852 5432
rect 108764 5312 108816 5364
rect 571892 5312 571944 5364
rect 17224 5244 17276 5296
rect 90916 5244 90968 5296
rect 101588 5244 101640 5296
rect 571984 5244 572036 5296
rect 87328 5176 87380 5228
rect 572076 5176 572128 5228
rect 80244 5108 80296 5160
rect 572168 5108 572220 5160
rect 24860 5040 24912 5092
rect 49608 5040 49660 5092
rect 69480 5040 69532 5092
rect 572260 5040 572312 5092
rect 48228 4972 48280 5024
rect 572352 4972 572404 5024
rect 24124 4904 24176 4956
rect 24860 4904 24912 4956
rect 26700 4904 26752 4956
rect 572444 4904 572496 4956
rect 21916 4836 21968 4888
rect 572536 4836 572588 4888
rect 17224 4768 17276 4820
rect 572628 4768 572680 4820
rect 572 4700 624 4752
rect 389180 4700 389232 4752
rect 65984 4632 66036 4684
rect 454040 4632 454092 4684
rect 62396 4564 62448 4616
rect 444380 4564 444432 4616
rect 83832 4496 83884 4548
rect 462320 4496 462372 4548
rect 58808 4428 58860 4480
rect 436100 4428 436152 4480
rect 51632 4360 51684 4412
rect 426440 4360 426492 4412
rect 112352 4292 112404 4344
rect 471980 4292 472032 4344
rect 29092 4224 29144 4276
rect 119436 4224 119488 4276
rect 17132 4088 17184 4140
rect 55220 4088 55272 4140
rect 63592 4088 63644 4140
rect 64788 4088 64840 4140
rect 68284 4088 68336 4140
rect 75460 4088 75512 4140
rect 252560 4088 252612 4140
rect 21732 4020 21784 4072
rect 76656 4020 76708 4072
rect 17408 3952 17460 4004
rect 84936 4020 84988 4072
rect 92112 4020 92164 4072
rect 270500 4020 270552 4072
rect 79048 3952 79100 4004
rect 79968 3952 80020 4004
rect 82636 3952 82688 4004
rect 17500 3884 17552 3936
rect 88524 3884 88576 3936
rect 89720 3884 89772 3936
rect 289820 3952 289872 4004
rect 97908 3884 97960 3936
rect 307760 3884 307812 3936
rect 17592 3816 17644 3868
rect 86132 3816 86184 3868
rect 86868 3816 86920 3868
rect 93308 3816 93360 3868
rect 93768 3816 93820 3868
rect 103980 3816 104032 3868
rect 325700 3816 325752 3868
rect 17684 3748 17736 3800
rect 102784 3748 102836 3800
rect 343640 3748 343692 3800
rect 19524 3680 19576 3732
rect 113548 3680 113600 3732
rect 114468 3680 114520 3732
rect 114744 3680 114796 3732
rect 115848 3680 115900 3732
rect 121828 3680 121880 3732
rect 122748 3680 122800 3732
rect 124220 3680 124272 3732
rect 125416 3680 125468 3732
rect 362960 3680 363012 3732
rect 21548 3612 21600 3664
rect 12440 3544 12492 3596
rect 13636 3544 13688 3596
rect 18328 3544 18380 3596
rect 19156 3544 19208 3596
rect 20720 3544 20772 3596
rect 21824 3544 21876 3596
rect 24308 3544 24360 3596
rect 24768 3544 24820 3596
rect 34980 3612 35032 3664
rect 499580 3612 499632 3664
rect 30288 3544 30340 3596
rect 33876 3544 33928 3596
rect 34428 3544 34480 3596
rect 42156 3544 42208 3596
rect 42708 3544 42760 3596
rect 43352 3544 43404 3596
rect 44088 3544 44140 3596
rect 46940 3544 46992 3596
rect 48136 3544 48188 3596
rect 50528 3544 50580 3596
rect 50988 3544 51040 3596
rect 517520 3544 517572 3596
rect 7656 3476 7708 3528
rect 8208 3476 8260 3528
rect 8852 3476 8904 3528
rect 9588 3476 9640 3528
rect 10048 3476 10100 3528
rect 10968 3476 11020 3528
rect 11244 3476 11296 3528
rect 554780 3476 554832 3528
rect 2872 3408 2924 3460
rect 14464 3408 14516 3460
rect 16028 3408 16080 3460
rect 563060 3408 563112 3460
rect 21272 3340 21324 3392
rect 60004 3340 60056 3392
rect 71872 3340 71924 3392
rect 73068 3340 73120 3392
rect 234620 3340 234672 3392
rect 17868 3272 17920 3324
rect 25504 3272 25556 3324
rect 56416 3272 56468 3324
rect 61200 3272 61252 3324
rect 215300 3272 215352 3324
rect 22008 3204 22060 3256
rect 52828 3204 52880 3256
rect 54024 3204 54076 3256
rect 197360 3204 197412 3256
rect 19248 3136 19300 3188
rect 36176 3136 36228 3188
rect 151820 3136 151872 3188
rect 29092 3068 29144 3120
rect 133880 3068 133932 3120
rect 17776 3000 17828 3052
rect 120632 3000 120684 3052
rect 17316 2932 17368 2984
rect 23112 2932 23164 2984
rect 24860 2932 24912 2984
rect 94504 2932 94556 2984
rect 96896 2932 96948 2984
rect 97908 2932 97960 2984
rect 111156 2932 111208 2984
rect 118240 2932 118292 2984
rect 33140 2864 33192 2916
rect 98092 2864 98144 2916
rect 115940 2864 115992 2916
rect 21456 2796 21508 2848
rect 49332 2796 49384 2848
rect 45744 2728 45796 2780
rect 49608 2728 49660 2780
rect 105176 2796 105228 2848
rect 5264 552 5316 604
rect 5448 552 5500 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 40512 700466 40540 703520
rect 105464 700670 105492 703520
rect 170324 700738 170352 703520
rect 135168 700732 135220 700738
rect 135168 700674 135220 700680
rect 170312 700732 170364 700738
rect 170312 700674 170364 700680
rect 105452 700664 105504 700670
rect 105452 700606 105504 700612
rect 106188 700664 106240 700670
rect 106188 700606 106240 700612
rect 118608 700664 118660 700670
rect 118608 700606 118660 700612
rect 100668 700596 100720 700602
rect 100668 700538 100720 700544
rect 82728 700528 82780 700534
rect 82728 700470 82780 700476
rect 40500 700460 40552 700466
rect 40500 700402 40552 700408
rect 41328 700460 41380 700466
rect 41328 700402 41380 700408
rect 64788 700460 64840 700466
rect 64788 700402 64840 700408
rect 28908 700324 28960 700330
rect 28908 700266 28960 700272
rect 21824 686792 21876 686798
rect 21824 686734 21876 686740
rect 21548 686588 21600 686594
rect 21548 686530 21600 686536
rect 9588 686452 9640 686458
rect 9588 686394 9640 686400
rect 6828 669384 6880 669390
rect 6828 669326 6880 669332
rect 3422 667992 3478 668001
rect 3422 667927 3424 667936
rect 3476 667927 3478 667936
rect 3424 667898 3476 667904
rect 5448 643136 5500 643142
rect 5448 643078 5500 643084
rect 3422 610464 3478 610473
rect 3422 610399 3478 610408
rect 3436 610026 3464 610399
rect 3424 610020 3476 610026
rect 3424 609962 3476 609968
rect 3146 553072 3202 553081
rect 3146 553007 3202 553016
rect 3160 552090 3188 553007
rect 3148 552084 3200 552090
rect 3148 552026 3200 552032
rect 3422 495544 3478 495553
rect 3422 495479 3478 495488
rect 3330 323096 3386 323105
rect 3330 323031 3386 323040
rect 3344 322998 3372 323031
rect 3332 322992 3384 322998
rect 3332 322934 3384 322940
rect 3332 108996 3384 109002
rect 3332 108938 3384 108944
rect 3344 107681 3372 108938
rect 3330 107672 3386 107681
rect 3330 107607 3386 107616
rect 3332 64864 3384 64870
rect 3332 64806 3384 64812
rect 3344 64569 3372 64806
rect 3330 64560 3386 64569
rect 3330 64495 3386 64504
rect 3148 22092 3200 22098
rect 3148 22034 3200 22040
rect 3160 21457 3188 22034
rect 3146 21448 3202 21457
rect 3146 21383 3202 21392
rect 3436 17746 3464 495479
rect 3514 438016 3570 438025
rect 3514 437951 3570 437960
rect 3528 437510 3556 437951
rect 3516 437504 3568 437510
rect 3516 437446 3568 437452
rect 3514 380624 3570 380633
rect 3514 380559 3570 380568
rect 3528 60722 3556 380559
rect 3606 280120 3662 280129
rect 3606 280055 3662 280064
rect 3620 113150 3648 280055
rect 3698 237008 3754 237017
rect 3698 236943 3754 236952
rect 3712 140758 3740 236943
rect 3882 193896 3938 193905
rect 3882 193831 3938 193840
rect 3792 191888 3844 191894
rect 3792 191830 3844 191836
rect 3804 150793 3832 191830
rect 3896 167006 3924 193831
rect 3884 167000 3936 167006
rect 3884 166942 3936 166948
rect 3790 150784 3846 150793
rect 3790 150719 3846 150728
rect 3700 140752 3752 140758
rect 3700 140694 3752 140700
rect 3608 113144 3660 113150
rect 3608 113086 3660 113092
rect 3516 60716 3568 60722
rect 3516 60658 3568 60664
rect 3424 17740 3476 17746
rect 3424 17682 3476 17688
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 1676 5500 1728 5506
rect 1676 5442 1728 5448
rect 572 4752 624 4758
rect 572 4694 624 4700
rect 584 480 612 4694
rect 1688 480 1716 5442
rect 2872 3460 2924 3466
rect 2872 3402 2924 3408
rect 2884 480 2912 3402
rect 4080 480 4108 6122
rect 5460 610 5488 643078
rect 6840 626 6868 669326
rect 7564 437504 7616 437510
rect 7564 437446 7616 437452
rect 7576 34474 7604 437446
rect 8208 324352 8260 324358
rect 8208 324294 8260 324300
rect 7564 34468 7616 34474
rect 7564 34410 7616 34416
rect 8220 3534 8248 324294
rect 9600 3534 9628 686394
rect 13728 686384 13780 686390
rect 13728 686326 13780 686332
rect 13636 351960 13688 351966
rect 13636 351902 13688 351908
rect 10324 322992 10376 322998
rect 10324 322934 10376 322940
rect 10336 86630 10364 322934
rect 11704 271924 11756 271930
rect 11704 271866 11756 271872
rect 10324 86624 10376 86630
rect 10324 86566 10376 86572
rect 11716 22098 11744 271866
rect 11796 218068 11848 218074
rect 11796 218010 11848 218016
rect 11808 109002 11836 218010
rect 11796 108996 11848 109002
rect 11796 108938 11848 108944
rect 11704 22092 11756 22098
rect 11704 22034 11756 22040
rect 10968 17536 11020 17542
rect 10968 17478 11020 17484
rect 10980 3534 11008 17478
rect 13648 3602 13676 351902
rect 12440 3596 12492 3602
rect 12440 3538 12492 3544
rect 13636 3596 13688 3602
rect 13636 3538 13688 3544
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8852 3528 8904 3534
rect 8852 3470 8904 3476
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 5264 604 5316 610
rect 5264 546 5316 552
rect 5448 604 5500 610
rect 5448 546 5500 552
rect 6472 598 6868 626
rect 5276 480 5304 546
rect 6472 480 6500 598
rect 7668 480 7696 3470
rect 8864 480 8892 3470
rect 10060 480 10088 3470
rect 11256 480 11284 3470
rect 12452 480 12480 3538
rect 13740 3482 13768 686326
rect 21364 686316 21416 686322
rect 21364 686258 21416 686264
rect 21272 686044 21324 686050
rect 21272 685986 21324 685992
rect 17866 670576 17922 670585
rect 17866 670511 17922 670520
rect 17880 669390 17908 670511
rect 17868 669384 17920 669390
rect 17868 669326 17920 669332
rect 19984 667956 20036 667962
rect 19984 667898 20036 667904
rect 17866 644056 17922 644065
rect 17866 643991 17922 644000
rect 17880 643142 17908 643991
rect 17868 643136 17920 643142
rect 17868 643078 17920 643084
rect 17866 617536 17922 617545
rect 17866 617471 17922 617480
rect 15844 610020 15896 610026
rect 15844 609962 15896 609968
rect 14464 298172 14516 298178
rect 14464 298114 14516 298120
rect 13648 3454 13768 3482
rect 14476 3466 14504 298114
rect 14556 245676 14608 245682
rect 14556 245618 14608 245624
rect 14568 64870 14596 245618
rect 14556 64864 14608 64870
rect 14556 64806 14608 64812
rect 15856 17814 15884 609962
rect 17774 590880 17830 590889
rect 17774 590815 17830 590824
rect 17682 564360 17738 564369
rect 17682 564295 17738 564304
rect 17590 537840 17646 537849
rect 17590 537775 17646 537784
rect 17498 511320 17554 511329
rect 17498 511255 17554 511264
rect 17406 484664 17462 484673
rect 17406 484599 17462 484608
rect 17314 431624 17370 431633
rect 17314 431559 17370 431568
rect 17222 404968 17278 404977
rect 17222 404903 17278 404912
rect 17130 378448 17186 378457
rect 17130 378383 17186 378392
rect 17040 351960 17092 351966
rect 17038 351928 17040 351937
rect 17092 351928 17094 351937
rect 17038 351863 17094 351872
rect 17038 325408 17094 325417
rect 17038 325343 17094 325352
rect 17052 324358 17080 325343
rect 17040 324352 17092 324358
rect 17040 324294 17092 324300
rect 17038 298752 17094 298761
rect 17038 298687 17094 298696
rect 17052 298178 17080 298687
rect 17040 298172 17092 298178
rect 17040 298114 17092 298120
rect 17038 272232 17094 272241
rect 17038 272167 17094 272176
rect 17052 271930 17080 272167
rect 17040 271924 17092 271930
rect 17040 271866 17092 271872
rect 17038 245712 17094 245721
rect 17038 245647 17040 245656
rect 17092 245647 17094 245656
rect 17040 245618 17092 245624
rect 17038 219056 17094 219065
rect 17038 218991 17094 219000
rect 17052 218074 17080 218991
rect 17040 218068 17092 218074
rect 17040 218010 17092 218016
rect 17038 192536 17094 192545
rect 17038 192471 17094 192480
rect 17052 191894 17080 192471
rect 17040 191888 17092 191894
rect 17040 191830 17092 191836
rect 17040 167000 17092 167006
rect 17040 166942 17092 166948
rect 17052 166025 17080 166942
rect 17038 166016 17094 166025
rect 17038 165951 17094 165960
rect 16764 140752 16816 140758
rect 16764 140694 16816 140700
rect 16776 139505 16804 140694
rect 16762 139496 16818 139505
rect 16762 139431 16818 139440
rect 17040 113144 17092 113150
rect 17040 113086 17092 113092
rect 17052 112849 17080 113086
rect 17038 112840 17094 112849
rect 17038 112775 17094 112784
rect 17040 86624 17092 86630
rect 17040 86566 17092 86572
rect 17052 86329 17080 86566
rect 17038 86320 17094 86329
rect 17038 86255 17094 86264
rect 16948 60716 17000 60722
rect 16948 60658 17000 60664
rect 16960 59809 16988 60658
rect 16946 59800 17002 59809
rect 16946 59735 17002 59744
rect 17040 34468 17092 34474
rect 17040 34410 17092 34416
rect 17052 33289 17080 34410
rect 17038 33280 17094 33289
rect 17038 33215 17094 33224
rect 15844 17808 15896 17814
rect 15844 17750 15896 17756
rect 15108 17332 15160 17338
rect 15108 17274 15160 17280
rect 15120 3482 15148 17274
rect 17144 4146 17172 378383
rect 17236 5302 17264 404903
rect 17224 5296 17276 5302
rect 17224 5238 17276 5244
rect 17224 4820 17276 4826
rect 17224 4762 17276 4768
rect 17132 4140 17184 4146
rect 17132 4082 17184 4088
rect 14464 3460 14516 3466
rect 13648 480 13676 3454
rect 14464 3402 14516 3408
rect 14844 3454 15148 3482
rect 16028 3460 16080 3466
rect 14844 480 14872 3454
rect 16028 3402 16080 3408
rect 16040 480 16068 3402
rect 17236 480 17264 4762
rect 17328 2990 17356 431559
rect 17420 4010 17448 484599
rect 17408 4004 17460 4010
rect 17408 3946 17460 3952
rect 17512 3942 17540 511255
rect 17500 3936 17552 3942
rect 17500 3878 17552 3884
rect 17604 3874 17632 537775
rect 17592 3868 17644 3874
rect 17592 3810 17644 3816
rect 17696 3806 17724 564295
rect 17684 3800 17736 3806
rect 17684 3742 17736 3748
rect 17788 3058 17816 590815
rect 17880 3330 17908 617471
rect 18604 552084 18656 552090
rect 18604 552026 18656 552032
rect 18616 17882 18644 552026
rect 19246 458144 19302 458153
rect 19246 458079 19302 458088
rect 18604 17876 18656 17882
rect 18604 17818 18656 17824
rect 19154 17368 19210 17377
rect 19154 17303 19210 17312
rect 19168 3602 19196 17303
rect 18328 3596 18380 3602
rect 18328 3538 18380 3544
rect 19156 3596 19208 3602
rect 19156 3538 19208 3544
rect 17868 3324 17920 3330
rect 17868 3266 17920 3272
rect 17776 3052 17828 3058
rect 17776 2994 17828 3000
rect 17316 2984 17368 2990
rect 17316 2926 17368 2932
rect 18340 480 18368 3538
rect 19260 3194 19288 458079
rect 19996 20670 20024 667898
rect 19984 20664 20036 20670
rect 19984 20606 20036 20612
rect 19524 3732 19576 3738
rect 19524 3674 19576 3680
rect 19248 3188 19300 3194
rect 19248 3130 19300 3136
rect 19536 480 19564 3674
rect 20720 3596 20772 3602
rect 20720 3538 20772 3544
rect 20732 480 20760 3538
rect 21284 3398 21312 685986
rect 21376 20602 21404 686258
rect 21456 686180 21508 686186
rect 21456 686122 21508 686128
rect 21364 20596 21416 20602
rect 21364 20538 21416 20544
rect 21272 3392 21324 3398
rect 21272 3334 21324 3340
rect 21468 2854 21496 686122
rect 21560 3670 21588 686530
rect 21732 686520 21784 686526
rect 21732 686462 21784 686468
rect 21640 685976 21692 685982
rect 21640 685918 21692 685924
rect 21548 3664 21600 3670
rect 21548 3606 21600 3612
rect 21652 3505 21680 685918
rect 21744 4078 21772 686462
rect 21732 4072 21784 4078
rect 21732 4014 21784 4020
rect 21836 3602 21864 686734
rect 21916 686112 21968 686118
rect 21916 686054 21968 686060
rect 21928 5114 21956 686054
rect 28920 684162 28948 700266
rect 41340 686662 41368 700402
rect 46848 700392 46900 700398
rect 46848 700334 46900 700340
rect 41328 686656 41380 686662
rect 41328 686598 41380 686604
rect 28874 684134 28948 684162
rect 28874 683876 28902 684134
rect 46860 683890 46888 700334
rect 46552 683862 46888 683890
rect 64800 683754 64828 700402
rect 82740 687206 82768 700470
rect 82268 687200 82320 687206
rect 82268 687142 82320 687148
rect 82728 687200 82780 687206
rect 82728 687142 82780 687148
rect 82280 683890 82308 687142
rect 100680 686866 100708 700538
rect 99932 686860 99984 686866
rect 99932 686802 99984 686808
rect 100668 686860 100720 686866
rect 100668 686802 100720 686808
rect 99944 683890 99972 686802
rect 106200 686730 106228 700606
rect 118620 687138 118648 700606
rect 117688 687132 117740 687138
rect 117688 687074 117740 687080
rect 118608 687132 118660 687138
rect 118608 687074 118660 687080
rect 106188 686724 106240 686730
rect 106188 686666 106240 686672
rect 117700 683890 117728 687074
rect 135180 683890 135208 700674
rect 235184 700670 235212 703520
rect 235172 700664 235224 700670
rect 235172 700606 235224 700612
rect 300136 700602 300164 703520
rect 300124 700596 300176 700602
rect 300124 700538 300176 700544
rect 364996 700534 365024 703520
rect 364984 700528 365036 700534
rect 364984 700470 365036 700476
rect 429856 700466 429884 703520
rect 429844 700460 429896 700466
rect 429844 700402 429896 700408
rect 494808 700398 494836 703520
rect 494796 700392 494848 700398
rect 494796 700334 494848 700340
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 559748 686792 559800 686798
rect 559748 686734 559800 686740
rect 152464 686724 152516 686730
rect 152464 686666 152516 686672
rect 81972 683862 82308 683890
rect 99636 683862 99972 683890
rect 117392 683862 117728 683890
rect 135056 683862 135208 683890
rect 152476 683890 152504 686666
rect 170128 686656 170180 686662
rect 170128 686598 170180 686604
rect 170140 683890 170168 686598
rect 205640 686588 205692 686594
rect 205640 686530 205692 686536
rect 188528 686248 188580 686254
rect 188528 686190 188580 686196
rect 188540 683890 188568 686190
rect 152476 683862 152812 683890
rect 170140 683862 170476 683890
rect 188232 683862 188568 683890
rect 205652 683890 205680 686530
rect 276388 686520 276440 686526
rect 276388 686462 276440 686468
rect 223578 686352 223634 686361
rect 223578 686287 223634 686296
rect 223592 683890 223620 686287
rect 240966 686216 241022 686225
rect 240966 686151 241022 686160
rect 240980 683890 241008 686151
rect 258722 686080 258778 686089
rect 258722 686015 258778 686024
rect 258736 683890 258764 686015
rect 276400 683890 276428 686462
rect 364984 686452 365036 686458
rect 364984 686394 365036 686400
rect 347226 686080 347282 686089
rect 347226 686015 347282 686024
rect 347240 683890 347268 686015
rect 364996 683890 365024 686394
rect 382648 686384 382700 686390
rect 382648 686326 382700 686332
rect 382660 683890 382688 686326
rect 400404 686316 400456 686322
rect 400404 686258 400456 686264
rect 400416 683890 400444 686258
rect 542726 686216 542782 686225
rect 418160 686180 418212 686186
rect 542726 686151 542782 686160
rect 418160 686122 418212 686128
rect 418172 683890 418200 686122
rect 436100 686112 436152 686118
rect 436100 686054 436152 686060
rect 524970 686080 525026 686089
rect 436112 683890 436140 686054
rect 453488 686044 453540 686050
rect 524970 686015 525026 686024
rect 453488 685986 453540 685992
rect 453500 683890 453528 685986
rect 488908 685976 488960 685982
rect 471242 685944 471298 685953
rect 488908 685918 488960 685924
rect 507306 685944 507362 685953
rect 471242 685879 471298 685888
rect 471256 683890 471284 685879
rect 488920 683890 488948 685918
rect 507306 685879 507362 685888
rect 507320 683890 507348 685879
rect 524984 683890 525012 686015
rect 542740 683890 542768 686151
rect 205652 683862 205896 683890
rect 223592 683862 223652 683890
rect 240980 683862 241316 683890
rect 258736 683862 259072 683890
rect 276400 683862 276736 683890
rect 347240 683862 347576 683890
rect 364996 683862 365332 683890
rect 382660 683862 382996 683890
rect 400416 683862 400752 683890
rect 418172 683862 418416 683890
rect 436112 683862 436172 683890
rect 453500 683862 453836 683890
rect 471256 683862 471592 683890
rect 488920 683862 489256 683890
rect 507012 683862 507348 683890
rect 524676 683862 525012 683890
rect 542432 683862 542768 683890
rect 559760 683890 559788 686734
rect 580262 686352 580318 686361
rect 580262 686287 580318 686296
rect 567844 686248 567896 686254
rect 567844 686190 567896 686196
rect 559760 683862 560096 683890
rect 64216 683726 64828 683754
rect 293866 683768 293922 683777
rect 293922 683726 294492 683754
rect 293866 683703 293922 683712
rect 329746 683496 329802 683505
rect 329802 683454 329912 683482
rect 329746 683431 329802 683440
rect 311806 683360 311862 683369
rect 311862 683318 312156 683346
rect 311806 683295 311862 683304
rect 22374 682816 22430 682825
rect 22374 682751 22430 682760
rect 22282 682680 22338 682689
rect 22282 682615 22338 682624
rect 22296 19378 22324 682615
rect 22284 19372 22336 19378
rect 22284 19314 22336 19320
rect 22388 19310 22416 682751
rect 22558 682544 22614 682553
rect 22558 682479 22614 682488
rect 22466 682408 22522 682417
rect 22466 682343 22522 682352
rect 22376 19304 22428 19310
rect 22376 19246 22428 19252
rect 22480 18018 22508 682343
rect 22468 18012 22520 18018
rect 22468 17954 22520 17960
rect 22572 9654 22600 682479
rect 567856 669474 567884 686190
rect 567764 669446 567884 669474
rect 567764 661994 567792 669446
rect 567764 661978 567976 661994
rect 567764 661972 567988 661978
rect 567764 661966 567936 661972
rect 567936 661914 567988 661920
rect 567936 657008 567988 657014
rect 567856 656968 567936 656996
rect 567856 650162 567884 656968
rect 567936 656950 567988 656956
rect 567764 650134 567884 650162
rect 567764 642410 567792 650134
rect 567764 642394 567976 642410
rect 567764 642388 567988 642394
rect 567764 642382 567936 642388
rect 567936 642330 567988 642336
rect 567936 637696 567988 637702
rect 567856 637644 567936 637650
rect 567856 637638 567988 637644
rect 567856 637622 567976 637638
rect 567856 630578 567884 637622
rect 567764 630550 567884 630578
rect 567764 623098 567792 630550
rect 567764 623082 567976 623098
rect 567764 623076 567988 623082
rect 567764 623070 567936 623076
rect 567936 623018 567988 623024
rect 567936 618384 567988 618390
rect 567856 618332 567936 618338
rect 567856 618326 567988 618332
rect 567856 618310 567976 618326
rect 567856 613442 567884 618310
rect 567764 613414 567884 613442
rect 567764 607186 567792 613414
rect 567764 607170 567976 607186
rect 567764 607164 567988 607170
rect 567764 607158 567936 607164
rect 567936 607106 567988 607112
rect 571338 600944 571394 600953
rect 571338 600879 571394 600888
rect 567936 598936 567988 598942
rect 567856 598896 567936 598924
rect 567856 574682 567884 598896
rect 567936 598878 567988 598884
rect 567856 574654 567976 574682
rect 567948 572762 567976 574654
rect 567936 572756 567988 572762
rect 567936 572698 567988 572704
rect 567936 572620 567988 572626
rect 567936 572562 567988 572568
rect 567948 569922 567976 572562
rect 567856 569894 567976 569922
rect 567856 563258 567884 569894
rect 567856 563230 567976 563258
rect 567948 563174 567976 563230
rect 567936 563168 567988 563174
rect 567936 563110 567988 563116
rect 567936 560380 567988 560386
rect 567936 560322 567988 560328
rect 567948 553450 567976 560322
rect 567936 553444 567988 553450
rect 567936 553386 567988 553392
rect 567948 550662 567976 550693
rect 567936 550656 567988 550662
rect 567856 550604 567936 550610
rect 567856 550598 567988 550604
rect 567856 550582 567976 550598
rect 567856 536194 567884 550582
rect 567856 536166 567976 536194
rect 567948 534138 567976 536166
rect 567936 534132 567988 534138
rect 567936 534074 567988 534080
rect 567936 533996 567988 534002
rect 567936 533938 567988 533944
rect 567948 531298 567976 533938
rect 567856 531270 567976 531298
rect 567856 514842 567884 531270
rect 567856 514826 567976 514842
rect 567856 514820 567988 514826
rect 567856 514814 567936 514820
rect 567936 514762 567988 514768
rect 568028 514684 568080 514690
rect 568028 514626 568080 514632
rect 568040 505578 568068 514626
rect 568028 505572 568080 505578
rect 568028 505514 568080 505520
rect 568028 502444 568080 502450
rect 568028 502386 568080 502392
rect 568040 502314 568068 502386
rect 568028 502308 568080 502314
rect 568028 502250 568080 502256
rect 567936 495440 567988 495446
rect 567936 495382 567988 495388
rect 567948 492674 567976 495382
rect 567856 492646 567976 492674
rect 567856 487098 567884 492646
rect 567856 487082 567976 487098
rect 567856 487076 567988 487082
rect 567856 487070 567936 487076
rect 567936 487018 567988 487024
rect 571246 244760 571302 244769
rect 571246 244695 571302 244704
rect 571260 244390 571288 244695
rect 571248 244384 571300 244390
rect 571248 244326 571300 244332
rect 571248 221536 571300 221542
rect 571246 221504 571248 221513
rect 571300 221504 571302 221513
rect 571246 221439 571302 221448
rect 571246 197568 571302 197577
rect 571246 197503 571302 197512
rect 571260 197470 571288 197503
rect 571248 197464 571300 197470
rect 571248 197406 571300 197412
rect 571248 174208 571300 174214
rect 571246 174176 571248 174185
rect 571300 174176 571302 174185
rect 571246 174111 571302 174120
rect 571248 150408 571300 150414
rect 571246 150376 571248 150385
rect 571300 150376 571302 150385
rect 571246 150311 571302 150320
rect 571248 126744 571300 126750
rect 571246 126712 571248 126721
rect 571300 126712 571302 126721
rect 571246 126647 571302 126656
rect 571248 103080 571300 103086
rect 571246 103048 571248 103057
rect 571300 103048 571302 103057
rect 571246 102983 571302 102992
rect 571248 79280 571300 79286
rect 571246 79248 571248 79257
rect 571300 79248 571302 79257
rect 571246 79183 571302 79192
rect 571248 55344 571300 55350
rect 571246 55312 571248 55321
rect 571300 55312 571302 55321
rect 571246 55247 571302 55256
rect 24216 20664 24268 20670
rect 24268 20612 24564 20618
rect 24216 20606 24564 20612
rect 24228 20590 24564 20606
rect 27620 20596 27672 20602
rect 27620 20538 27672 20544
rect 24124 19304 24176 19310
rect 24124 19246 24176 19252
rect 24860 19304 24912 19310
rect 24860 19246 24912 19252
rect 22560 9648 22612 9654
rect 22560 9590 22612 9596
rect 21928 5086 22048 5114
rect 21916 4888 21968 4894
rect 21916 4830 21968 4836
rect 21824 3596 21876 3602
rect 21824 3538 21876 3544
rect 21638 3496 21694 3505
rect 21638 3431 21694 3440
rect 21456 2848 21508 2854
rect 21456 2790 21508 2796
rect 21928 480 21956 4830
rect 22020 3262 22048 5086
rect 24136 4962 24164 19246
rect 24768 17264 24820 17270
rect 24768 17206 24820 17212
rect 24124 4956 24176 4962
rect 24124 4898 24176 4904
rect 24780 3602 24808 17206
rect 24872 11014 24900 19246
rect 26148 17944 26200 17950
rect 26148 17886 26200 17892
rect 26160 15178 26188 17886
rect 26160 15150 26280 15178
rect 24860 11008 24912 11014
rect 24860 10950 24912 10956
rect 26252 10946 26280 15150
rect 26240 10940 26292 10946
rect 26240 10882 26292 10888
rect 24860 9648 24912 9654
rect 24860 9590 24912 9596
rect 24872 5098 24900 9590
rect 24860 5092 24912 5098
rect 24860 5034 24912 5040
rect 24860 4956 24912 4962
rect 24860 4898 24912 4904
rect 26700 4956 26752 4962
rect 26700 4898 26752 4904
rect 24308 3596 24360 3602
rect 24308 3538 24360 3544
rect 24768 3596 24820 3602
rect 24768 3538 24820 3544
rect 22008 3256 22060 3262
rect 22008 3198 22060 3204
rect 23112 2984 23164 2990
rect 23112 2926 23164 2932
rect 23124 480 23152 2926
rect 24320 480 24348 3538
rect 24872 2990 24900 4898
rect 25504 3324 25556 3330
rect 25504 3266 25556 3272
rect 24860 2984 24912 2990
rect 24860 2926 24912 2932
rect 25516 480 25544 3266
rect 26712 480 26740 4898
rect 27632 3346 27660 20538
rect 33336 20046 33672 20074
rect 42444 20046 42780 20074
rect 51644 20046 51980 20074
rect 61088 20046 61424 20074
rect 33336 17814 33364 20046
rect 42444 17882 42472 20046
rect 42432 17876 42484 17882
rect 42432 17818 42484 17824
rect 33324 17808 33376 17814
rect 33324 17750 33376 17756
rect 51644 17746 51672 20046
rect 61396 19310 61424 20046
rect 70228 20046 70288 20074
rect 79396 20046 79732 20074
rect 88596 20046 88932 20074
rect 61384 19304 61436 19310
rect 61384 19246 61436 19252
rect 70228 19242 70256 20046
rect 70216 19236 70268 19242
rect 70216 19178 70268 19184
rect 79704 19174 79732 20046
rect 79692 19168 79744 19174
rect 79692 19110 79744 19116
rect 88904 19106 88932 20046
rect 97368 20046 97704 20074
rect 106568 20046 106904 20074
rect 115952 20046 116012 20074
rect 124784 20046 125120 20074
rect 133892 20046 134320 20074
rect 143092 20046 143428 20074
rect 151832 20046 152628 20074
rect 161584 20046 161736 20074
rect 170600 20046 170936 20074
rect 179708 20046 180044 20074
rect 189092 20046 189244 20074
rect 197372 20046 198352 20074
rect 207216 20046 207552 20074
rect 215312 20046 216660 20074
rect 225432 20046 225768 20074
rect 234632 20046 234968 20074
rect 243740 20046 244076 20074
rect 252572 20046 253276 20074
rect 262232 20046 262384 20074
rect 270512 20046 271584 20074
rect 280356 20046 280692 20074
rect 289832 20046 289892 20074
rect 298664 20046 299000 20074
rect 307772 20046 308108 20074
rect 316972 20046 317308 20074
rect 325712 20046 326416 20074
rect 335464 20046 335616 20074
rect 343652 20046 344724 20074
rect 353588 20046 353924 20074
rect 362972 20046 363032 20074
rect 371896 20046 372232 20074
rect 381004 20046 381340 20074
rect 389192 20046 390540 20074
rect 398852 20046 399648 20074
rect 408512 20046 408756 20074
rect 417620 20046 417956 20074
rect 426452 20046 427064 20074
rect 436112 20046 436264 20074
rect 444392 20046 445372 20074
rect 454052 20046 454572 20074
rect 462332 20046 463680 20074
rect 471992 20046 472880 20074
rect 481652 20046 481988 20074
rect 490760 20046 491096 20074
rect 499592 20046 500296 20074
rect 509252 20046 509404 20074
rect 517532 20046 518604 20074
rect 527376 20046 527712 20074
rect 536852 20046 536912 20074
rect 545684 20046 546020 20074
rect 554792 20046 555220 20074
rect 563072 20046 564328 20074
rect 88892 19100 88944 19106
rect 88892 19042 88944 19048
rect 86868 17944 86920 17950
rect 86868 17886 86920 17892
rect 51632 17740 51684 17746
rect 51632 17682 51684 17688
rect 31666 17640 31722 17649
rect 31666 17575 31722 17584
rect 28816 11008 28868 11014
rect 28816 10950 28868 10956
rect 27712 10940 27764 10946
rect 27712 10882 27764 10888
rect 27724 8226 27752 10882
rect 28828 8362 28856 10950
rect 28816 8356 28868 8362
rect 28816 8298 28868 8304
rect 27712 8220 27764 8226
rect 27712 8162 27764 8168
rect 29092 8220 29144 8226
rect 29092 8162 29144 8168
rect 29104 4282 29132 8162
rect 29092 4276 29144 4282
rect 29092 4218 29144 4224
rect 30288 3596 30340 3602
rect 30288 3538 30340 3544
rect 27632 3318 27936 3346
rect 27908 480 27936 3318
rect 29092 3120 29144 3126
rect 29092 3062 29144 3068
rect 29104 480 29132 3062
rect 30300 480 30328 3538
rect 31680 3346 31708 17575
rect 64786 17504 64842 17513
rect 34428 17468 34480 17474
rect 64786 17439 64842 17448
rect 34428 17410 34480 17416
rect 33048 16652 33100 16658
rect 33048 16594 33100 16600
rect 33060 3346 33088 16594
rect 33140 8288 33192 8294
rect 33140 8230 33192 8236
rect 31496 3318 31708 3346
rect 32692 3318 33088 3346
rect 31496 480 31524 3318
rect 32692 480 32720 3318
rect 33152 2922 33180 8230
rect 34440 3602 34468 17410
rect 41328 17400 41380 17406
rect 41328 17342 41380 17348
rect 39948 16720 40000 16726
rect 39948 16662 40000 16668
rect 34980 3664 35032 3670
rect 34980 3606 35032 3612
rect 33876 3596 33928 3602
rect 33876 3538 33928 3544
rect 34428 3596 34480 3602
rect 34428 3538 34480 3544
rect 33140 2916 33192 2922
rect 33140 2858 33192 2864
rect 33888 480 33916 3538
rect 34992 480 35020 3606
rect 39960 3482 39988 16662
rect 41340 3482 41368 17342
rect 42706 17232 42762 17241
rect 42706 17167 42762 17176
rect 42720 3602 42748 17167
rect 64696 17060 64748 17066
rect 64696 17002 64748 17008
rect 57888 16992 57940 16998
rect 57888 16934 57940 16940
rect 50988 16924 51040 16930
rect 50988 16866 51040 16872
rect 48136 16856 48188 16862
rect 48136 16798 48188 16804
rect 44088 16788 44140 16794
rect 44088 16730 44140 16736
rect 44100 3602 44128 16730
rect 44546 3904 44602 3913
rect 44546 3839 44602 3848
rect 42156 3596 42208 3602
rect 42156 3538 42208 3544
rect 42708 3596 42760 3602
rect 42708 3538 42760 3544
rect 43352 3596 43404 3602
rect 43352 3538 43404 3544
rect 44088 3596 44140 3602
rect 44088 3538 44140 3544
rect 39776 3454 39988 3482
rect 40972 3454 41368 3482
rect 37370 3360 37426 3369
rect 37370 3295 37426 3304
rect 38566 3360 38622 3369
rect 38566 3295 38622 3304
rect 36176 3188 36228 3194
rect 36176 3130 36228 3136
rect 36188 480 36216 3130
rect 37384 480 37412 3295
rect 38580 480 38608 3295
rect 39776 480 39804 3454
rect 40972 480 41000 3454
rect 42168 480 42196 3538
rect 43364 480 43392 3538
rect 44560 480 44588 3839
rect 48148 3602 48176 16798
rect 49608 5092 49660 5098
rect 49608 5034 49660 5040
rect 48228 5024 48280 5030
rect 48228 4966 48280 4972
rect 46940 3596 46992 3602
rect 46940 3538 46992 3544
rect 48136 3596 48188 3602
rect 48136 3538 48188 3544
rect 45744 2780 45796 2786
rect 45744 2722 45796 2728
rect 45756 480 45784 2722
rect 46952 480 46980 3538
rect 48240 2530 48268 4966
rect 49332 2848 49384 2854
rect 49332 2790 49384 2796
rect 48148 2502 48268 2530
rect 48148 480 48176 2502
rect 49344 480 49372 2790
rect 49620 2786 49648 5034
rect 51000 3602 51028 16866
rect 51632 4412 51684 4418
rect 51632 4354 51684 4360
rect 50528 3596 50580 3602
rect 50528 3538 50580 3544
rect 50988 3596 51040 3602
rect 50988 3538 51040 3544
rect 49608 2780 49660 2786
rect 49608 2722 49660 2728
rect 50540 480 50568 3538
rect 51644 480 51672 4354
rect 55220 4140 55272 4146
rect 55220 4082 55272 4088
rect 52828 3256 52880 3262
rect 52828 3198 52880 3204
rect 54024 3256 54076 3262
rect 54024 3198 54076 3204
rect 52840 480 52868 3198
rect 54036 480 54064 3198
rect 55232 480 55260 4082
rect 57900 3482 57928 16934
rect 62396 4616 62448 4622
rect 62396 4558 62448 4564
rect 58808 4480 58860 4486
rect 58808 4422 58860 4428
rect 57624 3454 57928 3482
rect 56416 3324 56468 3330
rect 56416 3266 56468 3272
rect 56428 480 56456 3266
rect 57624 480 57652 3454
rect 58820 480 58848 4422
rect 60004 3392 60056 3398
rect 60004 3334 60056 3340
rect 60016 480 60044 3334
rect 61200 3324 61252 3330
rect 61200 3266 61252 3272
rect 61212 480 61240 3266
rect 62408 480 62436 4558
rect 63592 4140 63644 4146
rect 63592 4082 63644 4088
rect 63604 480 63632 4082
rect 64708 3482 64736 17002
rect 64800 4146 64828 17439
rect 79968 17196 80020 17202
rect 79968 17138 80020 17144
rect 73068 17128 73120 17134
rect 73068 17070 73120 17076
rect 67180 6248 67232 6254
rect 67180 6190 67232 6196
rect 65984 4684 66036 4690
rect 65984 4626 66036 4632
rect 64788 4140 64840 4146
rect 64788 4082 64840 4088
rect 64708 3454 64828 3482
rect 64800 480 64828 3454
rect 65996 480 66024 4626
rect 67192 480 67220 6190
rect 69480 5092 69532 5098
rect 69480 5034 69532 5040
rect 68284 4140 68336 4146
rect 68284 4082 68336 4088
rect 68296 480 68324 4082
rect 69492 480 69520 5034
rect 70674 3768 70730 3777
rect 70674 3703 70730 3712
rect 70688 480 70716 3703
rect 72974 3632 73030 3641
rect 72974 3567 73030 3576
rect 71872 3392 71924 3398
rect 71872 3334 71924 3340
rect 71884 480 71912 3334
rect 72988 3210 73016 3567
rect 73080 3398 73108 17070
rect 77852 6316 77904 6322
rect 77852 6258 77904 6264
rect 75460 4140 75512 4146
rect 75460 4082 75512 4088
rect 74262 3496 74318 3505
rect 74262 3431 74318 3440
rect 73068 3392 73120 3398
rect 73068 3334 73120 3340
rect 72988 3182 73108 3210
rect 73080 480 73108 3182
rect 74276 480 74304 3431
rect 75472 480 75500 4082
rect 76656 4072 76708 4078
rect 76656 4014 76708 4020
rect 76668 480 76696 4014
rect 77864 480 77892 6258
rect 79980 4010 80008 17138
rect 80244 5160 80296 5166
rect 80244 5102 80296 5108
rect 79048 4004 79100 4010
rect 79048 3946 79100 3952
rect 79968 4004 80020 4010
rect 79968 3946 80020 3952
rect 79060 480 79088 3946
rect 80256 480 80284 5102
rect 83832 4548 83884 4554
rect 83832 4490 83884 4496
rect 82636 4004 82688 4010
rect 82636 3946 82688 3952
rect 81438 3496 81494 3505
rect 81438 3431 81494 3440
rect 81452 480 81480 3431
rect 82648 480 82676 3946
rect 83844 480 83872 4490
rect 84936 4072 84988 4078
rect 84936 4014 84988 4020
rect 84948 480 84976 4014
rect 86880 3874 86908 17886
rect 93768 17876 93820 17882
rect 93768 17818 93820 17824
rect 90916 5296 90968 5302
rect 90916 5238 90968 5244
rect 87328 5228 87380 5234
rect 87328 5170 87380 5176
rect 86132 3868 86184 3874
rect 86132 3810 86184 3816
rect 86868 3868 86920 3874
rect 86868 3810 86920 3816
rect 86144 480 86172 3810
rect 87340 480 87368 5170
rect 88524 3936 88576 3942
rect 88524 3878 88576 3884
rect 89720 3936 89772 3942
rect 89720 3878 89772 3884
rect 88536 480 88564 3878
rect 89732 480 89760 3878
rect 90928 480 90956 5238
rect 92112 4072 92164 4078
rect 92112 4014 92164 4020
rect 92124 480 92152 4014
rect 93780 3874 93808 17818
rect 97368 17542 97396 20046
rect 100668 17808 100720 17814
rect 100668 17750 100720 17756
rect 97356 17536 97408 17542
rect 97356 17478 97408 17484
rect 97908 3936 97960 3942
rect 97908 3878 97960 3884
rect 93308 3868 93360 3874
rect 93308 3810 93360 3816
rect 93768 3868 93820 3874
rect 93768 3810 93820 3816
rect 93320 480 93348 3810
rect 95698 3632 95754 3641
rect 95698 3567 95754 3576
rect 94504 2984 94556 2990
rect 94504 2926 94556 2932
rect 94516 480 94544 2926
rect 95712 480 95740 3567
rect 97920 2990 97948 3878
rect 99286 3768 99342 3777
rect 99286 3703 99342 3712
rect 96896 2984 96948 2990
rect 96896 2926 96948 2932
rect 97908 2984 97960 2990
rect 97908 2926 97960 2932
rect 96908 480 96936 2926
rect 98092 2916 98144 2922
rect 98092 2858 98144 2864
rect 98104 480 98132 2858
rect 99300 480 99328 3703
rect 100680 3482 100708 17750
rect 106568 17338 106596 20046
rect 114466 19952 114522 19961
rect 114466 19887 114522 19896
rect 107568 17740 107620 17746
rect 107568 17682 107620 17688
rect 106556 17332 106608 17338
rect 106556 17274 106608 17280
rect 101588 5296 101640 5302
rect 101588 5238 101640 5244
rect 100496 3454 100708 3482
rect 100496 480 100524 3454
rect 101600 480 101628 5238
rect 106370 4040 106426 4049
rect 106370 3975 106426 3984
rect 103980 3868 104032 3874
rect 103980 3810 104032 3816
rect 102784 3800 102836 3806
rect 102784 3742 102836 3748
rect 102796 480 102824 3742
rect 103992 480 104020 3810
rect 105176 2848 105228 2854
rect 105176 2790 105228 2796
rect 105188 480 105216 2790
rect 106384 480 106412 3975
rect 107580 480 107608 17682
rect 108764 5364 108816 5370
rect 108764 5306 108816 5312
rect 108776 480 108804 5306
rect 112352 4344 112404 4350
rect 112352 4286 112404 4292
rect 109958 3904 110014 3913
rect 109958 3839 110014 3848
rect 109972 480 110000 3839
rect 111156 2984 111208 2990
rect 111156 2926 111208 2932
rect 111168 480 111196 2926
rect 112364 480 112392 4286
rect 114480 3738 114508 19887
rect 115848 17672 115900 17678
rect 115848 17614 115900 17620
rect 115860 3738 115888 17614
rect 113548 3732 113600 3738
rect 113548 3674 113600 3680
rect 114468 3732 114520 3738
rect 114468 3674 114520 3680
rect 114744 3732 114796 3738
rect 114744 3674 114796 3680
rect 115848 3732 115900 3738
rect 115848 3674 115900 3680
rect 113560 480 113588 3674
rect 114756 480 114784 3674
rect 115952 2922 115980 20046
rect 122748 17604 122800 17610
rect 122748 17546 122800 17552
rect 117136 17332 117188 17338
rect 117136 17274 117188 17280
rect 116032 5432 116084 5438
rect 116032 5374 116084 5380
rect 115940 2916 115992 2922
rect 115940 2858 115992 2864
rect 116044 2802 116072 5374
rect 115952 2774 116072 2802
rect 115952 480 115980 2774
rect 117148 480 117176 17274
rect 119436 4276 119488 4282
rect 119436 4218 119488 4224
rect 118240 2984 118292 2990
rect 118240 2926 118292 2932
rect 118252 480 118280 2926
rect 119448 480 119476 4218
rect 122760 3738 122788 17546
rect 124784 17270 124812 20046
rect 125508 17536 125560 17542
rect 125508 17478 125560 17484
rect 124772 17264 124824 17270
rect 124772 17206 124824 17212
rect 125416 17264 125468 17270
rect 125416 17206 125468 17212
rect 123024 6384 123076 6390
rect 123024 6326 123076 6332
rect 121828 3732 121880 3738
rect 121828 3674 121880 3680
rect 122748 3732 122800 3738
rect 122748 3674 122800 3680
rect 120632 3052 120684 3058
rect 120632 2994 120684 3000
rect 120644 480 120672 2994
rect 121840 480 121868 3674
rect 123036 480 123064 6326
rect 125428 3738 125456 17206
rect 124220 3732 124272 3738
rect 124220 3674 124272 3680
rect 125416 3732 125468 3738
rect 125416 3674 125468 3680
rect 124232 480 124260 3674
rect 125520 3482 125548 17478
rect 125428 3454 125548 3482
rect 125428 480 125456 3454
rect 133892 3126 133920 20046
rect 143092 16658 143120 20046
rect 143080 16652 143132 16658
rect 143080 16594 143132 16600
rect 151832 3194 151860 20046
rect 161584 16726 161612 20046
rect 170600 16794 170628 20046
rect 179708 16862 179736 20046
rect 189092 16930 189120 20046
rect 189080 16924 189132 16930
rect 189080 16866 189132 16872
rect 179696 16856 179748 16862
rect 179696 16798 179748 16804
rect 170588 16788 170640 16794
rect 170588 16730 170640 16736
rect 161572 16720 161624 16726
rect 161572 16662 161624 16668
rect 197372 3262 197400 20046
rect 207216 16998 207244 20046
rect 207204 16992 207256 16998
rect 207204 16934 207256 16940
rect 215312 3330 215340 20046
rect 225432 17066 225460 20046
rect 225420 17060 225472 17066
rect 225420 17002 225472 17008
rect 234632 3398 234660 20046
rect 243740 17134 243768 20046
rect 243728 17128 243780 17134
rect 243728 17070 243780 17076
rect 252572 4146 252600 20046
rect 262232 17202 262260 20046
rect 262220 17196 262272 17202
rect 262220 17138 262272 17144
rect 252560 4140 252612 4146
rect 252560 4082 252612 4088
rect 270512 4078 270540 20046
rect 280356 17950 280384 20046
rect 280344 17944 280396 17950
rect 280344 17886 280396 17892
rect 270500 4072 270552 4078
rect 270500 4014 270552 4020
rect 289832 4010 289860 20046
rect 298664 17882 298692 20046
rect 298652 17876 298704 17882
rect 298652 17818 298704 17824
rect 289820 4004 289872 4010
rect 289820 3946 289872 3952
rect 307772 3942 307800 20046
rect 316972 17814 317000 20046
rect 316960 17808 317012 17814
rect 316960 17750 317012 17756
rect 307760 3936 307812 3942
rect 307760 3878 307812 3884
rect 325712 3874 325740 20046
rect 335464 17746 335492 20046
rect 335452 17740 335504 17746
rect 335452 17682 335504 17688
rect 325700 3868 325752 3874
rect 325700 3810 325752 3816
rect 343652 3806 343680 20046
rect 353588 17678 353616 20046
rect 353576 17672 353628 17678
rect 353576 17614 353628 17620
rect 343640 3800 343692 3806
rect 343640 3742 343692 3748
rect 362972 3738 363000 20046
rect 371896 17610 371924 20046
rect 371884 17604 371936 17610
rect 371884 17546 371936 17552
rect 381004 17542 381032 20046
rect 380992 17536 381044 17542
rect 380992 17478 381044 17484
rect 389192 4758 389220 20046
rect 398852 5506 398880 20046
rect 408512 17474 408540 20046
rect 408500 17468 408552 17474
rect 408500 17410 408552 17416
rect 417620 17406 417648 20046
rect 417608 17400 417660 17406
rect 417608 17342 417660 17348
rect 398840 5500 398892 5506
rect 398840 5442 398892 5448
rect 389180 4752 389232 4758
rect 389180 4694 389232 4700
rect 426452 4418 426480 20046
rect 436112 4486 436140 20046
rect 444392 4622 444420 20046
rect 454052 4690 454080 20046
rect 454040 4684 454092 4690
rect 454040 4626 454092 4632
rect 444380 4616 444432 4622
rect 444380 4558 444432 4564
rect 462332 4554 462360 20046
rect 462320 4548 462372 4554
rect 462320 4490 462372 4496
rect 436100 4480 436152 4486
rect 436100 4422 436152 4428
rect 426440 4412 426492 4418
rect 426440 4354 426492 4360
rect 471992 4350 472020 20046
rect 481652 17377 481680 20046
rect 490760 17649 490788 20046
rect 490746 17640 490802 17649
rect 490746 17575 490802 17584
rect 481638 17368 481694 17377
rect 481638 17303 481694 17312
rect 471980 4344 472032 4350
rect 471980 4286 472032 4292
rect 362960 3732 363012 3738
rect 362960 3674 363012 3680
rect 499592 3670 499620 20046
rect 509252 17241 509280 20046
rect 509238 17232 509294 17241
rect 509238 17167 509294 17176
rect 499580 3664 499632 3670
rect 499580 3606 499632 3612
rect 517532 3602 517560 20046
rect 527376 17513 527404 20046
rect 527362 17504 527418 17513
rect 527362 17439 527418 17448
rect 536852 17338 536880 20046
rect 536840 17332 536892 17338
rect 536840 17274 536892 17280
rect 545684 17270 545712 20046
rect 545672 17264 545724 17270
rect 545672 17206 545724 17212
rect 517520 3596 517572 3602
rect 517520 3538 517572 3544
rect 554792 3534 554820 20046
rect 554780 3528 554832 3534
rect 554780 3470 554832 3476
rect 563072 3466 563100 20046
rect 571352 6322 571380 600879
rect 571430 577280 571486 577289
rect 571430 577215 571486 577224
rect 571340 6316 571392 6322
rect 571340 6258 571392 6264
rect 571444 6254 571472 577215
rect 571522 553480 571578 553489
rect 571522 553415 571578 553424
rect 571432 6248 571484 6254
rect 571432 6190 571484 6196
rect 563060 3460 563112 3466
rect 563060 3402 563112 3408
rect 234620 3392 234672 3398
rect 571536 3369 571564 553415
rect 571614 529816 571670 529825
rect 571614 529751 571670 529760
rect 571628 6186 571656 529751
rect 571706 506152 571762 506161
rect 571706 506087 571762 506096
rect 571720 6390 571748 506087
rect 579712 487144 579764 487150
rect 579712 487086 579764 487092
rect 579724 486849 579752 487086
rect 579710 486840 579766 486849
rect 579710 486775 579766 486784
rect 571798 482352 571854 482361
rect 571798 482287 571854 482296
rect 571708 6384 571760 6390
rect 571708 6326 571760 6332
rect 571616 6180 571668 6186
rect 571616 6122 571668 6128
rect 571812 5438 571840 482287
rect 571890 458688 571946 458697
rect 571890 458623 571946 458632
rect 571800 5432 571852 5438
rect 571800 5374 571852 5380
rect 571904 5370 571932 458623
rect 578882 439920 578938 439929
rect 578882 439855 578938 439864
rect 571982 435024 572038 435033
rect 571982 434959 572038 434968
rect 571892 5364 571944 5370
rect 571892 5306 571944 5312
rect 571996 5302 572024 434959
rect 572074 411224 572130 411233
rect 572074 411159 572130 411168
rect 571984 5296 572036 5302
rect 571984 5238 572036 5244
rect 572088 5234 572116 411159
rect 573364 392012 573416 392018
rect 573364 391954 573416 391960
rect 572166 387560 572222 387569
rect 572166 387495 572222 387504
rect 572076 5228 572128 5234
rect 572076 5170 572128 5176
rect 572180 5166 572208 387495
rect 572258 363896 572314 363905
rect 572258 363831 572314 363840
rect 572168 5160 572220 5166
rect 572168 5102 572220 5108
rect 572272 5098 572300 363831
rect 572350 340096 572406 340105
rect 572350 340031 572406 340040
rect 572260 5092 572312 5098
rect 572260 5034 572312 5040
rect 572364 5030 572392 340031
rect 572442 316432 572498 316441
rect 572442 316367 572498 316376
rect 572352 5024 572404 5030
rect 572352 4966 572404 4972
rect 572456 4962 572484 316367
rect 572534 292632 572590 292641
rect 572534 292567 572590 292576
rect 572444 4956 572496 4962
rect 572444 4898 572496 4904
rect 572548 4894 572576 292567
rect 572626 268968 572682 268977
rect 572626 268903 572682 268912
rect 572536 4888 572588 4894
rect 572536 4830 572588 4836
rect 572640 4826 572668 268903
rect 573376 221542 573404 391954
rect 577504 345568 577556 345574
rect 577504 345510 577556 345516
rect 574744 298172 574796 298178
rect 574744 298114 574796 298120
rect 573364 221536 573416 221542
rect 573364 221478 573416 221484
rect 573364 204332 573416 204338
rect 573364 204274 573416 204280
rect 573376 126750 573404 204274
rect 574756 174214 574784 298114
rect 576124 251252 576176 251258
rect 576124 251194 576176 251200
rect 574744 174208 574796 174214
rect 574744 174150 574796 174156
rect 574744 157412 574796 157418
rect 574744 157354 574796 157360
rect 573364 126744 573416 126750
rect 573364 126686 573416 126692
rect 573364 110492 573416 110498
rect 573364 110434 573416 110440
rect 573376 79286 573404 110434
rect 574756 103086 574784 157354
rect 576136 150414 576164 251194
rect 577516 197470 577544 345510
rect 578896 244390 578924 439855
rect 579618 393000 579674 393009
rect 579618 392935 579674 392944
rect 579632 392018 579660 392935
rect 579620 392012 579672 392018
rect 579620 391954 579672 391960
rect 579618 346080 579674 346089
rect 579618 346015 579674 346024
rect 579632 345574 579660 346015
rect 579620 345568 579672 345574
rect 579620 345510 579672 345516
rect 579618 299160 579674 299169
rect 579618 299095 579674 299104
rect 579632 298178 579660 299095
rect 579620 298172 579672 298178
rect 579620 298114 579672 298120
rect 579618 252240 579674 252249
rect 579618 252175 579674 252184
rect 579632 251258 579660 252175
rect 579620 251252 579672 251258
rect 579620 251194 579672 251200
rect 578884 244384 578936 244390
rect 578884 244326 578936 244332
rect 579618 205320 579674 205329
rect 579618 205255 579674 205264
rect 579632 204338 579660 205255
rect 579620 204332 579672 204338
rect 579620 204274 579672 204280
rect 577504 197464 577556 197470
rect 577504 197406 577556 197412
rect 579618 158400 579674 158409
rect 579618 158335 579674 158344
rect 579632 157418 579660 158335
rect 579620 157412 579672 157418
rect 579620 157354 579672 157360
rect 576124 150408 576176 150414
rect 576124 150350 576176 150356
rect 579618 111480 579674 111489
rect 579618 111415 579674 111424
rect 579632 110498 579660 111415
rect 579620 110492 579672 110498
rect 579620 110434 579672 110440
rect 574744 103080 574796 103086
rect 574744 103022 574796 103028
rect 573364 79280 573416 79286
rect 573364 79222 573416 79228
rect 580170 64560 580226 64569
rect 580170 64495 580226 64504
rect 580184 63578 580212 64495
rect 577412 63572 577464 63578
rect 577412 63514 577464 63520
rect 580172 63572 580224 63578
rect 580172 63514 580224 63520
rect 577424 55350 577452 63514
rect 577412 55344 577464 55350
rect 577412 55286 577464 55292
rect 573362 31920 573418 31929
rect 573362 31855 573418 31864
rect 573376 17950 573404 31855
rect 580276 19106 580304 686287
rect 580354 639432 580410 639441
rect 580354 639367 580410 639376
rect 580368 19174 580396 639367
rect 580446 592512 580502 592521
rect 580446 592447 580502 592456
rect 580460 19242 580488 592447
rect 580538 545592 580594 545601
rect 580538 545527 580594 545536
rect 580552 19310 580580 545527
rect 580540 19304 580592 19310
rect 580540 19246 580592 19252
rect 580448 19236 580500 19242
rect 580448 19178 580500 19184
rect 580356 19168 580408 19174
rect 580356 19110 580408 19116
rect 580264 19100 580316 19106
rect 580264 19042 580316 19048
rect 573364 17944 573416 17950
rect 573364 17886 573416 17892
rect 579804 17944 579856 17950
rect 579804 17886 579856 17892
rect 579816 17649 579844 17886
rect 579802 17640 579858 17649
rect 579802 17575 579858 17584
rect 572628 4820 572680 4826
rect 572628 4762 572680 4768
rect 234620 3334 234672 3340
rect 571522 3360 571578 3369
rect 215300 3324 215352 3330
rect 571522 3295 571578 3304
rect 215300 3266 215352 3272
rect 197360 3256 197412 3262
rect 197360 3198 197412 3204
rect 151820 3188 151872 3194
rect 151820 3130 151872 3136
rect 133880 3120 133932 3126
rect 133880 3062 133932 3068
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 667956 3478 667992
rect 3422 667936 3424 667956
rect 3424 667936 3476 667956
rect 3476 667936 3478 667956
rect 3422 610408 3478 610464
rect 3146 553016 3202 553072
rect 3422 495488 3478 495544
rect 3330 323040 3386 323096
rect 3330 107616 3386 107672
rect 3330 64504 3386 64560
rect 3146 21392 3202 21448
rect 3514 437960 3570 438016
rect 3514 380568 3570 380624
rect 3606 280064 3662 280120
rect 3698 236952 3754 237008
rect 3882 193840 3938 193896
rect 3790 150728 3846 150784
rect 17866 670520 17922 670576
rect 17866 644000 17922 644056
rect 17866 617480 17922 617536
rect 17774 590824 17830 590880
rect 17682 564304 17738 564360
rect 17590 537784 17646 537840
rect 17498 511264 17554 511320
rect 17406 484608 17462 484664
rect 17314 431568 17370 431624
rect 17222 404912 17278 404968
rect 17130 378392 17186 378448
rect 17038 351908 17040 351928
rect 17040 351908 17092 351928
rect 17092 351908 17094 351928
rect 17038 351872 17094 351908
rect 17038 325352 17094 325408
rect 17038 298696 17094 298752
rect 17038 272176 17094 272232
rect 17038 245676 17094 245712
rect 17038 245656 17040 245676
rect 17040 245656 17092 245676
rect 17092 245656 17094 245676
rect 17038 219000 17094 219056
rect 17038 192480 17094 192536
rect 17038 165960 17094 166016
rect 16762 139440 16818 139496
rect 17038 112784 17094 112840
rect 17038 86264 17094 86320
rect 16946 59744 17002 59800
rect 17038 33224 17094 33280
rect 19246 458088 19302 458144
rect 19154 17312 19210 17368
rect 223578 686296 223634 686352
rect 240966 686160 241022 686216
rect 258722 686024 258778 686080
rect 347226 686024 347282 686080
rect 542726 686160 542782 686216
rect 524970 686024 525026 686080
rect 471242 685888 471298 685944
rect 507306 685888 507362 685944
rect 580262 686296 580318 686352
rect 293866 683712 293922 683768
rect 329746 683440 329802 683496
rect 311806 683304 311862 683360
rect 22374 682760 22430 682816
rect 22282 682624 22338 682680
rect 22558 682488 22614 682544
rect 22466 682352 22522 682408
rect 571338 600888 571394 600944
rect 571246 244704 571302 244760
rect 571246 221484 571248 221504
rect 571248 221484 571300 221504
rect 571300 221484 571302 221504
rect 571246 221448 571302 221484
rect 571246 197512 571302 197568
rect 571246 174156 571248 174176
rect 571248 174156 571300 174176
rect 571300 174156 571302 174176
rect 571246 174120 571302 174156
rect 571246 150356 571248 150376
rect 571248 150356 571300 150376
rect 571300 150356 571302 150376
rect 571246 150320 571302 150356
rect 571246 126692 571248 126712
rect 571248 126692 571300 126712
rect 571300 126692 571302 126712
rect 571246 126656 571302 126692
rect 571246 103028 571248 103048
rect 571248 103028 571300 103048
rect 571300 103028 571302 103048
rect 571246 102992 571302 103028
rect 571246 79228 571248 79248
rect 571248 79228 571300 79248
rect 571300 79228 571302 79248
rect 571246 79192 571302 79228
rect 571246 55292 571248 55312
rect 571248 55292 571300 55312
rect 571300 55292 571302 55312
rect 571246 55256 571302 55292
rect 21638 3440 21694 3496
rect 31666 17584 31722 17640
rect 64786 17448 64842 17504
rect 42706 17176 42762 17232
rect 44546 3848 44602 3904
rect 37370 3304 37426 3360
rect 38566 3304 38622 3360
rect 70674 3712 70730 3768
rect 72974 3576 73030 3632
rect 74262 3440 74318 3496
rect 81438 3440 81494 3496
rect 95698 3576 95754 3632
rect 99286 3712 99342 3768
rect 114466 19896 114522 19952
rect 106370 3984 106426 4040
rect 109958 3848 110014 3904
rect 490746 17584 490802 17640
rect 481638 17312 481694 17368
rect 509238 17176 509294 17232
rect 527362 17448 527418 17504
rect 571430 577224 571486 577280
rect 571522 553424 571578 553480
rect 571614 529760 571670 529816
rect 571706 506096 571762 506152
rect 579710 486784 579766 486840
rect 571798 482296 571854 482352
rect 571890 458632 571946 458688
rect 578882 439864 578938 439920
rect 571982 434968 572038 435024
rect 572074 411168 572130 411224
rect 572166 387504 572222 387560
rect 572258 363840 572314 363896
rect 572350 340040 572406 340096
rect 572442 316376 572498 316432
rect 572534 292576 572590 292632
rect 572626 268912 572682 268968
rect 579618 392944 579674 393000
rect 579618 346024 579674 346080
rect 579618 299104 579674 299160
rect 579618 252184 579674 252240
rect 579618 205264 579674 205320
rect 579618 158344 579674 158400
rect 579618 111424 579674 111480
rect 580170 64504 580226 64560
rect 573362 31864 573418 31920
rect 580354 639376 580410 639432
rect 580446 592456 580502 592512
rect 580538 545536 580594 545592
rect 579802 17584 579858 17640
rect 571522 3304 571578 3360
<< metal3 >>
rect 583520 697900 584960 698140
rect -960 696540 480 696780
rect 23238 686292 23244 686356
rect 23308 686354 23314 686356
rect 223573 686354 223639 686357
rect 23308 686352 223639 686354
rect 23308 686296 223578 686352
rect 223634 686296 223639 686352
rect 23308 686294 223639 686296
rect 23308 686292 23314 686294
rect 223573 686291 223639 686294
rect 580257 686354 580323 686357
rect 583520 686354 584960 686444
rect 580257 686352 584960 686354
rect 580257 686296 580262 686352
rect 580318 686296 584960 686352
rect 580257 686294 584960 686296
rect 580257 686291 580323 686294
rect 23054 686156 23060 686220
rect 23124 686218 23130 686220
rect 240961 686218 241027 686221
rect 23124 686216 241027 686218
rect 23124 686160 240966 686216
rect 241022 686160 241027 686216
rect 23124 686158 241027 686160
rect 23124 686156 23130 686158
rect 240961 686155 241027 686158
rect 542721 686218 542787 686221
rect 561622 686218 561628 686220
rect 542721 686216 561628 686218
rect 542721 686160 542726 686216
rect 542782 686160 561628 686216
rect 542721 686158 561628 686160
rect 542721 686155 542787 686158
rect 561622 686156 561628 686158
rect 561692 686156 561698 686220
rect 583520 686204 584960 686294
rect 23606 686020 23612 686084
rect 23676 686082 23682 686084
rect 258717 686082 258783 686085
rect 23676 686080 258783 686082
rect 23676 686024 258722 686080
rect 258778 686024 258783 686080
rect 23676 686022 258783 686024
rect 23676 686020 23682 686022
rect 258717 686019 258783 686022
rect 337326 686020 337332 686084
rect 337396 686082 337402 686084
rect 347221 686082 347287 686085
rect 337396 686080 347287 686082
rect 337396 686024 347226 686080
rect 347282 686024 347287 686080
rect 337396 686022 347287 686024
rect 337396 686020 337402 686022
rect 347221 686019 347287 686022
rect 524965 686082 525031 686085
rect 563278 686082 563284 686084
rect 524965 686080 563284 686082
rect 524965 686024 524970 686080
rect 525026 686024 563284 686080
rect 524965 686022 563284 686024
rect 524965 686019 525031 686022
rect 563278 686020 563284 686022
rect 563348 686020 563354 686084
rect 22870 685884 22876 685948
rect 22940 685946 22946 685948
rect 471237 685946 471303 685949
rect 22940 685944 471303 685946
rect 22940 685888 471242 685944
rect 471298 685888 471303 685944
rect 22940 685886 471303 685888
rect 22940 685884 22946 685886
rect 471237 685883 471303 685886
rect 507301 685946 507367 685949
rect 563094 685946 563100 685948
rect 507301 685944 563100 685946
rect 507301 685888 507306 685944
rect 507362 685888 563100 685944
rect 507301 685886 563100 685888
rect 507301 685883 507367 685886
rect 563094 685884 563100 685886
rect 563164 685884 563170 685948
rect 284886 683708 284892 683772
rect 284956 683770 284962 683772
rect 293861 683770 293927 683773
rect 284956 683768 293927 683770
rect 284956 683712 293866 683768
rect 293922 683712 293927 683768
rect 284956 683710 293927 683712
rect 284956 683708 284962 683710
rect 293861 683707 293927 683710
rect 323158 683436 323164 683500
rect 323228 683498 323234 683500
rect 329741 683498 329807 683501
rect 323228 683496 329807 683498
rect 323228 683440 329746 683496
rect 329802 683440 329807 683496
rect 323228 683438 329807 683440
rect 323228 683436 323234 683438
rect 329741 683435 329807 683438
rect 311801 683364 311867 683365
rect 311750 683362 311756 683364
rect 311710 683302 311756 683362
rect 311820 683360 311867 683364
rect 311862 683304 311867 683360
rect 311750 683300 311756 683302
rect 311820 683300 311867 683304
rect 311801 683299 311867 683300
rect 22369 682818 22435 682821
rect 284886 682818 284892 682820
rect 22369 682816 284892 682818
rect 22369 682760 22374 682816
rect 22430 682760 284892 682816
rect 22369 682758 284892 682760
rect 22369 682755 22435 682758
rect 284886 682756 284892 682758
rect 284956 682756 284962 682820
rect 22277 682682 22343 682685
rect 311750 682682 311756 682684
rect 22277 682680 311756 682682
rect 22277 682624 22282 682680
rect 22338 682624 311756 682680
rect 22277 682622 311756 682624
rect 22277 682619 22343 682622
rect 311750 682620 311756 682622
rect 311820 682620 311826 682684
rect 22553 682546 22619 682549
rect 323158 682546 323164 682548
rect 22553 682544 323164 682546
rect 22553 682488 22558 682544
rect 22614 682488 323164 682544
rect 22553 682486 323164 682488
rect 22553 682483 22619 682486
rect 323158 682484 323164 682486
rect 323228 682484 323234 682548
rect 22461 682410 22527 682413
rect 337326 682410 337332 682412
rect 22461 682408 337332 682410
rect -960 682124 480 682364
rect 22461 682352 22466 682408
rect 22522 682352 337332 682408
rect 22461 682350 337332 682352
rect 22461 682347 22527 682350
rect 337326 682348 337332 682350
rect 337396 682348 337402 682412
rect 583520 674508 584960 674748
rect 571374 672074 571380 672076
rect 568836 672014 571380 672074
rect 571374 672012 571380 672014
rect 571444 672012 571450 672076
rect 17861 670578 17927 670581
rect 17861 670576 20148 670578
rect 17861 670520 17866 670576
rect 17922 670520 20148 670576
rect 17861 670518 20148 670520
rect 17861 670515 17927 670518
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 583520 662676 584960 662916
rect -960 653428 480 653668
rect 583520 650980 584960 651220
rect 571558 648410 571564 648412
rect 568836 648350 571564 648410
rect 571558 648348 571564 648350
rect 571628 648348 571634 648412
rect 17861 644058 17927 644061
rect 17861 644056 20148 644058
rect 17861 644000 17866 644056
rect 17922 644000 20148 644056
rect 17861 643998 20148 644000
rect 17861 643995 17927 643998
rect 580349 639434 580415 639437
rect 583520 639434 584960 639524
rect 580349 639432 584960 639434
rect 580349 639376 580354 639432
rect 580410 639376 584960 639432
rect 580349 639374 584960 639376
rect 580349 639371 580415 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 583520 627588 584960 627828
rect -960 624732 480 624972
rect 571742 624610 571748 624612
rect 568836 624550 571748 624610
rect 571742 624548 571748 624550
rect 571812 624548 571818 624612
rect 17861 617538 17927 617541
rect 17861 617536 20148 617538
rect 17861 617480 17866 617536
rect 17922 617480 20148 617536
rect 17861 617478 20148 617480
rect 17861 617475 17927 617478
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3417 610466 3483 610469
rect -960 610464 3483 610466
rect -960 610408 3422 610464
rect 3478 610408 3483 610464
rect -960 610406 3483 610408
rect -960 610316 480 610406
rect 3417 610403 3483 610406
rect 583520 604060 584960 604300
rect 571333 600946 571399 600949
rect 568836 600944 571399 600946
rect 568836 600888 571338 600944
rect 571394 600888 571399 600944
rect 568836 600886 571399 600888
rect 571333 600883 571399 600886
rect -960 595900 480 596140
rect 580441 592514 580507 592517
rect 583520 592514 584960 592604
rect 580441 592512 584960 592514
rect 580441 592456 580446 592512
rect 580502 592456 584960 592512
rect 580441 592454 584960 592456
rect 580441 592451 580507 592454
rect 583520 592364 584960 592454
rect 17769 590882 17835 590885
rect 17769 590880 20148 590882
rect 17769 590824 17774 590880
rect 17830 590824 20148 590880
rect 17769 590822 20148 590824
rect 17769 590819 17835 590822
rect -960 581620 480 581860
rect 583520 580668 584960 580908
rect 571425 577282 571491 577285
rect 568836 577280 571491 577282
rect 568836 577224 571430 577280
rect 571486 577224 571491 577280
rect 568836 577222 571491 577224
rect 571425 577219 571491 577222
rect 583520 568836 584960 569076
rect -960 567204 480 567444
rect 17677 564362 17743 564365
rect 17677 564360 20148 564362
rect 17677 564304 17682 564360
rect 17738 564304 20148 564360
rect 17677 564302 20148 564304
rect 17677 564299 17743 564302
rect 583520 557140 584960 557380
rect 571517 553482 571583 553485
rect 568836 553480 571583 553482
rect 568836 553424 571522 553480
rect 571578 553424 571583 553480
rect 568836 553422 571583 553424
rect 571517 553419 571583 553422
rect -960 553074 480 553164
rect 3141 553074 3207 553077
rect -960 553072 3207 553074
rect -960 553016 3146 553072
rect 3202 553016 3207 553072
rect -960 553014 3207 553016
rect -960 552924 480 553014
rect 3141 553011 3207 553014
rect 580533 545594 580599 545597
rect 583520 545594 584960 545684
rect 580533 545592 584960 545594
rect 580533 545536 580538 545592
rect 580594 545536 584960 545592
rect 580533 545534 584960 545536
rect 580533 545531 580599 545534
rect 583520 545444 584960 545534
rect -960 538508 480 538748
rect 17585 537842 17651 537845
rect 17585 537840 20148 537842
rect 17585 537784 17590 537840
rect 17646 537784 20148 537840
rect 17585 537782 20148 537784
rect 17585 537779 17651 537782
rect 583520 533748 584960 533988
rect 571609 529818 571675 529821
rect 568836 529816 571675 529818
rect 568836 529760 571614 529816
rect 571670 529760 571675 529816
rect 568836 529758 571675 529760
rect 571609 529755 571675 529758
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 17493 511322 17559 511325
rect 17493 511320 20148 511322
rect 17493 511264 17498 511320
rect 17554 511264 20148 511320
rect 17493 511262 20148 511264
rect 17493 511259 17559 511262
rect 583520 510220 584960 510460
rect -960 509812 480 510052
rect 571701 506154 571767 506157
rect 568836 506152 571767 506154
rect 568836 506096 571706 506152
rect 571762 506096 571767 506152
rect 568836 506094 571767 506096
rect 571701 506091 571767 506094
rect 583520 498524 584960 498764
rect -960 495546 480 495636
rect 3417 495546 3483 495549
rect -960 495544 3483 495546
rect -960 495488 3422 495544
rect 3478 495488 3483 495544
rect -960 495486 3483 495488
rect -960 495396 480 495486
rect 3417 495483 3483 495486
rect 579705 486842 579771 486845
rect 583520 486842 584960 486932
rect 579705 486840 584960 486842
rect 579705 486784 579710 486840
rect 579766 486784 584960 486840
rect 579705 486782 584960 486784
rect 579705 486779 579771 486782
rect 583520 486692 584960 486782
rect 17401 484666 17467 484669
rect 17401 484664 20148 484666
rect 17401 484608 17406 484664
rect 17462 484608 20148 484664
rect 17401 484606 20148 484608
rect 17401 484603 17467 484606
rect 571793 482354 571859 482357
rect 568836 482352 571859 482354
rect 568836 482296 571798 482352
rect 571854 482296 571859 482352
rect 568836 482294 571859 482296
rect 571793 482291 571859 482294
rect -960 480980 480 481220
rect 583520 474996 584960 475236
rect -960 466700 480 466940
rect 583520 463300 584960 463540
rect 571885 458690 571951 458693
rect 568836 458688 571951 458690
rect 568836 458632 571890 458688
rect 571946 458632 571951 458688
rect 568836 458630 571951 458632
rect 571885 458627 571951 458630
rect 19241 458146 19307 458149
rect 19241 458144 20148 458146
rect 19241 458088 19246 458144
rect 19302 458088 20148 458144
rect 19241 458086 20148 458088
rect 19241 458083 19307 458086
rect -960 452284 480 452524
rect 583520 451604 584960 451844
rect 578877 439922 578943 439925
rect 583520 439922 584960 440012
rect 578877 439920 584960 439922
rect 578877 439864 578882 439920
rect 578938 439864 584960 439920
rect 578877 439862 584960 439864
rect 578877 439859 578943 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 3509 438018 3575 438021
rect -960 438016 3575 438018
rect -960 437960 3514 438016
rect 3570 437960 3575 438016
rect -960 437958 3575 437960
rect -960 437868 480 437958
rect 3509 437955 3575 437958
rect 571977 435026 572043 435029
rect 568836 435024 572043 435026
rect 568836 434968 571982 435024
rect 572038 434968 572043 435024
rect 568836 434966 572043 434968
rect 571977 434963 572043 434966
rect 17309 431626 17375 431629
rect 17309 431624 20148 431626
rect 17309 431568 17314 431624
rect 17370 431568 20148 431624
rect 17309 431566 20148 431568
rect 17309 431563 17375 431566
rect 583520 428076 584960 428316
rect -960 423588 480 423828
rect 583520 416380 584960 416620
rect 572069 411226 572135 411229
rect 568836 411224 572135 411226
rect 568836 411168 572074 411224
rect 572130 411168 572135 411224
rect 568836 411166 572135 411168
rect 572069 411163 572135 411166
rect -960 409172 480 409412
rect 17217 404970 17283 404973
rect 17217 404968 20148 404970
rect 17217 404912 17222 404968
rect 17278 404912 20148 404968
rect 17217 404910 20148 404912
rect 17217 404907 17283 404910
rect 583520 404684 584960 404924
rect -960 394892 480 395132
rect 579613 393002 579679 393005
rect 583520 393002 584960 393092
rect 579613 393000 584960 393002
rect 579613 392944 579618 393000
rect 579674 392944 584960 393000
rect 579613 392942 584960 392944
rect 579613 392939 579679 392942
rect 583520 392852 584960 392942
rect 572161 387562 572227 387565
rect 568836 387560 572227 387562
rect 568836 387504 572166 387560
rect 572222 387504 572227 387560
rect 568836 387502 572227 387504
rect 572161 387499 572227 387502
rect 583520 381156 584960 381396
rect -960 380626 480 380716
rect 3509 380626 3575 380629
rect -960 380624 3575 380626
rect -960 380568 3514 380624
rect 3570 380568 3575 380624
rect -960 380566 3575 380568
rect -960 380476 480 380566
rect 3509 380563 3575 380566
rect 17125 378450 17191 378453
rect 17125 378448 20148 378450
rect 17125 378392 17130 378448
rect 17186 378392 20148 378448
rect 17125 378390 20148 378392
rect 17125 378387 17191 378390
rect 583520 369460 584960 369700
rect -960 366060 480 366300
rect 572253 363898 572319 363901
rect 568836 363896 572319 363898
rect 568836 363840 572258 363896
rect 572314 363840 572319 363896
rect 568836 363838 572319 363840
rect 572253 363835 572319 363838
rect 583520 357764 584960 358004
rect -960 351780 480 352020
rect 17033 351930 17099 351933
rect 17033 351928 20148 351930
rect 17033 351872 17038 351928
rect 17094 351872 20148 351928
rect 17033 351870 20148 351872
rect 17033 351867 17099 351870
rect 579613 346082 579679 346085
rect 583520 346082 584960 346172
rect 579613 346080 584960 346082
rect 579613 346024 579618 346080
rect 579674 346024 584960 346080
rect 579613 346022 584960 346024
rect 579613 346019 579679 346022
rect 583520 345932 584960 346022
rect 572345 340098 572411 340101
rect 568836 340096 572411 340098
rect 568836 340040 572350 340096
rect 572406 340040 572411 340096
rect 568836 340038 572411 340040
rect 572345 340035 572411 340038
rect -960 337364 480 337604
rect 583520 334236 584960 334476
rect 17033 325410 17099 325413
rect 17033 325408 20148 325410
rect 17033 325352 17038 325408
rect 17094 325352 20148 325408
rect 17033 325350 20148 325352
rect 17033 325347 17099 325350
rect -960 323098 480 323188
rect 3325 323098 3391 323101
rect -960 323096 3391 323098
rect -960 323040 3330 323096
rect 3386 323040 3391 323096
rect -960 323038 3391 323040
rect -960 322948 480 323038
rect 3325 323035 3391 323038
rect 583520 322540 584960 322780
rect 572437 316434 572503 316437
rect 568836 316432 572503 316434
rect 568836 316376 572442 316432
rect 572498 316376 572503 316432
rect 568836 316374 572503 316376
rect 572437 316371 572503 316374
rect 583520 310708 584960 310948
rect -960 308668 480 308908
rect 579613 299162 579679 299165
rect 583520 299162 584960 299252
rect 579613 299160 584960 299162
rect 579613 299104 579618 299160
rect 579674 299104 584960 299160
rect 579613 299102 584960 299104
rect 579613 299099 579679 299102
rect 583520 299012 584960 299102
rect 17033 298754 17099 298757
rect 17033 298752 20148 298754
rect 17033 298696 17038 298752
rect 17094 298696 20148 298752
rect 17033 298694 20148 298696
rect 17033 298691 17099 298694
rect -960 294252 480 294492
rect 572529 292634 572595 292637
rect 568836 292632 572595 292634
rect 568836 292576 572534 292632
rect 572590 292576 572595 292632
rect 568836 292574 572595 292576
rect 572529 292571 572595 292574
rect 583520 287316 584960 287556
rect -960 280122 480 280212
rect 3601 280122 3667 280125
rect -960 280120 3667 280122
rect -960 280064 3606 280120
rect 3662 280064 3667 280120
rect -960 280062 3667 280064
rect -960 279972 480 280062
rect 3601 280059 3667 280062
rect 583520 275620 584960 275860
rect 17033 272234 17099 272237
rect 17033 272232 20148 272234
rect 17033 272176 17038 272232
rect 17094 272176 20148 272232
rect 17033 272174 20148 272176
rect 17033 272171 17099 272174
rect 572621 268970 572687 268973
rect 568836 268968 572687 268970
rect 568836 268912 572626 268968
rect 572682 268912 572687 268968
rect 568836 268910 572687 268912
rect 572621 268907 572687 268910
rect -960 265556 480 265796
rect 583520 263788 584960 264028
rect 579613 252242 579679 252245
rect 583520 252242 584960 252332
rect 579613 252240 584960 252242
rect 579613 252184 579618 252240
rect 579674 252184 584960 252240
rect 579613 252182 584960 252184
rect 579613 252179 579679 252182
rect 583520 252092 584960 252182
rect -960 251140 480 251380
rect 17033 245714 17099 245717
rect 17033 245712 20148 245714
rect 17033 245656 17038 245712
rect 17094 245656 20148 245712
rect 17033 245654 20148 245656
rect 17033 245651 17099 245654
rect 568806 244762 568866 245276
rect 571241 244762 571307 244765
rect 568806 244760 571307 244762
rect 568806 244704 571246 244760
rect 571302 244704 571307 244760
rect 568806 244702 571307 244704
rect 571241 244699 571307 244702
rect 583520 240396 584960 240636
rect -960 237010 480 237100
rect 3693 237010 3759 237013
rect -960 237008 3759 237010
rect -960 236952 3698 237008
rect 3754 236952 3759 237008
rect -960 236950 3759 236952
rect -960 236860 480 236950
rect 3693 236947 3759 236950
rect 583520 228700 584960 228940
rect -960 222444 480 222684
rect 571241 221506 571307 221509
rect 568836 221504 571307 221506
rect 568836 221448 571246 221504
rect 571302 221448 571307 221504
rect 568836 221446 571307 221448
rect 571241 221443 571307 221446
rect 17033 219058 17099 219061
rect 17033 219056 20148 219058
rect 17033 219000 17038 219056
rect 17094 219000 20148 219056
rect 17033 218998 20148 219000
rect 17033 218995 17099 218998
rect 583520 216868 584960 217108
rect -960 208028 480 208268
rect 579613 205322 579679 205325
rect 583520 205322 584960 205412
rect 579613 205320 584960 205322
rect 579613 205264 579618 205320
rect 579674 205264 584960 205320
rect 579613 205262 584960 205264
rect 579613 205259 579679 205262
rect 583520 205172 584960 205262
rect 568806 197570 568866 197812
rect 571241 197570 571307 197573
rect 568806 197568 571307 197570
rect 568806 197512 571246 197568
rect 571302 197512 571307 197568
rect 568806 197510 571307 197512
rect 571241 197507 571307 197510
rect -960 193898 480 193988
rect 3877 193898 3943 193901
rect -960 193896 3943 193898
rect -960 193840 3882 193896
rect 3938 193840 3943 193896
rect -960 193838 3943 193840
rect -960 193748 480 193838
rect 3877 193835 3943 193838
rect 583520 193476 584960 193716
rect 17033 192538 17099 192541
rect 17033 192536 20148 192538
rect 17033 192480 17038 192536
rect 17094 192480 20148 192536
rect 17033 192478 20148 192480
rect 17033 192475 17099 192478
rect 583520 181780 584960 182020
rect -960 179332 480 179572
rect 571241 174178 571307 174181
rect 568836 174176 571307 174178
rect 568836 174120 571246 174176
rect 571302 174120 571307 174176
rect 568836 174118 571307 174120
rect 571241 174115 571307 174118
rect 583520 169948 584960 170188
rect 17033 166018 17099 166021
rect 17033 166016 20148 166018
rect 17033 165960 17038 166016
rect 17094 165960 20148 166016
rect 17033 165958 20148 165960
rect 17033 165955 17099 165958
rect -960 164916 480 165156
rect 579613 158402 579679 158405
rect 583520 158402 584960 158492
rect 579613 158400 584960 158402
rect 579613 158344 579618 158400
rect 579674 158344 584960 158400
rect 579613 158342 584960 158344
rect 579613 158339 579679 158342
rect 583520 158252 584960 158342
rect -960 150786 480 150876
rect 3785 150786 3851 150789
rect -960 150784 3851 150786
rect -960 150728 3790 150784
rect 3846 150728 3851 150784
rect -960 150726 3851 150728
rect -960 150636 480 150726
rect 3785 150723 3851 150726
rect 571241 150378 571307 150381
rect 568836 150376 571307 150378
rect 568836 150320 571246 150376
rect 571302 150320 571307 150376
rect 568836 150318 571307 150320
rect 571241 150315 571307 150318
rect 583520 146556 584960 146796
rect 16757 139498 16823 139501
rect 16757 139496 20148 139498
rect 16757 139440 16762 139496
rect 16818 139440 20148 139496
rect 16757 139438 20148 139440
rect 16757 139435 16823 139438
rect -960 136220 480 136460
rect 583520 134724 584960 134964
rect 571241 126714 571307 126717
rect 568836 126712 571307 126714
rect 568836 126656 571246 126712
rect 571302 126656 571307 126712
rect 568836 126654 571307 126656
rect 571241 126651 571307 126654
rect 583520 123028 584960 123268
rect -960 121940 480 122180
rect 17033 112842 17099 112845
rect 17033 112840 20148 112842
rect 17033 112784 17038 112840
rect 17094 112784 20148 112840
rect 17033 112782 20148 112784
rect 17033 112779 17099 112782
rect 579613 111482 579679 111485
rect 583520 111482 584960 111572
rect 579613 111480 584960 111482
rect 579613 111424 579618 111480
rect 579674 111424 584960 111480
rect 579613 111422 584960 111424
rect 579613 111419 579679 111422
rect 583520 111332 584960 111422
rect -960 107674 480 107764
rect 3325 107674 3391 107677
rect -960 107672 3391 107674
rect -960 107616 3330 107672
rect 3386 107616 3391 107672
rect -960 107614 3391 107616
rect -960 107524 480 107614
rect 3325 107611 3391 107614
rect 571241 103050 571307 103053
rect 568836 103048 571307 103050
rect 568836 102992 571246 103048
rect 571302 102992 571307 103048
rect 568836 102990 571307 102992
rect 571241 102987 571307 102990
rect 583520 99636 584960 99876
rect -960 93108 480 93348
rect 583520 87804 584960 88044
rect 17033 86322 17099 86325
rect 17033 86320 20148 86322
rect 17033 86264 17038 86320
rect 17094 86264 20148 86320
rect 17033 86262 20148 86264
rect 17033 86259 17099 86262
rect 571241 79250 571307 79253
rect 568836 79248 571307 79250
rect 568836 79192 571246 79248
rect 571302 79192 571307 79248
rect 568836 79190 571307 79192
rect 571241 79187 571307 79190
rect -960 78828 480 79068
rect 583520 76108 584960 76348
rect -960 64562 480 64652
rect 3325 64562 3391 64565
rect -960 64560 3391 64562
rect -960 64504 3330 64560
rect 3386 64504 3391 64560
rect -960 64502 3391 64504
rect -960 64412 480 64502
rect 3325 64499 3391 64502
rect 580165 64562 580231 64565
rect 583520 64562 584960 64652
rect 580165 64560 584960 64562
rect 580165 64504 580170 64560
rect 580226 64504 584960 64560
rect 580165 64502 584960 64504
rect 580165 64499 580231 64502
rect 583520 64412 584960 64502
rect 16941 59802 17007 59805
rect 16941 59800 20148 59802
rect 16941 59744 16946 59800
rect 17002 59744 20148 59800
rect 16941 59742 20148 59744
rect 16941 59739 17007 59742
rect 568622 55314 568682 55556
rect 571241 55314 571307 55317
rect 568622 55312 571307 55314
rect 568622 55256 571246 55312
rect 571302 55256 571307 55312
rect 568622 55254 571307 55256
rect 571241 55251 571307 55254
rect 583520 52716 584960 52956
rect -960 49996 480 50236
rect 583520 40884 584960 41124
rect -960 35716 480 35956
rect 17033 33282 17099 33285
rect 17033 33280 20148 33282
rect 17033 33224 17038 33280
rect 17094 33224 20148 33280
rect 17033 33222 20148 33224
rect 17033 33219 17099 33222
rect 573357 31922 573423 31925
rect 568836 31920 573423 31922
rect 568836 31864 573362 31920
rect 573418 31864 573423 31920
rect 568836 31862 573423 31864
rect 573357 31859 573423 31862
rect 583520 29188 584960 29428
rect -960 21450 480 21540
rect 3141 21450 3207 21453
rect -960 21448 3207 21450
rect -960 21392 3146 21448
rect 3202 21392 3207 21448
rect -960 21390 3207 21392
rect -960 21300 480 21390
rect 3141 21387 3207 21390
rect 114461 19954 114527 19957
rect 561622 19954 561628 19956
rect 114461 19952 561628 19954
rect 114461 19896 114466 19952
rect 114522 19896 561628 19952
rect 114461 19894 561628 19896
rect 114461 19891 114527 19894
rect 561622 19892 561628 19894
rect 561692 19892 561698 19956
rect 31661 17642 31727 17645
rect 490741 17642 490807 17645
rect 31661 17640 490807 17642
rect 31661 17584 31666 17640
rect 31722 17584 490746 17640
rect 490802 17584 490807 17640
rect 31661 17582 490807 17584
rect 31661 17579 31727 17582
rect 490741 17579 490807 17582
rect 579797 17642 579863 17645
rect 583520 17642 584960 17732
rect 579797 17640 584960 17642
rect 579797 17584 579802 17640
rect 579858 17584 584960 17640
rect 579797 17582 584960 17584
rect 579797 17579 579863 17582
rect 64781 17506 64847 17509
rect 527357 17506 527423 17509
rect 64781 17504 527423 17506
rect 64781 17448 64786 17504
rect 64842 17448 527362 17504
rect 527418 17448 527423 17504
rect 583520 17492 584960 17582
rect 64781 17446 527423 17448
rect 64781 17443 64847 17446
rect 527357 17443 527423 17446
rect 19149 17370 19215 17373
rect 481633 17370 481699 17373
rect 19149 17368 481699 17370
rect 19149 17312 19154 17368
rect 19210 17312 481638 17368
rect 481694 17312 481699 17368
rect 19149 17310 481699 17312
rect 19149 17307 19215 17310
rect 481633 17307 481699 17310
rect 42701 17234 42767 17237
rect 509233 17234 509299 17237
rect 42701 17232 509299 17234
rect 42701 17176 42706 17232
rect 42762 17176 509238 17232
rect 509294 17176 509299 17232
rect 42701 17174 509299 17176
rect 42701 17171 42767 17174
rect 509233 17171 509299 17174
rect -960 7020 480 7260
rect 583520 5796 584960 6036
rect 106365 4042 106431 4045
rect 563278 4042 563284 4044
rect 106365 4040 563284 4042
rect 106365 3984 106370 4040
rect 106426 3984 563284 4040
rect 106365 3982 563284 3984
rect 106365 3979 106431 3982
rect 563278 3980 563284 3982
rect 563348 3980 563354 4044
rect 23054 3844 23060 3908
rect 23124 3906 23130 3908
rect 44541 3906 44607 3909
rect 23124 3904 44607 3906
rect 23124 3848 44546 3904
rect 44602 3848 44607 3904
rect 23124 3846 44607 3848
rect 23124 3844 23130 3846
rect 44541 3843 44607 3846
rect 109953 3906 110019 3909
rect 571374 3906 571380 3908
rect 109953 3904 571380 3906
rect 109953 3848 109958 3904
rect 110014 3848 571380 3904
rect 109953 3846 571380 3848
rect 109953 3843 110019 3846
rect 571374 3844 571380 3846
rect 571444 3844 571450 3908
rect 22870 3708 22876 3772
rect 22940 3770 22946 3772
rect 70669 3770 70735 3773
rect 22940 3768 70735 3770
rect 22940 3712 70674 3768
rect 70730 3712 70735 3768
rect 22940 3710 70735 3712
rect 22940 3708 22946 3710
rect 70669 3707 70735 3710
rect 99281 3770 99347 3773
rect 563094 3770 563100 3772
rect 99281 3768 563100 3770
rect 99281 3712 99286 3768
rect 99342 3712 563100 3768
rect 99281 3710 563100 3712
rect 99281 3707 99347 3710
rect 563094 3708 563100 3710
rect 563164 3708 563170 3772
rect 23606 3572 23612 3636
rect 23676 3634 23682 3636
rect 72969 3634 73035 3637
rect 23676 3632 73035 3634
rect 23676 3576 72974 3632
rect 73030 3576 73035 3632
rect 23676 3574 73035 3576
rect 23676 3572 23682 3574
rect 72969 3571 73035 3574
rect 95693 3634 95759 3637
rect 571558 3634 571564 3636
rect 95693 3632 571564 3634
rect 95693 3576 95698 3632
rect 95754 3576 571564 3632
rect 95693 3574 571564 3576
rect 95693 3571 95759 3574
rect 571558 3572 571564 3574
rect 571628 3572 571634 3636
rect 21633 3498 21699 3501
rect 74257 3498 74323 3501
rect 21633 3496 74323 3498
rect 21633 3440 21638 3496
rect 21694 3440 74262 3496
rect 74318 3440 74323 3496
rect 21633 3438 74323 3440
rect 21633 3435 21699 3438
rect 74257 3435 74323 3438
rect 81433 3498 81499 3501
rect 571742 3498 571748 3500
rect 81433 3496 571748 3498
rect 81433 3440 81438 3496
rect 81494 3440 571748 3496
rect 81433 3438 571748 3440
rect 81433 3435 81499 3438
rect 571742 3436 571748 3438
rect 571812 3436 571818 3500
rect 23238 3300 23244 3364
rect 23308 3362 23314 3364
rect 37365 3362 37431 3365
rect 23308 3360 37431 3362
rect 23308 3304 37370 3360
rect 37426 3304 37431 3360
rect 23308 3302 37431 3304
rect 23308 3300 23314 3302
rect 37365 3299 37431 3302
rect 38561 3362 38627 3365
rect 571517 3362 571583 3365
rect 38561 3360 571583 3362
rect 38561 3304 38566 3360
rect 38622 3304 571522 3360
rect 571578 3304 571583 3360
rect 38561 3302 571583 3304
rect 38561 3299 38627 3302
rect 571517 3299 571583 3302
<< via3 >>
rect 23244 686292 23308 686356
rect 23060 686156 23124 686220
rect 561628 686156 561692 686220
rect 23612 686020 23676 686084
rect 337332 686020 337396 686084
rect 563284 686020 563348 686084
rect 22876 685884 22940 685948
rect 563100 685884 563164 685948
rect 284892 683708 284956 683772
rect 323164 683436 323228 683500
rect 311756 683360 311820 683364
rect 311756 683304 311806 683360
rect 311806 683304 311820 683360
rect 311756 683300 311820 683304
rect 284892 682756 284956 682820
rect 311756 682620 311820 682684
rect 323164 682484 323228 682548
rect 337332 682348 337396 682412
rect 571380 672012 571444 672076
rect 571564 648348 571628 648412
rect 571748 624548 571812 624612
rect 561628 19892 561692 19956
rect 563284 3980 563348 4044
rect 23060 3844 23124 3908
rect 571380 3844 571444 3908
rect 22876 3708 22940 3772
rect 563100 3708 563164 3772
rect 23612 3572 23676 3636
rect 571564 3572 571628 3636
rect 571748 3436 571812 3500
rect 23244 3300 23308 3364
<< metal4 >>
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 668454 -2336 705222
rect -2936 668218 -2754 668454
rect -2518 668218 -2336 668454
rect -2936 668134 -2336 668218
rect -2936 667898 -2754 668134
rect -2518 667898 -2336 668134
rect -2936 632454 -2336 667898
rect -2936 632218 -2754 632454
rect -2518 632218 -2336 632454
rect -2936 632134 -2336 632218
rect -2936 631898 -2754 632134
rect -2518 631898 -2336 632134
rect -2936 596454 -2336 631898
rect -2936 596218 -2754 596454
rect -2518 596218 -2336 596454
rect -2936 596134 -2336 596218
rect -2936 595898 -2754 596134
rect -2518 595898 -2336 596134
rect -2936 560454 -2336 595898
rect -2936 560218 -2754 560454
rect -2518 560218 -2336 560454
rect -2936 560134 -2336 560218
rect -2936 559898 -2754 560134
rect -2518 559898 -2336 560134
rect -2936 524454 -2336 559898
rect -2936 524218 -2754 524454
rect -2518 524218 -2336 524454
rect -2936 524134 -2336 524218
rect -2936 523898 -2754 524134
rect -2518 523898 -2336 524134
rect -2936 488454 -2336 523898
rect -2936 488218 -2754 488454
rect -2518 488218 -2336 488454
rect -2936 488134 -2336 488218
rect -2936 487898 -2754 488134
rect -2518 487898 -2336 488134
rect -2936 452454 -2336 487898
rect -2936 452218 -2754 452454
rect -2518 452218 -2336 452454
rect -2936 452134 -2336 452218
rect -2936 451898 -2754 452134
rect -2518 451898 -2336 452134
rect -2936 416454 -2336 451898
rect -2936 416218 -2754 416454
rect -2518 416218 -2336 416454
rect -2936 416134 -2336 416218
rect -2936 415898 -2754 416134
rect -2518 415898 -2336 416134
rect -2936 380454 -2336 415898
rect -2936 380218 -2754 380454
rect -2518 380218 -2336 380454
rect -2936 380134 -2336 380218
rect -2936 379898 -2754 380134
rect -2518 379898 -2336 380134
rect -2936 344454 -2336 379898
rect -2936 344218 -2754 344454
rect -2518 344218 -2336 344454
rect -2936 344134 -2336 344218
rect -2936 343898 -2754 344134
rect -2518 343898 -2336 344134
rect -2936 308454 -2336 343898
rect -2936 308218 -2754 308454
rect -2518 308218 -2336 308454
rect -2936 308134 -2336 308218
rect -2936 307898 -2754 308134
rect -2518 307898 -2336 308134
rect -2936 272454 -2336 307898
rect -2936 272218 -2754 272454
rect -2518 272218 -2336 272454
rect -2936 272134 -2336 272218
rect -2936 271898 -2754 272134
rect -2518 271898 -2336 272134
rect -2936 236454 -2336 271898
rect -2936 236218 -2754 236454
rect -2518 236218 -2336 236454
rect -2936 236134 -2336 236218
rect -2936 235898 -2754 236134
rect -2518 235898 -2336 236134
rect -2936 200454 -2336 235898
rect -2936 200218 -2754 200454
rect -2518 200218 -2336 200454
rect -2936 200134 -2336 200218
rect -2936 199898 -2754 200134
rect -2518 199898 -2336 200134
rect -2936 164454 -2336 199898
rect -2936 164218 -2754 164454
rect -2518 164218 -2336 164454
rect -2936 164134 -2336 164218
rect -2936 163898 -2754 164134
rect -2518 163898 -2336 164134
rect -2936 128454 -2336 163898
rect -2936 128218 -2754 128454
rect -2518 128218 -2336 128454
rect -2936 128134 -2336 128218
rect -2936 127898 -2754 128134
rect -2518 127898 -2336 128134
rect -2936 92454 -2336 127898
rect -2936 92218 -2754 92454
rect -2518 92218 -2336 92454
rect -2936 92134 -2336 92218
rect -2936 91898 -2754 92134
rect -2518 91898 -2336 92134
rect -2936 56454 -2336 91898
rect -2936 56218 -2754 56454
rect -2518 56218 -2336 56454
rect -2936 56134 -2336 56218
rect -2936 55898 -2754 56134
rect -2518 55898 -2336 56134
rect -2936 20454 -2336 55898
rect -2936 20218 -2754 20454
rect -2518 20218 -2336 20454
rect -2936 20134 -2336 20218
rect -2936 19898 -2754 20134
rect -2518 19898 -2336 20134
rect -2936 -1286 -2336 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect 37072 704838 37672 705800
rect 37072 704602 37254 704838
rect 37490 704602 37672 704838
rect 37072 704518 37672 704602
rect 37072 704282 37254 704518
rect 37490 704282 37672 704518
rect 37072 686454 37672 704282
rect 23243 686356 23309 686357
rect 23243 686292 23244 686356
rect 23308 686292 23309 686356
rect 23243 686291 23309 686292
rect -1996 686134 -1396 686218
rect 23059 686220 23125 686221
rect 23059 686156 23060 686220
rect 23124 686156 23125 686220
rect 23059 686155 23125 686156
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect 22875 685948 22941 685949
rect 22875 685884 22876 685948
rect 22940 685884 22941 685948
rect 22875 685883 22941 685884
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect 22878 3773 22938 685883
rect 23062 3909 23122 686155
rect 23059 3908 23125 3909
rect 23059 3844 23060 3908
rect 23124 3844 23125 3908
rect 23059 3843 23125 3844
rect 22875 3772 22941 3773
rect 22875 3708 22876 3772
rect 22940 3708 22941 3772
rect 22875 3707 22941 3708
rect 23246 3365 23306 686291
rect 37072 686218 37254 686454
rect 37490 686218 37672 686454
rect 37072 686134 37672 686218
rect 23611 686084 23677 686085
rect 23611 686020 23612 686084
rect 23676 686020 23677 686084
rect 23611 686019 23677 686020
rect 23614 3637 23674 686019
rect 37072 685898 37254 686134
rect 37490 685898 37672 686134
rect 23611 3636 23677 3637
rect 23611 3572 23612 3636
rect 23676 3572 23677 3636
rect 23611 3571 23677 3572
rect 23243 3364 23309 3365
rect 23243 3300 23244 3364
rect 23308 3300 23309 3364
rect 23243 3299 23309 3300
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 37072 2454 37672 685898
rect 37072 2218 37254 2454
rect 37490 2218 37672 2454
rect 37072 2134 37672 2218
rect 37072 1898 37254 2134
rect 37490 1898 37672 2134
rect 37072 -346 37672 1898
rect 37072 -582 37254 -346
rect 37490 -582 37672 -346
rect 37072 -666 37672 -582
rect 37072 -902 37254 -666
rect 37490 -902 37672 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 37072 -1864 37672 -902
rect 110943 705778 111543 705800
rect 110943 705542 111125 705778
rect 111361 705542 111543 705778
rect 110943 705458 111543 705542
rect 110943 705222 111125 705458
rect 111361 705222 111543 705458
rect 110943 -1286 111543 705222
rect 110943 -1522 111125 -1286
rect 111361 -1522 111543 -1286
rect 110943 -1606 111543 -1522
rect 110943 -1842 111125 -1606
rect 111361 -1842 111543 -1606
rect 110943 -1864 111543 -1842
rect 184814 704838 185414 705800
rect 184814 704602 184996 704838
rect 185232 704602 185414 704838
rect 184814 704518 185414 704602
rect 184814 704282 184996 704518
rect 185232 704282 185414 704518
rect 184814 686454 185414 704282
rect 184814 686218 184996 686454
rect 185232 686218 185414 686454
rect 184814 686134 185414 686218
rect 184814 685898 184996 686134
rect 185232 685898 185414 686134
rect 184814 2454 185414 685898
rect 184814 2218 184996 2454
rect 185232 2218 185414 2454
rect 184814 2134 185414 2218
rect 184814 1898 184996 2134
rect 185232 1898 185414 2134
rect 184814 -346 185414 1898
rect 184814 -582 184996 -346
rect 185232 -582 185414 -346
rect 184814 -666 185414 -582
rect 184814 -902 184996 -666
rect 185232 -902 185414 -666
rect 184814 -1864 185414 -902
rect 258685 705778 259285 705800
rect 258685 705542 258867 705778
rect 259103 705542 259285 705778
rect 258685 705458 259285 705542
rect 258685 705222 258867 705458
rect 259103 705222 259285 705458
rect 258685 -1286 259285 705222
rect 332556 704838 333156 705800
rect 332556 704602 332738 704838
rect 332974 704602 333156 704838
rect 332556 704518 333156 704602
rect 332556 704282 332738 704518
rect 332974 704282 333156 704518
rect 332556 686454 333156 704282
rect 332556 686218 332738 686454
rect 332974 686218 333156 686454
rect 332556 686134 333156 686218
rect 332556 685898 332738 686134
rect 332974 685898 333156 686134
rect 406427 705778 407027 705800
rect 406427 705542 406609 705778
rect 406845 705542 407027 705778
rect 406427 705458 407027 705542
rect 406427 705222 406609 705458
rect 406845 705222 407027 705458
rect 337331 686084 337397 686085
rect 337331 686020 337332 686084
rect 337396 686020 337397 686084
rect 337331 686019 337397 686020
rect 284891 683772 284957 683773
rect 284891 683708 284892 683772
rect 284956 683708 284957 683772
rect 284891 683707 284957 683708
rect 284894 682821 284954 683707
rect 323163 683500 323229 683501
rect 323163 683436 323164 683500
rect 323228 683436 323229 683500
rect 323163 683435 323229 683436
rect 311755 683364 311821 683365
rect 311755 683300 311756 683364
rect 311820 683300 311821 683364
rect 311755 683299 311821 683300
rect 284891 682820 284957 682821
rect 284891 682756 284892 682820
rect 284956 682756 284957 682820
rect 284891 682755 284957 682756
rect 311758 682685 311818 683299
rect 311755 682684 311821 682685
rect 311755 682620 311756 682684
rect 311820 682620 311821 682684
rect 311755 682619 311821 682620
rect 323166 682549 323226 683435
rect 323163 682548 323229 682549
rect 323163 682484 323164 682548
rect 323228 682484 323229 682548
rect 323163 682483 323229 682484
rect 258685 -1522 258867 -1286
rect 259103 -1522 259285 -1286
rect 258685 -1606 259285 -1522
rect 258685 -1842 258867 -1606
rect 259103 -1842 259285 -1606
rect 258685 -1864 259285 -1842
rect 332556 2454 333156 685898
rect 337334 682413 337394 686019
rect 337331 682412 337397 682413
rect 337331 682348 337332 682412
rect 337396 682348 337397 682412
rect 337331 682347 337397 682348
rect 332556 2218 332738 2454
rect 332974 2218 333156 2454
rect 332556 2134 333156 2218
rect 332556 1898 332738 2134
rect 332974 1898 333156 2134
rect 332556 -346 333156 1898
rect 332556 -582 332738 -346
rect 332974 -582 333156 -346
rect 332556 -666 333156 -582
rect 332556 -902 332738 -666
rect 332974 -902 333156 -666
rect 332556 -1864 333156 -902
rect 406427 -1286 407027 705222
rect 406427 -1522 406609 -1286
rect 406845 -1522 407027 -1286
rect 406427 -1606 407027 -1522
rect 406427 -1842 406609 -1606
rect 406845 -1842 407027 -1606
rect 406427 -1864 407027 -1842
rect 480298 704838 480898 705800
rect 480298 704602 480480 704838
rect 480716 704602 480898 704838
rect 480298 704518 480898 704602
rect 480298 704282 480480 704518
rect 480716 704282 480898 704518
rect 480298 686454 480898 704282
rect 480298 686218 480480 686454
rect 480716 686218 480898 686454
rect 480298 686134 480898 686218
rect 480298 685898 480480 686134
rect 480716 685898 480898 686134
rect 480298 2454 480898 685898
rect 480298 2218 480480 2454
rect 480716 2218 480898 2454
rect 480298 2134 480898 2218
rect 480298 1898 480480 2134
rect 480716 1898 480898 2134
rect 480298 -346 480898 1898
rect 480298 -582 480480 -346
rect 480716 -582 480898 -346
rect 480298 -666 480898 -582
rect 480298 -902 480480 -666
rect 480716 -902 480898 -666
rect 480298 -1864 480898 -902
rect 554169 705778 554769 705800
rect 554169 705542 554351 705778
rect 554587 705542 554769 705778
rect 554169 705458 554769 705542
rect 554169 705222 554351 705458
rect 554587 705222 554769 705458
rect 554169 -1286 554769 705222
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 561627 686220 561693 686221
rect 561627 686156 561628 686220
rect 561692 686156 561693 686220
rect 561627 686155 561693 686156
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 561630 19957 561690 686155
rect 585320 686134 585920 686218
rect 563283 686084 563349 686085
rect 563283 686020 563284 686084
rect 563348 686020 563349 686084
rect 563283 686019 563349 686020
rect 563099 685948 563165 685949
rect 563099 685884 563100 685948
rect 563164 685884 563165 685948
rect 563099 685883 563165 685884
rect 561627 19956 561693 19957
rect 561627 19892 561628 19956
rect 561692 19892 561693 19956
rect 561627 19891 561693 19892
rect 563102 3773 563162 685883
rect 563286 4045 563346 686019
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 571379 672076 571445 672077
rect 571379 672012 571380 672076
rect 571444 672012 571445 672076
rect 571379 672011 571445 672012
rect 563283 4044 563349 4045
rect 563283 3980 563284 4044
rect 563348 3980 563349 4044
rect 563283 3979 563349 3980
rect 571382 3909 571442 672011
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 571563 648412 571629 648413
rect 571563 648348 571564 648412
rect 571628 648348 571629 648412
rect 571563 648347 571629 648348
rect 571379 3908 571445 3909
rect 571379 3844 571380 3908
rect 571444 3844 571445 3908
rect 571379 3843 571445 3844
rect 563099 3772 563165 3773
rect 563099 3708 563100 3772
rect 563164 3708 563165 3772
rect 563099 3707 563165 3708
rect 571566 3637 571626 648347
rect 571747 624612 571813 624613
rect 571747 624548 571748 624612
rect 571812 624548 571813 624612
rect 571747 624547 571813 624548
rect 571563 3636 571629 3637
rect 571563 3572 571564 3636
rect 571628 3572 571629 3636
rect 571563 3571 571629 3572
rect 571750 3501 571810 624547
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 571747 3500 571813 3501
rect 571747 3436 571748 3500
rect 571812 3436 571813 3500
rect 571747 3435 571813 3436
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 668454 586860 705222
rect 586260 668218 586442 668454
rect 586678 668218 586860 668454
rect 586260 668134 586860 668218
rect 586260 667898 586442 668134
rect 586678 667898 586860 668134
rect 586260 632454 586860 667898
rect 586260 632218 586442 632454
rect 586678 632218 586860 632454
rect 586260 632134 586860 632218
rect 586260 631898 586442 632134
rect 586678 631898 586860 632134
rect 586260 596454 586860 631898
rect 586260 596218 586442 596454
rect 586678 596218 586860 596454
rect 586260 596134 586860 596218
rect 586260 595898 586442 596134
rect 586678 595898 586860 596134
rect 586260 560454 586860 595898
rect 586260 560218 586442 560454
rect 586678 560218 586860 560454
rect 586260 560134 586860 560218
rect 586260 559898 586442 560134
rect 586678 559898 586860 560134
rect 586260 524454 586860 559898
rect 586260 524218 586442 524454
rect 586678 524218 586860 524454
rect 586260 524134 586860 524218
rect 586260 523898 586442 524134
rect 586678 523898 586860 524134
rect 586260 488454 586860 523898
rect 586260 488218 586442 488454
rect 586678 488218 586860 488454
rect 586260 488134 586860 488218
rect 586260 487898 586442 488134
rect 586678 487898 586860 488134
rect 586260 452454 586860 487898
rect 586260 452218 586442 452454
rect 586678 452218 586860 452454
rect 586260 452134 586860 452218
rect 586260 451898 586442 452134
rect 586678 451898 586860 452134
rect 586260 416454 586860 451898
rect 586260 416218 586442 416454
rect 586678 416218 586860 416454
rect 586260 416134 586860 416218
rect 586260 415898 586442 416134
rect 586678 415898 586860 416134
rect 586260 380454 586860 415898
rect 586260 380218 586442 380454
rect 586678 380218 586860 380454
rect 586260 380134 586860 380218
rect 586260 379898 586442 380134
rect 586678 379898 586860 380134
rect 586260 344454 586860 379898
rect 586260 344218 586442 344454
rect 586678 344218 586860 344454
rect 586260 344134 586860 344218
rect 586260 343898 586442 344134
rect 586678 343898 586860 344134
rect 586260 308454 586860 343898
rect 586260 308218 586442 308454
rect 586678 308218 586860 308454
rect 586260 308134 586860 308218
rect 586260 307898 586442 308134
rect 586678 307898 586860 308134
rect 586260 272454 586860 307898
rect 586260 272218 586442 272454
rect 586678 272218 586860 272454
rect 586260 272134 586860 272218
rect 586260 271898 586442 272134
rect 586678 271898 586860 272134
rect 586260 236454 586860 271898
rect 586260 236218 586442 236454
rect 586678 236218 586860 236454
rect 586260 236134 586860 236218
rect 586260 235898 586442 236134
rect 586678 235898 586860 236134
rect 586260 200454 586860 235898
rect 586260 200218 586442 200454
rect 586678 200218 586860 200454
rect 586260 200134 586860 200218
rect 586260 199898 586442 200134
rect 586678 199898 586860 200134
rect 586260 164454 586860 199898
rect 586260 164218 586442 164454
rect 586678 164218 586860 164454
rect 586260 164134 586860 164218
rect 586260 163898 586442 164134
rect 586678 163898 586860 164134
rect 586260 128454 586860 163898
rect 586260 128218 586442 128454
rect 586678 128218 586860 128454
rect 586260 128134 586860 128218
rect 586260 127898 586442 128134
rect 586678 127898 586860 128134
rect 586260 92454 586860 127898
rect 586260 92218 586442 92454
rect 586678 92218 586860 92454
rect 586260 92134 586860 92218
rect 586260 91898 586442 92134
rect 586678 91898 586860 92134
rect 586260 56454 586860 91898
rect 586260 56218 586442 56454
rect 586678 56218 586860 56454
rect 586260 56134 586860 56218
rect 586260 55898 586442 56134
rect 586678 55898 586860 56134
rect 586260 20454 586860 55898
rect 586260 20218 586442 20454
rect 586678 20218 586860 20454
rect 586260 20134 586860 20218
rect 586260 19898 586442 20134
rect 586678 19898 586860 20134
rect 554169 -1522 554351 -1286
rect 554587 -1522 554769 -1286
rect 554169 -1606 554769 -1522
rect 554169 -1842 554351 -1606
rect 554587 -1842 554769 -1606
rect 554169 -1864 554769 -1842
rect 586260 -1286 586860 19898
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
<< via4 >>
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 668218 -2518 668454
rect -2754 667898 -2518 668134
rect -2754 632218 -2518 632454
rect -2754 631898 -2518 632134
rect -2754 596218 -2518 596454
rect -2754 595898 -2518 596134
rect -2754 560218 -2518 560454
rect -2754 559898 -2518 560134
rect -2754 524218 -2518 524454
rect -2754 523898 -2518 524134
rect -2754 488218 -2518 488454
rect -2754 487898 -2518 488134
rect -2754 452218 -2518 452454
rect -2754 451898 -2518 452134
rect -2754 416218 -2518 416454
rect -2754 415898 -2518 416134
rect -2754 380218 -2518 380454
rect -2754 379898 -2518 380134
rect -2754 344218 -2518 344454
rect -2754 343898 -2518 344134
rect -2754 308218 -2518 308454
rect -2754 307898 -2518 308134
rect -2754 272218 -2518 272454
rect -2754 271898 -2518 272134
rect -2754 236218 -2518 236454
rect -2754 235898 -2518 236134
rect -2754 200218 -2518 200454
rect -2754 199898 -2518 200134
rect -2754 164218 -2518 164454
rect -2754 163898 -2518 164134
rect -2754 128218 -2518 128454
rect -2754 127898 -2518 128134
rect -2754 92218 -2518 92454
rect -2754 91898 -2518 92134
rect -2754 56218 -2518 56454
rect -2754 55898 -2518 56134
rect -2754 20218 -2518 20454
rect -2754 19898 -2518 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect 37254 704602 37490 704838
rect 37254 704282 37490 704518
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect 37254 686218 37490 686454
rect 37254 685898 37490 686134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 37254 2218 37490 2454
rect 37254 1898 37490 2134
rect 37254 -582 37490 -346
rect 37254 -902 37490 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 111125 705542 111361 705778
rect 111125 705222 111361 705458
rect 111125 -1522 111361 -1286
rect 111125 -1842 111361 -1606
rect 184996 704602 185232 704838
rect 184996 704282 185232 704518
rect 184996 686218 185232 686454
rect 184996 685898 185232 686134
rect 184996 2218 185232 2454
rect 184996 1898 185232 2134
rect 184996 -582 185232 -346
rect 184996 -902 185232 -666
rect 258867 705542 259103 705778
rect 258867 705222 259103 705458
rect 332738 704602 332974 704838
rect 332738 704282 332974 704518
rect 332738 686218 332974 686454
rect 332738 685898 332974 686134
rect 406609 705542 406845 705778
rect 406609 705222 406845 705458
rect 258867 -1522 259103 -1286
rect 258867 -1842 259103 -1606
rect 332738 2218 332974 2454
rect 332738 1898 332974 2134
rect 332738 -582 332974 -346
rect 332738 -902 332974 -666
rect 406609 -1522 406845 -1286
rect 406609 -1842 406845 -1606
rect 480480 704602 480716 704838
rect 480480 704282 480716 704518
rect 480480 686218 480716 686454
rect 480480 685898 480716 686134
rect 480480 2218 480716 2454
rect 480480 1898 480716 2134
rect 480480 -582 480716 -346
rect 480480 -902 480716 -666
rect 554351 705542 554587 705778
rect 554351 705222 554587 705458
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 668218 586678 668454
rect 586442 667898 586678 668134
rect 586442 632218 586678 632454
rect 586442 631898 586678 632134
rect 586442 596218 586678 596454
rect 586442 595898 586678 596134
rect 586442 560218 586678 560454
rect 586442 559898 586678 560134
rect 586442 524218 586678 524454
rect 586442 523898 586678 524134
rect 586442 488218 586678 488454
rect 586442 487898 586678 488134
rect 586442 452218 586678 452454
rect 586442 451898 586678 452134
rect 586442 416218 586678 416454
rect 586442 415898 586678 416134
rect 586442 380218 586678 380454
rect 586442 379898 586678 380134
rect 586442 344218 586678 344454
rect 586442 343898 586678 344134
rect 586442 308218 586678 308454
rect 586442 307898 586678 308134
rect 586442 272218 586678 272454
rect 586442 271898 586678 272134
rect 586442 236218 586678 236454
rect 586442 235898 586678 236134
rect 586442 200218 586678 200454
rect 586442 199898 586678 200134
rect 586442 164218 586678 164454
rect 586442 163898 586678 164134
rect 586442 128218 586678 128454
rect 586442 127898 586678 128134
rect 586442 92218 586678 92454
rect 586442 91898 586678 92134
rect 586442 56218 586678 56454
rect 586442 55898 586678 56134
rect 586442 20218 586678 20454
rect 586442 19898 586678 20134
rect 554351 -1522 554587 -1286
rect 554351 -1842 554587 -1606
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
<< metal5 >>
rect -2936 705800 -2336 705802
rect 110943 705800 111543 705802
rect 258685 705800 259285 705802
rect 406427 705800 407027 705802
rect 554169 705800 554769 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 111125 705778
rect 111361 705542 258867 705778
rect 259103 705542 406609 705778
rect 406845 705542 554351 705778
rect 554587 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 111125 705458
rect 111361 705222 258867 705458
rect 259103 705222 406609 705458
rect 406845 705222 554351 705458
rect 554587 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 110943 705198 111543 705200
rect 258685 705198 259285 705200
rect 406427 705198 407027 705200
rect 554169 705198 554769 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 37072 704860 37672 704862
rect 184814 704860 185414 704862
rect 332556 704860 333156 704862
rect 480298 704860 480898 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 37254 704838
rect 37490 704602 184996 704838
rect 185232 704602 332738 704838
rect 332974 704602 480480 704838
rect 480716 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 37254 704518
rect 37490 704282 184996 704518
rect 185232 704282 332738 704518
rect 332974 704282 480480 704518
rect 480716 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 37072 704258 37672 704260
rect 184814 704258 185414 704260
rect 332556 704258 333156 704260
rect 480298 704258 480898 704260
rect 585320 704258 585920 704260
rect -1996 686476 -1396 686478
rect 37072 686476 37672 686478
rect 184814 686476 185414 686478
rect 332556 686476 333156 686478
rect 480298 686476 480898 686478
rect 585320 686476 585920 686478
rect -2936 686454 586860 686476
rect -2936 686218 -1814 686454
rect -1578 686218 37254 686454
rect 37490 686218 184996 686454
rect 185232 686218 332738 686454
rect 332974 686218 480480 686454
rect 480716 686218 585502 686454
rect 585738 686218 586860 686454
rect -2936 686134 586860 686218
rect -2936 685898 -1814 686134
rect -1578 685898 37254 686134
rect 37490 685898 184996 686134
rect 185232 685898 332738 686134
rect 332974 685898 480480 686134
rect 480716 685898 585502 686134
rect 585738 685898 586860 686134
rect -2936 685876 586860 685898
rect -1996 685874 -1396 685876
rect 37072 685874 37672 685876
rect 184814 685874 185414 685876
rect 332556 685874 333156 685876
rect 480298 685874 480898 685876
rect 585320 685874 585920 685876
rect -2936 668476 -2336 668478
rect 586260 668476 586860 668478
rect -2936 668454 20000 668476
rect -2936 668218 -2754 668454
rect -2518 668218 20000 668454
rect -2936 668134 20000 668218
rect -2936 667898 -2754 668134
rect -2518 667898 20000 668134
rect -2936 667876 20000 667898
rect 569000 668454 586860 668476
rect 569000 668218 586442 668454
rect 586678 668218 586860 668454
rect 569000 668134 586860 668218
rect 569000 667898 586442 668134
rect 586678 667898 586860 668134
rect 569000 667876 586860 667898
rect -2936 667874 -2336 667876
rect 586260 667874 586860 667876
rect -1996 650476 -1396 650478
rect 585320 650476 585920 650478
rect -2936 650454 20000 650476
rect -2936 650218 -1814 650454
rect -1578 650218 20000 650454
rect -2936 650134 20000 650218
rect -2936 649898 -1814 650134
rect -1578 649898 20000 650134
rect -2936 649876 20000 649898
rect 569000 650454 586860 650476
rect 569000 650218 585502 650454
rect 585738 650218 586860 650454
rect 569000 650134 586860 650218
rect 569000 649898 585502 650134
rect 585738 649898 586860 650134
rect 569000 649876 586860 649898
rect -1996 649874 -1396 649876
rect 585320 649874 585920 649876
rect -2936 632476 -2336 632478
rect 586260 632476 586860 632478
rect -2936 632454 20000 632476
rect -2936 632218 -2754 632454
rect -2518 632218 20000 632454
rect -2936 632134 20000 632218
rect -2936 631898 -2754 632134
rect -2518 631898 20000 632134
rect -2936 631876 20000 631898
rect 569000 632454 586860 632476
rect 569000 632218 586442 632454
rect 586678 632218 586860 632454
rect 569000 632134 586860 632218
rect 569000 631898 586442 632134
rect 586678 631898 586860 632134
rect 569000 631876 586860 631898
rect -2936 631874 -2336 631876
rect 586260 631874 586860 631876
rect -1996 614476 -1396 614478
rect 585320 614476 585920 614478
rect -2936 614454 20000 614476
rect -2936 614218 -1814 614454
rect -1578 614218 20000 614454
rect -2936 614134 20000 614218
rect -2936 613898 -1814 614134
rect -1578 613898 20000 614134
rect -2936 613876 20000 613898
rect 569000 614454 586860 614476
rect 569000 614218 585502 614454
rect 585738 614218 586860 614454
rect 569000 614134 586860 614218
rect 569000 613898 585502 614134
rect 585738 613898 586860 614134
rect 569000 613876 586860 613898
rect -1996 613874 -1396 613876
rect 585320 613874 585920 613876
rect -2936 596476 -2336 596478
rect 586260 596476 586860 596478
rect -2936 596454 20000 596476
rect -2936 596218 -2754 596454
rect -2518 596218 20000 596454
rect -2936 596134 20000 596218
rect -2936 595898 -2754 596134
rect -2518 595898 20000 596134
rect -2936 595876 20000 595898
rect 569000 596454 586860 596476
rect 569000 596218 586442 596454
rect 586678 596218 586860 596454
rect 569000 596134 586860 596218
rect 569000 595898 586442 596134
rect 586678 595898 586860 596134
rect 569000 595876 586860 595898
rect -2936 595874 -2336 595876
rect 586260 595874 586860 595876
rect -1996 578476 -1396 578478
rect 585320 578476 585920 578478
rect -2936 578454 20000 578476
rect -2936 578218 -1814 578454
rect -1578 578218 20000 578454
rect -2936 578134 20000 578218
rect -2936 577898 -1814 578134
rect -1578 577898 20000 578134
rect -2936 577876 20000 577898
rect 569000 578454 586860 578476
rect 569000 578218 585502 578454
rect 585738 578218 586860 578454
rect 569000 578134 586860 578218
rect 569000 577898 585502 578134
rect 585738 577898 586860 578134
rect 569000 577876 586860 577898
rect -1996 577874 -1396 577876
rect 585320 577874 585920 577876
rect -2936 560476 -2336 560478
rect 586260 560476 586860 560478
rect -2936 560454 20000 560476
rect -2936 560218 -2754 560454
rect -2518 560218 20000 560454
rect -2936 560134 20000 560218
rect -2936 559898 -2754 560134
rect -2518 559898 20000 560134
rect -2936 559876 20000 559898
rect 569000 560454 586860 560476
rect 569000 560218 586442 560454
rect 586678 560218 586860 560454
rect 569000 560134 586860 560218
rect 569000 559898 586442 560134
rect 586678 559898 586860 560134
rect 569000 559876 586860 559898
rect -2936 559874 -2336 559876
rect 586260 559874 586860 559876
rect -1996 542476 -1396 542478
rect 585320 542476 585920 542478
rect -2936 542454 20000 542476
rect -2936 542218 -1814 542454
rect -1578 542218 20000 542454
rect -2936 542134 20000 542218
rect -2936 541898 -1814 542134
rect -1578 541898 20000 542134
rect -2936 541876 20000 541898
rect 569000 542454 586860 542476
rect 569000 542218 585502 542454
rect 585738 542218 586860 542454
rect 569000 542134 586860 542218
rect 569000 541898 585502 542134
rect 585738 541898 586860 542134
rect 569000 541876 586860 541898
rect -1996 541874 -1396 541876
rect 585320 541874 585920 541876
rect -2936 524476 -2336 524478
rect 586260 524476 586860 524478
rect -2936 524454 20000 524476
rect -2936 524218 -2754 524454
rect -2518 524218 20000 524454
rect -2936 524134 20000 524218
rect -2936 523898 -2754 524134
rect -2518 523898 20000 524134
rect -2936 523876 20000 523898
rect 569000 524454 586860 524476
rect 569000 524218 586442 524454
rect 586678 524218 586860 524454
rect 569000 524134 586860 524218
rect 569000 523898 586442 524134
rect 586678 523898 586860 524134
rect 569000 523876 586860 523898
rect -2936 523874 -2336 523876
rect 586260 523874 586860 523876
rect -1996 506476 -1396 506478
rect 585320 506476 585920 506478
rect -2936 506454 20000 506476
rect -2936 506218 -1814 506454
rect -1578 506218 20000 506454
rect -2936 506134 20000 506218
rect -2936 505898 -1814 506134
rect -1578 505898 20000 506134
rect -2936 505876 20000 505898
rect 569000 506454 586860 506476
rect 569000 506218 585502 506454
rect 585738 506218 586860 506454
rect 569000 506134 586860 506218
rect 569000 505898 585502 506134
rect 585738 505898 586860 506134
rect 569000 505876 586860 505898
rect -1996 505874 -1396 505876
rect 585320 505874 585920 505876
rect -2936 488476 -2336 488478
rect 586260 488476 586860 488478
rect -2936 488454 20000 488476
rect -2936 488218 -2754 488454
rect -2518 488218 20000 488454
rect -2936 488134 20000 488218
rect -2936 487898 -2754 488134
rect -2518 487898 20000 488134
rect -2936 487876 20000 487898
rect 569000 488454 586860 488476
rect 569000 488218 586442 488454
rect 586678 488218 586860 488454
rect 569000 488134 586860 488218
rect 569000 487898 586442 488134
rect 586678 487898 586860 488134
rect 569000 487876 586860 487898
rect -2936 487874 -2336 487876
rect 586260 487874 586860 487876
rect -1996 470476 -1396 470478
rect 585320 470476 585920 470478
rect -2936 470454 20000 470476
rect -2936 470218 -1814 470454
rect -1578 470218 20000 470454
rect -2936 470134 20000 470218
rect -2936 469898 -1814 470134
rect -1578 469898 20000 470134
rect -2936 469876 20000 469898
rect 569000 470454 586860 470476
rect 569000 470218 585502 470454
rect 585738 470218 586860 470454
rect 569000 470134 586860 470218
rect 569000 469898 585502 470134
rect 585738 469898 586860 470134
rect 569000 469876 586860 469898
rect -1996 469874 -1396 469876
rect 585320 469874 585920 469876
rect -2936 452476 -2336 452478
rect 586260 452476 586860 452478
rect -2936 452454 20000 452476
rect -2936 452218 -2754 452454
rect -2518 452218 20000 452454
rect -2936 452134 20000 452218
rect -2936 451898 -2754 452134
rect -2518 451898 20000 452134
rect -2936 451876 20000 451898
rect 569000 452454 586860 452476
rect 569000 452218 586442 452454
rect 586678 452218 586860 452454
rect 569000 452134 586860 452218
rect 569000 451898 586442 452134
rect 586678 451898 586860 452134
rect 569000 451876 586860 451898
rect -2936 451874 -2336 451876
rect 586260 451874 586860 451876
rect -1996 434476 -1396 434478
rect 585320 434476 585920 434478
rect -2936 434454 20000 434476
rect -2936 434218 -1814 434454
rect -1578 434218 20000 434454
rect -2936 434134 20000 434218
rect -2936 433898 -1814 434134
rect -1578 433898 20000 434134
rect -2936 433876 20000 433898
rect 569000 434454 586860 434476
rect 569000 434218 585502 434454
rect 585738 434218 586860 434454
rect 569000 434134 586860 434218
rect 569000 433898 585502 434134
rect 585738 433898 586860 434134
rect 569000 433876 586860 433898
rect -1996 433874 -1396 433876
rect 585320 433874 585920 433876
rect -2936 416476 -2336 416478
rect 586260 416476 586860 416478
rect -2936 416454 20000 416476
rect -2936 416218 -2754 416454
rect -2518 416218 20000 416454
rect -2936 416134 20000 416218
rect -2936 415898 -2754 416134
rect -2518 415898 20000 416134
rect -2936 415876 20000 415898
rect 569000 416454 586860 416476
rect 569000 416218 586442 416454
rect 586678 416218 586860 416454
rect 569000 416134 586860 416218
rect 569000 415898 586442 416134
rect 586678 415898 586860 416134
rect 569000 415876 586860 415898
rect -2936 415874 -2336 415876
rect 586260 415874 586860 415876
rect -1996 398476 -1396 398478
rect 585320 398476 585920 398478
rect -2936 398454 20000 398476
rect -2936 398218 -1814 398454
rect -1578 398218 20000 398454
rect -2936 398134 20000 398218
rect -2936 397898 -1814 398134
rect -1578 397898 20000 398134
rect -2936 397876 20000 397898
rect 569000 398454 586860 398476
rect 569000 398218 585502 398454
rect 585738 398218 586860 398454
rect 569000 398134 586860 398218
rect 569000 397898 585502 398134
rect 585738 397898 586860 398134
rect 569000 397876 586860 397898
rect -1996 397874 -1396 397876
rect 585320 397874 585920 397876
rect -2936 380476 -2336 380478
rect 586260 380476 586860 380478
rect -2936 380454 20000 380476
rect -2936 380218 -2754 380454
rect -2518 380218 20000 380454
rect -2936 380134 20000 380218
rect -2936 379898 -2754 380134
rect -2518 379898 20000 380134
rect -2936 379876 20000 379898
rect 569000 380454 586860 380476
rect 569000 380218 586442 380454
rect 586678 380218 586860 380454
rect 569000 380134 586860 380218
rect 569000 379898 586442 380134
rect 586678 379898 586860 380134
rect 569000 379876 586860 379898
rect -2936 379874 -2336 379876
rect 586260 379874 586860 379876
rect -1996 362476 -1396 362478
rect 585320 362476 585920 362478
rect -2936 362454 20000 362476
rect -2936 362218 -1814 362454
rect -1578 362218 20000 362454
rect -2936 362134 20000 362218
rect -2936 361898 -1814 362134
rect -1578 361898 20000 362134
rect -2936 361876 20000 361898
rect 569000 362454 586860 362476
rect 569000 362218 585502 362454
rect 585738 362218 586860 362454
rect 569000 362134 586860 362218
rect 569000 361898 585502 362134
rect 585738 361898 586860 362134
rect 569000 361876 586860 361898
rect -1996 361874 -1396 361876
rect 585320 361874 585920 361876
rect -2936 344476 -2336 344478
rect 586260 344476 586860 344478
rect -2936 344454 20000 344476
rect -2936 344218 -2754 344454
rect -2518 344218 20000 344454
rect -2936 344134 20000 344218
rect -2936 343898 -2754 344134
rect -2518 343898 20000 344134
rect -2936 343876 20000 343898
rect 569000 344454 586860 344476
rect 569000 344218 586442 344454
rect 586678 344218 586860 344454
rect 569000 344134 586860 344218
rect 569000 343898 586442 344134
rect 586678 343898 586860 344134
rect 569000 343876 586860 343898
rect -2936 343874 -2336 343876
rect 586260 343874 586860 343876
rect -1996 326476 -1396 326478
rect 585320 326476 585920 326478
rect -2936 326454 20000 326476
rect -2936 326218 -1814 326454
rect -1578 326218 20000 326454
rect -2936 326134 20000 326218
rect -2936 325898 -1814 326134
rect -1578 325898 20000 326134
rect -2936 325876 20000 325898
rect 569000 326454 586860 326476
rect 569000 326218 585502 326454
rect 585738 326218 586860 326454
rect 569000 326134 586860 326218
rect 569000 325898 585502 326134
rect 585738 325898 586860 326134
rect 569000 325876 586860 325898
rect -1996 325874 -1396 325876
rect 585320 325874 585920 325876
rect -2936 308476 -2336 308478
rect 586260 308476 586860 308478
rect -2936 308454 20000 308476
rect -2936 308218 -2754 308454
rect -2518 308218 20000 308454
rect -2936 308134 20000 308218
rect -2936 307898 -2754 308134
rect -2518 307898 20000 308134
rect -2936 307876 20000 307898
rect 569000 308454 586860 308476
rect 569000 308218 586442 308454
rect 586678 308218 586860 308454
rect 569000 308134 586860 308218
rect 569000 307898 586442 308134
rect 586678 307898 586860 308134
rect 569000 307876 586860 307898
rect -2936 307874 -2336 307876
rect 586260 307874 586860 307876
rect -1996 290476 -1396 290478
rect 585320 290476 585920 290478
rect -2936 290454 20000 290476
rect -2936 290218 -1814 290454
rect -1578 290218 20000 290454
rect -2936 290134 20000 290218
rect -2936 289898 -1814 290134
rect -1578 289898 20000 290134
rect -2936 289876 20000 289898
rect 569000 290454 586860 290476
rect 569000 290218 585502 290454
rect 585738 290218 586860 290454
rect 569000 290134 586860 290218
rect 569000 289898 585502 290134
rect 585738 289898 586860 290134
rect 569000 289876 586860 289898
rect -1996 289874 -1396 289876
rect 585320 289874 585920 289876
rect -2936 272476 -2336 272478
rect 586260 272476 586860 272478
rect -2936 272454 20000 272476
rect -2936 272218 -2754 272454
rect -2518 272218 20000 272454
rect -2936 272134 20000 272218
rect -2936 271898 -2754 272134
rect -2518 271898 20000 272134
rect -2936 271876 20000 271898
rect 569000 272454 586860 272476
rect 569000 272218 586442 272454
rect 586678 272218 586860 272454
rect 569000 272134 586860 272218
rect 569000 271898 586442 272134
rect 586678 271898 586860 272134
rect 569000 271876 586860 271898
rect -2936 271874 -2336 271876
rect 586260 271874 586860 271876
rect -1996 254476 -1396 254478
rect 585320 254476 585920 254478
rect -2936 254454 20000 254476
rect -2936 254218 -1814 254454
rect -1578 254218 20000 254454
rect -2936 254134 20000 254218
rect -2936 253898 -1814 254134
rect -1578 253898 20000 254134
rect -2936 253876 20000 253898
rect 569000 254454 586860 254476
rect 569000 254218 585502 254454
rect 585738 254218 586860 254454
rect 569000 254134 586860 254218
rect 569000 253898 585502 254134
rect 585738 253898 586860 254134
rect 569000 253876 586860 253898
rect -1996 253874 -1396 253876
rect 585320 253874 585920 253876
rect -2936 236476 -2336 236478
rect 586260 236476 586860 236478
rect -2936 236454 20000 236476
rect -2936 236218 -2754 236454
rect -2518 236218 20000 236454
rect -2936 236134 20000 236218
rect -2936 235898 -2754 236134
rect -2518 235898 20000 236134
rect -2936 235876 20000 235898
rect 569000 236454 586860 236476
rect 569000 236218 586442 236454
rect 586678 236218 586860 236454
rect 569000 236134 586860 236218
rect 569000 235898 586442 236134
rect 586678 235898 586860 236134
rect 569000 235876 586860 235898
rect -2936 235874 -2336 235876
rect 586260 235874 586860 235876
rect -1996 218476 -1396 218478
rect 585320 218476 585920 218478
rect -2936 218454 20000 218476
rect -2936 218218 -1814 218454
rect -1578 218218 20000 218454
rect -2936 218134 20000 218218
rect -2936 217898 -1814 218134
rect -1578 217898 20000 218134
rect -2936 217876 20000 217898
rect 569000 218454 586860 218476
rect 569000 218218 585502 218454
rect 585738 218218 586860 218454
rect 569000 218134 586860 218218
rect 569000 217898 585502 218134
rect 585738 217898 586860 218134
rect 569000 217876 586860 217898
rect -1996 217874 -1396 217876
rect 585320 217874 585920 217876
rect -2936 200476 -2336 200478
rect 586260 200476 586860 200478
rect -2936 200454 20000 200476
rect -2936 200218 -2754 200454
rect -2518 200218 20000 200454
rect -2936 200134 20000 200218
rect -2936 199898 -2754 200134
rect -2518 199898 20000 200134
rect -2936 199876 20000 199898
rect 569000 200454 586860 200476
rect 569000 200218 586442 200454
rect 586678 200218 586860 200454
rect 569000 200134 586860 200218
rect 569000 199898 586442 200134
rect 586678 199898 586860 200134
rect 569000 199876 586860 199898
rect -2936 199874 -2336 199876
rect 586260 199874 586860 199876
rect -1996 182476 -1396 182478
rect 585320 182476 585920 182478
rect -2936 182454 20000 182476
rect -2936 182218 -1814 182454
rect -1578 182218 20000 182454
rect -2936 182134 20000 182218
rect -2936 181898 -1814 182134
rect -1578 181898 20000 182134
rect -2936 181876 20000 181898
rect 569000 182454 586860 182476
rect 569000 182218 585502 182454
rect 585738 182218 586860 182454
rect 569000 182134 586860 182218
rect 569000 181898 585502 182134
rect 585738 181898 586860 182134
rect 569000 181876 586860 181898
rect -1996 181874 -1396 181876
rect 585320 181874 585920 181876
rect -2936 164476 -2336 164478
rect 586260 164476 586860 164478
rect -2936 164454 20000 164476
rect -2936 164218 -2754 164454
rect -2518 164218 20000 164454
rect -2936 164134 20000 164218
rect -2936 163898 -2754 164134
rect -2518 163898 20000 164134
rect -2936 163876 20000 163898
rect 569000 164454 586860 164476
rect 569000 164218 586442 164454
rect 586678 164218 586860 164454
rect 569000 164134 586860 164218
rect 569000 163898 586442 164134
rect 586678 163898 586860 164134
rect 569000 163876 586860 163898
rect -2936 163874 -2336 163876
rect 586260 163874 586860 163876
rect -1996 146476 -1396 146478
rect 585320 146476 585920 146478
rect -2936 146454 20000 146476
rect -2936 146218 -1814 146454
rect -1578 146218 20000 146454
rect -2936 146134 20000 146218
rect -2936 145898 -1814 146134
rect -1578 145898 20000 146134
rect -2936 145876 20000 145898
rect 569000 146454 586860 146476
rect 569000 146218 585502 146454
rect 585738 146218 586860 146454
rect 569000 146134 586860 146218
rect 569000 145898 585502 146134
rect 585738 145898 586860 146134
rect 569000 145876 586860 145898
rect -1996 145874 -1396 145876
rect 585320 145874 585920 145876
rect -2936 128476 -2336 128478
rect 586260 128476 586860 128478
rect -2936 128454 20000 128476
rect -2936 128218 -2754 128454
rect -2518 128218 20000 128454
rect -2936 128134 20000 128218
rect -2936 127898 -2754 128134
rect -2518 127898 20000 128134
rect -2936 127876 20000 127898
rect 569000 128454 586860 128476
rect 569000 128218 586442 128454
rect 586678 128218 586860 128454
rect 569000 128134 586860 128218
rect 569000 127898 586442 128134
rect 586678 127898 586860 128134
rect 569000 127876 586860 127898
rect -2936 127874 -2336 127876
rect 586260 127874 586860 127876
rect -1996 110476 -1396 110478
rect 585320 110476 585920 110478
rect -2936 110454 20000 110476
rect -2936 110218 -1814 110454
rect -1578 110218 20000 110454
rect -2936 110134 20000 110218
rect -2936 109898 -1814 110134
rect -1578 109898 20000 110134
rect -2936 109876 20000 109898
rect 569000 110454 586860 110476
rect 569000 110218 585502 110454
rect 585738 110218 586860 110454
rect 569000 110134 586860 110218
rect 569000 109898 585502 110134
rect 585738 109898 586860 110134
rect 569000 109876 586860 109898
rect -1996 109874 -1396 109876
rect 585320 109874 585920 109876
rect -2936 92476 -2336 92478
rect 586260 92476 586860 92478
rect -2936 92454 20000 92476
rect -2936 92218 -2754 92454
rect -2518 92218 20000 92454
rect -2936 92134 20000 92218
rect -2936 91898 -2754 92134
rect -2518 91898 20000 92134
rect -2936 91876 20000 91898
rect 569000 92454 586860 92476
rect 569000 92218 586442 92454
rect 586678 92218 586860 92454
rect 569000 92134 586860 92218
rect 569000 91898 586442 92134
rect 586678 91898 586860 92134
rect 569000 91876 586860 91898
rect -2936 91874 -2336 91876
rect 586260 91874 586860 91876
rect -1996 74476 -1396 74478
rect 585320 74476 585920 74478
rect -2936 74454 20000 74476
rect -2936 74218 -1814 74454
rect -1578 74218 20000 74454
rect -2936 74134 20000 74218
rect -2936 73898 -1814 74134
rect -1578 73898 20000 74134
rect -2936 73876 20000 73898
rect 569000 74454 586860 74476
rect 569000 74218 585502 74454
rect 585738 74218 586860 74454
rect 569000 74134 586860 74218
rect 569000 73898 585502 74134
rect 585738 73898 586860 74134
rect 569000 73876 586860 73898
rect -1996 73874 -1396 73876
rect 585320 73874 585920 73876
rect -2936 56476 -2336 56478
rect 586260 56476 586860 56478
rect -2936 56454 20000 56476
rect -2936 56218 -2754 56454
rect -2518 56218 20000 56454
rect -2936 56134 20000 56218
rect -2936 55898 -2754 56134
rect -2518 55898 20000 56134
rect -2936 55876 20000 55898
rect 569000 56454 586860 56476
rect 569000 56218 586442 56454
rect 586678 56218 586860 56454
rect 569000 56134 586860 56218
rect 569000 55898 586442 56134
rect 586678 55898 586860 56134
rect 569000 55876 586860 55898
rect -2936 55874 -2336 55876
rect 586260 55874 586860 55876
rect -1996 38476 -1396 38478
rect 585320 38476 585920 38478
rect -2936 38454 20000 38476
rect -2936 38218 -1814 38454
rect -1578 38218 20000 38454
rect -2936 38134 20000 38218
rect -2936 37898 -1814 38134
rect -1578 37898 20000 38134
rect -2936 37876 20000 37898
rect 569000 38454 586860 38476
rect 569000 38218 585502 38454
rect 585738 38218 586860 38454
rect 569000 38134 586860 38218
rect 569000 37898 585502 38134
rect 585738 37898 586860 38134
rect 569000 37876 586860 37898
rect -1996 37874 -1396 37876
rect 585320 37874 585920 37876
rect -2936 20476 -2336 20478
rect 586260 20476 586860 20478
rect -2936 20454 20000 20476
rect -2936 20218 -2754 20454
rect -2518 20218 20000 20454
rect -2936 20134 20000 20218
rect -2936 19898 -2754 20134
rect -2518 19898 20000 20134
rect -2936 19876 20000 19898
rect 569000 20454 586860 20476
rect 569000 20218 586442 20454
rect 586678 20218 586860 20454
rect 569000 20134 586860 20218
rect 569000 19898 586442 20134
rect 586678 19898 586860 20134
rect 569000 19876 586860 19898
rect -2936 19874 -2336 19876
rect 586260 19874 586860 19876
rect -1996 2476 -1396 2478
rect 37072 2476 37672 2478
rect 184814 2476 185414 2478
rect 332556 2476 333156 2478
rect 480298 2476 480898 2478
rect 585320 2476 585920 2478
rect -2936 2454 586860 2476
rect -2936 2218 -1814 2454
rect -1578 2218 37254 2454
rect 37490 2218 184996 2454
rect 185232 2218 332738 2454
rect 332974 2218 480480 2454
rect 480716 2218 585502 2454
rect 585738 2218 586860 2454
rect -2936 2134 586860 2218
rect -2936 1898 -1814 2134
rect -1578 1898 37254 2134
rect 37490 1898 184996 2134
rect 185232 1898 332738 2134
rect 332974 1898 480480 2134
rect 480716 1898 585502 2134
rect 585738 1898 586860 2134
rect -2936 1876 586860 1898
rect -1996 1874 -1396 1876
rect 37072 1874 37672 1876
rect 184814 1874 185414 1876
rect 332556 1874 333156 1876
rect 480298 1874 480898 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 37072 -324 37672 -322
rect 184814 -324 185414 -322
rect 332556 -324 333156 -322
rect 480298 -324 480898 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 37254 -346
rect 37490 -582 184996 -346
rect 185232 -582 332738 -346
rect 332974 -582 480480 -346
rect 480716 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 37254 -666
rect 37490 -902 184996 -666
rect 185232 -902 332738 -666
rect 332974 -902 480480 -666
rect 480716 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 37072 -926 37672 -924
rect 184814 -926 185414 -924
rect 332556 -926 333156 -924
rect 480298 -926 480898 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 110943 -1264 111543 -1262
rect 258685 -1264 259285 -1262
rect 406427 -1264 407027 -1262
rect 554169 -1264 554769 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 111125 -1286
rect 111361 -1522 258867 -1286
rect 259103 -1522 406609 -1286
rect 406845 -1522 554351 -1286
rect 554587 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 111125 -1606
rect 111361 -1842 258867 -1606
rect 259103 -1842 406609 -1606
rect 406845 -1842 554351 -1606
rect 554587 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 110943 -1866 111543 -1864
rect 258685 -1866 259285 -1864
rect 406427 -1866 407027 -1864
rect 554169 -1866 554769 -1864
rect 586260 -1866 586860 -1864
use fpga  fpga250
timestamp 1608322654
transform 1 0 20000 0 1 20000
box 0 0 549000 664000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 637 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>

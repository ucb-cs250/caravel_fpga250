VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga
  CLASS BLOCK ;
  FOREIGN fpga ;
  ORIGIN -0.005 0.000 ;
  SIZE 3843.105 BY 3888.080 ;
  PIN gpio_east[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 3789.690 74.080 3793.690 74.680 ;
    END
  END gpio_east[0]
  PIN gpio_east[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 3789.690 133.920 3793.690 134.520 ;
    END
  END gpio_east[1]
  PIN gpio_east[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 3789.690 194.440 3793.690 195.040 ;
    END
  END gpio_east[2]
  PIN gpio_east[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 3789.690 254.960 3793.690 255.560 ;
    END
  END gpio_east[3]
  PIN gpio_east[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 3789.690 314.800 3793.690 315.400 ;
    END
  END gpio_east[4]
  PIN gpio_east[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 3789.690 375.320 3793.690 375.920 ;
    END
  END gpio_east[5]
  PIN gpio_east[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 3789.690 435.840 3793.690 436.440 ;
    END
  END gpio_east[6]
  PIN gpio_east[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 3789.690 495.680 3793.690 496.280 ;
    END
  END gpio_east[7]
  PIN gpio_east[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 3789.690 556.200 3793.690 556.800 ;
    END
  END gpio_east[8]
  PIN gpio_east[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 3789.690 616.720 3793.690 617.320 ;
    END
  END gpio_east[9]
  PIN gpio_north[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 748.980 3840.120 749.260 3844.120 ;
    END
  END gpio_north[0]
  PIN gpio_north[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 859.380 3840.120 859.660 3844.120 ;
    END
  END gpio_north[1]
  PIN gpio_north[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 970.240 3840.120 970.520 3844.120 ;
    END
  END gpio_north[2]
  PIN gpio_north[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1081.100 3840.120 1081.380 3844.120 ;
    END
  END gpio_north[3]
  PIN gpio_north[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1191.500 3840.120 1191.780 3844.120 ;
    END
  END gpio_north[4]
  PIN gpio_north[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1302.360 3840.120 1302.640 3844.120 ;
    END
  END gpio_north[5]
  PIN gpio_north[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1413.220 3840.120 1413.500 3844.120 ;
    END
  END gpio_north[6]
  PIN gpio_north[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1523.620 3840.120 1523.900 3844.120 ;
    END
  END gpio_north[7]
  PIN gpio_north[8]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1634.480 3840.120 1634.760 3844.120 ;
    END
  END gpio_north[8]
  PIN gpio_north[9]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1745.340 3840.120 1745.620 3844.120 ;
    END
  END gpio_north[9]
  PIN gpio_south[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 755.420 44.120 755.700 48.120 ;
    END
  END gpio_south[0]
  PIN gpio_south[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 879.160 44.120 879.440 48.120 ;
    END
  END gpio_south[1]
  PIN gpio_south[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1003.360 44.120 1003.640 48.120 ;
    END
  END gpio_south[2]
  PIN gpio_south[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1127.100 44.120 1127.380 48.120 ;
    END
  END gpio_south[3]
  PIN gpio_south[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1251.300 44.120 1251.580 48.120 ;
    END
  END gpio_south[4]
  PIN gpio_south[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1375.040 44.120 1375.320 48.120 ;
    END
  END gpio_south[5]
  PIN gpio_south[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1499.240 44.120 1499.520 48.120 ;
    END
  END gpio_south[6]
  PIN gpio_south[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1622.980 44.120 1623.260 48.120 ;
    END
  END gpio_south[7]
  PIN gpio_west[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 693.690 111.480 697.690 112.080 ;
    END
  END gpio_west[0]
  PIN gpio_west[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 693.690 246.800 697.690 247.400 ;
    END
  END gpio_west[1]
  PIN gpio_west[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 693.690 382.800 697.690 383.400 ;
    END
  END gpio_west[2]
  PIN gpio_west[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 693.690 518.120 697.690 518.720 ;
    END
  END gpio_west[3]
  PIN gpio_west[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 693.690 654.120 697.690 654.720 ;
    END
  END gpio_west[4]
  PIN gpio_west[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 693.690 789.440 697.690 790.040 ;
    END
  END gpio_west[5]
  PIN gpio_west[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 693.690 925.440 697.690 926.040 ;
    END
  END gpio_west[6]
  PIN gpio_west[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 693.690 1061.440 697.690 1062.040 ;
    END
  END gpio_west[7]
  PIN gpio_west[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 693.690 1196.760 697.690 1197.360 ;
    END
  END gpio_west[8]
  PIN gpio_west[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 693.690 1332.760 697.690 1333.360 ;
    END
  END gpio_west[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1855.740 3840.120 1856.020 3844.120 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1747.180 44.120 1747.460 48.120 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1966.600 3840.120 1966.880 3844.120 ;
    END
  END wbs_ack_o
  PIN wbs_addr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3789.690 2607.080 3793.690 2607.680 ;
    END
  END wbs_addr_i[0]
  PIN wbs_addr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3789.690 2727.440 3793.690 2728.040 ;
    END
  END wbs_addr_i[10]
  PIN wbs_addr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3789.690 2787.960 3793.690 2788.560 ;
    END
  END wbs_addr_i[11]
  PIN wbs_addr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2519.980 3840.120 2520.260 3844.120 ;
    END
  END wbs_addr_i[12]
  PIN wbs_addr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1995.120 44.120 1995.400 48.120 ;
    END
  END wbs_addr_i[13]
  PIN wbs_addr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2119.320 44.120 2119.600 48.120 ;
    END
  END wbs_addr_i[14]
  PIN wbs_addr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 693.690 1875.400 697.690 1876.000 ;
    END
  END wbs_addr_i[15]
  PIN wbs_addr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2630.840 3840.120 2631.120 3844.120 ;
    END
  END wbs_addr_i[16]
  PIN wbs_addr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3789.690 2848.480 3793.690 2849.080 ;
    END
  END wbs_addr_i[17]
  PIN wbs_addr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2741.700 3840.120 2741.980 3844.120 ;
    END
  END wbs_addr_i[18]
  PIN wbs_addr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2852.100 3840.120 2852.380 3844.120 ;
    END
  END wbs_addr_i[19]
  PIN wbs_addr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 693.690 1468.080 697.690 1468.680 ;
    END
  END wbs_addr_i[1]
  PIN wbs_addr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2243.060 44.120 2243.340 48.120 ;
    END
  END wbs_addr_i[20]
  PIN wbs_addr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2367.260 44.120 2367.540 48.120 ;
    END
  END wbs_addr_i[21]
  PIN wbs_addr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3789.690 2908.320 3793.690 2908.920 ;
    END
  END wbs_addr_i[22]
  PIN wbs_addr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2962.960 3840.120 2963.240 3844.120 ;
    END
  END wbs_addr_i[23]
  PIN wbs_addr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3073.820 3840.120 3074.100 3844.120 ;
    END
  END wbs_addr_i[24]
  PIN wbs_addr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3184.220 3840.120 3184.500 3844.120 ;
    END
  END wbs_addr_i[25]
  PIN wbs_addr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2491.000 44.120 2491.280 48.120 ;
    END
  END wbs_addr_i[26]
  PIN wbs_addr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 693.690 2011.400 697.690 2012.000 ;
    END
  END wbs_addr_i[27]
  PIN wbs_addr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 693.690 2146.720 697.690 2147.320 ;
    END
  END wbs_addr_i[28]
  PIN wbs_addr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3789.690 2968.840 3793.690 2969.440 ;
    END
  END wbs_addr_i[29]
  PIN wbs_addr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3789.690 2667.600 3793.690 2668.200 ;
    END
  END wbs_addr_i[2]
  PIN wbs_addr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 693.690 2282.720 697.690 2283.320 ;
    END
  END wbs_addr_i[30]
  PIN wbs_addr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3789.690 3029.360 3793.690 3029.960 ;
    END
  END wbs_addr_i[31]
  PIN wbs_addr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 693.690 1604.080 697.690 1604.680 ;
    END
  END wbs_addr_i[3]
  PIN wbs_addr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2077.460 3840.120 2077.740 3844.120 ;
    END
  END wbs_addr_i[4]
  PIN wbs_addr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 693.690 1739.400 697.690 1740.000 ;
    END
  END wbs_addr_i[5]
  PIN wbs_addr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2187.860 3840.120 2188.140 3844.120 ;
    END
  END wbs_addr_i[6]
  PIN wbs_addr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2298.720 3840.120 2299.000 3844.120 ;
    END
  END wbs_addr_i[7]
  PIN wbs_addr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2409.580 3840.120 2409.860 3844.120 ;
    END
  END wbs_addr_i[8]
  PIN wbs_addr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1871.380 44.120 1871.660 48.120 ;
    END
  END wbs_addr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 693.690 2418.040 697.690 2418.640 ;
    END
  END wbs_cyc_i
  PIN wbs_data_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2615.200 44.120 2615.480 48.120 ;
    END
  END wbs_data_i[0]
  PIN wbs_data_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 693.690 2825.360 697.690 2825.960 ;
    END
  END wbs_data_i[10]
  PIN wbs_data_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3111.080 44.120 3111.360 48.120 ;
    END
  END wbs_data_i[11]
  PIN wbs_data_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3789.690 3330.600 3793.690 3331.200 ;
    END
  END wbs_data_i[12]
  PIN wbs_data_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3295.080 3840.120 3295.360 3844.120 ;
    END
  END wbs_data_i[13]
  PIN wbs_data_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3405.940 3840.120 3406.220 3844.120 ;
    END
  END wbs_data_i[14]
  PIN wbs_data_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3789.690 3391.120 3793.690 3391.720 ;
    END
  END wbs_data_i[15]
  PIN wbs_data_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3235.280 44.120 3235.560 48.120 ;
    END
  END wbs_data_i[16]
  PIN wbs_data_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3516.340 3840.120 3516.620 3844.120 ;
    END
  END wbs_data_i[17]
  PIN wbs_data_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3359.020 44.120 3359.300 48.120 ;
    END
  END wbs_data_i[18]
  PIN wbs_data_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 693.690 2961.360 697.690 2961.960 ;
    END
  END wbs_data_i[19]
  PIN wbs_data_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3789.690 3089.200 3793.690 3089.800 ;
    END
  END wbs_data_i[1]
  PIN wbs_data_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3789.690 3451.640 3793.690 3452.240 ;
    END
  END wbs_data_i[20]
  PIN wbs_data_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3789.690 3511.480 3793.690 3512.080 ;
    END
  END wbs_data_i[21]
  PIN wbs_data_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 693.690 3096.680 697.690 3097.280 ;
    END
  END wbs_data_i[22]
  PIN wbs_data_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 693.690 3232.680 697.690 3233.280 ;
    END
  END wbs_data_i[23]
  PIN wbs_data_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 693.690 3368.000 697.690 3368.600 ;
    END
  END wbs_data_i[24]
  PIN wbs_data_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3483.220 44.120 3483.500 48.120 ;
    END
  END wbs_data_i[25]
  PIN wbs_data_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 693.690 3504.000 697.690 3504.600 ;
    END
  END wbs_data_i[26]
  PIN wbs_data_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 693.690 3639.320 697.690 3639.920 ;
    END
  END wbs_data_i[27]
  PIN wbs_data_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3627.200 3840.120 3627.480 3844.120 ;
    END
  END wbs_data_i[28]
  PIN wbs_data_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3789.690 3572.000 3793.690 3572.600 ;
    END
  END wbs_data_i[29]
  PIN wbs_data_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3789.690 3149.720 3793.690 3150.320 ;
    END
  END wbs_data_i[2]
  PIN wbs_data_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3606.960 44.120 3607.240 48.120 ;
    END
  END wbs_data_i[30]
  PIN wbs_data_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3789.690 3632.520 3793.690 3633.120 ;
    END
  END wbs_data_i[31]
  PIN wbs_data_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 693.690 2554.040 697.690 2554.640 ;
    END
  END wbs_data_i[3]
  PIN wbs_data_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 693.690 2689.360 697.690 2689.960 ;
    END
  END wbs_data_i[4]
  PIN wbs_data_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3789.690 3210.240 3793.690 3210.840 ;
    END
  END wbs_data_i[5]
  PIN wbs_data_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2738.940 44.120 2739.220 48.120 ;
    END
  END wbs_data_i[6]
  PIN wbs_data_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2863.140 44.120 2863.420 48.120 ;
    END
  END wbs_data_i[7]
  PIN wbs_data_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2987.340 44.120 2987.620 48.120 ;
    END
  END wbs_data_i[8]
  PIN wbs_data_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3789.690 3270.760 3793.690 3271.360 ;
    END
  END wbs_data_i[9]
  PIN wbs_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3789.690 676.560 3793.690 677.160 ;
    END
  END wbs_data_o[0]
  PIN wbs_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3789.690 1279.720 3793.690 1280.320 ;
    END
  END wbs_data_o[10]
  PIN wbs_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3789.690 1340.240 3793.690 1340.840 ;
    END
  END wbs_data_o[11]
  PIN wbs_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3789.690 1400.760 3793.690 1401.360 ;
    END
  END wbs_data_o[12]
  PIN wbs_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3789.690 1461.280 3793.690 1461.880 ;
    END
  END wbs_data_o[13]
  PIN wbs_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3789.690 1521.120 3793.690 1521.720 ;
    END
  END wbs_data_o[14]
  PIN wbs_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3789.690 1581.640 3793.690 1582.240 ;
    END
  END wbs_data_o[15]
  PIN wbs_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3789.690 1642.160 3793.690 1642.760 ;
    END
  END wbs_data_o[16]
  PIN wbs_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3789.690 1702.000 3793.690 1702.600 ;
    END
  END wbs_data_o[17]
  PIN wbs_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3789.690 1762.520 3793.690 1763.120 ;
    END
  END wbs_data_o[18]
  PIN wbs_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3789.690 1823.040 3793.690 1823.640 ;
    END
  END wbs_data_o[19]
  PIN wbs_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3789.690 737.080 3793.690 737.680 ;
    END
  END wbs_data_o[1]
  PIN wbs_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3789.690 1882.880 3793.690 1883.480 ;
    END
  END wbs_data_o[20]
  PIN wbs_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3789.690 1943.400 3793.690 1944.000 ;
    END
  END wbs_data_o[21]
  PIN wbs_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3789.690 2003.920 3793.690 2004.520 ;
    END
  END wbs_data_o[22]
  PIN wbs_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3789.690 2064.440 3793.690 2065.040 ;
    END
  END wbs_data_o[23]
  PIN wbs_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3789.690 2124.280 3793.690 2124.880 ;
    END
  END wbs_data_o[24]
  PIN wbs_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3789.690 2184.800 3793.690 2185.400 ;
    END
  END wbs_data_o[25]
  PIN wbs_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3789.690 2245.320 3793.690 2245.920 ;
    END
  END wbs_data_o[26]
  PIN wbs_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3789.690 2305.160 3793.690 2305.760 ;
    END
  END wbs_data_o[27]
  PIN wbs_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3789.690 2365.680 3793.690 2366.280 ;
    END
  END wbs_data_o[28]
  PIN wbs_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3789.690 2426.200 3793.690 2426.800 ;
    END
  END wbs_data_o[29]
  PIN wbs_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3789.690 797.600 3793.690 798.200 ;
    END
  END wbs_data_o[2]
  PIN wbs_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3789.690 2486.040 3793.690 2486.640 ;
    END
  END wbs_data_o[30]
  PIN wbs_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3789.690 2546.560 3793.690 2547.160 ;
    END
  END wbs_data_o[31]
  PIN wbs_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3789.690 858.120 3793.690 858.720 ;
    END
  END wbs_data_o[3]
  PIN wbs_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3789.690 917.960 3793.690 918.560 ;
    END
  END wbs_data_o[4]
  PIN wbs_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3789.690 978.480 3793.690 979.080 ;
    END
  END wbs_data_o[5]
  PIN wbs_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3789.690 1039.000 3793.690 1039.600 ;
    END
  END wbs_data_o[6]
  PIN wbs_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3789.690 1098.840 3793.690 1099.440 ;
    END
  END wbs_data_o[7]
  PIN wbs_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3789.690 1159.360 3793.690 1159.960 ;
    END
  END wbs_data_o[8]
  PIN wbs_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3789.690 1219.880 3793.690 1220.480 ;
    END
  END wbs_data_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3789.690 3692.360 3793.690 3692.960 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3789.690 3752.880 3793.690 3753.480 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3789.690 3813.400 3793.690 3814.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3738.060 3840.120 3738.340 3844.120 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 693.690 3775.320 697.690 3775.920 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3731.160 44.120 3731.440 48.120 ;
    END
  END wbs_we_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 669.210 25.000 3818.110 45.000 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 644.210 0.000 3843.110 20.000 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 699.210 54.915 3788.110 3833.165 ;
      LAYER met1 ;
        RECT 699.210 54.760 3788.110 3833.320 ;
      LAYER met2 ;
        RECT 708.040 3839.840 748.700 3840.120 ;
        RECT 749.540 3839.840 859.100 3840.120 ;
        RECT 859.940 3839.840 969.960 3840.120 ;
        RECT 970.800 3839.840 1080.820 3840.120 ;
        RECT 1081.660 3839.840 1191.220 3840.120 ;
        RECT 1192.060 3839.840 1302.080 3840.120 ;
        RECT 1302.920 3839.840 1412.940 3840.120 ;
        RECT 1413.780 3839.840 1523.340 3840.120 ;
        RECT 1524.180 3839.840 1634.200 3840.120 ;
        RECT 1635.040 3839.840 1745.060 3840.120 ;
        RECT 1745.900 3839.840 1855.460 3840.120 ;
        RECT 1856.300 3839.840 1966.320 3840.120 ;
        RECT 1967.160 3839.840 2077.180 3840.120 ;
        RECT 2078.020 3839.840 2187.580 3840.120 ;
        RECT 2188.420 3839.840 2298.440 3840.120 ;
        RECT 2299.280 3839.840 2409.300 3840.120 ;
        RECT 2410.140 3839.840 2519.700 3840.120 ;
        RECT 2520.540 3839.840 2630.560 3840.120 ;
        RECT 2631.400 3839.840 2741.420 3840.120 ;
        RECT 2742.260 3839.840 2851.820 3840.120 ;
        RECT 2852.660 3839.840 2962.680 3840.120 ;
        RECT 2963.520 3839.840 3073.540 3840.120 ;
        RECT 3074.380 3839.840 3183.940 3840.120 ;
        RECT 3184.780 3839.840 3294.800 3840.120 ;
        RECT 3295.640 3839.840 3405.660 3840.120 ;
        RECT 3406.500 3839.840 3516.060 3840.120 ;
        RECT 3516.900 3839.840 3626.920 3840.120 ;
        RECT 3627.760 3839.840 3737.780 3840.120 ;
        RECT 3738.620 3839.840 3777.900 3840.120 ;
        RECT 708.040 48.400 3777.900 3839.840 ;
        RECT 708.040 48.120 755.140 48.400 ;
        RECT 755.980 48.120 878.880 48.400 ;
        RECT 879.720 48.120 1003.080 48.400 ;
        RECT 1003.920 48.120 1126.820 48.400 ;
        RECT 1127.660 48.120 1251.020 48.400 ;
        RECT 1251.860 48.120 1374.760 48.400 ;
        RECT 1375.600 48.120 1498.960 48.400 ;
        RECT 1499.800 48.120 1622.700 48.400 ;
        RECT 1623.540 48.120 1746.900 48.400 ;
        RECT 1747.740 48.120 1871.100 48.400 ;
        RECT 1871.940 48.120 1994.840 48.400 ;
        RECT 1995.680 48.120 2119.040 48.400 ;
        RECT 2119.880 48.120 2242.780 48.400 ;
        RECT 2243.620 48.120 2366.980 48.400 ;
        RECT 2367.820 48.120 2490.720 48.400 ;
        RECT 2491.560 48.120 2614.920 48.400 ;
        RECT 2615.760 48.120 2738.660 48.400 ;
        RECT 2739.500 48.120 2862.860 48.400 ;
        RECT 2863.700 48.120 2987.060 48.400 ;
        RECT 2987.900 48.120 3110.800 48.400 ;
        RECT 3111.640 48.120 3235.000 48.400 ;
        RECT 3235.840 48.120 3358.740 48.400 ;
        RECT 3359.580 48.120 3482.940 48.400 ;
        RECT 3483.780 48.120 3606.680 48.400 ;
        RECT 3607.520 48.120 3730.880 48.400 ;
        RECT 3731.720 48.120 3777.900 48.400 ;
      LAYER met3 ;
        RECT 697.690 3814.400 3789.690 3833.245 ;
        RECT 697.690 3813.000 3789.290 3814.400 ;
        RECT 697.690 3776.320 3789.690 3813.000 ;
        RECT 698.090 3774.920 3789.690 3776.320 ;
        RECT 697.690 3753.880 3789.690 3774.920 ;
        RECT 697.690 3752.480 3789.290 3753.880 ;
        RECT 697.690 3693.360 3789.690 3752.480 ;
        RECT 697.690 3691.960 3789.290 3693.360 ;
        RECT 697.690 3640.320 3789.690 3691.960 ;
        RECT 698.090 3638.920 3789.690 3640.320 ;
        RECT 697.690 3633.520 3789.690 3638.920 ;
        RECT 697.690 3632.120 3789.290 3633.520 ;
        RECT 697.690 3573.000 3789.690 3632.120 ;
        RECT 697.690 3571.600 3789.290 3573.000 ;
        RECT 697.690 3512.480 3789.690 3571.600 ;
        RECT 697.690 3511.080 3789.290 3512.480 ;
        RECT 697.690 3505.000 3789.690 3511.080 ;
        RECT 698.090 3503.600 3789.690 3505.000 ;
        RECT 697.690 3452.640 3789.690 3503.600 ;
        RECT 697.690 3451.240 3789.290 3452.640 ;
        RECT 697.690 3392.120 3789.690 3451.240 ;
        RECT 697.690 3390.720 3789.290 3392.120 ;
        RECT 697.690 3369.000 3789.690 3390.720 ;
        RECT 698.090 3367.600 3789.690 3369.000 ;
        RECT 697.690 3331.600 3789.690 3367.600 ;
        RECT 697.690 3330.200 3789.290 3331.600 ;
        RECT 697.690 3271.760 3789.690 3330.200 ;
        RECT 697.690 3270.360 3789.290 3271.760 ;
        RECT 697.690 3233.680 3789.690 3270.360 ;
        RECT 698.090 3232.280 3789.690 3233.680 ;
        RECT 697.690 3211.240 3789.690 3232.280 ;
        RECT 697.690 3209.840 3789.290 3211.240 ;
        RECT 697.690 3150.720 3789.690 3209.840 ;
        RECT 697.690 3149.320 3789.290 3150.720 ;
        RECT 697.690 3097.680 3789.690 3149.320 ;
        RECT 698.090 3096.280 3789.690 3097.680 ;
        RECT 697.690 3090.200 3789.690 3096.280 ;
        RECT 697.690 3088.800 3789.290 3090.200 ;
        RECT 697.690 3030.360 3789.690 3088.800 ;
        RECT 697.690 3028.960 3789.290 3030.360 ;
        RECT 697.690 2969.840 3789.690 3028.960 ;
        RECT 697.690 2968.440 3789.290 2969.840 ;
        RECT 697.690 2962.360 3789.690 2968.440 ;
        RECT 698.090 2960.960 3789.690 2962.360 ;
        RECT 697.690 2909.320 3789.690 2960.960 ;
        RECT 697.690 2907.920 3789.290 2909.320 ;
        RECT 697.690 2849.480 3789.690 2907.920 ;
        RECT 697.690 2848.080 3789.290 2849.480 ;
        RECT 697.690 2826.360 3789.690 2848.080 ;
        RECT 698.090 2824.960 3789.690 2826.360 ;
        RECT 697.690 2788.960 3789.690 2824.960 ;
        RECT 697.690 2787.560 3789.290 2788.960 ;
        RECT 697.690 2728.440 3789.690 2787.560 ;
        RECT 697.690 2727.040 3789.290 2728.440 ;
        RECT 697.690 2690.360 3789.690 2727.040 ;
        RECT 698.090 2688.960 3789.690 2690.360 ;
        RECT 697.690 2668.600 3789.690 2688.960 ;
        RECT 697.690 2667.200 3789.290 2668.600 ;
        RECT 697.690 2608.080 3789.690 2667.200 ;
        RECT 697.690 2606.680 3789.290 2608.080 ;
        RECT 697.690 2555.040 3789.690 2606.680 ;
        RECT 698.090 2553.640 3789.690 2555.040 ;
        RECT 697.690 2547.560 3789.690 2553.640 ;
        RECT 697.690 2546.160 3789.290 2547.560 ;
        RECT 697.690 2487.040 3789.690 2546.160 ;
        RECT 697.690 2485.640 3789.290 2487.040 ;
        RECT 697.690 2427.200 3789.690 2485.640 ;
        RECT 697.690 2425.800 3789.290 2427.200 ;
        RECT 697.690 2419.040 3789.690 2425.800 ;
        RECT 698.090 2417.640 3789.690 2419.040 ;
        RECT 697.690 2366.680 3789.690 2417.640 ;
        RECT 697.690 2365.280 3789.290 2366.680 ;
        RECT 697.690 2306.160 3789.690 2365.280 ;
        RECT 697.690 2304.760 3789.290 2306.160 ;
        RECT 697.690 2283.720 3789.690 2304.760 ;
        RECT 698.090 2282.320 3789.690 2283.720 ;
        RECT 697.690 2246.320 3789.690 2282.320 ;
        RECT 697.690 2244.920 3789.290 2246.320 ;
        RECT 697.690 2185.800 3789.690 2244.920 ;
        RECT 697.690 2184.400 3789.290 2185.800 ;
        RECT 697.690 2147.720 3789.690 2184.400 ;
        RECT 698.090 2146.320 3789.690 2147.720 ;
        RECT 697.690 2125.280 3789.690 2146.320 ;
        RECT 697.690 2123.880 3789.290 2125.280 ;
        RECT 697.690 2065.440 3789.690 2123.880 ;
        RECT 697.690 2064.040 3789.290 2065.440 ;
        RECT 697.690 2012.400 3789.690 2064.040 ;
        RECT 698.090 2011.000 3789.690 2012.400 ;
        RECT 697.690 2004.920 3789.690 2011.000 ;
        RECT 697.690 2003.520 3789.290 2004.920 ;
        RECT 697.690 1944.400 3789.690 2003.520 ;
        RECT 697.690 1943.000 3789.290 1944.400 ;
        RECT 697.690 1883.880 3789.690 1943.000 ;
        RECT 697.690 1882.480 3789.290 1883.880 ;
        RECT 697.690 1876.400 3789.690 1882.480 ;
        RECT 698.090 1875.000 3789.690 1876.400 ;
        RECT 697.690 1824.040 3789.690 1875.000 ;
        RECT 697.690 1822.640 3789.290 1824.040 ;
        RECT 697.690 1763.520 3789.690 1822.640 ;
        RECT 697.690 1762.120 3789.290 1763.520 ;
        RECT 697.690 1740.400 3789.690 1762.120 ;
        RECT 698.090 1739.000 3789.690 1740.400 ;
        RECT 697.690 1703.000 3789.690 1739.000 ;
        RECT 697.690 1701.600 3789.290 1703.000 ;
        RECT 697.690 1643.160 3789.690 1701.600 ;
        RECT 697.690 1641.760 3789.290 1643.160 ;
        RECT 697.690 1605.080 3789.690 1641.760 ;
        RECT 698.090 1603.680 3789.690 1605.080 ;
        RECT 697.690 1582.640 3789.690 1603.680 ;
        RECT 697.690 1581.240 3789.290 1582.640 ;
        RECT 697.690 1522.120 3789.690 1581.240 ;
        RECT 697.690 1520.720 3789.290 1522.120 ;
        RECT 697.690 1469.080 3789.690 1520.720 ;
        RECT 698.090 1467.680 3789.690 1469.080 ;
        RECT 697.690 1462.280 3789.690 1467.680 ;
        RECT 697.690 1460.880 3789.290 1462.280 ;
        RECT 697.690 1401.760 3789.690 1460.880 ;
        RECT 697.690 1400.360 3789.290 1401.760 ;
        RECT 697.690 1341.240 3789.690 1400.360 ;
        RECT 697.690 1339.840 3789.290 1341.240 ;
        RECT 697.690 1333.760 3789.690 1339.840 ;
        RECT 698.090 1332.360 3789.690 1333.760 ;
        RECT 697.690 1280.720 3789.690 1332.360 ;
        RECT 697.690 1279.320 3789.290 1280.720 ;
        RECT 697.690 1220.880 3789.690 1279.320 ;
        RECT 697.690 1219.480 3789.290 1220.880 ;
        RECT 697.690 1197.760 3789.690 1219.480 ;
        RECT 698.090 1196.360 3789.690 1197.760 ;
        RECT 697.690 1160.360 3789.690 1196.360 ;
        RECT 697.690 1158.960 3789.290 1160.360 ;
        RECT 697.690 1099.840 3789.690 1158.960 ;
        RECT 697.690 1098.440 3789.290 1099.840 ;
        RECT 697.690 1062.440 3789.690 1098.440 ;
        RECT 698.090 1061.040 3789.690 1062.440 ;
        RECT 697.690 1040.000 3789.690 1061.040 ;
        RECT 697.690 1038.600 3789.290 1040.000 ;
        RECT 697.690 979.480 3789.690 1038.600 ;
        RECT 697.690 978.080 3789.290 979.480 ;
        RECT 697.690 926.440 3789.690 978.080 ;
        RECT 698.090 925.040 3789.690 926.440 ;
        RECT 697.690 918.960 3789.690 925.040 ;
        RECT 697.690 917.560 3789.290 918.960 ;
        RECT 697.690 859.120 3789.690 917.560 ;
        RECT 697.690 857.720 3789.290 859.120 ;
        RECT 697.690 798.600 3789.690 857.720 ;
        RECT 697.690 797.200 3789.290 798.600 ;
        RECT 697.690 790.440 3789.690 797.200 ;
        RECT 698.090 789.040 3789.690 790.440 ;
        RECT 697.690 738.080 3789.690 789.040 ;
        RECT 697.690 736.680 3789.290 738.080 ;
        RECT 697.690 677.560 3789.690 736.680 ;
        RECT 697.690 676.160 3789.290 677.560 ;
        RECT 697.690 655.120 3789.690 676.160 ;
        RECT 698.090 653.720 3789.690 655.120 ;
        RECT 697.690 617.720 3789.690 653.720 ;
        RECT 697.690 616.320 3789.290 617.720 ;
        RECT 697.690 557.200 3789.690 616.320 ;
        RECT 697.690 555.800 3789.290 557.200 ;
        RECT 697.690 519.120 3789.690 555.800 ;
        RECT 698.090 517.720 3789.690 519.120 ;
        RECT 697.690 496.680 3789.690 517.720 ;
        RECT 697.690 495.280 3789.290 496.680 ;
        RECT 697.690 436.840 3789.690 495.280 ;
        RECT 697.690 435.440 3789.290 436.840 ;
        RECT 697.690 383.800 3789.690 435.440 ;
        RECT 698.090 382.400 3789.690 383.800 ;
        RECT 697.690 376.320 3789.690 382.400 ;
        RECT 697.690 374.920 3789.290 376.320 ;
        RECT 697.690 315.800 3789.690 374.920 ;
        RECT 697.690 314.400 3789.290 315.800 ;
        RECT 697.690 255.960 3789.690 314.400 ;
        RECT 697.690 254.560 3789.290 255.960 ;
        RECT 697.690 247.800 3789.690 254.560 ;
        RECT 698.090 246.400 3789.690 247.800 ;
        RECT 697.690 195.440 3789.690 246.400 ;
        RECT 697.690 194.040 3789.290 195.440 ;
        RECT 697.690 134.920 3789.690 194.040 ;
        RECT 697.690 133.520 3789.290 134.920 ;
        RECT 697.690 112.480 3789.690 133.520 ;
        RECT 698.090 111.080 3789.690 112.480 ;
        RECT 697.690 75.080 3789.690 111.080 ;
        RECT 697.690 73.680 3789.290 75.080 ;
        RECT 697.690 54.835 3789.690 73.680 ;
      LAYER met4 ;
        RECT 644.210 0.000 3843.110 3888.080 ;
      LAYER met5 ;
        RECT 0.005 70.610 3843.110 3888.080 ;
  END
END fpga
END LIBRARY


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2884.510 90.040 2897.690 90.250 ;
        RECT 2881.000 89.950 2897.690 90.040 ;
        RECT 2881.000 89.440 2885.000 89.950 ;
        RECT 2897.390 88.890 2897.690 89.950 ;
        RECT 2897.390 88.590 2898.610 88.890 ;
        RECT 2898.310 88.210 2898.610 88.590 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2898.310 87.910 2924.800 88.210 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1076.010 3444.780 1076.330 3444.840 ;
        RECT 2880.590 3444.780 2880.910 3444.840 ;
        RECT 1076.010 3444.640 2880.910 3444.780 ;
        RECT 1076.010 3444.580 1076.330 3444.640 ;
        RECT 2880.590 3444.580 2880.910 3444.640 ;
        RECT 2880.590 2435.660 2880.910 2435.720 ;
        RECT 2898.070 2435.660 2898.390 2435.720 ;
        RECT 2880.590 2435.520 2898.390 2435.660 ;
        RECT 2880.590 2435.460 2880.910 2435.520 ;
        RECT 2898.070 2435.460 2898.390 2435.520 ;
      LAYER via ;
        RECT 1076.040 3444.580 1076.300 3444.840 ;
        RECT 2880.620 3444.580 2880.880 3444.840 ;
        RECT 2880.620 2435.460 2880.880 2435.720 ;
        RECT 2898.100 2435.460 2898.360 2435.720 ;
      LAYER met2 ;
        RECT 1076.040 3444.550 1076.300 3444.870 ;
        RECT 2880.620 3444.550 2880.880 3444.870 ;
        RECT 1076.100 3435.000 1076.240 3444.550 ;
        RECT 1076.070 3431.000 1076.350 3435.000 ;
        RECT 2880.680 2435.750 2880.820 3444.550 ;
        RECT 2880.620 2435.430 2880.880 2435.750 ;
        RECT 2898.100 2435.430 2898.360 2435.750 ;
        RECT 2898.160 2434.245 2898.300 2435.430 ;
        RECT 2898.090 2433.875 2898.370 2434.245 ;
      LAYER via2 ;
        RECT 2898.090 2433.920 2898.370 2434.200 ;
      LAYER met3 ;
        RECT 2898.065 2434.210 2898.395 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2898.065 2433.910 2924.800 2434.210 ;
        RECT 2898.065 2433.895 2898.395 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 263.650 34.240 263.970 34.300 ;
        RECT 2902.670 34.240 2902.990 34.300 ;
        RECT 263.650 34.100 2902.990 34.240 ;
        RECT 263.650 34.040 263.970 34.100 ;
        RECT 2902.670 34.040 2902.990 34.100 ;
      LAYER via ;
        RECT 263.680 34.040 263.940 34.300 ;
        RECT 2902.700 34.040 2902.960 34.300 ;
      LAYER met2 ;
        RECT 2902.690 2669.155 2902.970 2669.525 ;
        RECT 263.710 35.000 263.990 39.000 ;
        RECT 263.740 34.330 263.880 35.000 ;
        RECT 2902.760 34.330 2902.900 2669.155 ;
        RECT 263.680 34.010 263.940 34.330 ;
        RECT 2902.700 34.010 2902.960 34.330 ;
      LAYER via2 ;
        RECT 2902.690 2669.200 2902.970 2669.480 ;
      LAYER met3 ;
        RECT 2902.665 2669.490 2902.995 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2902.665 2669.190 2924.800 2669.490 ;
        RECT 2902.665 2669.175 2902.995 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 314.710 33.900 315.030 33.960 ;
        RECT 2902.210 33.900 2902.530 33.960 ;
        RECT 314.710 33.760 2902.530 33.900 ;
        RECT 314.710 33.700 315.030 33.760 ;
        RECT 2902.210 33.700 2902.530 33.760 ;
      LAYER via ;
        RECT 314.740 33.700 315.000 33.960 ;
        RECT 2902.240 33.700 2902.500 33.960 ;
      LAYER met2 ;
        RECT 2902.230 2903.755 2902.510 2904.125 ;
        RECT 314.770 35.000 315.050 39.000 ;
        RECT 314.800 33.990 314.940 35.000 ;
        RECT 2902.300 33.990 2902.440 2903.755 ;
        RECT 314.740 33.670 315.000 33.990 ;
        RECT 2902.240 33.670 2902.500 33.990 ;
      LAYER via2 ;
        RECT 2902.230 2903.800 2902.510 2904.080 ;
      LAYER met3 ;
        RECT 2902.205 2904.090 2902.535 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2902.205 2903.790 2924.800 2904.090 ;
        RECT 2902.205 2903.775 2902.535 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 365.310 33.560 365.630 33.620 ;
        RECT 2901.750 33.560 2902.070 33.620 ;
        RECT 365.310 33.420 2902.070 33.560 ;
        RECT 365.310 33.360 365.630 33.420 ;
        RECT 2901.750 33.360 2902.070 33.420 ;
      LAYER via ;
        RECT 365.340 33.360 365.600 33.620 ;
        RECT 2901.780 33.360 2902.040 33.620 ;
      LAYER met2 ;
        RECT 2901.770 3138.355 2902.050 3138.725 ;
        RECT 365.370 35.000 365.650 39.000 ;
        RECT 365.400 33.650 365.540 35.000 ;
        RECT 2901.840 33.650 2901.980 3138.355 ;
        RECT 365.340 33.330 365.600 33.650 ;
        RECT 2901.780 33.330 2902.040 33.650 ;
      LAYER via2 ;
        RECT 2901.770 3138.400 2902.050 3138.680 ;
      LAYER met3 ;
        RECT 2901.745 3138.690 2902.075 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2901.745 3138.390 2924.800 3138.690 ;
        RECT 2901.745 3138.375 2902.075 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 416.370 33.220 416.690 33.280 ;
        RECT 2901.290 33.220 2901.610 33.280 ;
        RECT 416.370 33.080 2901.610 33.220 ;
        RECT 416.370 33.020 416.690 33.080 ;
        RECT 2901.290 33.020 2901.610 33.080 ;
      LAYER via ;
        RECT 416.400 33.020 416.660 33.280 ;
        RECT 2901.320 33.020 2901.580 33.280 ;
      LAYER met2 ;
        RECT 2901.310 3372.955 2901.590 3373.325 ;
        RECT 416.430 35.000 416.710 39.000 ;
        RECT 416.460 33.310 416.600 35.000 ;
        RECT 2901.380 33.310 2901.520 3372.955 ;
        RECT 416.400 32.990 416.660 33.310 ;
        RECT 2901.320 32.990 2901.580 33.310 ;
      LAYER via2 ;
        RECT 2901.310 3373.000 2901.590 3373.280 ;
      LAYER met3 ;
        RECT 2901.285 3373.290 2901.615 3373.305 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2901.285 3372.990 2924.800 3373.290 ;
        RECT 2901.285 3372.975 2901.615 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 96.210 3501.560 96.530 3501.620 ;
        RECT 2798.250 3501.560 2798.570 3501.620 ;
        RECT 96.210 3501.420 2798.570 3501.560 ;
        RECT 96.210 3501.360 96.530 3501.420 ;
        RECT 2798.250 3501.360 2798.570 3501.420 ;
        RECT 89.770 3449.880 90.090 3449.940 ;
        RECT 96.210 3449.880 96.530 3449.940 ;
        RECT 89.770 3449.740 96.530 3449.880 ;
        RECT 89.770 3449.680 90.090 3449.740 ;
        RECT 96.210 3449.680 96.530 3449.740 ;
      LAYER via ;
        RECT 96.240 3501.360 96.500 3501.620 ;
        RECT 2798.280 3501.360 2798.540 3501.620 ;
        RECT 89.800 3449.680 90.060 3449.940 ;
        RECT 96.240 3449.680 96.500 3449.940 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3501.650 2798.480 3517.600 ;
        RECT 96.240 3501.330 96.500 3501.650 ;
        RECT 2798.280 3501.330 2798.540 3501.650 ;
        RECT 96.300 3449.970 96.440 3501.330 ;
        RECT 89.800 3449.650 90.060 3449.970 ;
        RECT 96.240 3449.650 96.500 3449.970 ;
        RECT 89.860 3435.000 90.000 3449.650 ;
        RECT 89.830 3431.000 90.110 3435.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 199.710 3501.900 200.030 3501.960 ;
        RECT 2473.950 3501.900 2474.270 3501.960 ;
        RECT 199.710 3501.760 2474.270 3501.900 ;
        RECT 199.710 3501.700 200.030 3501.760 ;
        RECT 2473.950 3501.700 2474.270 3501.760 ;
      LAYER via ;
        RECT 199.740 3501.700 200.000 3501.960 ;
        RECT 2473.980 3501.700 2474.240 3501.960 ;
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3501.990 2474.180 3517.600 ;
        RECT 199.740 3501.670 200.000 3501.990 ;
        RECT 2473.980 3501.670 2474.240 3501.990 ;
        RECT 199.310 3434.410 199.590 3435.000 ;
        RECT 199.800 3434.410 199.940 3501.670 ;
        RECT 199.310 3434.270 199.940 3434.410 ;
        RECT 199.310 3431.000 199.590 3434.270 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 310.110 3502.240 310.430 3502.300 ;
        RECT 2149.190 3502.240 2149.510 3502.300 ;
        RECT 310.110 3502.100 2149.510 3502.240 ;
        RECT 310.110 3502.040 310.430 3502.100 ;
        RECT 2149.190 3502.040 2149.510 3502.100 ;
      LAYER via ;
        RECT 310.140 3502.040 310.400 3502.300 ;
        RECT 2149.220 3502.040 2149.480 3502.300 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3502.330 2149.420 3517.600 ;
        RECT 310.140 3502.010 310.400 3502.330 ;
        RECT 2149.220 3502.010 2149.480 3502.330 ;
        RECT 308.790 3434.410 309.070 3435.000 ;
        RECT 310.200 3434.410 310.340 3502.010 ;
        RECT 308.790 3434.270 310.340 3434.410 ;
        RECT 308.790 3431.000 309.070 3434.270 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 420.510 3502.580 420.830 3502.640 ;
        RECT 1824.890 3502.580 1825.210 3502.640 ;
        RECT 420.510 3502.440 1825.210 3502.580 ;
        RECT 420.510 3502.380 420.830 3502.440 ;
        RECT 1824.890 3502.380 1825.210 3502.440 ;
      LAYER via ;
        RECT 420.540 3502.380 420.800 3502.640 ;
        RECT 1824.920 3502.380 1825.180 3502.640 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3502.670 1825.120 3517.600 ;
        RECT 420.540 3502.350 420.800 3502.670 ;
        RECT 1824.920 3502.350 1825.180 3502.670 ;
        RECT 418.270 3434.410 418.550 3435.000 ;
        RECT 420.600 3434.410 420.740 3502.350 ;
        RECT 418.270 3434.270 420.740 3434.410 ;
        RECT 418.270 3431.000 418.550 3434.270 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 530.910 3502.920 531.230 3502.980 ;
        RECT 1500.590 3502.920 1500.910 3502.980 ;
        RECT 530.910 3502.780 1500.910 3502.920 ;
        RECT 530.910 3502.720 531.230 3502.780 ;
        RECT 1500.590 3502.720 1500.910 3502.780 ;
      LAYER via ;
        RECT 530.940 3502.720 531.200 3502.980 ;
        RECT 1500.620 3502.720 1500.880 3502.980 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3503.010 1500.820 3517.600 ;
        RECT 530.940 3502.690 531.200 3503.010 ;
        RECT 1500.620 3502.690 1500.880 3503.010 ;
        RECT 531.000 3435.090 531.140 3502.690 ;
        RECT 528.210 3434.410 528.490 3435.000 ;
        RECT 529.620 3434.950 531.140 3435.090 ;
        RECT 529.620 3434.410 529.760 3434.950 ;
        RECT 528.210 3434.270 529.760 3434.410 ;
        RECT 528.210 3431.000 528.490 3434.270 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2895.310 199.820 2895.630 199.880 ;
        RECT 2903.130 199.820 2903.450 199.880 ;
        RECT 2895.310 199.680 2903.450 199.820 ;
        RECT 2895.310 199.620 2895.630 199.680 ;
        RECT 2903.130 199.620 2903.450 199.680 ;
      LAYER via ;
        RECT 2895.340 199.620 2895.600 199.880 ;
        RECT 2903.160 199.620 2903.420 199.880 ;
      LAYER met2 ;
        RECT 2903.150 322.475 2903.430 322.845 ;
        RECT 2903.220 199.910 2903.360 322.475 ;
        RECT 2895.340 199.765 2895.600 199.910 ;
        RECT 2895.330 199.395 2895.610 199.765 ;
        RECT 2903.160 199.590 2903.420 199.910 ;
      LAYER via2 ;
        RECT 2903.150 322.520 2903.430 322.800 ;
        RECT 2895.330 199.440 2895.610 199.720 ;
      LAYER met3 ;
        RECT 2903.125 322.810 2903.455 322.825 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2903.125 322.510 2924.800 322.810 ;
        RECT 2903.125 322.495 2903.455 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
        RECT 2895.305 199.730 2895.635 199.745 ;
        RECT 2884.510 199.520 2895.635 199.730 ;
        RECT 2881.000 199.430 2895.635 199.520 ;
        RECT 2881.000 198.920 2885.000 199.430 ;
        RECT 2895.305 199.415 2895.635 199.430 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 641.310 3503.260 641.630 3503.320 ;
        RECT 1175.830 3503.260 1176.150 3503.320 ;
        RECT 641.310 3503.120 1176.150 3503.260 ;
        RECT 641.310 3503.060 641.630 3503.120 ;
        RECT 1175.830 3503.060 1176.150 3503.120 ;
        RECT 637.630 3447.840 637.950 3447.900 ;
        RECT 641.310 3447.840 641.630 3447.900 ;
        RECT 637.630 3447.700 641.630 3447.840 ;
        RECT 637.630 3447.640 637.950 3447.700 ;
        RECT 641.310 3447.640 641.630 3447.700 ;
      LAYER via ;
        RECT 641.340 3503.060 641.600 3503.320 ;
        RECT 1175.860 3503.060 1176.120 3503.320 ;
        RECT 637.660 3447.640 637.920 3447.900 ;
        RECT 641.340 3447.640 641.600 3447.900 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3503.350 1176.060 3517.600 ;
        RECT 641.340 3503.030 641.600 3503.350 ;
        RECT 1175.860 3503.030 1176.120 3503.350 ;
        RECT 641.400 3447.930 641.540 3503.030 ;
        RECT 637.660 3447.610 637.920 3447.930 ;
        RECT 641.340 3447.610 641.600 3447.930 ;
        RECT 637.720 3435.000 637.860 3447.610 ;
        RECT 637.690 3431.000 637.970 3435.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 751.710 3503.600 752.030 3503.660 ;
        RECT 851.530 3503.600 851.850 3503.660 ;
        RECT 751.710 3503.460 851.850 3503.600 ;
        RECT 751.710 3503.400 752.030 3503.460 ;
        RECT 851.530 3503.400 851.850 3503.460 ;
        RECT 747.110 3447.840 747.430 3447.900 ;
        RECT 751.710 3447.840 752.030 3447.900 ;
        RECT 747.110 3447.700 752.030 3447.840 ;
        RECT 747.110 3447.640 747.430 3447.700 ;
        RECT 751.710 3447.640 752.030 3447.700 ;
      LAYER via ;
        RECT 751.740 3503.400 752.000 3503.660 ;
        RECT 851.560 3503.400 851.820 3503.660 ;
        RECT 747.140 3447.640 747.400 3447.900 ;
        RECT 751.740 3447.640 752.000 3447.900 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3503.690 851.760 3517.600 ;
        RECT 751.740 3503.370 752.000 3503.690 ;
        RECT 851.560 3503.370 851.820 3503.690 ;
        RECT 751.800 3447.930 751.940 3503.370 ;
        RECT 747.140 3447.610 747.400 3447.930 ;
        RECT 751.740 3447.610 752.000 3447.930 ;
        RECT 747.200 3435.000 747.340 3447.610 ;
        RECT 747.170 3431.000 747.450 3435.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 527.230 3498.500 527.550 3498.560 ;
        RECT 530.450 3498.500 530.770 3498.560 ;
        RECT 527.230 3498.360 530.770 3498.500 ;
        RECT 527.230 3498.300 527.550 3498.360 ;
        RECT 530.450 3498.300 530.770 3498.360 ;
        RECT 530.450 3446.820 530.770 3446.880 ;
        RECT 857.050 3446.820 857.370 3446.880 ;
        RECT 530.450 3446.680 857.370 3446.820 ;
        RECT 530.450 3446.620 530.770 3446.680 ;
        RECT 857.050 3446.620 857.370 3446.680 ;
      LAYER via ;
        RECT 527.260 3498.300 527.520 3498.560 ;
        RECT 530.480 3498.300 530.740 3498.560 ;
        RECT 530.480 3446.620 530.740 3446.880 ;
        RECT 857.080 3446.620 857.340 3446.880 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3498.590 527.460 3517.600 ;
        RECT 527.260 3498.270 527.520 3498.590 ;
        RECT 530.480 3498.270 530.740 3498.590 ;
        RECT 530.540 3446.910 530.680 3498.270 ;
        RECT 530.480 3446.590 530.740 3446.910 ;
        RECT 857.080 3446.590 857.340 3446.910 ;
        RECT 857.140 3435.000 857.280 3446.590 ;
        RECT 857.110 3431.000 857.390 3435.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 202.470 3502.240 202.790 3502.300 ;
        RECT 206.610 3502.240 206.930 3502.300 ;
        RECT 202.470 3502.100 206.930 3502.240 ;
        RECT 202.470 3502.040 202.790 3502.100 ;
        RECT 206.610 3502.040 206.930 3502.100 ;
        RECT 206.610 3446.480 206.930 3446.540 ;
        RECT 966.530 3446.480 966.850 3446.540 ;
        RECT 206.610 3446.340 966.850 3446.480 ;
        RECT 206.610 3446.280 206.930 3446.340 ;
        RECT 966.530 3446.280 966.850 3446.340 ;
      LAYER via ;
        RECT 202.500 3502.040 202.760 3502.300 ;
        RECT 206.640 3502.040 206.900 3502.300 ;
        RECT 206.640 3446.280 206.900 3446.540 ;
        RECT 966.560 3446.280 966.820 3446.540 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3502.330 202.700 3517.600 ;
        RECT 202.500 3502.010 202.760 3502.330 ;
        RECT 206.640 3502.010 206.900 3502.330 ;
        RECT 206.700 3446.570 206.840 3502.010 ;
        RECT 206.640 3446.250 206.900 3446.570 ;
        RECT 966.560 3446.250 966.820 3446.570 ;
        RECT 966.620 3435.000 966.760 3446.250 ;
        RECT 966.590 3431.000 966.870 3435.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.630 3408.740 16.950 3408.800 ;
        RECT 30.890 3408.740 31.210 3408.800 ;
        RECT 16.630 3408.600 31.210 3408.740 ;
        RECT 16.630 3408.540 16.950 3408.600 ;
        RECT 30.890 3408.540 31.210 3408.600 ;
        RECT 30.890 27.440 31.210 27.500 ;
        RECT 60.330 27.440 60.650 27.500 ;
        RECT 30.890 27.300 60.650 27.440 ;
        RECT 30.890 27.240 31.210 27.300 ;
        RECT 60.330 27.240 60.650 27.300 ;
      LAYER via ;
        RECT 16.660 3408.540 16.920 3408.800 ;
        RECT 30.920 3408.540 31.180 3408.800 ;
        RECT 30.920 27.240 31.180 27.500 ;
        RECT 60.360 27.240 60.620 27.500 ;
      LAYER met2 ;
        RECT 16.650 3411.035 16.930 3411.405 ;
        RECT 16.720 3408.830 16.860 3411.035 ;
        RECT 16.660 3408.510 16.920 3408.830 ;
        RECT 30.920 3408.510 31.180 3408.830 ;
        RECT 30.980 27.530 31.120 3408.510 ;
        RECT 60.390 35.000 60.670 39.000 ;
        RECT 60.420 27.530 60.560 35.000 ;
        RECT 30.920 27.210 31.180 27.530 ;
        RECT 60.360 27.210 60.620 27.530 ;
      LAYER via2 ;
        RECT 16.650 3411.080 16.930 3411.360 ;
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 16.625 3411.370 16.955 3411.385 ;
        RECT -4.800 3411.070 16.955 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 16.625 3411.055 16.955 3411.070 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 15.710 3121.100 16.030 3121.160 ;
        RECT 31.350 3121.100 31.670 3121.160 ;
        RECT 15.710 3120.960 31.670 3121.100 ;
        RECT 15.710 3120.900 16.030 3120.960 ;
        RECT 31.350 3120.900 31.670 3120.960 ;
        RECT 31.350 23.700 31.670 23.760 ;
        RECT 110.930 23.700 111.250 23.760 ;
        RECT 31.350 23.560 111.250 23.700 ;
        RECT 31.350 23.500 31.670 23.560 ;
        RECT 110.930 23.500 111.250 23.560 ;
      LAYER via ;
        RECT 15.740 3120.900 16.000 3121.160 ;
        RECT 31.380 3120.900 31.640 3121.160 ;
        RECT 31.380 23.500 31.640 23.760 ;
        RECT 110.960 23.500 111.220 23.760 ;
      LAYER met2 ;
        RECT 15.730 3124.075 16.010 3124.445 ;
        RECT 15.800 3121.190 15.940 3124.075 ;
        RECT 15.740 3120.870 16.000 3121.190 ;
        RECT 31.380 3120.870 31.640 3121.190 ;
        RECT 31.440 23.790 31.580 3120.870 ;
        RECT 110.990 35.000 111.270 39.000 ;
        RECT 111.020 23.790 111.160 35.000 ;
        RECT 31.380 23.470 31.640 23.790 ;
        RECT 110.960 23.470 111.220 23.790 ;
      LAYER via2 ;
        RECT 15.730 3124.120 16.010 3124.400 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 15.705 3124.410 16.035 3124.425 ;
        RECT -4.800 3124.110 16.035 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 15.705 3124.095 16.035 3124.110 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 20.310 2836.520 20.630 2836.580 ;
        RECT 37.790 2836.520 38.110 2836.580 ;
        RECT 20.310 2836.380 38.110 2836.520 ;
        RECT 20.310 2836.320 20.630 2836.380 ;
        RECT 37.790 2836.320 38.110 2836.380 ;
        RECT 37.790 27.100 38.110 27.160 ;
        RECT 161.990 27.100 162.310 27.160 ;
        RECT 37.790 26.960 162.310 27.100 ;
        RECT 37.790 26.900 38.110 26.960 ;
        RECT 161.990 26.900 162.310 26.960 ;
      LAYER via ;
        RECT 20.340 2836.320 20.600 2836.580 ;
        RECT 37.820 2836.320 38.080 2836.580 ;
        RECT 37.820 26.900 38.080 27.160 ;
        RECT 162.020 26.900 162.280 27.160 ;
      LAYER met2 ;
        RECT 20.330 2836.435 20.610 2836.805 ;
        RECT 20.340 2836.290 20.600 2836.435 ;
        RECT 37.820 2836.290 38.080 2836.610 ;
        RECT 37.880 27.190 38.020 2836.290 ;
        RECT 162.050 35.000 162.330 39.000 ;
        RECT 162.080 27.190 162.220 35.000 ;
        RECT 37.820 26.870 38.080 27.190 ;
        RECT 162.020 26.870 162.280 27.190 ;
      LAYER via2 ;
        RECT 20.330 2836.480 20.610 2836.760 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 20.305 2836.770 20.635 2836.785 ;
        RECT -4.800 2836.470 20.635 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 20.305 2836.455 20.635 2836.470 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 25.740 17.410 25.800 ;
        RECT 212.590 25.740 212.910 25.800 ;
        RECT 17.090 25.600 212.910 25.740 ;
        RECT 17.090 25.540 17.410 25.600 ;
        RECT 212.590 25.540 212.910 25.600 ;
      LAYER via ;
        RECT 17.120 25.540 17.380 25.800 ;
        RECT 212.620 25.540 212.880 25.800 ;
      LAYER met2 ;
        RECT 17.110 2549.475 17.390 2549.845 ;
        RECT 17.180 25.830 17.320 2549.475 ;
        RECT 212.650 35.000 212.930 39.000 ;
        RECT 212.680 25.830 212.820 35.000 ;
        RECT 17.120 25.510 17.380 25.830 ;
        RECT 212.620 25.510 212.880 25.830 ;
      LAYER via2 ;
        RECT 17.110 2549.520 17.390 2549.800 ;
      LAYER met3 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 17.085 2549.810 17.415 2549.825 ;
        RECT -4.800 2549.510 17.415 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 17.085 2549.495 17.415 2549.510 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.570 2261.835 17.850 2262.205 ;
        RECT 17.640 93.005 17.780 2261.835 ;
        RECT 17.570 92.635 17.850 93.005 ;
      LAYER via2 ;
        RECT 17.570 2261.880 17.850 2262.160 ;
        RECT 17.570 92.680 17.850 92.960 ;
      LAYER met3 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 17.545 2262.170 17.875 2262.185 ;
        RECT -4.800 2261.870 17.875 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 17.545 2261.855 17.875 2261.870 ;
        RECT 17.545 92.970 17.875 92.985 ;
        RECT 17.545 92.670 35.570 92.970 ;
        RECT 17.545 92.655 17.875 92.670 ;
        RECT 35.270 90.040 35.570 92.670 ;
        RECT 35.000 89.440 39.000 90.040 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.030 1974.875 18.310 1975.245 ;
        RECT 18.100 199.765 18.240 1974.875 ;
        RECT 18.030 199.395 18.310 199.765 ;
      LAYER via2 ;
        RECT 18.030 1974.920 18.310 1975.200 ;
        RECT 18.030 199.440 18.310 199.720 ;
      LAYER met3 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 18.005 1975.210 18.335 1975.225 ;
        RECT -4.800 1974.910 18.335 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 18.005 1974.895 18.335 1974.910 ;
        RECT 18.005 199.730 18.335 199.745 ;
        RECT 18.005 199.520 35.570 199.730 ;
        RECT 18.005 199.430 39.000 199.520 ;
        RECT 18.005 199.415 18.335 199.430 ;
        RECT 35.000 198.920 39.000 199.430 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2895.310 309.980 2895.630 310.040 ;
        RECT 2904.050 309.980 2904.370 310.040 ;
        RECT 2895.310 309.840 2904.370 309.980 ;
        RECT 2895.310 309.780 2895.630 309.840 ;
        RECT 2904.050 309.780 2904.370 309.840 ;
      LAYER via ;
        RECT 2895.340 309.780 2895.600 310.040 ;
        RECT 2904.080 309.780 2904.340 310.040 ;
      LAYER met2 ;
        RECT 2904.070 557.075 2904.350 557.445 ;
        RECT 2904.140 310.070 2904.280 557.075 ;
        RECT 2895.340 309.925 2895.600 310.070 ;
        RECT 2895.330 309.555 2895.610 309.925 ;
        RECT 2904.080 309.750 2904.340 310.070 ;
      LAYER via2 ;
        RECT 2904.070 557.120 2904.350 557.400 ;
        RECT 2895.330 309.600 2895.610 309.880 ;
      LAYER met3 ;
        RECT 2904.045 557.410 2904.375 557.425 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2904.045 557.110 2924.800 557.410 ;
        RECT 2904.045 557.095 2904.375 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
        RECT 2895.305 309.890 2895.635 309.905 ;
        RECT 2884.510 309.590 2895.635 309.890 ;
        RECT 2884.510 309.000 2884.810 309.590 ;
        RECT 2895.305 309.575 2895.635 309.590 ;
        RECT 2881.000 308.400 2885.000 309.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 1687.235 18.770 1687.605 ;
        RECT 18.560 310.605 18.700 1687.235 ;
        RECT 18.490 310.235 18.770 310.605 ;
      LAYER via2 ;
        RECT 18.490 1687.280 18.770 1687.560 ;
        RECT 18.490 310.280 18.770 310.560 ;
      LAYER met3 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 18.465 1687.570 18.795 1687.585 ;
        RECT -4.800 1687.270 18.795 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
        RECT 18.465 1687.255 18.795 1687.270 ;
        RECT 18.465 310.570 18.795 310.585 ;
        RECT 18.465 310.270 35.570 310.570 ;
        RECT 18.465 310.255 18.795 310.270 ;
        RECT 35.270 309.000 35.570 310.270 ;
        RECT 35.000 308.400 39.000 309.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.950 1471.675 19.230 1472.045 ;
        RECT 19.020 420.765 19.160 1471.675 ;
        RECT 18.950 420.395 19.230 420.765 ;
      LAYER via2 ;
        RECT 18.950 1471.720 19.230 1472.000 ;
        RECT 18.950 420.440 19.230 420.720 ;
      LAYER met3 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 18.925 1472.010 19.255 1472.025 ;
        RECT -4.800 1471.710 19.255 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 18.925 1471.695 19.255 1471.710 ;
        RECT 18.925 420.730 19.255 420.745 ;
        RECT 18.925 420.430 35.570 420.730 ;
        RECT 18.925 420.415 19.255 420.430 ;
        RECT 35.270 418.480 35.570 420.430 ;
        RECT 35.000 417.880 39.000 418.480 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.870 1256.115 20.150 1256.485 ;
        RECT 19.940 530.245 20.080 1256.115 ;
        RECT 19.870 529.875 20.150 530.245 ;
      LAYER via2 ;
        RECT 19.870 1256.160 20.150 1256.440 ;
        RECT 19.870 529.920 20.150 530.200 ;
      LAYER met3 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 19.845 1256.450 20.175 1256.465 ;
        RECT -4.800 1256.150 20.175 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 19.845 1256.135 20.175 1256.150 ;
        RECT 19.845 530.210 20.175 530.225 ;
        RECT 19.845 529.910 35.570 530.210 ;
        RECT 19.845 529.895 20.175 529.910 ;
        RECT 35.270 528.640 35.570 529.910 ;
        RECT 35.000 528.040 39.000 528.640 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.630 641.480 16.950 641.540 ;
        RECT 20.770 641.480 21.090 641.540 ;
        RECT 16.630 641.340 21.090 641.480 ;
        RECT 16.630 641.280 16.950 641.340 ;
        RECT 20.770 641.280 21.090 641.340 ;
      LAYER via ;
        RECT 16.660 641.280 16.920 641.540 ;
        RECT 20.800 641.280 21.060 641.540 ;
      LAYER met2 ;
        RECT 16.650 1040.555 16.930 1040.925 ;
        RECT 16.720 641.570 16.860 1040.555 ;
        RECT 16.660 641.250 16.920 641.570 ;
        RECT 20.800 641.250 21.060 641.570 ;
        RECT 20.860 641.085 21.000 641.250 ;
        RECT 20.790 640.715 21.070 641.085 ;
      LAYER via2 ;
        RECT 16.650 1040.600 16.930 1040.880 ;
        RECT 20.790 640.760 21.070 641.040 ;
      LAYER met3 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 16.625 1040.890 16.955 1040.905 ;
        RECT -4.800 1040.590 16.955 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
        RECT 16.625 1040.575 16.955 1040.590 ;
        RECT 20.765 641.050 21.095 641.065 ;
        RECT 20.765 640.750 35.570 641.050 ;
        RECT 20.765 640.735 21.095 640.750 ;
        RECT 35.270 638.120 35.570 640.750 ;
        RECT 35.000 637.520 39.000 638.120 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.550 824.995 23.830 825.365 ;
        RECT 23.620 750.565 23.760 824.995 ;
        RECT 23.550 750.195 23.830 750.565 ;
      LAYER via2 ;
        RECT 23.550 825.040 23.830 825.320 ;
        RECT 23.550 750.240 23.830 750.520 ;
      LAYER met3 ;
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 23.525 825.330 23.855 825.345 ;
        RECT -4.800 825.030 23.855 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
        RECT 23.525 825.015 23.855 825.030 ;
        RECT 23.525 750.530 23.855 750.545 ;
        RECT 23.525 750.230 35.570 750.530 ;
        RECT 23.525 750.215 23.855 750.230 ;
        RECT 35.270 747.600 35.570 750.230 ;
        RECT 35.000 747.000 39.000 747.600 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.170 855.680 16.490 855.740 ;
        RECT 23.530 855.680 23.850 855.740 ;
        RECT 16.170 855.540 23.850 855.680 ;
        RECT 16.170 855.480 16.490 855.540 ;
        RECT 23.530 855.480 23.850 855.540 ;
      LAYER via ;
        RECT 16.200 855.480 16.460 855.740 ;
        RECT 23.560 855.480 23.820 855.740 ;
      LAYER met2 ;
        RECT 16.200 855.450 16.460 855.770 ;
        RECT 23.550 855.595 23.830 855.965 ;
        RECT 23.560 855.450 23.820 855.595 ;
        RECT 16.260 610.485 16.400 855.450 ;
        RECT 16.190 610.115 16.470 610.485 ;
      LAYER via2 ;
        RECT 23.550 855.640 23.830 855.920 ;
        RECT 16.190 610.160 16.470 610.440 ;
      LAYER met3 ;
        RECT 35.000 857.160 39.000 857.760 ;
        RECT 23.525 855.930 23.855 855.945 ;
        RECT 35.270 855.930 35.570 857.160 ;
        RECT 23.525 855.630 35.570 855.930 ;
        RECT 23.525 855.615 23.855 855.630 ;
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 16.165 610.450 16.495 610.465 ;
        RECT -4.800 610.150 16.495 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 16.165 610.135 16.495 610.150 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.330 966.435 20.610 966.805 ;
        RECT 20.400 394.925 20.540 966.435 ;
        RECT 20.330 394.555 20.610 394.925 ;
      LAYER via2 ;
        RECT 20.330 966.480 20.610 966.760 ;
        RECT 20.330 394.600 20.610 394.880 ;
      LAYER met3 ;
        RECT 20.305 966.770 20.635 966.785 ;
        RECT 35.000 966.770 39.000 967.240 ;
        RECT 20.305 966.640 39.000 966.770 ;
        RECT 20.305 966.470 35.570 966.640 ;
        RECT 20.305 966.455 20.635 966.470 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 20.305 394.890 20.635 394.905 ;
        RECT -4.800 394.590 20.635 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 20.305 394.575 20.635 394.590 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.410 1076.595 19.690 1076.965 ;
        RECT 19.480 179.365 19.620 1076.595 ;
        RECT 19.410 178.995 19.690 179.365 ;
      LAYER via2 ;
        RECT 19.410 1076.640 19.690 1076.920 ;
        RECT 19.410 179.040 19.690 179.320 ;
      LAYER met3 ;
        RECT 19.385 1076.930 19.715 1076.945 ;
        RECT 19.385 1076.720 35.570 1076.930 ;
        RECT 19.385 1076.630 39.000 1076.720 ;
        RECT 19.385 1076.615 19.715 1076.630 ;
        RECT 35.000 1076.120 39.000 1076.630 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 19.385 179.330 19.715 179.345 ;
        RECT -4.800 179.030 19.715 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 19.385 179.015 19.715 179.030 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2895.310 420.820 2895.630 420.880 ;
        RECT 2903.590 420.820 2903.910 420.880 ;
        RECT 2895.310 420.680 2903.910 420.820 ;
        RECT 2895.310 420.620 2895.630 420.680 ;
        RECT 2903.590 420.620 2903.910 420.680 ;
      LAYER via ;
        RECT 2895.340 420.620 2895.600 420.880 ;
        RECT 2903.620 420.620 2903.880 420.880 ;
      LAYER met2 ;
        RECT 2903.610 791.675 2903.890 792.045 ;
        RECT 2903.680 420.910 2903.820 791.675 ;
        RECT 2895.340 420.765 2895.600 420.910 ;
        RECT 2895.330 420.395 2895.610 420.765 ;
        RECT 2903.620 420.590 2903.880 420.910 ;
      LAYER via2 ;
        RECT 2903.610 791.720 2903.890 792.000 ;
        RECT 2895.330 420.440 2895.610 420.720 ;
      LAYER met3 ;
        RECT 2903.585 792.010 2903.915 792.025 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2903.585 791.710 2924.800 792.010 ;
        RECT 2903.585 791.695 2903.915 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
        RECT 2895.305 420.730 2895.635 420.745 ;
        RECT 2884.510 420.430 2895.635 420.730 ;
        RECT 2884.510 418.480 2884.810 420.430 ;
        RECT 2895.305 420.415 2895.635 420.430 ;
        RECT 2881.000 417.880 2885.000 418.480 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2895.310 530.980 2895.630 531.040 ;
        RECT 2903.130 530.980 2903.450 531.040 ;
        RECT 2895.310 530.840 2903.450 530.980 ;
        RECT 2895.310 530.780 2895.630 530.840 ;
        RECT 2903.130 530.780 2903.450 530.840 ;
      LAYER via ;
        RECT 2895.340 530.780 2895.600 531.040 ;
        RECT 2903.160 530.780 2903.420 531.040 ;
      LAYER met2 ;
        RECT 2903.150 1026.275 2903.430 1026.645 ;
        RECT 2903.220 531.070 2903.360 1026.275 ;
        RECT 2895.340 530.925 2895.600 531.070 ;
        RECT 2895.330 530.555 2895.610 530.925 ;
        RECT 2903.160 530.750 2903.420 531.070 ;
      LAYER via2 ;
        RECT 2903.150 1026.320 2903.430 1026.600 ;
        RECT 2895.330 530.600 2895.610 530.880 ;
      LAYER met3 ;
        RECT 2903.125 1026.610 2903.455 1026.625 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2903.125 1026.310 2924.800 1026.610 ;
        RECT 2903.125 1026.295 2903.455 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
        RECT 2895.305 530.890 2895.635 530.905 ;
        RECT 2884.510 530.590 2895.635 530.890 ;
        RECT 2884.510 528.640 2884.810 530.590 ;
        RECT 2895.305 530.575 2895.635 530.590 ;
        RECT 2881.000 528.040 2885.000 528.640 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2895.310 639.780 2895.630 639.840 ;
        RECT 2900.830 639.780 2901.150 639.840 ;
        RECT 2895.310 639.640 2901.150 639.780 ;
        RECT 2895.310 639.580 2895.630 639.640 ;
        RECT 2900.830 639.580 2901.150 639.640 ;
      LAYER via ;
        RECT 2895.340 639.580 2895.600 639.840 ;
        RECT 2900.860 639.580 2901.120 639.840 ;
      LAYER met2 ;
        RECT 2900.850 1260.875 2901.130 1261.245 ;
        RECT 2900.920 639.870 2901.060 1260.875 ;
        RECT 2895.340 639.725 2895.600 639.870 ;
        RECT 2895.330 639.355 2895.610 639.725 ;
        RECT 2900.860 639.550 2901.120 639.870 ;
      LAYER via2 ;
        RECT 2900.850 1260.920 2901.130 1261.200 ;
        RECT 2895.330 639.400 2895.610 639.680 ;
      LAYER met3 ;
        RECT 2900.825 1261.210 2901.155 1261.225 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2900.825 1260.910 2924.800 1261.210 ;
        RECT 2900.825 1260.895 2901.155 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
        RECT 2895.305 639.690 2895.635 639.705 ;
        RECT 2884.510 639.390 2895.635 639.690 ;
        RECT 2884.510 638.120 2884.810 639.390 ;
        RECT 2895.305 639.375 2895.635 639.390 ;
        RECT 2881.000 637.520 2885.000 638.120 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2895.310 750.620 2895.630 750.680 ;
        RECT 2904.510 750.620 2904.830 750.680 ;
        RECT 2895.310 750.480 2904.830 750.620 ;
        RECT 2895.310 750.420 2895.630 750.480 ;
        RECT 2904.510 750.420 2904.830 750.480 ;
      LAYER via ;
        RECT 2895.340 750.420 2895.600 750.680 ;
        RECT 2904.540 750.420 2904.800 750.680 ;
      LAYER met2 ;
        RECT 2904.530 1495.475 2904.810 1495.845 ;
        RECT 2904.600 750.710 2904.740 1495.475 ;
        RECT 2895.340 750.565 2895.600 750.710 ;
        RECT 2895.330 750.195 2895.610 750.565 ;
        RECT 2904.540 750.390 2904.800 750.710 ;
      LAYER via2 ;
        RECT 2904.530 1495.520 2904.810 1495.800 ;
        RECT 2895.330 750.240 2895.610 750.520 ;
      LAYER met3 ;
        RECT 2904.505 1495.810 2904.835 1495.825 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2904.505 1495.510 2924.800 1495.810 ;
        RECT 2904.505 1495.495 2904.835 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
        RECT 2895.305 750.530 2895.635 750.545 ;
        RECT 2884.510 750.230 2895.635 750.530 ;
        RECT 2884.510 747.600 2884.810 750.230 ;
        RECT 2895.305 750.215 2895.635 750.230 ;
        RECT 2881.000 747.000 2885.000 747.600 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2895.310 860.780 2895.630 860.840 ;
        RECT 2904.050 860.780 2904.370 860.840 ;
        RECT 2895.310 860.640 2904.370 860.780 ;
        RECT 2895.310 860.580 2895.630 860.640 ;
        RECT 2904.050 860.580 2904.370 860.640 ;
      LAYER via ;
        RECT 2895.340 860.580 2895.600 860.840 ;
        RECT 2904.080 860.580 2904.340 860.840 ;
      LAYER met2 ;
        RECT 2904.070 1730.075 2904.350 1730.445 ;
        RECT 2904.140 860.870 2904.280 1730.075 ;
        RECT 2895.340 860.725 2895.600 860.870 ;
        RECT 2895.330 860.355 2895.610 860.725 ;
        RECT 2904.080 860.550 2904.340 860.870 ;
      LAYER via2 ;
        RECT 2904.070 1730.120 2904.350 1730.400 ;
        RECT 2895.330 860.400 2895.610 860.680 ;
      LAYER met3 ;
        RECT 2904.045 1730.410 2904.375 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2904.045 1730.110 2924.800 1730.410 ;
        RECT 2904.045 1730.095 2904.375 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
        RECT 2895.305 860.690 2895.635 860.705 ;
        RECT 2884.510 860.390 2895.635 860.690 ;
        RECT 2884.510 857.760 2884.810 860.390 ;
        RECT 2895.305 860.375 2895.635 860.390 ;
        RECT 2881.000 857.160 2885.000 857.760 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2895.310 970.260 2895.630 970.320 ;
        RECT 2903.590 970.260 2903.910 970.320 ;
        RECT 2895.310 970.120 2903.910 970.260 ;
        RECT 2895.310 970.060 2895.630 970.120 ;
        RECT 2903.590 970.060 2903.910 970.120 ;
      LAYER via ;
        RECT 2895.340 970.060 2895.600 970.320 ;
        RECT 2903.620 970.060 2903.880 970.320 ;
      LAYER met2 ;
        RECT 2903.610 1964.675 2903.890 1965.045 ;
        RECT 2903.680 970.350 2903.820 1964.675 ;
        RECT 2895.340 970.205 2895.600 970.350 ;
        RECT 2895.330 969.835 2895.610 970.205 ;
        RECT 2903.620 970.030 2903.880 970.350 ;
      LAYER via2 ;
        RECT 2903.610 1964.720 2903.890 1965.000 ;
        RECT 2895.330 969.880 2895.610 970.160 ;
      LAYER met3 ;
        RECT 2903.585 1965.010 2903.915 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2903.585 1964.710 2924.800 1965.010 ;
        RECT 2903.585 1964.695 2903.915 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
        RECT 2895.305 970.170 2895.635 970.185 ;
        RECT 2884.510 969.870 2895.635 970.170 ;
        RECT 2884.510 967.240 2884.810 969.870 ;
        RECT 2895.305 969.855 2895.635 969.870 ;
        RECT 2881.000 966.640 2885.000 967.240 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2895.310 1081.780 2895.630 1081.840 ;
        RECT 2903.130 1081.780 2903.450 1081.840 ;
        RECT 2895.310 1081.640 2903.450 1081.780 ;
        RECT 2895.310 1081.580 2895.630 1081.640 ;
        RECT 2903.130 1081.580 2903.450 1081.640 ;
      LAYER via ;
        RECT 2895.340 1081.580 2895.600 1081.840 ;
        RECT 2903.160 1081.580 2903.420 1081.840 ;
      LAYER met2 ;
        RECT 2903.150 2199.275 2903.430 2199.645 ;
        RECT 2903.220 1081.870 2903.360 2199.275 ;
        RECT 2895.340 1081.550 2895.600 1081.870 ;
        RECT 2903.160 1081.550 2903.420 1081.870 ;
        RECT 2895.400 1079.685 2895.540 1081.550 ;
        RECT 2895.330 1079.315 2895.610 1079.685 ;
      LAYER via2 ;
        RECT 2903.150 2199.320 2903.430 2199.600 ;
        RECT 2895.330 1079.360 2895.610 1079.640 ;
      LAYER met3 ;
        RECT 2903.125 2199.610 2903.455 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2903.125 2199.310 2924.800 2199.610 ;
        RECT 2903.125 2199.295 2903.455 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
        RECT 2895.305 1079.650 2895.635 1079.665 ;
        RECT 2884.510 1079.350 2895.635 1079.650 ;
        RECT 2884.510 1076.720 2884.810 1079.350 ;
        RECT 2895.305 1079.335 2895.635 1079.350 ;
        RECT 2881.000 1076.120 2885.000 1076.720 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 204.420 2924.800 205.620 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2551.100 2924.800 2552.300 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2785.700 2924.800 2786.900 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3020.300 2924.800 3021.500 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3254.900 2924.800 3256.100 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3489.500 2924.800 3490.700 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 439.020 2924.800 440.220 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 3267.140 2.400 3268.340 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2979.500 2.400 2980.700 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2692.540 2.400 2693.740 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2404.900 2.400 2406.100 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2117.940 2.400 2119.140 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1830.300 2.400 1831.500 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 673.620 2924.800 674.820 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1543.340 2.400 1544.540 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1327.780 2.400 1328.980 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1112.220 2.400 1113.420 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 896.660 2.400 897.860 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 681.100 2.400 682.300 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 465.540 2.400 466.740 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 249.980 2.400 251.180 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 35.100 2.400 36.300 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 908.900 2924.800 910.100 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1143.500 2924.800 1144.700 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1378.100 2924.800 1379.300 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1612.700 2924.800 1613.900 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1847.300 2924.800 1848.500 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2081.900 2924.800 2083.100 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2316.500 2924.800 2317.700 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 145.940 2924.800 147.140 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2492.620 2924.800 2493.820 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2727.220 2924.800 2728.420 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2961.820 2924.800 2963.020 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3196.420 2924.800 3197.620 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3431.020 2924.800 3432.220 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 380.540 2924.800 381.740 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 3339.220 2.400 3340.420 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 3051.580 2.400 3052.780 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2764.620 2.400 2765.820 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2476.980 2.400 2478.180 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2189.340 2.400 2190.540 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1902.380 2.400 1903.580 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 615.140 2924.800 616.340 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1614.740 2.400 1615.940 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1399.860 2.400 1401.060 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1184.300 2.400 1185.500 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 968.740 2.400 969.940 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 753.180 2.400 754.380 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 537.620 2.400 538.820 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 322.060 2.400 323.260 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 106.500 2.400 107.700 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 849.740 2924.800 850.940 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1084.340 2924.800 1085.540 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1318.940 2924.800 1320.140 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1553.540 2924.800 1554.740 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1788.820 2924.800 1790.020 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2023.420 2924.800 2024.620 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2258.020 2924.800 2259.220 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 674.310 -4.800 674.870 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2879.745 1062.925 2879.915 1104.915 ;
        RECT 2880.665 1007.505 2880.835 1062.415 ;
        RECT 2881.125 931.345 2881.295 959.055 ;
        RECT 2880.205 96.645 2880.375 120.955 ;
      LAYER mcon ;
        RECT 2879.745 1104.745 2879.915 1104.915 ;
        RECT 2880.665 1062.245 2880.835 1062.415 ;
        RECT 2881.125 958.885 2881.295 959.055 ;
        RECT 2880.205 120.785 2880.375 120.955 ;
      LAYER met1 ;
        RECT 2880.130 1171.540 2880.450 1171.600 ;
        RECT 2881.970 1171.540 2882.290 1171.600 ;
        RECT 2880.130 1171.400 2882.290 1171.540 ;
        RECT 2880.130 1171.340 2880.450 1171.400 ;
        RECT 2881.970 1171.340 2882.290 1171.400 ;
        RECT 2879.670 1104.900 2879.990 1104.960 ;
        RECT 2879.475 1104.760 2879.990 1104.900 ;
        RECT 2879.670 1104.700 2879.990 1104.760 ;
        RECT 2879.685 1063.080 2879.975 1063.125 ;
        RECT 2880.590 1063.080 2880.910 1063.140 ;
        RECT 2879.685 1062.940 2880.910 1063.080 ;
        RECT 2879.685 1062.895 2879.975 1062.940 ;
        RECT 2880.590 1062.880 2880.910 1062.940 ;
        RECT 2880.590 1062.400 2880.910 1062.460 ;
        RECT 2880.395 1062.260 2880.910 1062.400 ;
        RECT 2880.590 1062.200 2880.910 1062.260 ;
        RECT 2880.605 1007.660 2880.895 1007.705 ;
        RECT 2881.050 1007.660 2881.370 1007.720 ;
        RECT 2880.605 1007.520 2881.370 1007.660 ;
        RECT 2880.605 1007.475 2880.895 1007.520 ;
        RECT 2881.050 1007.460 2881.370 1007.520 ;
        RECT 2881.050 959.040 2881.370 959.100 ;
        RECT 2880.855 958.900 2881.370 959.040 ;
        RECT 2881.050 958.840 2881.370 958.900 ;
        RECT 2881.050 931.500 2881.370 931.560 ;
        RECT 2880.855 931.360 2881.370 931.500 ;
        RECT 2881.050 931.300 2881.370 931.360 ;
        RECT 2881.510 428.100 2881.830 428.360 ;
        RECT 2881.600 427.680 2881.740 428.100 ;
        RECT 2881.510 427.420 2881.830 427.680 ;
        RECT 2881.050 289.920 2881.370 289.980 ;
        RECT 2881.510 289.920 2881.830 289.980 ;
        RECT 2881.050 289.780 2881.830 289.920 ;
        RECT 2881.050 289.720 2881.370 289.780 ;
        RECT 2881.510 289.720 2881.830 289.780 ;
        RECT 2880.145 120.940 2880.435 120.985 ;
        RECT 2881.050 120.940 2881.370 121.000 ;
        RECT 2880.145 120.800 2881.370 120.940 ;
        RECT 2880.145 120.755 2880.435 120.800 ;
        RECT 2881.050 120.740 2881.370 120.800 ;
        RECT 2880.130 96.800 2880.450 96.860 ;
        RECT 2879.935 96.660 2880.450 96.800 ;
        RECT 2880.130 96.600 2880.450 96.660 ;
        RECT 2.830 37.980 3.150 38.040 ;
        RECT 2878.750 37.980 2879.070 38.040 ;
        RECT 2.830 37.840 2879.070 37.980 ;
        RECT 2.830 37.780 3.150 37.840 ;
        RECT 2878.750 37.780 2879.070 37.840 ;
      LAYER via ;
        RECT 2880.160 1171.340 2880.420 1171.600 ;
        RECT 2882.000 1171.340 2882.260 1171.600 ;
        RECT 2879.700 1104.700 2879.960 1104.960 ;
        RECT 2880.620 1062.880 2880.880 1063.140 ;
        RECT 2880.620 1062.200 2880.880 1062.460 ;
        RECT 2881.080 1007.460 2881.340 1007.720 ;
        RECT 2881.080 958.840 2881.340 959.100 ;
        RECT 2881.080 931.300 2881.340 931.560 ;
        RECT 2881.540 428.100 2881.800 428.360 ;
        RECT 2881.540 427.420 2881.800 427.680 ;
        RECT 2881.080 289.720 2881.340 289.980 ;
        RECT 2881.540 289.720 2881.800 289.980 ;
        RECT 2881.080 120.740 2881.340 121.000 ;
        RECT 2880.160 96.600 2880.420 96.860 ;
        RECT 2.860 37.780 3.120 38.040 ;
        RECT 2878.780 37.780 2879.040 38.040 ;
      LAYER met2 ;
        RECT 2881.990 1182.675 2882.270 1183.045 ;
        RECT 2882.060 1171.630 2882.200 1182.675 ;
        RECT 2880.160 1171.310 2880.420 1171.630 ;
        RECT 2882.000 1171.310 2882.260 1171.630 ;
        RECT 2880.220 1125.810 2880.360 1171.310 ;
        RECT 2879.760 1125.670 2880.360 1125.810 ;
        RECT 2879.760 1104.990 2879.900 1125.670 ;
        RECT 2879.700 1104.670 2879.960 1104.990 ;
        RECT 2880.620 1062.850 2880.880 1063.170 ;
        RECT 2880.680 1062.490 2880.820 1062.850 ;
        RECT 2880.620 1062.170 2880.880 1062.490 ;
        RECT 2881.080 1007.430 2881.340 1007.750 ;
        RECT 2881.140 959.130 2881.280 1007.430 ;
        RECT 2881.080 958.810 2881.340 959.130 ;
        RECT 2881.080 931.270 2881.340 931.590 ;
        RECT 2881.140 683.810 2881.280 931.270 ;
        RECT 2880.680 683.670 2881.280 683.810 ;
        RECT 2880.680 641.650 2880.820 683.670 ;
        RECT 2880.680 641.510 2881.280 641.650 ;
        RECT 2881.140 545.260 2881.280 641.510 ;
        RECT 2881.140 545.120 2881.740 545.260 ;
        RECT 2881.600 428.390 2881.740 545.120 ;
        RECT 2881.540 428.070 2881.800 428.390 ;
        RECT 2881.540 427.450 2881.800 427.710 ;
        RECT 2881.140 427.390 2881.800 427.450 ;
        RECT 2881.140 427.310 2881.740 427.390 ;
        RECT 2881.140 397.530 2881.280 427.310 ;
        RECT 2881.140 397.390 2881.740 397.530 ;
        RECT 2881.600 290.010 2881.740 397.390 ;
        RECT 2881.080 289.690 2881.340 290.010 ;
        RECT 2881.540 289.690 2881.800 290.010 ;
        RECT 2881.140 121.030 2881.280 289.690 ;
        RECT 2881.080 120.710 2881.340 121.030 ;
        RECT 2880.160 96.570 2880.420 96.890 ;
        RECT 2880.220 58.210 2880.360 96.570 ;
        RECT 2878.840 58.070 2880.360 58.210 ;
        RECT 2878.840 38.070 2878.980 58.070 ;
        RECT 2.860 37.750 3.120 38.070 ;
        RECT 2878.780 37.750 2879.040 38.070 ;
        RECT 2.920 2.400 3.060 37.750 ;
        RECT 2.710 -4.800 3.270 2.400 ;
      LAYER via2 ;
        RECT 2881.990 1182.720 2882.270 1183.000 ;
      LAYER met3 ;
        RECT 2881.000 1185.600 2885.000 1186.200 ;
        RECT 2881.750 1183.025 2882.050 1185.600 ;
        RECT 2881.750 1182.710 2882.295 1183.025 ;
        RECT 2881.965 1182.695 2882.295 1182.710 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2879.745 962.625 2879.915 994.415 ;
        RECT 2879.745 869.805 2879.915 914.855 ;
        RECT 2879.745 803.845 2879.915 853.655 ;
        RECT 2879.745 752.165 2879.915 767.295 ;
        RECT 2879.745 721.905 2879.915 746.895 ;
        RECT 2879.745 662.745 2879.915 704.735 ;
        RECT 2879.745 592.705 2879.915 660.535 ;
        RECT 2880.665 512.125 2880.835 544.255 ;
        RECT 2881.125 351.645 2881.295 469.115 ;
        RECT 2879.745 289.085 2879.915 316.795 ;
        RECT 2880.205 196.945 2880.375 258.995 ;
        RECT 2879.745 101.405 2879.915 186.235 ;
      LAYER mcon ;
        RECT 2879.745 994.245 2879.915 994.415 ;
        RECT 2879.745 914.685 2879.915 914.855 ;
        RECT 2879.745 853.485 2879.915 853.655 ;
        RECT 2879.745 767.125 2879.915 767.295 ;
        RECT 2879.745 746.725 2879.915 746.895 ;
        RECT 2879.745 704.565 2879.915 704.735 ;
        RECT 2879.745 660.365 2879.915 660.535 ;
        RECT 2880.665 544.085 2880.835 544.255 ;
        RECT 2881.125 468.945 2881.295 469.115 ;
        RECT 2879.745 316.625 2879.915 316.795 ;
        RECT 2880.205 258.825 2880.375 258.995 ;
        RECT 2879.745 186.065 2879.915 186.235 ;
      LAYER met1 ;
        RECT 2879.670 1208.600 2879.990 1208.660 ;
        RECT 2881.510 1208.600 2881.830 1208.660 ;
        RECT 2879.670 1208.460 2881.830 1208.600 ;
        RECT 2879.670 1208.400 2879.990 1208.460 ;
        RECT 2881.510 1208.400 2881.830 1208.460 ;
        RECT 2879.670 1183.440 2879.990 1183.500 ;
        RECT 2881.050 1183.440 2881.370 1183.500 ;
        RECT 2879.670 1183.300 2881.370 1183.440 ;
        RECT 2879.670 1183.240 2879.990 1183.300 ;
        RECT 2881.050 1183.240 2881.370 1183.300 ;
        RECT 2881.050 1087.560 2881.370 1087.620 ;
        RECT 2881.970 1087.560 2882.290 1087.620 ;
        RECT 2881.050 1087.420 2882.290 1087.560 ;
        RECT 2881.050 1087.360 2881.370 1087.420 ;
        RECT 2881.970 1087.360 2882.290 1087.420 ;
        RECT 2879.685 994.400 2879.975 994.445 ;
        RECT 2881.510 994.400 2881.830 994.460 ;
        RECT 2879.685 994.260 2881.830 994.400 ;
        RECT 2879.685 994.215 2879.975 994.260 ;
        RECT 2881.510 994.200 2881.830 994.260 ;
        RECT 2879.685 962.780 2879.975 962.825 ;
        RECT 2880.590 962.780 2880.910 962.840 ;
        RECT 2879.685 962.640 2880.910 962.780 ;
        RECT 2879.685 962.595 2879.975 962.640 ;
        RECT 2880.590 962.580 2880.910 962.640 ;
        RECT 2879.685 914.840 2879.975 914.885 ;
        RECT 2880.130 914.840 2880.450 914.900 ;
        RECT 2879.685 914.700 2880.450 914.840 ;
        RECT 2879.685 914.655 2879.975 914.700 ;
        RECT 2880.130 914.640 2880.450 914.700 ;
        RECT 2879.670 869.960 2879.990 870.020 ;
        RECT 2879.475 869.820 2879.990 869.960 ;
        RECT 2879.670 869.760 2879.990 869.820 ;
        RECT 2879.670 853.640 2879.990 853.700 ;
        RECT 2879.475 853.500 2879.990 853.640 ;
        RECT 2879.670 853.440 2879.990 853.500 ;
        RECT 2879.670 804.000 2879.990 804.060 ;
        RECT 2879.475 803.860 2879.990 804.000 ;
        RECT 2879.670 803.800 2879.990 803.860 ;
        RECT 2879.670 767.280 2879.990 767.340 ;
        RECT 2879.475 767.140 2879.990 767.280 ;
        RECT 2879.670 767.080 2879.990 767.140 ;
        RECT 2879.670 752.320 2879.990 752.380 ;
        RECT 2879.475 752.180 2879.990 752.320 ;
        RECT 2879.670 752.120 2879.990 752.180 ;
        RECT 2879.670 746.880 2879.990 746.940 ;
        RECT 2879.475 746.740 2879.990 746.880 ;
        RECT 2879.670 746.680 2879.990 746.740 ;
        RECT 2879.670 722.060 2879.990 722.120 ;
        RECT 2879.475 721.920 2879.990 722.060 ;
        RECT 2879.670 721.860 2879.990 721.920 ;
        RECT 2879.670 704.720 2879.990 704.780 ;
        RECT 2879.475 704.580 2879.990 704.720 ;
        RECT 2879.670 704.520 2879.990 704.580 ;
        RECT 2879.670 662.900 2879.990 662.960 ;
        RECT 2879.475 662.760 2879.990 662.900 ;
        RECT 2879.670 662.700 2879.990 662.760 ;
        RECT 2879.670 660.520 2879.990 660.580 ;
        RECT 2879.475 660.380 2879.990 660.520 ;
        RECT 2879.670 660.320 2879.990 660.380 ;
        RECT 2879.685 592.860 2879.975 592.905 ;
        RECT 2880.590 592.860 2880.910 592.920 ;
        RECT 2879.685 592.720 2880.910 592.860 ;
        RECT 2879.685 592.675 2879.975 592.720 ;
        RECT 2880.590 592.660 2880.910 592.720 ;
        RECT 2880.590 544.240 2880.910 544.300 ;
        RECT 2880.395 544.100 2880.910 544.240 ;
        RECT 2880.590 544.040 2880.910 544.100 ;
        RECT 2879.670 512.280 2879.990 512.340 ;
        RECT 2880.605 512.280 2880.895 512.325 ;
        RECT 2879.670 512.140 2880.895 512.280 ;
        RECT 2879.670 512.080 2879.990 512.140 ;
        RECT 2880.605 512.095 2880.895 512.140 ;
        RECT 2879.670 502.220 2879.990 502.480 ;
        RECT 2879.760 501.800 2879.900 502.220 ;
        RECT 2879.670 501.540 2879.990 501.800 ;
        RECT 2879.670 469.100 2879.990 469.160 ;
        RECT 2881.065 469.100 2881.355 469.145 ;
        RECT 2879.670 468.960 2881.355 469.100 ;
        RECT 2879.670 468.900 2879.990 468.960 ;
        RECT 2881.065 468.915 2881.355 468.960 ;
        RECT 2879.670 351.800 2879.990 351.860 ;
        RECT 2881.065 351.800 2881.355 351.845 ;
        RECT 2879.670 351.660 2881.355 351.800 ;
        RECT 2879.670 351.600 2879.990 351.660 ;
        RECT 2881.065 351.615 2881.355 351.660 ;
        RECT 2879.670 316.780 2879.990 316.840 ;
        RECT 2879.475 316.640 2879.990 316.780 ;
        RECT 2879.670 316.580 2879.990 316.640 ;
        RECT 2879.685 289.240 2879.975 289.285 ;
        RECT 2880.590 289.240 2880.910 289.300 ;
        RECT 2879.685 289.100 2880.910 289.240 ;
        RECT 2879.685 289.055 2879.975 289.100 ;
        RECT 2880.590 289.040 2880.910 289.100 ;
        RECT 2880.145 258.980 2880.435 259.025 ;
        RECT 2880.590 258.980 2880.910 259.040 ;
        RECT 2880.145 258.840 2880.910 258.980 ;
        RECT 2880.145 258.795 2880.435 258.840 ;
        RECT 2880.590 258.780 2880.910 258.840 ;
        RECT 2879.670 197.100 2879.990 197.160 ;
        RECT 2880.145 197.100 2880.435 197.145 ;
        RECT 2879.670 196.960 2880.435 197.100 ;
        RECT 2879.670 196.900 2879.990 196.960 ;
        RECT 2880.145 196.915 2880.435 196.960 ;
        RECT 2879.670 186.220 2879.990 186.280 ;
        RECT 2879.475 186.080 2879.990 186.220 ;
        RECT 2879.670 186.020 2879.990 186.080 ;
        RECT 2879.670 101.560 2879.990 101.620 ;
        RECT 2879.475 101.420 2879.990 101.560 ;
        RECT 2879.670 101.360 2879.990 101.420 ;
        RECT 2879.670 86.260 2879.990 86.320 ;
        RECT 2881.510 86.260 2881.830 86.320 ;
        RECT 2879.670 86.120 2881.830 86.260 ;
        RECT 2879.670 86.060 2879.990 86.120 ;
        RECT 2881.510 86.060 2881.830 86.120 ;
        RECT 8.350 38.320 8.670 38.380 ;
        RECT 2881.510 38.320 2881.830 38.380 ;
        RECT 8.350 38.180 2881.830 38.320 ;
        RECT 8.350 38.120 8.670 38.180 ;
        RECT 2881.510 38.120 2881.830 38.180 ;
      LAYER via ;
        RECT 2879.700 1208.400 2879.960 1208.660 ;
        RECT 2881.540 1208.400 2881.800 1208.660 ;
        RECT 2879.700 1183.240 2879.960 1183.500 ;
        RECT 2881.080 1183.240 2881.340 1183.500 ;
        RECT 2881.080 1087.360 2881.340 1087.620 ;
        RECT 2882.000 1087.360 2882.260 1087.620 ;
        RECT 2881.540 994.200 2881.800 994.460 ;
        RECT 2880.620 962.580 2880.880 962.840 ;
        RECT 2880.160 914.640 2880.420 914.900 ;
        RECT 2879.700 869.760 2879.960 870.020 ;
        RECT 2879.700 853.440 2879.960 853.700 ;
        RECT 2879.700 803.800 2879.960 804.060 ;
        RECT 2879.700 767.080 2879.960 767.340 ;
        RECT 2879.700 752.120 2879.960 752.380 ;
        RECT 2879.700 746.680 2879.960 746.940 ;
        RECT 2879.700 721.860 2879.960 722.120 ;
        RECT 2879.700 704.520 2879.960 704.780 ;
        RECT 2879.700 662.700 2879.960 662.960 ;
        RECT 2879.700 660.320 2879.960 660.580 ;
        RECT 2880.620 592.660 2880.880 592.920 ;
        RECT 2880.620 544.040 2880.880 544.300 ;
        RECT 2879.700 512.080 2879.960 512.340 ;
        RECT 2879.700 502.220 2879.960 502.480 ;
        RECT 2879.700 501.540 2879.960 501.800 ;
        RECT 2879.700 468.900 2879.960 469.160 ;
        RECT 2879.700 351.600 2879.960 351.860 ;
        RECT 2879.700 316.580 2879.960 316.840 ;
        RECT 2880.620 289.040 2880.880 289.300 ;
        RECT 2880.620 258.780 2880.880 259.040 ;
        RECT 2879.700 196.900 2879.960 197.160 ;
        RECT 2879.700 186.020 2879.960 186.280 ;
        RECT 2879.700 101.360 2879.960 101.620 ;
        RECT 2879.700 86.060 2879.960 86.320 ;
        RECT 2881.540 86.060 2881.800 86.320 ;
        RECT 8.380 38.120 8.640 38.380 ;
        RECT 2881.540 38.120 2881.800 38.380 ;
      LAYER met2 ;
        RECT 2881.530 1292.835 2881.810 1293.205 ;
        RECT 2881.600 1208.690 2881.740 1292.835 ;
        RECT 2879.700 1208.370 2879.960 1208.690 ;
        RECT 2881.540 1208.370 2881.800 1208.690 ;
        RECT 2879.760 1183.530 2879.900 1208.370 ;
        RECT 2879.700 1183.210 2879.960 1183.530 ;
        RECT 2881.080 1183.210 2881.340 1183.530 ;
        RECT 2881.140 1087.650 2881.280 1183.210 ;
        RECT 2881.080 1087.330 2881.340 1087.650 ;
        RECT 2882.000 1087.330 2882.260 1087.650 ;
        RECT 2882.060 1086.370 2882.200 1087.330 ;
        RECT 2881.600 1086.230 2882.200 1086.370 ;
        RECT 2881.600 994.490 2881.740 1086.230 ;
        RECT 2881.540 994.170 2881.800 994.490 ;
        RECT 2880.620 962.550 2880.880 962.870 ;
        RECT 2880.680 930.650 2880.820 962.550 ;
        RECT 2880.220 930.510 2880.820 930.650 ;
        RECT 2880.220 914.930 2880.360 930.510 ;
        RECT 2880.160 914.610 2880.420 914.930 ;
        RECT 2879.700 869.730 2879.960 870.050 ;
        RECT 2879.760 853.730 2879.900 869.730 ;
        RECT 2879.700 853.410 2879.960 853.730 ;
        RECT 2879.700 803.770 2879.960 804.090 ;
        RECT 2879.760 767.370 2879.900 803.770 ;
        RECT 2879.700 767.050 2879.960 767.370 ;
        RECT 2879.700 752.090 2879.960 752.410 ;
        RECT 2879.760 746.970 2879.900 752.090 ;
        RECT 2879.700 746.650 2879.960 746.970 ;
        RECT 2879.700 721.830 2879.960 722.150 ;
        RECT 2879.760 704.810 2879.900 721.830 ;
        RECT 2879.700 704.490 2879.960 704.810 ;
        RECT 2879.700 662.670 2879.960 662.990 ;
        RECT 2879.760 660.610 2879.900 662.670 ;
        RECT 2879.700 660.290 2879.960 660.610 ;
        RECT 2880.620 592.630 2880.880 592.950 ;
        RECT 2880.680 544.330 2880.820 592.630 ;
        RECT 2880.620 544.010 2880.880 544.330 ;
        RECT 2879.700 512.050 2879.960 512.370 ;
        RECT 2879.760 502.510 2879.900 512.050 ;
        RECT 2879.700 502.190 2879.960 502.510 ;
        RECT 2879.700 501.510 2879.960 501.830 ;
        RECT 2879.760 469.190 2879.900 501.510 ;
        RECT 2879.700 468.870 2879.960 469.190 ;
        RECT 2879.700 351.570 2879.960 351.890 ;
        RECT 2879.760 316.870 2879.900 351.570 ;
        RECT 2879.700 316.550 2879.960 316.870 ;
        RECT 2880.620 289.010 2880.880 289.330 ;
        RECT 2880.680 259.070 2880.820 289.010 ;
        RECT 2880.620 258.750 2880.880 259.070 ;
        RECT 2879.700 196.870 2879.960 197.190 ;
        RECT 2879.760 186.310 2879.900 196.870 ;
        RECT 2879.700 185.990 2879.960 186.310 ;
        RECT 2879.700 101.330 2879.960 101.650 ;
        RECT 2879.760 86.350 2879.900 101.330 ;
        RECT 2879.700 86.030 2879.960 86.350 ;
        RECT 2881.540 86.030 2881.800 86.350 ;
        RECT 2881.600 38.410 2881.740 86.030 ;
        RECT 8.380 38.090 8.640 38.410 ;
        RECT 2881.540 38.090 2881.800 38.410 ;
        RECT 8.440 2.400 8.580 38.090 ;
        RECT 8.230 -4.800 8.790 2.400 ;
      LAYER via2 ;
        RECT 2881.530 1292.880 2881.810 1293.160 ;
      LAYER met3 ;
        RECT 2881.000 1295.760 2885.000 1296.360 ;
        RECT 2881.750 1293.185 2882.050 1295.760 ;
        RECT 2881.505 1292.870 2882.050 1293.185 ;
        RECT 2881.505 1292.855 2881.835 1292.870 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 45.610 3446.140 45.930 3446.200 ;
        RECT 1185.950 3446.140 1186.270 3446.200 ;
        RECT 45.610 3446.000 1186.270 3446.140 ;
        RECT 45.610 3445.940 45.930 3446.000 ;
        RECT 1185.950 3445.940 1186.270 3446.000 ;
        RECT 45.610 19.280 45.930 19.340 ;
        RECT 44.780 19.140 45.930 19.280 ;
        RECT 14.330 18.940 14.650 19.000 ;
        RECT 44.780 18.940 44.920 19.140 ;
        RECT 45.610 19.080 45.930 19.140 ;
        RECT 14.330 18.800 44.920 18.940 ;
        RECT 14.330 18.740 14.650 18.800 ;
      LAYER via ;
        RECT 45.640 3445.940 45.900 3446.200 ;
        RECT 1185.980 3445.940 1186.240 3446.200 ;
        RECT 14.360 18.740 14.620 19.000 ;
        RECT 45.640 19.080 45.900 19.340 ;
      LAYER met2 ;
        RECT 45.640 3445.910 45.900 3446.230 ;
        RECT 1185.980 3445.910 1186.240 3446.230 ;
        RECT 45.700 19.370 45.840 3445.910 ;
        RECT 1186.040 3435.000 1186.180 3445.910 ;
        RECT 1186.010 3431.000 1186.290 3435.000 ;
        RECT 45.640 19.050 45.900 19.370 ;
        RECT 14.360 18.710 14.620 19.030 ;
        RECT 14.420 2.400 14.560 18.710 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 45.150 3445.800 45.470 3445.860 ;
        RECT 1295.430 3445.800 1295.750 3445.860 ;
        RECT 45.150 3445.660 1295.750 3445.800 ;
        RECT 45.150 3445.600 45.470 3445.660 ;
        RECT 1295.430 3445.600 1295.750 3445.660 ;
        RECT 38.250 17.240 38.570 17.300 ;
        RECT 45.150 17.240 45.470 17.300 ;
        RECT 38.250 17.100 45.470 17.240 ;
        RECT 38.250 17.040 38.570 17.100 ;
        RECT 45.150 17.040 45.470 17.100 ;
      LAYER via ;
        RECT 45.180 3445.600 45.440 3445.860 ;
        RECT 1295.460 3445.600 1295.720 3445.860 ;
        RECT 38.280 17.040 38.540 17.300 ;
        RECT 45.180 17.040 45.440 17.300 ;
      LAYER met2 ;
        RECT 45.180 3445.570 45.440 3445.890 ;
        RECT 1295.460 3445.570 1295.720 3445.890 ;
        RECT 45.240 17.330 45.380 3445.570 ;
        RECT 1295.520 3435.000 1295.660 3445.570 ;
        RECT 1295.490 3431.000 1295.770 3435.000 ;
        RECT 38.280 17.010 38.540 17.330 ;
        RECT 45.180 17.010 45.440 17.330 ;
        RECT 38.340 2.400 38.480 17.010 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 48.830 3445.120 49.150 3445.180 ;
        RECT 1514.850 3445.120 1515.170 3445.180 ;
        RECT 48.830 3444.980 1515.170 3445.120 ;
        RECT 48.830 3444.920 49.150 3444.980 ;
        RECT 1514.850 3444.920 1515.170 3444.980 ;
        RECT 48.830 15.200 49.150 15.260 ;
        RECT 240.650 15.200 240.970 15.260 ;
        RECT 48.830 15.060 240.970 15.200 ;
        RECT 48.830 15.000 49.150 15.060 ;
        RECT 240.650 15.000 240.970 15.060 ;
      LAYER via ;
        RECT 48.860 3444.920 49.120 3445.180 ;
        RECT 1514.880 3444.920 1515.140 3445.180 ;
        RECT 48.860 15.000 49.120 15.260 ;
        RECT 240.680 15.000 240.940 15.260 ;
      LAYER met2 ;
        RECT 48.860 3444.890 49.120 3445.210 ;
        RECT 1514.880 3444.890 1515.140 3445.210 ;
        RECT 48.920 15.290 49.060 3444.890 ;
        RECT 1514.940 3435.000 1515.080 3444.890 ;
        RECT 1514.910 3431.000 1515.190 3435.000 ;
        RECT 48.860 14.970 49.120 15.290 ;
        RECT 240.680 14.970 240.940 15.290 ;
        RECT 240.740 2.400 240.880 14.970 ;
        RECT 240.530 -4.800 241.090 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 258.130 25.740 258.450 25.800 ;
        RECT 2197.950 25.740 2198.270 25.800 ;
        RECT 258.130 25.600 2198.270 25.740 ;
        RECT 258.130 25.540 258.450 25.600 ;
        RECT 2197.950 25.540 2198.270 25.600 ;
      LAYER via ;
        RECT 258.160 25.540 258.420 25.800 ;
        RECT 2197.980 25.540 2198.240 25.800 ;
      LAYER met2 ;
        RECT 2198.010 35.000 2198.290 39.000 ;
        RECT 2198.040 25.830 2198.180 35.000 ;
        RECT 258.160 25.510 258.420 25.830 ;
        RECT 2197.980 25.510 2198.240 25.830 ;
        RECT 258.220 2.400 258.360 25.510 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 276.070 25.400 276.390 25.460 ;
        RECT 2248.550 25.400 2248.870 25.460 ;
        RECT 276.070 25.260 2248.870 25.400 ;
        RECT 276.070 25.200 276.390 25.260 ;
        RECT 2248.550 25.200 2248.870 25.260 ;
      LAYER via ;
        RECT 276.100 25.200 276.360 25.460 ;
        RECT 2248.580 25.200 2248.840 25.460 ;
      LAYER met2 ;
        RECT 2248.610 35.000 2248.890 39.000 ;
        RECT 2248.640 25.490 2248.780 35.000 ;
        RECT 276.100 25.170 276.360 25.490 ;
        RECT 2248.580 25.170 2248.840 25.490 ;
        RECT 276.160 2.400 276.300 25.170 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2879.745 1393.745 2879.915 1495.915 ;
        RECT 2879.745 1313.505 2879.915 1365.015 ;
        RECT 2879.745 1245.505 2879.915 1288.175 ;
        RECT 2881.585 993.565 2881.755 996.455 ;
        RECT 2881.125 603.585 2881.295 652.715 ;
        RECT 2879.745 360.825 2879.915 406.895 ;
        RECT 2881.585 286.365 2881.755 294.015 ;
      LAYER mcon ;
        RECT 2879.745 1495.745 2879.915 1495.915 ;
        RECT 2879.745 1364.845 2879.915 1365.015 ;
        RECT 2879.745 1288.005 2879.915 1288.175 ;
        RECT 2881.585 996.285 2881.755 996.455 ;
        RECT 2881.125 652.545 2881.295 652.715 ;
        RECT 2879.745 406.725 2879.915 406.895 ;
        RECT 2881.585 293.845 2881.755 294.015 ;
      LAYER met1 ;
        RECT 2879.670 1539.080 2879.990 1539.140 ;
        RECT 2881.510 1539.080 2881.830 1539.140 ;
        RECT 2879.670 1538.940 2881.830 1539.080 ;
        RECT 2879.670 1538.880 2879.990 1538.940 ;
        RECT 2881.510 1538.880 2881.830 1538.940 ;
        RECT 2879.670 1495.900 2879.990 1495.960 ;
        RECT 2879.475 1495.760 2879.990 1495.900 ;
        RECT 2879.670 1495.700 2879.990 1495.760 ;
        RECT 2879.670 1393.900 2879.990 1393.960 ;
        RECT 2879.475 1393.760 2879.990 1393.900 ;
        RECT 2879.670 1393.700 2879.990 1393.760 ;
        RECT 2879.670 1365.000 2879.990 1365.060 ;
        RECT 2879.475 1364.860 2879.990 1365.000 ;
        RECT 2879.670 1364.800 2879.990 1364.860 ;
        RECT 2879.670 1313.660 2879.990 1313.720 ;
        RECT 2879.475 1313.520 2879.990 1313.660 ;
        RECT 2879.670 1313.460 2879.990 1313.520 ;
        RECT 2879.670 1288.160 2879.990 1288.220 ;
        RECT 2879.475 1288.020 2879.990 1288.160 ;
        RECT 2879.670 1287.960 2879.990 1288.020 ;
        RECT 2879.670 1245.660 2879.990 1245.720 ;
        RECT 2879.475 1245.520 2879.990 1245.660 ;
        RECT 2879.670 1245.460 2879.990 1245.520 ;
        RECT 2879.670 1175.280 2879.990 1175.340 ;
        RECT 2881.510 1175.280 2881.830 1175.340 ;
        RECT 2879.670 1175.140 2881.830 1175.280 ;
        RECT 2879.670 1175.080 2879.990 1175.140 ;
        RECT 2881.510 1175.080 2881.830 1175.140 ;
        RECT 2879.670 1013.780 2879.990 1013.840 ;
        RECT 2881.050 1013.780 2881.370 1013.840 ;
        RECT 2879.670 1013.640 2881.370 1013.780 ;
        RECT 2879.670 1013.580 2879.990 1013.640 ;
        RECT 2881.050 1013.580 2881.370 1013.640 ;
        RECT 2879.670 996.440 2879.990 996.500 ;
        RECT 2881.525 996.440 2881.815 996.485 ;
        RECT 2879.670 996.300 2881.815 996.440 ;
        RECT 2879.670 996.240 2879.990 996.300 ;
        RECT 2881.525 996.255 2881.815 996.300 ;
        RECT 2881.510 993.720 2881.830 993.780 ;
        RECT 2881.315 993.580 2881.830 993.720 ;
        RECT 2881.510 993.520 2881.830 993.580 ;
        RECT 2879.670 924.700 2879.990 924.760 ;
        RECT 2881.510 924.700 2881.830 924.760 ;
        RECT 2879.670 924.560 2881.830 924.700 ;
        RECT 2879.670 924.500 2879.990 924.560 ;
        RECT 2881.510 924.500 2881.830 924.560 ;
        RECT 2879.670 916.880 2879.990 916.940 ;
        RECT 2881.510 916.880 2881.830 916.940 ;
        RECT 2879.670 916.740 2881.830 916.880 ;
        RECT 2879.670 916.680 2879.990 916.740 ;
        RECT 2881.510 916.680 2881.830 916.740 ;
        RECT 2880.130 722.740 2880.450 722.800 ;
        RECT 2881.510 722.740 2881.830 722.800 ;
        RECT 2880.130 722.600 2881.830 722.740 ;
        RECT 2880.130 722.540 2880.450 722.600 ;
        RECT 2881.510 722.540 2881.830 722.600 ;
        RECT 2880.130 685.340 2880.450 685.400 ;
        RECT 2879.760 685.200 2880.450 685.340 ;
        RECT 2879.760 685.060 2879.900 685.200 ;
        RECT 2880.130 685.140 2880.450 685.200 ;
        RECT 2879.670 684.800 2879.990 685.060 ;
        RECT 2879.670 652.700 2879.990 652.760 ;
        RECT 2881.065 652.700 2881.355 652.745 ;
        RECT 2879.670 652.560 2881.355 652.700 ;
        RECT 2879.670 652.500 2879.990 652.560 ;
        RECT 2881.065 652.515 2881.355 652.560 ;
        RECT 2881.065 603.740 2881.355 603.785 ;
        RECT 2881.510 603.740 2881.830 603.800 ;
        RECT 2881.065 603.600 2881.830 603.740 ;
        RECT 2881.065 603.555 2881.355 603.600 ;
        RECT 2881.510 603.540 2881.830 603.600 ;
        RECT 2879.670 520.780 2879.990 520.840 ;
        RECT 2881.970 520.780 2882.290 520.840 ;
        RECT 2879.670 520.640 2882.290 520.780 ;
        RECT 2879.670 520.580 2879.990 520.640 ;
        RECT 2881.970 520.580 2882.290 520.640 ;
        RECT 2879.670 406.880 2879.990 406.940 ;
        RECT 2879.475 406.740 2879.990 406.880 ;
        RECT 2879.670 406.680 2879.990 406.740 ;
        RECT 2879.670 360.980 2879.990 361.040 ;
        RECT 2879.475 360.840 2879.990 360.980 ;
        RECT 2879.670 360.780 2879.990 360.840 ;
        RECT 2879.670 294.000 2879.990 294.060 ;
        RECT 2881.525 294.000 2881.815 294.045 ;
        RECT 2879.670 293.860 2881.815 294.000 ;
        RECT 2879.670 293.800 2879.990 293.860 ;
        RECT 2881.525 293.815 2881.815 293.860 ;
        RECT 2881.510 286.520 2881.830 286.580 ;
        RECT 2881.315 286.380 2881.830 286.520 ;
        RECT 2881.510 286.320 2881.830 286.380 ;
        RECT 2880.130 143.380 2880.450 143.440 ;
        RECT 2881.510 143.380 2881.830 143.440 ;
        RECT 2880.130 143.240 2881.830 143.380 ;
        RECT 2880.130 143.180 2880.450 143.240 ;
        RECT 2881.510 143.180 2881.830 143.240 ;
        RECT 2880.130 107.000 2880.450 107.060 ;
        RECT 2881.510 107.000 2881.830 107.060 ;
        RECT 2880.130 106.860 2881.830 107.000 ;
        RECT 2880.130 106.800 2880.450 106.860 ;
        RECT 2881.510 106.800 2881.830 106.860 ;
        RECT 294.010 38.660 294.330 38.720 ;
        RECT 2881.050 38.660 2881.370 38.720 ;
        RECT 294.010 38.520 2881.370 38.660 ;
        RECT 294.010 38.460 294.330 38.520 ;
        RECT 2881.050 38.460 2881.370 38.520 ;
      LAYER via ;
        RECT 2879.700 1538.880 2879.960 1539.140 ;
        RECT 2881.540 1538.880 2881.800 1539.140 ;
        RECT 2879.700 1495.700 2879.960 1495.960 ;
        RECT 2879.700 1393.700 2879.960 1393.960 ;
        RECT 2879.700 1364.800 2879.960 1365.060 ;
        RECT 2879.700 1313.460 2879.960 1313.720 ;
        RECT 2879.700 1287.960 2879.960 1288.220 ;
        RECT 2879.700 1245.460 2879.960 1245.720 ;
        RECT 2879.700 1175.080 2879.960 1175.340 ;
        RECT 2881.540 1175.080 2881.800 1175.340 ;
        RECT 2879.700 1013.580 2879.960 1013.840 ;
        RECT 2881.080 1013.580 2881.340 1013.840 ;
        RECT 2879.700 996.240 2879.960 996.500 ;
        RECT 2881.540 993.520 2881.800 993.780 ;
        RECT 2879.700 924.500 2879.960 924.760 ;
        RECT 2881.540 924.500 2881.800 924.760 ;
        RECT 2879.700 916.680 2879.960 916.940 ;
        RECT 2881.540 916.680 2881.800 916.940 ;
        RECT 2880.160 722.540 2880.420 722.800 ;
        RECT 2881.540 722.540 2881.800 722.800 ;
        RECT 2880.160 685.140 2880.420 685.400 ;
        RECT 2879.700 684.800 2879.960 685.060 ;
        RECT 2879.700 652.500 2879.960 652.760 ;
        RECT 2881.540 603.540 2881.800 603.800 ;
        RECT 2879.700 520.580 2879.960 520.840 ;
        RECT 2882.000 520.580 2882.260 520.840 ;
        RECT 2879.700 406.680 2879.960 406.940 ;
        RECT 2879.700 360.780 2879.960 361.040 ;
        RECT 2879.700 293.800 2879.960 294.060 ;
        RECT 2881.540 286.320 2881.800 286.580 ;
        RECT 2880.160 143.180 2880.420 143.440 ;
        RECT 2881.540 143.180 2881.800 143.440 ;
        RECT 2880.160 106.800 2880.420 107.060 ;
        RECT 2881.540 106.800 2881.800 107.060 ;
        RECT 294.040 38.460 294.300 38.720 ;
        RECT 2881.080 38.460 2881.340 38.720 ;
      LAYER met2 ;
        RECT 2881.530 1621.955 2881.810 1622.325 ;
        RECT 2881.600 1539.170 2881.740 1621.955 ;
        RECT 2879.700 1538.850 2879.960 1539.170 ;
        RECT 2881.540 1538.850 2881.800 1539.170 ;
        RECT 2879.760 1495.990 2879.900 1538.850 ;
        RECT 2879.700 1495.670 2879.960 1495.990 ;
        RECT 2879.700 1393.900 2879.960 1393.990 ;
        RECT 2879.300 1393.760 2879.960 1393.900 ;
        RECT 2879.300 1365.170 2879.440 1393.760 ;
        RECT 2879.700 1393.670 2879.960 1393.760 ;
        RECT 2879.300 1365.090 2879.900 1365.170 ;
        RECT 2879.300 1365.030 2879.960 1365.090 ;
        RECT 2879.700 1364.770 2879.960 1365.030 ;
        RECT 2879.700 1313.430 2879.960 1313.750 ;
        RECT 2879.760 1311.450 2879.900 1313.430 ;
        RECT 2879.300 1311.310 2879.900 1311.450 ;
        RECT 2879.300 1288.330 2879.440 1311.310 ;
        RECT 2879.300 1288.250 2879.900 1288.330 ;
        RECT 2879.300 1288.190 2879.960 1288.250 ;
        RECT 2879.700 1287.930 2879.960 1288.190 ;
        RECT 2879.700 1245.430 2879.960 1245.750 ;
        RECT 2879.760 1231.890 2879.900 1245.430 ;
        RECT 2879.300 1231.750 2879.900 1231.890 ;
        RECT 2879.300 1175.450 2879.440 1231.750 ;
        RECT 2879.300 1175.370 2879.900 1175.450 ;
        RECT 2879.300 1175.310 2879.960 1175.370 ;
        RECT 2879.700 1175.050 2879.960 1175.310 ;
        RECT 2881.540 1175.050 2881.800 1175.370 ;
        RECT 2881.600 1087.050 2881.740 1175.050 ;
        RECT 2881.140 1086.910 2881.740 1087.050 ;
        RECT 2881.140 1013.870 2881.280 1086.910 ;
        RECT 2879.700 1013.550 2879.960 1013.870 ;
        RECT 2881.080 1013.550 2881.340 1013.870 ;
        RECT 2879.760 996.530 2879.900 1013.550 ;
        RECT 2879.700 996.210 2879.960 996.530 ;
        RECT 2881.540 993.490 2881.800 993.810 ;
        RECT 2881.600 924.790 2881.740 993.490 ;
        RECT 2879.700 924.530 2879.960 924.790 ;
        RECT 2879.300 924.470 2879.960 924.530 ;
        RECT 2881.540 924.470 2881.800 924.790 ;
        RECT 2879.300 924.390 2879.900 924.470 ;
        RECT 2879.300 917.050 2879.440 924.390 ;
        RECT 2879.300 916.970 2879.900 917.050 ;
        RECT 2879.300 916.910 2879.960 916.970 ;
        RECT 2879.700 916.650 2879.960 916.910 ;
        RECT 2881.540 916.650 2881.800 916.970 ;
        RECT 2881.600 722.830 2881.740 916.650 ;
        RECT 2880.160 722.570 2880.420 722.830 ;
        RECT 2879.300 722.510 2880.420 722.570 ;
        RECT 2881.540 722.510 2881.800 722.830 ;
        RECT 2879.300 722.430 2880.360 722.510 ;
        RECT 2879.300 702.170 2879.440 722.430 ;
        RECT 2879.300 702.030 2880.360 702.170 ;
        RECT 2880.220 685.430 2880.360 702.030 ;
        RECT 2880.160 685.110 2880.420 685.430 ;
        RECT 2879.700 684.770 2879.960 685.090 ;
        RECT 2879.760 684.490 2879.900 684.770 ;
        RECT 2879.300 684.350 2879.900 684.490 ;
        RECT 2879.300 659.840 2879.440 684.350 ;
        RECT 2879.300 659.700 2879.900 659.840 ;
        RECT 2879.760 652.790 2879.900 659.700 ;
        RECT 2879.700 652.470 2879.960 652.790 ;
        RECT 2881.540 603.510 2881.800 603.830 ;
        RECT 2881.600 545.600 2881.740 603.510 ;
        RECT 2881.600 545.460 2882.200 545.600 ;
        RECT 2882.060 520.870 2882.200 545.460 ;
        RECT 2879.700 520.610 2879.960 520.870 ;
        RECT 2879.300 520.550 2879.960 520.610 ;
        RECT 2882.000 520.550 2882.260 520.870 ;
        RECT 2879.300 520.470 2879.900 520.550 ;
        RECT 2879.300 467.570 2879.440 520.470 ;
        RECT 2879.300 467.430 2880.820 467.570 ;
        RECT 2880.680 443.090 2880.820 467.430 ;
        RECT 2879.300 442.950 2880.820 443.090 ;
        RECT 2879.300 406.880 2879.440 442.950 ;
        RECT 2879.700 406.880 2879.960 406.970 ;
        RECT 2879.300 406.740 2879.960 406.880 ;
        RECT 2879.700 406.650 2879.960 406.740 ;
        RECT 2879.700 360.810 2879.960 361.070 ;
        RECT 2879.300 360.750 2879.960 360.810 ;
        RECT 2879.300 360.670 2879.900 360.750 ;
        RECT 2879.300 294.000 2879.440 360.670 ;
        RECT 2879.700 294.000 2879.960 294.090 ;
        RECT 2879.300 293.860 2879.960 294.000 ;
        RECT 2879.700 293.770 2879.960 293.860 ;
        RECT 2881.540 286.290 2881.800 286.610 ;
        RECT 2881.600 143.470 2881.740 286.290 ;
        RECT 2880.160 143.150 2880.420 143.470 ;
        RECT 2881.540 143.150 2881.800 143.470 ;
        RECT 2880.220 107.090 2880.360 143.150 ;
        RECT 2880.160 106.770 2880.420 107.090 ;
        RECT 2881.540 106.770 2881.800 107.090 ;
        RECT 2881.600 101.730 2881.740 106.770 ;
        RECT 2881.140 101.590 2881.740 101.730 ;
        RECT 2881.140 38.750 2881.280 101.590 ;
        RECT 294.040 38.430 294.300 38.750 ;
        RECT 2881.080 38.430 2881.340 38.750 ;
        RECT 294.100 2.400 294.240 38.430 ;
        RECT 293.890 -4.800 294.450 2.400 ;
      LAYER via2 ;
        RECT 2881.530 1622.000 2881.810 1622.280 ;
      LAYER met3 ;
        RECT 2881.000 1624.880 2885.000 1625.480 ;
        RECT 2881.750 1622.305 2882.050 1624.880 ;
        RECT 2881.505 1621.990 2882.050 1622.305 ;
        RECT 2881.505 1621.975 2881.835 1621.990 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 311.950 25.060 312.270 25.120 ;
        RECT 2299.610 25.060 2299.930 25.120 ;
        RECT 311.950 24.920 2299.930 25.060 ;
        RECT 311.950 24.860 312.270 24.920 ;
        RECT 2299.610 24.860 2299.930 24.920 ;
      LAYER via ;
        RECT 311.980 24.860 312.240 25.120 ;
        RECT 2299.640 24.860 2299.900 25.120 ;
      LAYER met2 ;
        RECT 2299.670 35.000 2299.950 39.000 ;
        RECT 2299.700 25.150 2299.840 35.000 ;
        RECT 311.980 24.830 312.240 25.150 ;
        RECT 2299.640 24.830 2299.900 25.150 ;
        RECT 312.040 2.400 312.180 24.830 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 32.270 31.860 32.590 31.920 ;
        RECT 329.890 31.860 330.210 31.920 ;
        RECT 32.270 31.720 330.210 31.860 ;
        RECT 32.270 31.660 32.590 31.720 ;
        RECT 329.890 31.660 330.210 31.720 ;
      LAYER via ;
        RECT 32.300 31.660 32.560 31.920 ;
        RECT 329.920 31.660 330.180 31.920 ;
      LAYER met2 ;
        RECT 32.290 1621.955 32.570 1622.325 ;
        RECT 32.360 31.950 32.500 1621.955 ;
        RECT 32.300 31.630 32.560 31.950 ;
        RECT 329.920 31.630 330.180 31.950 ;
        RECT 329.980 2.400 330.120 31.630 ;
        RECT 329.770 -4.800 330.330 2.400 ;
      LAYER via2 ;
        RECT 32.290 1622.000 32.570 1622.280 ;
      LAYER met3 ;
        RECT 35.000 1624.880 39.000 1625.480 ;
        RECT 32.265 1622.290 32.595 1622.305 ;
        RECT 35.270 1622.290 35.570 1624.880 ;
        RECT 32.265 1621.990 35.570 1622.290 ;
        RECT 32.265 1621.975 32.595 1621.990 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2880.205 1531.785 2880.375 1579.895 ;
        RECT 2880.205 1351.585 2880.375 1361.615 ;
        RECT 2880.205 1215.585 2880.375 1287.495 ;
        RECT 2880.205 1079.925 2880.375 1087.575 ;
        RECT 2880.665 685.865 2880.835 748.595 ;
        RECT 2880.205 521.305 2880.375 570.095 ;
        RECT 2880.205 373.745 2880.375 397.375 ;
        RECT 2880.205 289.935 2880.375 337.875 ;
        RECT 2880.205 289.765 2880.835 289.935 ;
        RECT 2880.665 286.535 2880.835 289.765 ;
        RECT 2879.745 286.365 2880.835 286.535 ;
        RECT 2879.745 217.345 2879.915 286.365 ;
        RECT 2880.205 169.065 2880.375 176.715 ;
        RECT 347.445 37.485 347.615 39.015 ;
      LAYER mcon ;
        RECT 2880.205 1579.725 2880.375 1579.895 ;
        RECT 2880.205 1361.445 2880.375 1361.615 ;
        RECT 2880.205 1287.325 2880.375 1287.495 ;
        RECT 2880.205 1087.405 2880.375 1087.575 ;
        RECT 2880.665 748.425 2880.835 748.595 ;
        RECT 2880.205 569.925 2880.375 570.095 ;
        RECT 2880.205 397.205 2880.375 397.375 ;
        RECT 2880.205 337.705 2880.375 337.875 ;
        RECT 2880.205 176.545 2880.375 176.715 ;
        RECT 347.445 38.845 347.615 39.015 ;
      LAYER met1 ;
        RECT 2880.590 1628.500 2880.910 1628.560 ;
        RECT 2881.050 1628.500 2881.370 1628.560 ;
        RECT 2880.590 1628.360 2881.370 1628.500 ;
        RECT 2880.590 1628.300 2880.910 1628.360 ;
        RECT 2881.050 1628.300 2881.370 1628.360 ;
        RECT 2880.145 1579.880 2880.435 1579.925 ;
        RECT 2880.590 1579.880 2880.910 1579.940 ;
        RECT 2880.145 1579.740 2880.910 1579.880 ;
        RECT 2880.145 1579.695 2880.435 1579.740 ;
        RECT 2880.590 1579.680 2880.910 1579.740 ;
        RECT 2880.130 1531.940 2880.450 1532.000 ;
        RECT 2879.935 1531.800 2880.450 1531.940 ;
        RECT 2880.130 1531.740 2880.450 1531.800 ;
        RECT 2880.130 1432.120 2880.450 1432.380 ;
        RECT 2880.220 1431.360 2880.360 1432.120 ;
        RECT 2880.130 1431.100 2880.450 1431.360 ;
        RECT 2880.130 1361.600 2880.450 1361.660 ;
        RECT 2880.130 1361.460 2880.645 1361.600 ;
        RECT 2880.130 1361.400 2880.450 1361.460 ;
        RECT 2880.130 1351.740 2880.450 1351.800 ;
        RECT 2880.130 1351.600 2880.645 1351.740 ;
        RECT 2880.130 1351.540 2880.450 1351.600 ;
        RECT 2879.670 1287.480 2879.990 1287.540 ;
        RECT 2880.145 1287.480 2880.435 1287.525 ;
        RECT 2879.670 1287.340 2880.435 1287.480 ;
        RECT 2879.670 1287.280 2879.990 1287.340 ;
        RECT 2880.145 1287.295 2880.435 1287.340 ;
        RECT 2880.130 1215.740 2880.450 1215.800 ;
        RECT 2879.935 1215.600 2880.450 1215.740 ;
        RECT 2880.130 1215.540 2880.450 1215.600 ;
        RECT 2880.130 1207.040 2880.450 1207.300 ;
        RECT 2880.220 1206.220 2880.360 1207.040 ;
        RECT 2880.590 1206.220 2880.910 1206.280 ;
        RECT 2880.220 1206.080 2880.910 1206.220 ;
        RECT 2880.590 1206.020 2880.910 1206.080 ;
        RECT 2880.130 1087.560 2880.450 1087.620 ;
        RECT 2879.935 1087.420 2880.450 1087.560 ;
        RECT 2880.130 1087.360 2880.450 1087.420 ;
        RECT 2879.670 1080.080 2879.990 1080.140 ;
        RECT 2880.145 1080.080 2880.435 1080.125 ;
        RECT 2879.670 1079.940 2880.435 1080.080 ;
        RECT 2879.670 1079.880 2879.990 1079.940 ;
        RECT 2880.145 1079.895 2880.435 1079.940 ;
        RECT 2880.130 748.580 2880.450 748.640 ;
        RECT 2880.605 748.580 2880.895 748.625 ;
        RECT 2880.130 748.440 2880.895 748.580 ;
        RECT 2880.130 748.380 2880.450 748.440 ;
        RECT 2880.605 748.395 2880.895 748.440 ;
        RECT 2879.670 686.020 2879.990 686.080 ;
        RECT 2880.605 686.020 2880.895 686.065 ;
        RECT 2879.670 685.880 2880.895 686.020 ;
        RECT 2879.670 685.820 2879.990 685.880 ;
        RECT 2880.605 685.835 2880.895 685.880 ;
        RECT 2879.670 608.160 2879.990 608.220 ;
        RECT 2880.590 608.160 2880.910 608.220 ;
        RECT 2879.670 608.020 2880.910 608.160 ;
        RECT 2879.670 607.960 2879.990 608.020 ;
        RECT 2880.590 607.960 2880.910 608.020 ;
        RECT 2879.670 570.080 2879.990 570.140 ;
        RECT 2880.145 570.080 2880.435 570.125 ;
        RECT 2879.670 569.940 2880.435 570.080 ;
        RECT 2879.670 569.880 2879.990 569.940 ;
        RECT 2880.145 569.895 2880.435 569.940 ;
        RECT 2879.670 521.460 2879.990 521.520 ;
        RECT 2880.145 521.460 2880.435 521.505 ;
        RECT 2879.670 521.320 2880.435 521.460 ;
        RECT 2879.670 521.260 2879.990 521.320 ;
        RECT 2880.145 521.275 2880.435 521.320 ;
        RECT 2879.670 397.360 2879.990 397.420 ;
        RECT 2880.145 397.360 2880.435 397.405 ;
        RECT 2879.670 397.220 2880.435 397.360 ;
        RECT 2879.670 397.160 2879.990 397.220 ;
        RECT 2880.145 397.175 2880.435 397.220 ;
        RECT 2880.130 373.900 2880.450 373.960 ;
        RECT 2879.935 373.760 2880.450 373.900 ;
        RECT 2880.130 373.700 2880.450 373.760 ;
        RECT 2880.130 337.860 2880.450 337.920 ;
        RECT 2879.935 337.720 2880.450 337.860 ;
        RECT 2880.130 337.660 2880.450 337.720 ;
        RECT 2879.670 217.500 2879.990 217.560 ;
        RECT 2879.475 217.360 2879.990 217.500 ;
        RECT 2879.670 217.300 2879.990 217.360 ;
        RECT 2879.670 176.700 2879.990 176.760 ;
        RECT 2880.145 176.700 2880.435 176.745 ;
        RECT 2879.670 176.560 2880.435 176.700 ;
        RECT 2879.670 176.500 2879.990 176.560 ;
        RECT 2880.145 176.515 2880.435 176.560 ;
        RECT 2879.670 169.220 2879.990 169.280 ;
        RECT 2880.145 169.220 2880.435 169.265 ;
        RECT 2879.670 169.080 2880.435 169.220 ;
        RECT 2879.670 169.020 2879.990 169.080 ;
        RECT 2880.145 169.035 2880.435 169.080 ;
        RECT 2879.670 102.920 2879.990 102.980 ;
        RECT 2880.590 102.920 2880.910 102.980 ;
        RECT 2879.670 102.780 2880.910 102.920 ;
        RECT 2879.670 102.720 2879.990 102.780 ;
        RECT 2880.590 102.720 2880.910 102.780 ;
        RECT 347.385 39.000 347.675 39.045 ;
        RECT 2880.590 39.000 2880.910 39.060 ;
        RECT 347.385 38.860 2880.910 39.000 ;
        RECT 347.385 38.815 347.675 38.860 ;
        RECT 2880.590 38.800 2880.910 38.860 ;
        RECT 347.370 37.640 347.690 37.700 ;
        RECT 347.175 37.500 347.690 37.640 ;
        RECT 347.370 37.440 347.690 37.500 ;
      LAYER via ;
        RECT 2880.620 1628.300 2880.880 1628.560 ;
        RECT 2881.080 1628.300 2881.340 1628.560 ;
        RECT 2880.620 1579.680 2880.880 1579.940 ;
        RECT 2880.160 1531.740 2880.420 1532.000 ;
        RECT 2880.160 1432.120 2880.420 1432.380 ;
        RECT 2880.160 1431.100 2880.420 1431.360 ;
        RECT 2880.160 1361.400 2880.420 1361.660 ;
        RECT 2880.160 1351.540 2880.420 1351.800 ;
        RECT 2879.700 1287.280 2879.960 1287.540 ;
        RECT 2880.160 1215.540 2880.420 1215.800 ;
        RECT 2880.160 1207.040 2880.420 1207.300 ;
        RECT 2880.620 1206.020 2880.880 1206.280 ;
        RECT 2880.160 1087.360 2880.420 1087.620 ;
        RECT 2879.700 1079.880 2879.960 1080.140 ;
        RECT 2880.160 748.380 2880.420 748.640 ;
        RECT 2879.700 685.820 2879.960 686.080 ;
        RECT 2879.700 607.960 2879.960 608.220 ;
        RECT 2880.620 607.960 2880.880 608.220 ;
        RECT 2879.700 569.880 2879.960 570.140 ;
        RECT 2879.700 521.260 2879.960 521.520 ;
        RECT 2879.700 397.160 2879.960 397.420 ;
        RECT 2880.160 373.700 2880.420 373.960 ;
        RECT 2880.160 337.660 2880.420 337.920 ;
        RECT 2879.700 217.300 2879.960 217.560 ;
        RECT 2879.700 176.500 2879.960 176.760 ;
        RECT 2879.700 169.020 2879.960 169.280 ;
        RECT 2879.700 102.720 2879.960 102.980 ;
        RECT 2880.620 102.720 2880.880 102.980 ;
        RECT 2880.620 38.800 2880.880 39.060 ;
        RECT 347.400 37.440 347.660 37.700 ;
      LAYER met2 ;
        RECT 2881.530 1731.690 2881.810 1731.805 ;
        RECT 2881.140 1731.550 2881.810 1731.690 ;
        RECT 2881.140 1628.590 2881.280 1731.550 ;
        RECT 2881.530 1731.435 2881.810 1731.550 ;
        RECT 2880.620 1628.270 2880.880 1628.590 ;
        RECT 2881.080 1628.270 2881.340 1628.590 ;
        RECT 2880.680 1579.970 2880.820 1628.270 ;
        RECT 2880.620 1579.650 2880.880 1579.970 ;
        RECT 2880.160 1531.710 2880.420 1532.030 ;
        RECT 2880.220 1432.410 2880.360 1531.710 ;
        RECT 2880.160 1432.090 2880.420 1432.410 ;
        RECT 2880.160 1431.070 2880.420 1431.390 ;
        RECT 2880.220 1361.690 2880.360 1431.070 ;
        RECT 2880.160 1361.370 2880.420 1361.690 ;
        RECT 2880.160 1351.510 2880.420 1351.830 ;
        RECT 2880.220 1314.170 2880.360 1351.510 ;
        RECT 2878.840 1314.030 2880.360 1314.170 ;
        RECT 2878.840 1287.650 2878.980 1314.030 ;
        RECT 2878.840 1287.570 2879.900 1287.650 ;
        RECT 2878.840 1287.510 2879.960 1287.570 ;
        RECT 2879.700 1287.250 2879.960 1287.510 ;
        RECT 2880.160 1215.510 2880.420 1215.830 ;
        RECT 2880.220 1207.330 2880.360 1215.510 ;
        RECT 2880.160 1207.010 2880.420 1207.330 ;
        RECT 2880.620 1205.990 2880.880 1206.310 ;
        RECT 2880.680 1125.130 2880.820 1205.990 ;
        RECT 2880.220 1124.990 2880.820 1125.130 ;
        RECT 2880.220 1087.650 2880.360 1124.990 ;
        RECT 2880.160 1087.330 2880.420 1087.650 ;
        RECT 2879.700 1079.850 2879.960 1080.170 ;
        RECT 2879.760 1078.210 2879.900 1079.850 ;
        RECT 2877.460 1078.070 2879.900 1078.210 ;
        RECT 2877.460 1077.530 2877.600 1078.070 ;
        RECT 2876.540 1077.390 2877.600 1077.530 ;
        RECT 2876.540 1019.730 2876.680 1077.390 ;
        RECT 2876.540 1019.590 2878.060 1019.730 ;
        RECT 2877.920 932.010 2878.060 1019.590 ;
        RECT 2876.540 931.870 2878.060 932.010 ;
        RECT 2876.540 887.130 2876.680 931.870 ;
        RECT 2876.540 886.990 2877.600 887.130 ;
        RECT 2877.460 885.090 2877.600 886.990 ;
        RECT 2877.460 884.950 2880.360 885.090 ;
        RECT 2880.220 876.930 2880.360 884.950 ;
        RECT 2877.460 876.790 2880.360 876.930 ;
        RECT 2877.460 826.610 2877.600 876.790 ;
        RECT 2877.460 826.470 2880.360 826.610 ;
        RECT 2880.220 748.670 2880.360 826.470 ;
        RECT 2880.160 748.350 2880.420 748.670 ;
        RECT 2879.700 685.850 2879.960 686.110 ;
        RECT 2878.840 685.790 2879.960 685.850 ;
        RECT 2878.840 685.710 2879.900 685.790 ;
        RECT 2878.840 640.970 2878.980 685.710 ;
        RECT 2878.840 640.830 2880.820 640.970 ;
        RECT 2880.680 608.250 2880.820 640.830 ;
        RECT 2879.700 608.160 2879.960 608.250 ;
        RECT 2874.700 608.020 2879.960 608.160 ;
        RECT 2874.700 570.250 2874.840 608.020 ;
        RECT 2879.700 607.930 2879.960 608.020 ;
        RECT 2880.620 607.930 2880.880 608.250 ;
        RECT 2874.700 570.170 2879.900 570.250 ;
        RECT 2874.700 570.110 2879.960 570.170 ;
        RECT 2879.700 569.850 2879.960 570.110 ;
        RECT 2879.700 521.290 2879.960 521.550 ;
        RECT 2878.840 521.230 2879.960 521.290 ;
        RECT 2878.840 521.150 2879.900 521.230 ;
        RECT 2878.840 466.890 2878.980 521.150 ;
        RECT 2878.840 466.750 2880.360 466.890 ;
        RECT 2880.220 452.610 2880.360 466.750 ;
        RECT 2878.840 452.470 2880.360 452.610 ;
        RECT 2878.840 397.530 2878.980 452.470 ;
        RECT 2878.840 397.450 2879.900 397.530 ;
        RECT 2878.840 397.390 2879.960 397.450 ;
        RECT 2879.700 397.130 2879.960 397.390 ;
        RECT 2880.160 373.670 2880.420 373.990 ;
        RECT 2880.220 337.950 2880.360 373.670 ;
        RECT 2880.160 337.630 2880.420 337.950 ;
        RECT 2879.700 217.500 2879.960 217.590 ;
        RECT 2878.840 217.360 2879.960 217.500 ;
        RECT 2878.840 207.810 2878.980 217.360 ;
        RECT 2879.700 217.270 2879.960 217.360 ;
        RECT 2877.460 207.670 2878.980 207.810 ;
        RECT 2877.460 186.050 2877.600 207.670 ;
        RECT 2877.460 185.910 2878.980 186.050 ;
        RECT 2878.840 184.690 2878.980 185.910 ;
        RECT 2878.840 184.550 2879.900 184.690 ;
        RECT 2879.760 176.790 2879.900 184.550 ;
        RECT 2879.700 176.470 2879.960 176.790 ;
        RECT 2879.700 169.220 2879.960 169.310 ;
        RECT 2879.300 169.080 2879.960 169.220 ;
        RECT 2879.300 105.130 2879.440 169.080 ;
        RECT 2879.700 168.990 2879.960 169.080 ;
        RECT 2879.300 104.990 2879.900 105.130 ;
        RECT 2879.760 103.010 2879.900 104.990 ;
        RECT 2879.700 102.690 2879.960 103.010 ;
        RECT 2880.620 102.690 2880.880 103.010 ;
        RECT 2880.680 39.090 2880.820 102.690 ;
        RECT 2880.620 38.770 2880.880 39.090 ;
        RECT 347.400 37.410 347.660 37.730 ;
        RECT 347.460 2.400 347.600 37.410 ;
        RECT 347.250 -4.800 347.810 2.400 ;
      LAYER via2 ;
        RECT 2881.530 1731.480 2881.810 1731.760 ;
      LAYER met3 ;
        RECT 2881.000 1734.360 2885.000 1734.960 ;
        RECT 2881.750 1731.785 2882.050 1734.360 ;
        RECT 2881.505 1731.470 2882.050 1731.785 ;
        RECT 2881.505 1731.455 2881.835 1731.470 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 365.310 31.860 365.630 31.920 ;
        RECT 2886.110 31.860 2886.430 31.920 ;
        RECT 365.310 31.720 2886.430 31.860 ;
        RECT 365.310 31.660 365.630 31.720 ;
        RECT 2886.110 31.660 2886.430 31.720 ;
      LAYER via ;
        RECT 365.340 31.660 365.600 31.920 ;
        RECT 2886.140 31.660 2886.400 31.920 ;
      LAYER met2 ;
        RECT 2886.130 1843.975 2886.410 1844.345 ;
        RECT 2886.200 31.950 2886.340 1843.975 ;
        RECT 365.340 31.630 365.600 31.950 ;
        RECT 2886.140 31.630 2886.400 31.950 ;
        RECT 365.400 2.400 365.540 31.630 ;
        RECT 365.190 -4.800 365.750 2.400 ;
      LAYER via2 ;
        RECT 2886.130 1844.020 2886.410 1844.300 ;
      LAYER met3 ;
        RECT 2881.000 1844.310 2885.000 1844.440 ;
        RECT 2886.105 1844.310 2886.435 1844.325 ;
        RECT 2881.000 1844.010 2886.435 1844.310 ;
        RECT 2881.000 1843.840 2885.000 1844.010 ;
        RECT 2886.105 1843.995 2886.435 1844.010 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 383.250 18.260 383.570 18.320 ;
        RECT 2350.210 18.260 2350.530 18.320 ;
        RECT 383.250 18.120 2350.530 18.260 ;
        RECT 383.250 18.060 383.570 18.120 ;
        RECT 2350.210 18.060 2350.530 18.120 ;
      LAYER via ;
        RECT 383.280 18.060 383.540 18.320 ;
        RECT 2350.240 18.060 2350.500 18.320 ;
      LAYER met2 ;
        RECT 2350.270 35.000 2350.550 39.000 ;
        RECT 2350.300 18.350 2350.440 35.000 ;
        RECT 383.280 18.030 383.540 18.350 ;
        RECT 2350.240 18.030 2350.500 18.350 ;
        RECT 383.340 2.400 383.480 18.030 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 401.190 24.720 401.510 24.780 ;
        RECT 2401.270 24.720 2401.590 24.780 ;
        RECT 401.190 24.580 2401.590 24.720 ;
        RECT 401.190 24.520 401.510 24.580 ;
        RECT 2401.270 24.520 2401.590 24.580 ;
      LAYER via ;
        RECT 401.220 24.520 401.480 24.780 ;
        RECT 2401.300 24.520 2401.560 24.780 ;
      LAYER met2 ;
        RECT 2401.330 35.000 2401.610 39.000 ;
        RECT 2401.360 24.810 2401.500 35.000 ;
        RECT 401.220 24.490 401.480 24.810 ;
        RECT 2401.300 24.490 2401.560 24.810 ;
        RECT 401.280 2.400 401.420 24.490 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 37.330 20.980 37.650 21.040 ;
        RECT 62.170 20.980 62.490 21.040 ;
        RECT 37.330 20.840 62.490 20.980 ;
        RECT 37.330 20.780 37.650 20.840 ;
        RECT 62.170 20.780 62.490 20.840 ;
      LAYER via ;
        RECT 37.360 20.780 37.620 21.040 ;
        RECT 62.200 20.780 62.460 21.040 ;
      LAYER met2 ;
        RECT 37.350 1182.675 37.630 1183.045 ;
        RECT 37.420 21.070 37.560 1182.675 ;
        RECT 37.360 20.750 37.620 21.070 ;
        RECT 62.200 20.750 62.460 21.070 ;
        RECT 62.260 2.400 62.400 20.750 ;
        RECT 62.050 -4.800 62.610 2.400 ;
      LAYER via2 ;
        RECT 37.350 1182.720 37.630 1183.000 ;
      LAYER met3 ;
        RECT 35.000 1185.600 39.000 1186.200 ;
        RECT 37.110 1183.025 37.410 1185.600 ;
        RECT 37.110 1182.710 37.655 1183.025 ;
        RECT 37.325 1182.695 37.655 1182.710 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 419.130 32.540 419.450 32.600 ;
        RECT 2885.650 32.540 2885.970 32.600 ;
        RECT 419.130 32.400 2885.970 32.540 ;
        RECT 419.130 32.340 419.450 32.400 ;
        RECT 2885.650 32.340 2885.970 32.400 ;
      LAYER via ;
        RECT 419.160 32.340 419.420 32.600 ;
        RECT 2885.680 32.340 2885.940 32.600 ;
      LAYER met2 ;
        RECT 2885.670 1953.455 2885.950 1953.825 ;
        RECT 2885.740 32.630 2885.880 1953.455 ;
        RECT 419.160 32.310 419.420 32.630 ;
        RECT 2885.680 32.310 2885.940 32.630 ;
        RECT 419.220 2.400 419.360 32.310 ;
        RECT 419.010 -4.800 419.570 2.400 ;
      LAYER via2 ;
        RECT 2885.670 1953.500 2885.950 1953.780 ;
      LAYER met3 ;
        RECT 2881.000 1953.790 2885.000 1953.920 ;
        RECT 2885.645 1953.790 2885.975 1953.805 ;
        RECT 2881.000 1953.490 2885.975 1953.790 ;
        RECT 2881.000 1953.320 2885.000 1953.490 ;
        RECT 2885.645 1953.475 2885.975 1953.490 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 436.610 17.920 436.930 17.980 ;
        RECT 2452.330 17.920 2452.650 17.980 ;
        RECT 436.610 17.780 2452.650 17.920 ;
        RECT 436.610 17.720 436.930 17.780 ;
        RECT 2452.330 17.720 2452.650 17.780 ;
      LAYER via ;
        RECT 436.640 17.720 436.900 17.980 ;
        RECT 2452.360 17.720 2452.620 17.980 ;
      LAYER met2 ;
        RECT 2452.390 35.000 2452.670 39.000 ;
        RECT 2452.420 18.010 2452.560 35.000 ;
        RECT 436.640 17.690 436.900 18.010 ;
        RECT 2452.360 17.690 2452.620 18.010 ;
        RECT 436.700 2.400 436.840 17.690 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 454.550 32.880 454.870 32.940 ;
        RECT 2885.190 32.880 2885.510 32.940 ;
        RECT 454.550 32.740 2885.510 32.880 ;
        RECT 454.550 32.680 454.870 32.740 ;
        RECT 2885.190 32.680 2885.510 32.740 ;
      LAYER via ;
        RECT 454.580 32.680 454.840 32.940 ;
        RECT 2885.220 32.680 2885.480 32.940 ;
      LAYER met2 ;
        RECT 2885.210 2062.595 2885.490 2062.965 ;
        RECT 2885.280 32.970 2885.420 2062.595 ;
        RECT 454.580 32.650 454.840 32.970 ;
        RECT 2885.220 32.650 2885.480 32.970 ;
        RECT 454.640 2.400 454.780 32.650 ;
        RECT 454.430 -4.800 454.990 2.400 ;
      LAYER via2 ;
        RECT 2885.210 2062.640 2885.490 2062.920 ;
      LAYER met3 ;
        RECT 2881.000 2063.480 2885.000 2064.080 ;
        RECT 2884.510 2062.930 2884.810 2063.480 ;
        RECT 2885.185 2062.930 2885.515 2062.945 ;
        RECT 2884.510 2062.630 2885.515 2062.930 ;
        RECT 2885.185 2062.615 2885.515 2062.630 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 472.490 30.500 472.810 30.560 ;
        RECT 2884.730 30.500 2885.050 30.560 ;
        RECT 472.490 30.360 2885.050 30.500 ;
        RECT 472.490 30.300 472.810 30.360 ;
        RECT 2884.730 30.300 2885.050 30.360 ;
      LAYER via ;
        RECT 472.520 30.300 472.780 30.560 ;
        RECT 2884.760 30.300 2885.020 30.560 ;
      LAYER met2 ;
        RECT 2884.750 2170.035 2885.030 2170.405 ;
        RECT 2884.820 30.590 2884.960 2170.035 ;
        RECT 472.520 30.270 472.780 30.590 ;
        RECT 2884.760 30.270 2885.020 30.590 ;
        RECT 472.580 2.400 472.720 30.270 ;
        RECT 472.370 -4.800 472.930 2.400 ;
      LAYER via2 ;
        RECT 2884.750 2170.080 2885.030 2170.360 ;
      LAYER met3 ;
        RECT 2881.000 2172.960 2885.000 2173.560 ;
        RECT 2884.510 2170.385 2884.810 2172.960 ;
        RECT 2884.510 2170.070 2885.055 2170.385 ;
        RECT 2884.725 2170.055 2885.055 2170.070 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 490.430 24.380 490.750 24.440 ;
        RECT 2502.930 24.380 2503.250 24.440 ;
        RECT 490.430 24.240 2503.250 24.380 ;
        RECT 490.430 24.180 490.750 24.240 ;
        RECT 2502.930 24.180 2503.250 24.240 ;
      LAYER via ;
        RECT 490.460 24.180 490.720 24.440 ;
        RECT 2502.960 24.180 2503.220 24.440 ;
      LAYER met2 ;
        RECT 2502.990 35.000 2503.270 39.000 ;
        RECT 2503.020 24.470 2503.160 35.000 ;
        RECT 490.460 24.150 490.720 24.470 ;
        RECT 2502.960 24.150 2503.220 24.470 ;
        RECT 490.520 2.400 490.660 24.150 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 507.910 30.160 508.230 30.220 ;
        RECT 2884.270 30.160 2884.590 30.220 ;
        RECT 507.910 30.020 2884.590 30.160 ;
        RECT 507.910 29.960 508.230 30.020 ;
        RECT 2884.270 29.960 2884.590 30.020 ;
      LAYER via ;
        RECT 507.940 29.960 508.200 30.220 ;
        RECT 2884.300 29.960 2884.560 30.220 ;
      LAYER met2 ;
        RECT 2884.290 2279.515 2884.570 2279.885 ;
        RECT 2884.360 30.250 2884.500 2279.515 ;
        RECT 507.940 29.930 508.200 30.250 ;
        RECT 2884.300 29.930 2884.560 30.250 ;
        RECT 508.000 2.400 508.140 29.930 ;
        RECT 507.790 -4.800 508.350 2.400 ;
      LAYER via2 ;
        RECT 2884.290 2279.560 2884.570 2279.840 ;
      LAYER met3 ;
        RECT 2881.000 2282.440 2885.000 2283.040 ;
        RECT 2884.510 2279.865 2884.810 2282.440 ;
        RECT 2884.265 2279.550 2884.810 2279.865 ;
        RECT 2884.265 2279.535 2884.595 2279.550 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 75.970 26.420 76.290 26.480 ;
        RECT 521.250 26.420 521.570 26.480 ;
        RECT 75.970 26.280 521.570 26.420 ;
        RECT 75.970 26.220 76.290 26.280 ;
        RECT 521.250 26.220 521.570 26.280 ;
        RECT 521.250 19.280 521.570 19.340 ;
        RECT 525.850 19.280 526.170 19.340 ;
        RECT 521.250 19.140 526.170 19.280 ;
        RECT 521.250 19.080 521.570 19.140 ;
        RECT 525.850 19.080 526.170 19.140 ;
      LAYER via ;
        RECT 76.000 26.220 76.260 26.480 ;
        RECT 521.280 26.220 521.540 26.480 ;
        RECT 521.280 19.080 521.540 19.340 ;
        RECT 525.880 19.080 526.140 19.340 ;
      LAYER met2 ;
        RECT 1622.970 3432.370 1623.250 3432.485 ;
        RECT 1624.390 3432.370 1624.670 3435.000 ;
        RECT 1622.970 3432.230 1624.670 3432.370 ;
        RECT 1622.970 3432.115 1623.250 3432.230 ;
        RECT 1624.390 3431.000 1624.670 3432.230 ;
        RECT 75.990 36.875 76.270 37.245 ;
        RECT 76.060 26.510 76.200 36.875 ;
        RECT 76.000 26.190 76.260 26.510 ;
        RECT 521.280 26.190 521.540 26.510 ;
        RECT 521.340 19.370 521.480 26.190 ;
        RECT 521.280 19.050 521.540 19.370 ;
        RECT 525.880 19.050 526.140 19.370 ;
        RECT 525.940 2.400 526.080 19.050 ;
        RECT 525.730 -4.800 526.290 2.400 ;
      LAYER via2 ;
        RECT 1622.970 3432.160 1623.250 3432.440 ;
        RECT 75.990 36.920 76.270 37.200 ;
      LAYER met3 ;
        RECT 831.950 3435.850 832.330 3435.860 ;
        RECT 888.070 3435.850 888.450 3435.860 ;
        RECT 831.950 3435.550 888.450 3435.850 ;
        RECT 831.950 3435.540 832.330 3435.550 ;
        RECT 888.070 3435.540 888.450 3435.550 ;
        RECT 1014.110 3435.850 1014.490 3435.860 ;
        RECT 1061.950 3435.850 1062.330 3435.860 ;
        RECT 1014.110 3435.550 1062.330 3435.850 ;
        RECT 1014.110 3435.540 1014.490 3435.550 ;
        RECT 1061.950 3435.540 1062.330 3435.550 ;
        RECT 1152.110 3435.850 1152.490 3435.860 ;
        RECT 1176.030 3435.850 1176.410 3435.860 ;
        RECT 1152.110 3435.550 1176.410 3435.850 ;
        RECT 1152.110 3435.540 1152.490 3435.550 ;
        RECT 1176.030 3435.540 1176.410 3435.550 ;
        RECT 50.870 3432.450 51.250 3432.460 ;
        RECT 62.830 3432.450 63.210 3432.460 ;
        RECT 50.870 3432.150 63.210 3432.450 ;
        RECT 50.870 3432.140 51.250 3432.150 ;
        RECT 62.830 3432.140 63.210 3432.150 ;
        RECT 475.910 3432.450 476.290 3432.460 ;
        RECT 499.830 3432.450 500.210 3432.460 ;
        RECT 475.910 3432.150 500.210 3432.450 ;
        RECT 475.910 3432.140 476.290 3432.150 ;
        RECT 499.830 3432.140 500.210 3432.150 ;
        RECT 1200.870 3432.450 1201.250 3432.460 ;
        RECT 1247.790 3432.450 1248.170 3432.460 ;
        RECT 1200.870 3432.150 1248.170 3432.450 ;
        RECT 1200.870 3432.140 1201.250 3432.150 ;
        RECT 1247.790 3432.140 1248.170 3432.150 ;
        RECT 1622.230 3432.450 1622.610 3432.460 ;
        RECT 1622.945 3432.450 1623.275 3432.465 ;
        RECT 1622.230 3432.150 1623.275 3432.450 ;
        RECT 1622.230 3432.140 1622.610 3432.150 ;
        RECT 1622.945 3432.135 1623.275 3432.150 ;
        RECT 911.070 3431.770 911.450 3431.780 ;
        RECT 931.310 3431.770 931.690 3431.780 ;
        RECT 911.070 3431.470 931.690 3431.770 ;
        RECT 911.070 3431.460 911.450 3431.470 ;
        RECT 931.310 3431.460 931.690 3431.470 ;
        RECT 50.870 37.210 51.250 37.220 ;
        RECT 75.965 37.210 76.295 37.225 ;
        RECT 50.870 36.910 76.295 37.210 ;
        RECT 50.870 36.900 51.250 36.910 ;
        RECT 75.965 36.895 76.295 36.910 ;
      LAYER via3 ;
        RECT 831.980 3435.540 832.300 3435.860 ;
        RECT 888.100 3435.540 888.420 3435.860 ;
        RECT 1014.140 3435.540 1014.460 3435.860 ;
        RECT 1061.980 3435.540 1062.300 3435.860 ;
        RECT 1152.140 3435.540 1152.460 3435.860 ;
        RECT 1176.060 3435.540 1176.380 3435.860 ;
        RECT 50.900 3432.140 51.220 3432.460 ;
        RECT 62.860 3432.140 63.180 3432.460 ;
        RECT 475.940 3432.140 476.260 3432.460 ;
        RECT 499.860 3432.140 500.180 3432.460 ;
        RECT 1200.900 3432.140 1201.220 3432.460 ;
        RECT 1247.820 3432.140 1248.140 3432.460 ;
        RECT 1622.260 3432.140 1622.580 3432.460 ;
        RECT 911.100 3431.460 911.420 3431.780 ;
        RECT 931.340 3431.460 931.660 3431.780 ;
        RECT 50.900 36.900 51.220 37.220 ;
      LAYER met4 ;
        RECT 831.975 3435.535 832.305 3435.865 ;
        RECT 888.095 3435.535 888.425 3435.865 ;
        RECT 831.990 3432.890 832.290 3435.535 ;
        RECT 50.895 3432.135 51.225 3432.465 ;
        RECT 50.910 37.225 51.210 3432.135 ;
        RECT 62.430 3431.710 63.610 3432.890 ;
        RECT 475.935 3432.135 476.265 3432.465 ;
        RECT 475.950 3429.490 476.250 3432.135 ;
        RECT 499.430 3431.710 500.610 3432.890 ;
        RECT 831.550 3431.710 832.730 3432.890 ;
        RECT 888.110 3429.490 888.410 3435.535 ;
        RECT 1013.710 3435.110 1014.890 3436.290 ;
        RECT 1061.975 3435.535 1062.305 3435.865 ;
        RECT 1061.990 3432.890 1062.290 3435.535 ;
        RECT 1151.710 3435.110 1152.890 3436.290 ;
        RECT 1176.055 3435.535 1176.385 3435.865 ;
        RECT 911.095 3431.455 911.425 3431.785 ;
        RECT 931.335 3431.455 931.665 3431.785 ;
        RECT 1061.550 3431.710 1062.730 3432.890 ;
        RECT 911.110 3429.490 911.410 3431.455 ;
        RECT 931.350 3429.490 931.650 3431.455 ;
        RECT 1176.070 3429.490 1176.370 3435.535 ;
        RECT 1200.895 3432.135 1201.225 3432.465 ;
        RECT 1200.910 3429.490 1201.210 3432.135 ;
        RECT 1247.390 3431.710 1248.570 3432.890 ;
        RECT 1621.830 3431.710 1623.010 3432.890 ;
        RECT 64.270 3429.050 65.450 3429.490 ;
        RECT 95.550 3429.050 96.730 3429.490 ;
        RECT 64.270 3428.750 96.730 3429.050 ;
        RECT 64.270 3428.310 65.450 3428.750 ;
        RECT 95.550 3428.310 96.730 3428.750 ;
        RECT 475.510 3428.310 476.690 3429.490 ;
        RECT 887.670 3428.310 888.850 3429.490 ;
        RECT 910.670 3428.310 911.850 3429.490 ;
        RECT 930.910 3428.310 932.090 3429.490 ;
        RECT 975.990 3429.050 977.170 3429.490 ;
        RECT 979.670 3429.050 980.850 3429.490 ;
        RECT 975.990 3428.750 980.850 3429.050 ;
        RECT 975.990 3428.310 977.170 3428.750 ;
        RECT 979.670 3428.310 980.850 3428.750 ;
        RECT 1175.630 3428.310 1176.810 3429.490 ;
        RECT 1200.470 3428.310 1201.650 3429.490 ;
        RECT 50.895 36.895 51.225 37.225 ;
      LAYER met5 ;
        RECT 979.460 3434.900 1015.100 3436.500 ;
        RECT 1122.980 3434.900 1153.100 3436.500 ;
        RECT 61.300 3431.500 63.820 3433.100 ;
        RECT 61.300 3429.700 62.900 3431.500 ;
        RECT 156.980 3429.700 159.500 3433.100 ;
        RECT 253.580 3429.700 256.100 3433.100 ;
        RECT 350.180 3429.700 352.700 3433.100 ;
        RECT 446.780 3429.700 449.300 3433.100 ;
        RECT 499.220 3431.500 545.900 3433.100 ;
        RECT 544.300 3429.700 545.900 3431.500 ;
        RECT 639.980 3429.700 642.500 3433.100 ;
        RECT 736.580 3429.700 739.100 3433.100 ;
        RECT 831.340 3429.700 832.940 3433.100 ;
        RECT 61.300 3428.100 65.660 3429.700 ;
        RECT 95.340 3428.100 476.900 3429.700 ;
        RECT 544.300 3428.100 832.940 3429.700 ;
        RECT 887.460 3428.100 912.060 3429.700 ;
        RECT 930.700 3428.100 977.380 3429.700 ;
        RECT 979.460 3428.100 981.060 3434.900 ;
        RECT 1122.980 3433.100 1124.580 3434.900 ;
        RECT 1061.340 3431.500 1077.660 3433.100 ;
        RECT 1076.060 3429.700 1077.660 3431.500 ;
        RECT 1121.140 3431.500 1124.580 3433.100 ;
        RECT 1247.180 3431.500 1270.860 3433.100 ;
        RECT 1121.140 3429.700 1122.740 3431.500 ;
        RECT 1269.260 3429.700 1270.860 3431.500 ;
        RECT 1316.180 3431.500 1367.460 3433.100 ;
        RECT 1316.180 3429.700 1317.780 3431.500 ;
        RECT 1076.060 3428.100 1122.740 3429.700 ;
        RECT 1175.420 3428.100 1201.860 3429.700 ;
        RECT 1269.260 3428.100 1317.780 3429.700 ;
        RECT 1365.860 3429.700 1367.460 3431.500 ;
        RECT 1412.780 3431.500 1464.060 3433.100 ;
        RECT 1412.780 3429.700 1414.380 3431.500 ;
        RECT 1365.860 3428.100 1414.380 3429.700 ;
        RECT 1462.460 3429.700 1464.060 3431.500 ;
        RECT 1509.380 3431.500 1560.660 3433.100 ;
        RECT 1509.380 3429.700 1510.980 3431.500 ;
        RECT 1462.460 3428.100 1510.980 3429.700 ;
        RECT 1559.060 3429.700 1560.660 3431.500 ;
        RECT 1604.140 3431.500 1623.220 3433.100 ;
        RECT 1604.140 3429.700 1605.740 3431.500 ;
        RECT 1559.060 3428.100 1605.740 3429.700 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 35.950 28.800 36.270 28.860 ;
        RECT 543.790 28.800 544.110 28.860 ;
        RECT 35.950 28.660 544.110 28.800 ;
        RECT 35.950 28.600 36.270 28.660 ;
        RECT 543.790 28.600 544.110 28.660 ;
      LAYER via ;
        RECT 35.980 28.600 36.240 28.860 ;
        RECT 543.820 28.600 544.080 28.860 ;
      LAYER met2 ;
        RECT 35.970 1732.115 36.250 1732.485 ;
        RECT 36.040 28.890 36.180 1732.115 ;
        RECT 35.980 28.570 36.240 28.890 ;
        RECT 543.820 28.570 544.080 28.890 ;
        RECT 543.880 2.400 544.020 28.570 ;
        RECT 543.670 -4.800 544.230 2.400 ;
      LAYER via2 ;
        RECT 35.970 1732.160 36.250 1732.440 ;
      LAYER met3 ;
        RECT 35.000 1734.360 39.000 1734.960 ;
        RECT 36.190 1732.465 36.490 1734.360 ;
        RECT 35.945 1732.150 36.490 1732.465 ;
        RECT 35.945 1732.135 36.275 1732.150 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 70.910 26.760 71.230 26.820 ;
        RECT 496.870 26.760 497.190 26.820 ;
        RECT 70.910 26.620 497.190 26.760 ;
        RECT 70.910 26.560 71.230 26.620 ;
        RECT 496.870 26.560 497.190 26.620 ;
        RECT 496.870 19.620 497.190 19.680 ;
        RECT 561.730 19.620 562.050 19.680 ;
        RECT 496.870 19.480 562.050 19.620 ;
        RECT 496.870 19.420 497.190 19.480 ;
        RECT 561.730 19.420 562.050 19.480 ;
      LAYER via ;
        RECT 70.940 26.560 71.200 26.820 ;
        RECT 496.900 26.560 497.160 26.820 ;
        RECT 496.900 19.420 497.160 19.680 ;
        RECT 561.760 19.420 562.020 19.680 ;
      LAYER met2 ;
        RECT 1733.830 3443.675 1734.110 3444.045 ;
        RECT 1733.900 3435.000 1734.040 3443.675 ;
        RECT 1733.870 3431.000 1734.150 3435.000 ;
        RECT 70.930 38.235 71.210 38.605 ;
        RECT 71.000 26.850 71.140 38.235 ;
        RECT 70.940 26.530 71.200 26.850 ;
        RECT 496.900 26.530 497.160 26.850 ;
        RECT 496.960 19.710 497.100 26.530 ;
        RECT 496.900 19.390 497.160 19.710 ;
        RECT 561.760 19.390 562.020 19.710 ;
        RECT 561.820 2.400 561.960 19.390 ;
        RECT 561.610 -4.800 562.170 2.400 ;
      LAYER via2 ;
        RECT 1733.830 3443.720 1734.110 3444.000 ;
        RECT 70.930 38.280 71.210 38.560 ;
      LAYER met3 ;
        RECT 1704.110 3444.010 1704.490 3444.020 ;
        RECT 1733.805 3444.010 1734.135 3444.025 ;
        RECT 1704.110 3443.710 1734.135 3444.010 ;
        RECT 1704.110 3443.700 1704.490 3443.710 ;
        RECT 1733.805 3443.695 1734.135 3443.710 ;
        RECT 469.470 3431.770 469.850 3431.780 ;
        RECT 516.390 3431.770 516.770 3431.780 ;
        RECT 469.470 3431.470 516.770 3431.770 ;
        RECT 469.470 3431.460 469.850 3431.470 ;
        RECT 516.390 3431.460 516.770 3431.470 ;
        RECT 541.230 3431.770 541.610 3431.780 ;
        RECT 565.150 3431.770 565.530 3431.780 ;
        RECT 541.230 3431.470 565.530 3431.770 ;
        RECT 541.230 3431.460 541.610 3431.470 ;
        RECT 565.150 3431.460 565.530 3431.470 ;
        RECT 1703.190 3431.770 1703.570 3431.780 ;
        RECT 1704.110 3431.770 1704.490 3431.780 ;
        RECT 1703.190 3431.470 1704.490 3431.770 ;
        RECT 1703.190 3431.460 1703.570 3431.470 ;
        RECT 1704.110 3431.460 1704.490 3431.470 ;
        RECT 52.710 38.570 53.090 38.580 ;
        RECT 70.905 38.570 71.235 38.585 ;
        RECT 52.710 38.270 71.235 38.570 ;
        RECT 52.710 38.260 53.090 38.270 ;
        RECT 70.905 38.255 71.235 38.270 ;
      LAYER via3 ;
        RECT 1704.140 3443.700 1704.460 3444.020 ;
        RECT 469.500 3431.460 469.820 3431.780 ;
        RECT 516.420 3431.460 516.740 3431.780 ;
        RECT 541.260 3431.460 541.580 3431.780 ;
        RECT 565.180 3431.460 565.500 3431.780 ;
        RECT 1703.220 3431.460 1703.540 3431.780 ;
        RECT 1704.140 3431.460 1704.460 3431.780 ;
        RECT 52.740 38.260 53.060 38.580 ;
      LAYER met4 ;
        RECT 1704.135 3443.695 1704.465 3444.025 ;
        RECT 1704.150 3431.785 1704.450 3443.695 ;
        RECT 469.495 3431.455 469.825 3431.785 ;
        RECT 516.415 3431.455 516.745 3431.785 ;
        RECT 541.255 3431.455 541.585 3431.785 ;
        RECT 565.175 3431.455 565.505 3431.785 ;
        RECT 1703.215 3431.455 1703.545 3431.785 ;
        RECT 1704.135 3431.455 1704.465 3431.785 ;
        RECT 469.510 3426.090 469.810 3431.455 ;
        RECT 516.430 3426.090 516.730 3431.455 ;
        RECT 541.270 3429.490 541.570 3431.455 ;
        RECT 540.830 3428.310 542.010 3429.490 ;
        RECT 565.190 3426.090 565.490 3431.455 ;
        RECT 1703.230 3429.490 1703.530 3431.455 ;
        RECT 835.230 3429.050 836.410 3429.490 ;
        RECT 820.950 3428.750 836.410 3429.050 ;
        RECT 820.950 3426.090 821.250 3428.750 ;
        RECT 835.230 3428.310 836.410 3428.750 ;
        RECT 1702.790 3428.310 1703.970 3429.490 ;
        RECT 469.070 3424.910 470.250 3426.090 ;
        RECT 515.990 3424.910 517.170 3426.090 ;
        RECT 564.750 3424.910 565.930 3426.090 ;
        RECT 820.510 3424.910 821.690 3426.090 ;
        RECT 52.310 3421.510 53.490 3422.690 ;
        RECT 52.750 38.585 53.050 3421.510 ;
        RECT 52.735 38.255 53.065 38.585 ;
      LAYER met5 ;
        RECT 516.700 3428.100 542.220 3429.700 ;
        RECT 835.020 3428.100 868.820 3429.700 ;
        RECT 516.700 3426.300 518.300 3428.100 ;
        RECT 61.300 3424.700 470.460 3426.300 ;
        RECT 61.300 3422.900 62.900 3424.700 ;
        RECT 52.100 3421.300 62.900 3422.900 ;
        RECT 156.980 3421.300 159.500 3424.700 ;
        RECT 253.580 3421.300 256.100 3424.700 ;
        RECT 350.180 3421.300 352.700 3424.700 ;
        RECT 446.780 3421.300 449.300 3424.700 ;
        RECT 515.780 3421.300 518.300 3426.300 ;
        RECT 564.540 3422.900 566.140 3426.300 ;
        RECT 612.380 3424.700 821.900 3426.300 ;
        RECT 612.380 3422.900 613.980 3424.700 ;
        RECT 564.540 3421.300 613.980 3422.900 ;
        RECT 736.580 3421.300 739.100 3424.700 ;
        RECT 867.220 3419.500 868.820 3428.100 ;
        RECT 984.060 3428.100 1027.060 3429.700 ;
        RECT 885.620 3424.700 929.540 3426.300 ;
        RECT 885.620 3422.900 887.220 3424.700 ;
        RECT 882.860 3421.300 887.220 3422.900 ;
        RECT 927.940 3422.900 929.540 3424.700 ;
        RECT 933.460 3424.700 967.260 3426.300 ;
        RECT 933.460 3422.900 935.060 3424.700 ;
        RECT 927.940 3421.300 935.060 3422.900 ;
        RECT 882.860 3419.500 884.460 3421.300 ;
        RECT 867.220 3417.900 884.460 3419.500 ;
        RECT 929.780 3417.900 932.300 3421.300 ;
        RECT 965.660 3419.500 967.260 3424.700 ;
        RECT 984.060 3419.500 985.660 3428.100 ;
        RECT 1025.460 3426.300 1027.060 3428.100 ;
        RECT 1610.580 3428.100 1704.180 3429.700 ;
        RECT 1025.460 3424.700 1028.900 3426.300 ;
        RECT 1027.300 3422.900 1028.900 3424.700 ;
        RECT 1076.060 3424.700 1124.580 3426.300 ;
        RECT 1076.060 3422.900 1077.660 3424.700 ;
        RECT 1027.300 3421.300 1077.660 3422.900 ;
        RECT 1122.980 3422.900 1124.580 3424.700 ;
        RECT 1172.660 3424.700 1221.180 3426.300 ;
        RECT 1172.660 3422.900 1174.260 3424.700 ;
        RECT 1122.980 3421.300 1174.260 3422.900 ;
        RECT 1219.580 3422.900 1221.180 3424.700 ;
        RECT 1302.380 3424.700 1317.780 3426.300 ;
        RECT 1219.580 3421.300 1257.060 3422.900 ;
        RECT 965.660 3417.900 985.660 3419.500 ;
        RECT 1255.460 3416.100 1257.060 3421.300 ;
        RECT 1302.380 3416.100 1303.980 3424.700 ;
        RECT 1316.180 3422.900 1317.780 3424.700 ;
        RECT 1398.980 3424.700 1414.380 3426.300 ;
        RECT 1316.180 3421.300 1353.660 3422.900 ;
        RECT 1255.460 3414.500 1303.980 3416.100 ;
        RECT 1352.060 3416.100 1353.660 3421.300 ;
        RECT 1398.980 3416.100 1400.580 3424.700 ;
        RECT 1412.780 3422.900 1414.380 3424.700 ;
        RECT 1495.580 3424.700 1510.980 3426.300 ;
        RECT 1412.780 3421.300 1450.260 3422.900 ;
        RECT 1352.060 3414.500 1400.580 3416.100 ;
        RECT 1448.660 3416.100 1450.260 3421.300 ;
        RECT 1495.580 3416.100 1497.180 3424.700 ;
        RECT 1509.380 3422.900 1510.980 3424.700 ;
        RECT 1592.180 3424.700 1605.740 3426.300 ;
        RECT 1509.380 3421.300 1546.860 3422.900 ;
        RECT 1448.660 3414.500 1497.180 3416.100 ;
        RECT 1545.260 3416.100 1546.860 3421.300 ;
        RECT 1592.180 3416.100 1593.780 3424.700 ;
        RECT 1604.140 3422.900 1605.740 3424.700 ;
        RECT 1610.580 3422.900 1612.180 3428.100 ;
        RECT 1604.140 3421.300 1612.180 3422.900 ;
        RECT 1545.260 3414.500 1593.780 3416.100 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 35.490 29.480 35.810 29.540 ;
        RECT 579.670 29.480 579.990 29.540 ;
        RECT 35.490 29.340 579.990 29.480 ;
        RECT 35.490 29.280 35.810 29.340 ;
        RECT 579.670 29.280 579.990 29.340 ;
      LAYER via ;
        RECT 35.520 29.280 35.780 29.540 ;
        RECT 579.700 29.280 579.960 29.540 ;
      LAYER met2 ;
        RECT 35.510 1842.275 35.790 1842.645 ;
        RECT 35.580 29.570 35.720 1842.275 ;
        RECT 35.520 29.250 35.780 29.570 ;
        RECT 579.700 29.250 579.960 29.570 ;
        RECT 579.760 2.400 579.900 29.250 ;
        RECT 579.550 -4.800 580.110 2.400 ;
      LAYER via2 ;
        RECT 35.510 1842.320 35.790 1842.600 ;
      LAYER met3 ;
        RECT 35.000 1843.840 39.000 1844.440 ;
        RECT 35.270 1842.625 35.570 1843.840 ;
        RECT 35.270 1842.310 35.815 1842.625 ;
        RECT 35.485 1842.295 35.815 1842.310 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 46.990 3445.460 47.310 3445.520 ;
        RECT 1404.910 3445.460 1405.230 3445.520 ;
        RECT 46.990 3445.320 1405.230 3445.460 ;
        RECT 46.990 3445.260 47.310 3445.320 ;
        RECT 1404.910 3445.260 1405.230 3445.320 ;
        RECT 46.990 38.660 47.310 38.720 ;
        RECT 86.090 38.660 86.410 38.720 ;
        RECT 46.990 38.520 86.410 38.660 ;
        RECT 46.990 38.460 47.310 38.520 ;
        RECT 86.090 38.460 86.410 38.520 ;
      LAYER via ;
        RECT 47.020 3445.260 47.280 3445.520 ;
        RECT 1404.940 3445.260 1405.200 3445.520 ;
        RECT 47.020 38.460 47.280 38.720 ;
        RECT 86.120 38.460 86.380 38.720 ;
      LAYER met2 ;
        RECT 47.020 3445.230 47.280 3445.550 ;
        RECT 1404.940 3445.230 1405.200 3445.550 ;
        RECT 47.080 38.750 47.220 3445.230 ;
        RECT 1405.000 3435.000 1405.140 3445.230 ;
        RECT 1404.970 3431.000 1405.250 3435.000 ;
        RECT 47.020 38.430 47.280 38.750 ;
        RECT 86.120 38.430 86.380 38.750 ;
        RECT 86.180 2.400 86.320 38.430 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 597.150 29.480 597.470 29.540 ;
        RECT 2893.930 29.480 2894.250 29.540 ;
        RECT 597.150 29.340 2894.250 29.480 ;
        RECT 597.150 29.280 597.470 29.340 ;
        RECT 2893.930 29.280 2894.250 29.340 ;
      LAYER via ;
        RECT 597.180 29.280 597.440 29.540 ;
        RECT 2893.960 29.280 2894.220 29.540 ;
      LAYER met2 ;
        RECT 2893.950 2389.675 2894.230 2390.045 ;
        RECT 2894.020 29.570 2894.160 2389.675 ;
        RECT 597.180 29.250 597.440 29.570 ;
        RECT 2893.960 29.250 2894.220 29.570 ;
        RECT 597.240 2.400 597.380 29.250 ;
        RECT 597.030 -4.800 597.590 2.400 ;
      LAYER via2 ;
        RECT 2893.950 2389.720 2894.230 2390.000 ;
      LAYER met3 ;
        RECT 2881.000 2392.600 2885.000 2393.200 ;
        RECT 2884.510 2390.010 2884.810 2392.600 ;
        RECT 2893.925 2390.010 2894.255 2390.025 ;
        RECT 2884.510 2389.710 2894.255 2390.010 ;
        RECT 2893.925 2389.695 2894.255 2389.710 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 46.530 3432.540 46.850 3432.600 ;
        RECT 1841.910 3432.540 1842.230 3432.600 ;
        RECT 46.530 3432.400 1842.230 3432.540 ;
        RECT 46.530 3432.340 46.850 3432.400 ;
        RECT 1841.910 3432.340 1842.230 3432.400 ;
        RECT 46.530 29.140 46.850 29.200 ;
        RECT 615.090 29.140 615.410 29.200 ;
        RECT 46.530 29.000 615.410 29.140 ;
        RECT 46.530 28.940 46.850 29.000 ;
        RECT 615.090 28.940 615.410 29.000 ;
      LAYER via ;
        RECT 46.560 3432.340 46.820 3432.600 ;
        RECT 1841.940 3432.340 1842.200 3432.600 ;
        RECT 46.560 28.940 46.820 29.200 ;
        RECT 615.120 28.940 615.380 29.200 ;
      LAYER met2 ;
        RECT 46.560 3432.310 46.820 3432.630 ;
        RECT 1841.940 3432.370 1842.200 3432.630 ;
        RECT 1843.350 3432.370 1843.630 3435.000 ;
        RECT 1841.940 3432.310 1843.630 3432.370 ;
        RECT 46.620 29.230 46.760 3432.310 ;
        RECT 1842.000 3432.230 1843.630 3432.310 ;
        RECT 1843.350 3431.000 1843.630 3432.230 ;
        RECT 46.560 28.910 46.820 29.230 ;
        RECT 615.120 28.910 615.380 29.230 ;
        RECT 615.180 2.400 615.320 28.910 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 109.550 30.840 109.870 30.900 ;
        RECT 2894.850 30.840 2895.170 30.900 ;
        RECT 109.550 30.700 2895.170 30.840 ;
        RECT 109.550 30.640 109.870 30.700 ;
        RECT 2894.850 30.640 2895.170 30.700 ;
      LAYER via ;
        RECT 109.580 30.640 109.840 30.900 ;
        RECT 2894.880 30.640 2895.140 30.900 ;
      LAYER met2 ;
        RECT 2894.870 1402.315 2895.150 1402.685 ;
        RECT 2894.940 30.930 2895.080 1402.315 ;
        RECT 109.580 30.610 109.840 30.930 ;
        RECT 2894.880 30.610 2895.140 30.930 ;
        RECT 109.640 2.400 109.780 30.610 ;
        RECT 109.430 -4.800 109.990 2.400 ;
      LAYER via2 ;
        RECT 2894.870 1402.360 2895.150 1402.640 ;
      LAYER met3 ;
        RECT 2881.000 1405.240 2885.000 1405.840 ;
        RECT 2884.510 1402.650 2884.810 1405.240 ;
        RECT 2894.845 1402.650 2895.175 1402.665 ;
        RECT 2884.510 1402.350 2895.175 1402.650 ;
        RECT 2894.845 1402.335 2895.175 1402.350 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 36.870 25.060 37.190 25.120 ;
        RECT 133.470 25.060 133.790 25.120 ;
        RECT 36.870 24.920 133.790 25.060 ;
        RECT 36.870 24.860 37.190 24.920 ;
        RECT 133.470 24.860 133.790 24.920 ;
      LAYER via ;
        RECT 36.900 24.860 37.160 25.120 ;
        RECT 133.500 24.860 133.760 25.120 ;
      LAYER met2 ;
        RECT 36.890 1292.835 37.170 1293.205 ;
        RECT 36.960 25.150 37.100 1292.835 ;
        RECT 36.900 24.830 37.160 25.150 ;
        RECT 133.500 24.830 133.760 25.150 ;
        RECT 133.560 2.400 133.700 24.830 ;
        RECT 133.350 -4.800 133.910 2.400 ;
      LAYER via2 ;
        RECT 36.890 1292.880 37.170 1293.160 ;
      LAYER met3 ;
        RECT 35.000 1295.760 39.000 1296.360 ;
        RECT 37.110 1293.185 37.410 1295.760 ;
        RECT 36.865 1292.870 37.410 1293.185 ;
        RECT 36.865 1292.855 37.195 1292.870 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 151.410 31.180 151.730 31.240 ;
        RECT 2894.390 31.180 2894.710 31.240 ;
        RECT 151.410 31.040 2894.710 31.180 ;
        RECT 151.410 30.980 151.730 31.040 ;
        RECT 2894.390 30.980 2894.710 31.040 ;
      LAYER via ;
        RECT 151.440 30.980 151.700 31.240 ;
        RECT 2894.420 30.980 2894.680 31.240 ;
      LAYER met2 ;
        RECT 2894.410 1513.155 2894.690 1513.525 ;
        RECT 2894.480 31.270 2894.620 1513.155 ;
        RECT 151.440 30.950 151.700 31.270 ;
        RECT 2894.420 30.950 2894.680 31.270 ;
        RECT 151.500 2.400 151.640 30.950 ;
        RECT 151.290 -4.800 151.850 2.400 ;
      LAYER via2 ;
        RECT 2894.410 1513.200 2894.690 1513.480 ;
      LAYER met3 ;
        RECT 2881.000 1514.720 2885.000 1515.320 ;
        RECT 2884.510 1513.490 2884.810 1514.720 ;
        RECT 2894.385 1513.490 2894.715 1513.505 ;
        RECT 2884.510 1513.190 2894.715 1513.490 ;
        RECT 2894.385 1513.175 2894.715 1513.190 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 36.410 24.720 36.730 24.780 ;
        RECT 169.350 24.720 169.670 24.780 ;
        RECT 36.410 24.580 169.670 24.720 ;
        RECT 36.410 24.520 36.730 24.580 ;
        RECT 169.350 24.520 169.670 24.580 ;
      LAYER via ;
        RECT 36.440 24.520 36.700 24.780 ;
        RECT 169.380 24.520 169.640 24.780 ;
      LAYER met2 ;
        RECT 36.430 1402.315 36.710 1402.685 ;
        RECT 36.500 24.810 36.640 1402.315 ;
        RECT 36.440 24.490 36.700 24.810 ;
        RECT 169.380 24.490 169.640 24.810 ;
        RECT 169.440 2.400 169.580 24.490 ;
        RECT 169.230 -4.800 169.790 2.400 ;
      LAYER via2 ;
        RECT 36.430 1402.360 36.710 1402.640 ;
      LAYER met3 ;
        RECT 35.000 1405.240 39.000 1405.840 ;
        RECT 36.190 1402.665 36.490 1405.240 ;
        RECT 36.190 1402.350 36.735 1402.665 ;
        RECT 36.405 1402.335 36.735 1402.350 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 186.830 18.940 187.150 19.000 ;
        RECT 2095.830 18.940 2096.150 19.000 ;
        RECT 186.830 18.800 2096.150 18.940 ;
        RECT 186.830 18.740 187.150 18.800 ;
        RECT 2095.830 18.740 2096.150 18.800 ;
      LAYER via ;
        RECT 186.860 18.740 187.120 19.000 ;
        RECT 2095.860 18.740 2096.120 19.000 ;
      LAYER met2 ;
        RECT 2095.890 35.000 2096.170 39.000 ;
        RECT 2095.920 19.030 2096.060 35.000 ;
        RECT 186.860 18.710 187.120 19.030 ;
        RECT 2095.860 18.710 2096.120 19.030 ;
        RECT 186.920 2.400 187.060 18.710 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 31.810 24.040 32.130 24.100 ;
        RECT 204.770 24.040 205.090 24.100 ;
        RECT 31.810 23.900 205.090 24.040 ;
        RECT 31.810 23.840 32.130 23.900 ;
        RECT 204.770 23.840 205.090 23.900 ;
      LAYER via ;
        RECT 31.840 23.840 32.100 24.100 ;
        RECT 204.800 23.840 205.060 24.100 ;
      LAYER met2 ;
        RECT 31.830 1513.155 32.110 1513.525 ;
        RECT 31.900 24.130 32.040 1513.155 ;
        RECT 31.840 23.810 32.100 24.130 ;
        RECT 204.800 23.810 205.060 24.130 ;
        RECT 204.860 2.400 205.000 23.810 ;
        RECT 204.650 -4.800 205.210 2.400 ;
      LAYER via2 ;
        RECT 31.830 1513.200 32.110 1513.480 ;
      LAYER met3 ;
        RECT 35.000 1514.720 39.000 1515.320 ;
        RECT 31.805 1513.490 32.135 1513.505 ;
        RECT 35.270 1513.490 35.570 1514.720 ;
        RECT 31.805 1513.190 35.570 1513.490 ;
        RECT 31.805 1513.175 32.135 1513.190 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 222.710 18.600 223.030 18.660 ;
        RECT 2146.890 18.600 2147.210 18.660 ;
        RECT 222.710 18.460 2147.210 18.600 ;
        RECT 222.710 18.400 223.030 18.460 ;
        RECT 2146.890 18.400 2147.210 18.460 ;
      LAYER via ;
        RECT 222.740 18.400 223.000 18.660 ;
        RECT 2146.920 18.400 2147.180 18.660 ;
      LAYER met2 ;
        RECT 2146.950 35.000 2147.230 39.000 ;
        RECT 2146.980 18.690 2147.120 35.000 ;
        RECT 222.740 18.370 223.000 18.690 ;
        RECT 2146.920 18.370 2147.180 18.690 ;
        RECT 222.800 2.400 222.940 18.370 ;
        RECT 222.590 -4.800 223.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 44.690 3444.440 45.010 3444.500 ;
        RECT 1953.230 3444.440 1953.550 3444.500 ;
        RECT 44.690 3444.300 1953.550 3444.440 ;
        RECT 44.690 3444.240 45.010 3444.300 ;
        RECT 1953.230 3444.240 1953.550 3444.300 ;
        RECT 20.310 15.540 20.630 15.600 ;
        RECT 44.690 15.540 45.010 15.600 ;
        RECT 20.310 15.400 45.010 15.540 ;
        RECT 20.310 15.340 20.630 15.400 ;
        RECT 44.690 15.340 45.010 15.400 ;
      LAYER via ;
        RECT 44.720 3444.240 44.980 3444.500 ;
        RECT 1953.260 3444.240 1953.520 3444.500 ;
        RECT 20.340 15.340 20.600 15.600 ;
        RECT 44.720 15.340 44.980 15.600 ;
      LAYER met2 ;
        RECT 44.720 3444.210 44.980 3444.530 ;
        RECT 1953.260 3444.210 1953.520 3444.530 ;
        RECT 44.780 15.630 44.920 3444.210 ;
        RECT 1953.320 3435.000 1953.460 3444.210 ;
        RECT 1953.290 3431.000 1953.570 3435.000 ;
        RECT 20.340 15.310 20.600 15.630 ;
        RECT 44.720 15.310 44.980 15.630 ;
        RECT 20.400 2.400 20.540 15.310 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2554.050 35.000 2554.330 39.000 ;
        RECT 2554.080 25.685 2554.220 35.000 ;
        RECT 44.250 25.315 44.530 25.685 ;
        RECT 2554.010 25.315 2554.290 25.685 ;
        RECT 44.320 2.400 44.460 25.315 ;
        RECT 44.110 -4.800 44.670 2.400 ;
      LAYER via2 ;
        RECT 44.250 25.360 44.530 25.640 ;
        RECT 2554.010 25.360 2554.290 25.640 ;
      LAYER met3 ;
        RECT 44.225 25.650 44.555 25.665 ;
        RECT 2553.985 25.650 2554.315 25.665 ;
        RECT 44.225 25.350 2554.315 25.650 ;
        RECT 44.225 25.335 44.555 25.350 ;
        RECT 2553.985 25.335 2554.315 25.350 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 48.370 3444.100 48.690 3444.160 ;
        RECT 2062.710 3444.100 2063.030 3444.160 ;
        RECT 48.370 3443.960 2063.030 3444.100 ;
        RECT 48.370 3443.900 48.690 3443.960 ;
        RECT 2062.710 3443.900 2063.030 3443.960 ;
        RECT 48.370 15.540 48.690 15.600 ;
        RECT 246.630 15.540 246.950 15.600 ;
        RECT 48.370 15.400 246.950 15.540 ;
        RECT 48.370 15.340 48.690 15.400 ;
        RECT 246.630 15.340 246.950 15.400 ;
      LAYER via ;
        RECT 48.400 3443.900 48.660 3444.160 ;
        RECT 2062.740 3443.900 2063.000 3444.160 ;
        RECT 48.400 15.340 48.660 15.600 ;
        RECT 246.660 15.340 246.920 15.600 ;
      LAYER met2 ;
        RECT 48.400 3443.870 48.660 3444.190 ;
        RECT 2062.740 3443.870 2063.000 3444.190 ;
        RECT 48.460 15.630 48.600 3443.870 ;
        RECT 2062.800 3435.000 2062.940 3443.870 ;
        RECT 2062.770 3431.000 2063.050 3435.000 ;
        RECT 48.400 15.310 48.660 15.630 ;
        RECT 246.660 15.310 246.920 15.630 ;
        RECT 246.720 2.400 246.860 15.310 ;
        RECT 246.510 -4.800 247.070 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 264.110 24.040 264.430 24.100 ;
        RECT 2757.770 24.040 2758.090 24.100 ;
        RECT 264.110 23.900 2758.090 24.040 ;
        RECT 264.110 23.840 264.430 23.900 ;
        RECT 2757.770 23.840 2758.090 23.900 ;
      LAYER via ;
        RECT 264.140 23.840 264.400 24.100 ;
        RECT 2757.800 23.840 2758.060 24.100 ;
      LAYER met2 ;
        RECT 2757.830 35.000 2758.110 39.000 ;
        RECT 2757.860 24.130 2758.000 35.000 ;
        RECT 264.140 23.810 264.400 24.130 ;
        RECT 2757.800 23.810 2758.060 24.130 ;
        RECT 264.200 2.400 264.340 23.810 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 47.910 3443.760 48.230 3443.820 ;
        RECT 2172.190 3443.760 2172.510 3443.820 ;
        RECT 47.910 3443.620 2172.510 3443.760 ;
        RECT 47.910 3443.560 48.230 3443.620 ;
        RECT 2172.190 3443.560 2172.510 3443.620 ;
        RECT 47.910 16.220 48.230 16.280 ;
        RECT 282.050 16.220 282.370 16.280 ;
        RECT 47.910 16.080 282.370 16.220 ;
        RECT 47.910 16.020 48.230 16.080 ;
        RECT 282.050 16.020 282.370 16.080 ;
      LAYER via ;
        RECT 47.940 3443.560 48.200 3443.820 ;
        RECT 2172.220 3443.560 2172.480 3443.820 ;
        RECT 47.940 16.020 48.200 16.280 ;
        RECT 282.080 16.020 282.340 16.280 ;
      LAYER met2 ;
        RECT 47.940 3443.530 48.200 3443.850 ;
        RECT 2172.220 3443.530 2172.480 3443.850 ;
        RECT 48.000 16.310 48.140 3443.530 ;
        RECT 2172.280 3435.000 2172.420 3443.530 ;
        RECT 2172.250 3431.000 2172.530 3435.000 ;
        RECT 47.940 15.990 48.200 16.310 ;
        RECT 282.080 15.990 282.340 16.310 ;
        RECT 282.140 2.400 282.280 15.990 ;
        RECT 281.930 -4.800 282.490 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 47.450 3447.160 47.770 3447.220 ;
        RECT 2282.130 3447.160 2282.450 3447.220 ;
        RECT 47.450 3447.020 2282.450 3447.160 ;
        RECT 47.450 3446.960 47.770 3447.020 ;
        RECT 2282.130 3446.960 2282.450 3447.020 ;
        RECT 47.450 16.560 47.770 16.620 ;
        RECT 299.990 16.560 300.310 16.620 ;
        RECT 47.450 16.420 300.310 16.560 ;
        RECT 47.450 16.360 47.770 16.420 ;
        RECT 299.990 16.360 300.310 16.420 ;
      LAYER via ;
        RECT 47.480 3446.960 47.740 3447.220 ;
        RECT 2282.160 3446.960 2282.420 3447.220 ;
        RECT 47.480 16.360 47.740 16.620 ;
        RECT 300.020 16.360 300.280 16.620 ;
      LAYER met2 ;
        RECT 47.480 3446.930 47.740 3447.250 ;
        RECT 2282.160 3446.930 2282.420 3447.250 ;
        RECT 47.540 16.650 47.680 3446.930 ;
        RECT 2282.220 3435.000 2282.360 3446.930 ;
        RECT 2282.190 3431.000 2282.470 3435.000 ;
        RECT 47.480 16.330 47.740 16.650 ;
        RECT 300.020 16.330 300.280 16.650 ;
        RECT 300.080 2.400 300.220 16.330 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 317.930 31.520 318.250 31.580 ;
        RECT 2893.010 31.520 2893.330 31.580 ;
        RECT 317.930 31.380 2893.330 31.520 ;
        RECT 317.930 31.320 318.250 31.380 ;
        RECT 2893.010 31.320 2893.330 31.380 ;
      LAYER via ;
        RECT 317.960 31.320 318.220 31.580 ;
        RECT 2893.040 31.320 2893.300 31.580 ;
      LAYER met2 ;
        RECT 2893.030 2719.475 2893.310 2719.845 ;
        RECT 2893.100 31.610 2893.240 2719.475 ;
        RECT 317.960 31.290 318.220 31.610 ;
        RECT 2893.040 31.290 2893.300 31.610 ;
        RECT 318.020 2.400 318.160 31.290 ;
        RECT 317.810 -4.800 318.370 2.400 ;
      LAYER via2 ;
        RECT 2893.030 2719.520 2893.310 2719.800 ;
      LAYER met3 ;
        RECT 2881.000 2721.040 2885.000 2721.640 ;
        RECT 2884.510 2719.810 2884.810 2721.040 ;
        RECT 2893.005 2719.810 2893.335 2719.825 ;
        RECT 2884.510 2719.510 2893.335 2719.810 ;
        RECT 2893.005 2719.495 2893.335 2719.510 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 34.570 24.380 34.890 24.440 ;
        RECT 335.870 24.380 336.190 24.440 ;
        RECT 34.570 24.240 336.190 24.380 ;
        RECT 34.570 24.180 34.890 24.240 ;
        RECT 335.870 24.180 336.190 24.240 ;
      LAYER via ;
        RECT 34.600 24.180 34.860 24.440 ;
        RECT 335.900 24.180 336.160 24.440 ;
      LAYER met2 ;
        RECT 34.590 2389.675 34.870 2390.045 ;
        RECT 34.660 24.470 34.800 2389.675 ;
        RECT 34.600 24.150 34.860 24.470 ;
        RECT 335.900 24.150 336.160 24.470 ;
        RECT 335.960 2.400 336.100 24.150 ;
        RECT 335.750 -4.800 336.310 2.400 ;
      LAYER via2 ;
        RECT 34.590 2389.720 34.870 2390.000 ;
      LAYER met3 ;
        RECT 35.000 2392.600 39.000 2393.200 ;
        RECT 34.565 2390.010 34.895 2390.025 ;
        RECT 35.270 2390.010 35.570 2392.600 ;
        RECT 34.565 2389.710 35.570 2390.010 ;
        RECT 34.565 2389.695 34.895 2389.710 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 24.910 16.900 25.230 16.960 ;
        RECT 353.350 16.900 353.670 16.960 ;
        RECT 24.910 16.760 353.670 16.900 ;
        RECT 24.910 16.700 25.230 16.760 ;
        RECT 353.350 16.700 353.670 16.760 ;
      LAYER via ;
        RECT 24.940 16.700 25.200 16.960 ;
        RECT 353.380 16.700 353.640 16.960 ;
      LAYER met2 ;
        RECT 25.390 2499.155 25.670 2499.525 ;
        RECT 25.460 27.610 25.600 2499.155 ;
        RECT 25.000 27.470 25.600 27.610 ;
        RECT 25.000 16.990 25.140 27.470 ;
        RECT 24.940 16.670 25.200 16.990 ;
        RECT 353.380 16.670 353.640 16.990 ;
        RECT 353.440 2.400 353.580 16.670 ;
        RECT 353.230 -4.800 353.790 2.400 ;
      LAYER via2 ;
        RECT 25.390 2499.200 25.670 2499.480 ;
      LAYER met3 ;
        RECT 35.000 2502.080 39.000 2502.680 ;
        RECT 25.365 2499.490 25.695 2499.505 ;
        RECT 35.270 2499.490 35.570 2502.080 ;
        RECT 25.365 2499.190 35.570 2499.490 ;
        RECT 25.365 2499.175 25.695 2499.190 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 25.370 18.260 25.690 18.320 ;
        RECT 371.290 18.260 371.610 18.320 ;
        RECT 25.370 18.120 371.610 18.260 ;
        RECT 25.370 18.060 25.690 18.120 ;
        RECT 371.290 18.060 371.610 18.120 ;
      LAYER via ;
        RECT 25.400 18.060 25.660 18.320 ;
        RECT 371.320 18.060 371.580 18.320 ;
      LAYER met2 ;
        RECT 25.850 2608.635 26.130 2609.005 ;
        RECT 25.920 26.930 26.060 2608.635 ;
        RECT 25.460 26.790 26.060 26.930 ;
        RECT 25.460 18.350 25.600 26.790 ;
        RECT 25.400 18.030 25.660 18.350 ;
        RECT 371.320 18.030 371.580 18.350 ;
        RECT 371.380 2.400 371.520 18.030 ;
        RECT 371.170 -4.800 371.730 2.400 ;
      LAYER via2 ;
        RECT 25.850 2608.680 26.130 2608.960 ;
      LAYER met3 ;
        RECT 35.000 2611.560 39.000 2612.160 ;
        RECT 25.825 2608.970 26.155 2608.985 ;
        RECT 35.270 2608.970 35.570 2611.560 ;
        RECT 25.825 2608.670 35.570 2608.970 ;
        RECT 25.825 2608.655 26.155 2608.670 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 389.230 32.200 389.550 32.260 ;
        RECT 2892.550 32.200 2892.870 32.260 ;
        RECT 389.230 32.060 2892.870 32.200 ;
        RECT 389.230 32.000 389.550 32.060 ;
        RECT 2892.550 32.000 2892.870 32.060 ;
      LAYER via ;
        RECT 389.260 32.000 389.520 32.260 ;
        RECT 2892.580 32.000 2892.840 32.260 ;
      LAYER met2 ;
        RECT 2892.570 2828.955 2892.850 2829.325 ;
        RECT 2892.640 32.290 2892.780 2828.955 ;
        RECT 389.260 31.970 389.520 32.290 ;
        RECT 2892.580 31.970 2892.840 32.290 ;
        RECT 389.320 2.400 389.460 31.970 ;
        RECT 389.110 -4.800 389.670 2.400 ;
      LAYER via2 ;
        RECT 2892.570 2829.000 2892.850 2829.280 ;
      LAYER met3 ;
        RECT 2881.000 2831.200 2885.000 2831.800 ;
        RECT 2884.510 2829.290 2884.810 2831.200 ;
        RECT 2892.545 2829.290 2892.875 2829.305 ;
        RECT 2884.510 2828.990 2892.875 2829.290 ;
        RECT 2892.545 2828.975 2892.875 2828.990 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 25.830 17.920 26.150 17.980 ;
        RECT 407.170 17.920 407.490 17.980 ;
        RECT 25.830 17.780 407.490 17.920 ;
        RECT 25.830 17.720 26.150 17.780 ;
        RECT 407.170 17.720 407.490 17.780 ;
      LAYER via ;
        RECT 25.860 17.720 26.120 17.980 ;
        RECT 407.200 17.720 407.460 17.980 ;
      LAYER met2 ;
        RECT 26.310 2719.475 26.590 2719.845 ;
        RECT 26.380 26.250 26.520 2719.475 ;
        RECT 25.920 26.110 26.520 26.250 ;
        RECT 25.920 18.010 26.060 26.110 ;
        RECT 25.860 17.690 26.120 18.010 ;
        RECT 407.200 17.690 407.460 18.010 ;
        RECT 407.260 2.400 407.400 17.690 ;
        RECT 407.050 -4.800 407.610 2.400 ;
      LAYER via2 ;
        RECT 26.310 2719.520 26.590 2719.800 ;
      LAYER met3 ;
        RECT 35.000 2721.040 39.000 2721.640 ;
        RECT 26.285 2719.810 26.615 2719.825 ;
        RECT 35.270 2719.810 35.570 2721.040 ;
        RECT 26.285 2719.510 35.570 2719.810 ;
        RECT 26.285 2719.495 26.615 2719.510 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 68.150 17.240 68.470 17.300 ;
        RECT 2605.050 17.240 2605.370 17.300 ;
        RECT 68.150 17.100 2605.370 17.240 ;
        RECT 68.150 17.040 68.470 17.100 ;
        RECT 2605.050 17.040 2605.370 17.100 ;
      LAYER via ;
        RECT 68.180 17.040 68.440 17.300 ;
        RECT 2605.080 17.040 2605.340 17.300 ;
      LAYER met2 ;
        RECT 2605.110 35.000 2605.390 39.000 ;
        RECT 2605.140 17.330 2605.280 35.000 ;
        RECT 68.180 17.010 68.440 17.330 ;
        RECT 2605.080 17.010 2605.340 17.330 ;
        RECT 68.240 2.400 68.380 17.010 ;
        RECT 68.030 -4.800 68.590 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2391.630 3442.995 2391.910 3443.365 ;
        RECT 2391.700 3435.000 2391.840 3442.995 ;
        RECT 2391.670 3431.000 2391.950 3435.000 ;
        RECT 424.670 37.555 424.950 37.925 ;
        RECT 424.740 2.400 424.880 37.555 ;
        RECT 424.530 -4.800 425.090 2.400 ;
      LAYER via2 ;
        RECT 2391.630 3443.040 2391.910 3443.320 ;
        RECT 424.670 37.600 424.950 37.880 ;
      LAYER met3 ;
        RECT 54.550 3443.330 54.930 3443.340 ;
        RECT 2391.605 3443.330 2391.935 3443.345 ;
        RECT 54.550 3443.030 2391.935 3443.330 ;
        RECT 54.550 3443.020 54.930 3443.030 ;
        RECT 2391.605 3443.015 2391.935 3443.030 ;
        RECT 54.550 37.890 54.930 37.900 ;
        RECT 424.645 37.890 424.975 37.905 ;
        RECT 54.550 37.590 424.975 37.890 ;
        RECT 54.550 37.580 54.930 37.590 ;
        RECT 424.645 37.575 424.975 37.590 ;
      LAYER via3 ;
        RECT 54.580 3443.020 54.900 3443.340 ;
        RECT 54.580 37.580 54.900 37.900 ;
      LAYER met4 ;
        RECT 54.575 3443.015 54.905 3443.345 ;
        RECT 54.590 37.905 54.890 3443.015 ;
        RECT 54.575 37.575 54.905 37.905 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 32.730 20.640 33.050 20.700 ;
        RECT 442.590 20.640 442.910 20.700 ;
        RECT 32.730 20.500 442.910 20.640 ;
        RECT 32.730 20.440 33.050 20.500 ;
        RECT 442.590 20.440 442.910 20.500 ;
      LAYER via ;
        RECT 32.760 20.440 33.020 20.700 ;
        RECT 442.620 20.440 442.880 20.700 ;
      LAYER met2 ;
        RECT 32.750 2831.335 33.030 2831.705 ;
        RECT 32.820 20.730 32.960 2831.335 ;
        RECT 32.760 20.410 33.020 20.730 ;
        RECT 442.620 20.410 442.880 20.730 ;
        RECT 442.680 2.400 442.820 20.410 ;
        RECT 442.470 -4.800 443.030 2.400 ;
      LAYER via2 ;
        RECT 32.750 2831.380 33.030 2831.660 ;
      LAYER met3 ;
        RECT 32.725 2831.670 33.055 2831.685 ;
        RECT 35.000 2831.670 39.000 2831.800 ;
        RECT 32.725 2831.370 39.000 2831.670 ;
        RECT 32.725 2831.355 33.055 2831.370 ;
        RECT 35.000 2831.200 39.000 2831.370 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 34.645 14.365 34.815 20.315 ;
        RECT 82.485 14.365 82.655 19.975 ;
      LAYER mcon ;
        RECT 34.645 20.145 34.815 20.315 ;
        RECT 82.485 19.805 82.655 19.975 ;
      LAYER met1 ;
        RECT 33.190 20.300 33.510 20.360 ;
        RECT 34.585 20.300 34.875 20.345 ;
        RECT 33.190 20.160 34.875 20.300 ;
        RECT 33.190 20.100 33.510 20.160 ;
        RECT 34.585 20.115 34.875 20.160 ;
        RECT 82.425 19.960 82.715 20.005 ;
        RECT 460.530 19.960 460.850 20.020 ;
        RECT 82.425 19.820 460.850 19.960 ;
        RECT 82.425 19.775 82.715 19.820 ;
        RECT 460.530 19.760 460.850 19.820 ;
        RECT 34.585 14.520 34.875 14.565 ;
        RECT 82.425 14.520 82.715 14.565 ;
        RECT 34.585 14.380 82.715 14.520 ;
        RECT 34.585 14.335 34.875 14.380 ;
        RECT 82.425 14.335 82.715 14.380 ;
      LAYER via ;
        RECT 33.220 20.100 33.480 20.360 ;
        RECT 460.560 19.760 460.820 20.020 ;
      LAYER met2 ;
        RECT 33.210 2940.815 33.490 2941.185 ;
        RECT 33.280 20.390 33.420 2940.815 ;
        RECT 33.220 20.070 33.480 20.390 ;
        RECT 460.560 19.730 460.820 20.050 ;
        RECT 460.620 2.400 460.760 19.730 ;
        RECT 460.410 -4.800 460.970 2.400 ;
      LAYER via2 ;
        RECT 33.210 2940.860 33.490 2941.140 ;
      LAYER met3 ;
        RECT 33.185 2941.150 33.515 2941.165 ;
        RECT 35.000 2941.150 39.000 2941.280 ;
        RECT 33.185 2940.850 39.000 2941.150 ;
        RECT 33.185 2940.835 33.515 2940.850 ;
        RECT 35.000 2940.680 39.000 2940.850 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 32.270 3007.880 32.590 3007.940 ;
        RECT 33.650 3007.880 33.970 3007.940 ;
        RECT 32.270 3007.740 33.970 3007.880 ;
        RECT 32.270 3007.680 32.590 3007.740 ;
        RECT 33.650 3007.680 33.970 3007.740 ;
        RECT 32.270 2959.600 32.590 2959.660 ;
        RECT 33.650 2959.600 33.970 2959.660 ;
        RECT 32.270 2959.460 33.970 2959.600 ;
        RECT 32.270 2959.400 32.590 2959.460 ;
        RECT 33.650 2959.400 33.970 2959.460 ;
        RECT 31.810 2911.320 32.130 2911.380 ;
        RECT 33.650 2911.320 33.970 2911.380 ;
        RECT 31.810 2911.180 33.970 2911.320 ;
        RECT 31.810 2911.120 32.130 2911.180 ;
        RECT 33.650 2911.120 33.970 2911.180 ;
        RECT 31.810 2862.360 32.130 2862.420 ;
        RECT 34.110 2862.360 34.430 2862.420 ;
        RECT 31.810 2862.220 34.430 2862.360 ;
        RECT 31.810 2862.160 32.130 2862.220 ;
        RECT 34.110 2862.160 34.430 2862.220 ;
        RECT 34.110 2816.120 34.430 2816.180 ;
        RECT 32.360 2815.980 34.430 2816.120 ;
        RECT 32.360 2815.500 32.500 2815.980 ;
        RECT 34.110 2815.920 34.430 2815.980 ;
        RECT 32.270 2815.240 32.590 2815.500 ;
        RECT 32.270 2767.160 32.590 2767.220 ;
        RECT 33.650 2767.160 33.970 2767.220 ;
        RECT 32.270 2767.020 33.970 2767.160 ;
        RECT 32.270 2766.960 32.590 2767.020 ;
        RECT 33.650 2766.960 33.970 2767.020 ;
        RECT 32.270 2670.600 32.590 2670.660 ;
        RECT 33.650 2670.600 33.970 2670.660 ;
        RECT 32.270 2670.460 33.970 2670.600 ;
        RECT 32.270 2670.400 32.590 2670.460 ;
        RECT 33.650 2670.400 33.970 2670.460 ;
        RECT 32.270 2574.040 32.590 2574.100 ;
        RECT 33.650 2574.040 33.970 2574.100 ;
        RECT 32.270 2573.900 33.970 2574.040 ;
        RECT 32.270 2573.840 32.590 2573.900 ;
        RECT 33.650 2573.840 33.970 2573.900 ;
        RECT 32.270 2477.480 32.590 2477.540 ;
        RECT 33.650 2477.480 33.970 2477.540 ;
        RECT 32.270 2477.340 33.970 2477.480 ;
        RECT 32.270 2477.280 32.590 2477.340 ;
        RECT 33.650 2477.280 33.970 2477.340 ;
        RECT 32.270 2380.580 32.590 2380.640 ;
        RECT 33.650 2380.580 33.970 2380.640 ;
        RECT 32.270 2380.440 33.970 2380.580 ;
        RECT 32.270 2380.380 32.590 2380.440 ;
        RECT 33.650 2380.380 33.970 2380.440 ;
        RECT 32.270 2284.020 32.590 2284.080 ;
        RECT 33.650 2284.020 33.970 2284.080 ;
        RECT 32.270 2283.880 33.970 2284.020 ;
        RECT 32.270 2283.820 32.590 2283.880 ;
        RECT 33.650 2283.820 33.970 2283.880 ;
        RECT 32.270 2187.460 32.590 2187.520 ;
        RECT 33.650 2187.460 33.970 2187.520 ;
        RECT 32.270 2187.320 33.970 2187.460 ;
        RECT 32.270 2187.260 32.590 2187.320 ;
        RECT 33.650 2187.260 33.970 2187.320 ;
        RECT 32.270 1994.340 32.590 1994.400 ;
        RECT 33.650 1994.340 33.970 1994.400 ;
        RECT 32.270 1994.200 33.970 1994.340 ;
        RECT 32.270 1994.140 32.590 1994.200 ;
        RECT 33.650 1994.140 33.970 1994.200 ;
        RECT 32.270 1945.720 32.590 1945.780 ;
        RECT 33.650 1945.720 33.970 1945.780 ;
        RECT 32.270 1945.580 33.970 1945.720 ;
        RECT 32.270 1945.520 32.590 1945.580 ;
        RECT 33.650 1945.520 33.970 1945.580 ;
        RECT 32.270 1897.780 32.590 1897.840 ;
        RECT 33.650 1897.780 33.970 1897.840 ;
        RECT 32.270 1897.640 33.970 1897.780 ;
        RECT 32.270 1897.580 32.590 1897.640 ;
        RECT 33.650 1897.580 33.970 1897.640 ;
        RECT 32.270 1849.160 32.590 1849.220 ;
        RECT 33.650 1849.160 33.970 1849.220 ;
        RECT 32.270 1849.020 33.970 1849.160 ;
        RECT 32.270 1848.960 32.590 1849.020 ;
        RECT 33.650 1848.960 33.970 1849.020 ;
        RECT 32.270 1801.220 32.590 1801.280 ;
        RECT 33.650 1801.220 33.970 1801.280 ;
        RECT 32.270 1801.080 33.970 1801.220 ;
        RECT 32.270 1801.020 32.590 1801.080 ;
        RECT 33.650 1801.020 33.970 1801.080 ;
        RECT 32.270 1752.600 32.590 1752.660 ;
        RECT 33.650 1752.600 33.970 1752.660 ;
        RECT 32.270 1752.460 33.970 1752.600 ;
        RECT 32.270 1752.400 32.590 1752.460 ;
        RECT 33.650 1752.400 33.970 1752.460 ;
        RECT 32.270 1704.660 32.590 1704.720 ;
        RECT 33.650 1704.660 33.970 1704.720 ;
        RECT 32.270 1704.520 33.970 1704.660 ;
        RECT 32.270 1704.460 32.590 1704.520 ;
        RECT 33.650 1704.460 33.970 1704.520 ;
        RECT 31.810 1656.040 32.130 1656.100 ;
        RECT 33.650 1656.040 33.970 1656.100 ;
        RECT 31.810 1655.900 33.970 1656.040 ;
        RECT 31.810 1655.840 32.130 1655.900 ;
        RECT 33.650 1655.840 33.970 1655.900 ;
        RECT 31.810 1608.100 32.130 1608.160 ;
        RECT 33.650 1608.100 33.970 1608.160 ;
        RECT 31.810 1607.960 33.970 1608.100 ;
        RECT 31.810 1607.900 32.130 1607.960 ;
        RECT 33.650 1607.900 33.970 1607.960 ;
        RECT 30.430 1559.140 30.750 1559.200 ;
        RECT 33.650 1559.140 33.970 1559.200 ;
        RECT 30.430 1559.000 33.970 1559.140 ;
        RECT 30.430 1558.940 30.750 1559.000 ;
        RECT 33.650 1558.940 33.970 1559.000 ;
        RECT 30.430 1511.200 30.750 1511.260 ;
        RECT 33.650 1511.200 33.970 1511.260 ;
        RECT 30.430 1511.060 33.970 1511.200 ;
        RECT 30.430 1511.000 30.750 1511.060 ;
        RECT 33.650 1511.000 33.970 1511.060 ;
        RECT 30.430 1462.580 30.750 1462.640 ;
        RECT 33.650 1462.580 33.970 1462.640 ;
        RECT 30.430 1462.440 33.970 1462.580 ;
        RECT 30.430 1462.380 30.750 1462.440 ;
        RECT 33.650 1462.380 33.970 1462.440 ;
        RECT 30.430 1414.640 30.750 1414.700 ;
        RECT 33.650 1414.640 33.970 1414.700 ;
        RECT 30.430 1414.500 33.970 1414.640 ;
        RECT 30.430 1414.440 30.750 1414.500 ;
        RECT 33.650 1414.440 33.970 1414.500 ;
        RECT 30.430 1366.020 30.750 1366.080 ;
        RECT 33.650 1366.020 33.970 1366.080 ;
        RECT 30.430 1365.880 33.970 1366.020 ;
        RECT 30.430 1365.820 30.750 1365.880 ;
        RECT 33.650 1365.820 33.970 1365.880 ;
        RECT 30.430 1318.080 30.750 1318.140 ;
        RECT 33.650 1318.080 33.970 1318.140 ;
        RECT 30.430 1317.940 33.970 1318.080 ;
        RECT 30.430 1317.880 30.750 1317.940 ;
        RECT 33.650 1317.880 33.970 1317.940 ;
        RECT 30.430 1269.460 30.750 1269.520 ;
        RECT 33.650 1269.460 33.970 1269.520 ;
        RECT 30.430 1269.320 33.970 1269.460 ;
        RECT 30.430 1269.260 30.750 1269.320 ;
        RECT 33.650 1269.260 33.970 1269.320 ;
        RECT 30.430 1221.520 30.750 1221.580 ;
        RECT 33.650 1221.520 33.970 1221.580 ;
        RECT 30.430 1221.380 33.970 1221.520 ;
        RECT 30.430 1221.320 30.750 1221.380 ;
        RECT 33.650 1221.320 33.970 1221.380 ;
        RECT 30.430 1172.900 30.750 1172.960 ;
        RECT 33.650 1172.900 33.970 1172.960 ;
        RECT 30.430 1172.760 33.970 1172.900 ;
        RECT 30.430 1172.700 30.750 1172.760 ;
        RECT 33.650 1172.700 33.970 1172.760 ;
        RECT 30.430 1124.960 30.750 1125.020 ;
        RECT 33.650 1124.960 33.970 1125.020 ;
        RECT 30.430 1124.820 33.970 1124.960 ;
        RECT 30.430 1124.760 30.750 1124.820 ;
        RECT 33.650 1124.760 33.970 1124.820 ;
        RECT 30.430 1076.340 30.750 1076.400 ;
        RECT 33.650 1076.340 33.970 1076.400 ;
        RECT 30.430 1076.200 33.970 1076.340 ;
        RECT 30.430 1076.140 30.750 1076.200 ;
        RECT 33.650 1076.140 33.970 1076.200 ;
        RECT 30.430 1028.400 30.750 1028.460 ;
        RECT 33.650 1028.400 33.970 1028.460 ;
        RECT 30.430 1028.260 33.970 1028.400 ;
        RECT 30.430 1028.200 30.750 1028.260 ;
        RECT 33.650 1028.200 33.970 1028.260 ;
        RECT 30.430 979.780 30.750 979.840 ;
        RECT 33.650 979.780 33.970 979.840 ;
        RECT 30.430 979.640 33.970 979.780 ;
        RECT 30.430 979.580 30.750 979.640 ;
        RECT 33.650 979.580 33.970 979.640 ;
        RECT 30.430 931.840 30.750 931.900 ;
        RECT 33.650 931.840 33.970 931.900 ;
        RECT 30.430 931.700 33.970 931.840 ;
        RECT 30.430 931.640 30.750 931.700 ;
        RECT 33.650 931.640 33.970 931.700 ;
        RECT 30.430 883.220 30.750 883.280 ;
        RECT 33.650 883.220 33.970 883.280 ;
        RECT 30.430 883.080 33.970 883.220 ;
        RECT 30.430 883.020 30.750 883.080 ;
        RECT 33.650 883.020 33.970 883.080 ;
        RECT 30.430 835.280 30.750 835.340 ;
        RECT 33.650 835.280 33.970 835.340 ;
        RECT 30.430 835.140 33.970 835.280 ;
        RECT 30.430 835.080 30.750 835.140 ;
        RECT 33.650 835.080 33.970 835.140 ;
        RECT 30.430 786.660 30.750 786.720 ;
        RECT 33.650 786.660 33.970 786.720 ;
        RECT 30.430 786.520 33.970 786.660 ;
        RECT 30.430 786.460 30.750 786.520 ;
        RECT 33.650 786.460 33.970 786.520 ;
        RECT 30.430 738.380 30.750 738.440 ;
        RECT 33.650 738.380 33.970 738.440 ;
        RECT 30.430 738.240 33.970 738.380 ;
        RECT 30.430 738.180 30.750 738.240 ;
        RECT 33.650 738.180 33.970 738.240 ;
        RECT 30.430 689.760 30.750 689.820 ;
        RECT 33.650 689.760 33.970 689.820 ;
        RECT 30.430 689.620 33.970 689.760 ;
        RECT 30.430 689.560 30.750 689.620 ;
        RECT 33.650 689.560 33.970 689.620 ;
        RECT 30.430 641.820 30.750 641.880 ;
        RECT 33.650 641.820 33.970 641.880 ;
        RECT 30.430 641.680 33.970 641.820 ;
        RECT 30.430 641.620 30.750 641.680 ;
        RECT 33.650 641.620 33.970 641.680 ;
        RECT 30.430 593.200 30.750 593.260 ;
        RECT 33.650 593.200 33.970 593.260 ;
        RECT 30.430 593.060 33.970 593.200 ;
        RECT 30.430 593.000 30.750 593.060 ;
        RECT 33.650 593.000 33.970 593.060 ;
        RECT 30.430 545.260 30.750 545.320 ;
        RECT 33.650 545.260 33.970 545.320 ;
        RECT 30.430 545.120 33.970 545.260 ;
        RECT 30.430 545.060 30.750 545.120 ;
        RECT 33.650 545.060 33.970 545.120 ;
        RECT 30.430 496.640 30.750 496.700 ;
        RECT 33.650 496.640 33.970 496.700 ;
        RECT 30.430 496.500 33.970 496.640 ;
        RECT 30.430 496.440 30.750 496.500 ;
        RECT 33.650 496.440 33.970 496.500 ;
        RECT 30.430 448.700 30.750 448.760 ;
        RECT 33.650 448.700 33.970 448.760 ;
        RECT 30.430 448.560 33.970 448.700 ;
        RECT 30.430 448.500 30.750 448.560 ;
        RECT 33.650 448.500 33.970 448.560 ;
        RECT 30.430 400.080 30.750 400.140 ;
        RECT 33.650 400.080 33.970 400.140 ;
        RECT 30.430 399.940 33.970 400.080 ;
        RECT 30.430 399.880 30.750 399.940 ;
        RECT 33.650 399.880 33.970 399.940 ;
        RECT 30.430 352.140 30.750 352.200 ;
        RECT 33.650 352.140 33.970 352.200 ;
        RECT 30.430 352.000 33.970 352.140 ;
        RECT 30.430 351.940 30.750 352.000 ;
        RECT 33.650 351.940 33.970 352.000 ;
        RECT 30.430 303.520 30.750 303.580 ;
        RECT 33.650 303.520 33.970 303.580 ;
        RECT 30.430 303.380 33.970 303.520 ;
        RECT 30.430 303.320 30.750 303.380 ;
        RECT 33.650 303.320 33.970 303.380 ;
        RECT 30.430 255.580 30.750 255.640 ;
        RECT 33.650 255.580 33.970 255.640 ;
        RECT 30.430 255.440 33.970 255.580 ;
        RECT 30.430 255.380 30.750 255.440 ;
        RECT 33.650 255.380 33.970 255.440 ;
        RECT 30.430 206.960 30.750 207.020 ;
        RECT 33.650 206.960 33.970 207.020 ;
        RECT 30.430 206.820 33.970 206.960 ;
        RECT 30.430 206.760 30.750 206.820 ;
        RECT 33.650 206.760 33.970 206.820 ;
        RECT 30.430 159.020 30.750 159.080 ;
        RECT 33.650 159.020 33.970 159.080 ;
        RECT 30.430 158.880 33.970 159.020 ;
        RECT 30.430 158.820 30.750 158.880 ;
        RECT 33.650 158.820 33.970 158.880 ;
        RECT 30.430 110.400 30.750 110.460 ;
        RECT 33.650 110.400 33.970 110.460 ;
        RECT 30.430 110.260 33.970 110.400 ;
        RECT 30.430 110.200 30.750 110.260 ;
        RECT 33.650 110.200 33.970 110.260 ;
        RECT 30.430 62.460 30.750 62.520 ;
        RECT 33.650 62.460 33.970 62.520 ;
        RECT 30.430 62.320 33.970 62.460 ;
        RECT 30.430 62.260 30.750 62.320 ;
        RECT 33.650 62.260 33.970 62.320 ;
        RECT 33.650 19.620 33.970 19.680 ;
        RECT 478.470 19.620 478.790 19.680 ;
        RECT 33.650 19.480 478.790 19.620 ;
        RECT 33.650 19.420 33.970 19.480 ;
        RECT 478.470 19.420 478.790 19.480 ;
      LAYER via ;
        RECT 32.300 3007.680 32.560 3007.940 ;
        RECT 33.680 3007.680 33.940 3007.940 ;
        RECT 32.300 2959.400 32.560 2959.660 ;
        RECT 33.680 2959.400 33.940 2959.660 ;
        RECT 31.840 2911.120 32.100 2911.380 ;
        RECT 33.680 2911.120 33.940 2911.380 ;
        RECT 31.840 2862.160 32.100 2862.420 ;
        RECT 34.140 2862.160 34.400 2862.420 ;
        RECT 34.140 2815.920 34.400 2816.180 ;
        RECT 32.300 2815.240 32.560 2815.500 ;
        RECT 32.300 2766.960 32.560 2767.220 ;
        RECT 33.680 2766.960 33.940 2767.220 ;
        RECT 32.300 2670.400 32.560 2670.660 ;
        RECT 33.680 2670.400 33.940 2670.660 ;
        RECT 32.300 2573.840 32.560 2574.100 ;
        RECT 33.680 2573.840 33.940 2574.100 ;
        RECT 32.300 2477.280 32.560 2477.540 ;
        RECT 33.680 2477.280 33.940 2477.540 ;
        RECT 32.300 2380.380 32.560 2380.640 ;
        RECT 33.680 2380.380 33.940 2380.640 ;
        RECT 32.300 2283.820 32.560 2284.080 ;
        RECT 33.680 2283.820 33.940 2284.080 ;
        RECT 32.300 2187.260 32.560 2187.520 ;
        RECT 33.680 2187.260 33.940 2187.520 ;
        RECT 32.300 1994.140 32.560 1994.400 ;
        RECT 33.680 1994.140 33.940 1994.400 ;
        RECT 32.300 1945.520 32.560 1945.780 ;
        RECT 33.680 1945.520 33.940 1945.780 ;
        RECT 32.300 1897.580 32.560 1897.840 ;
        RECT 33.680 1897.580 33.940 1897.840 ;
        RECT 32.300 1848.960 32.560 1849.220 ;
        RECT 33.680 1848.960 33.940 1849.220 ;
        RECT 32.300 1801.020 32.560 1801.280 ;
        RECT 33.680 1801.020 33.940 1801.280 ;
        RECT 32.300 1752.400 32.560 1752.660 ;
        RECT 33.680 1752.400 33.940 1752.660 ;
        RECT 32.300 1704.460 32.560 1704.720 ;
        RECT 33.680 1704.460 33.940 1704.720 ;
        RECT 31.840 1655.840 32.100 1656.100 ;
        RECT 33.680 1655.840 33.940 1656.100 ;
        RECT 31.840 1607.900 32.100 1608.160 ;
        RECT 33.680 1607.900 33.940 1608.160 ;
        RECT 30.460 1558.940 30.720 1559.200 ;
        RECT 33.680 1558.940 33.940 1559.200 ;
        RECT 30.460 1511.000 30.720 1511.260 ;
        RECT 33.680 1511.000 33.940 1511.260 ;
        RECT 30.460 1462.380 30.720 1462.640 ;
        RECT 33.680 1462.380 33.940 1462.640 ;
        RECT 30.460 1414.440 30.720 1414.700 ;
        RECT 33.680 1414.440 33.940 1414.700 ;
        RECT 30.460 1365.820 30.720 1366.080 ;
        RECT 33.680 1365.820 33.940 1366.080 ;
        RECT 30.460 1317.880 30.720 1318.140 ;
        RECT 33.680 1317.880 33.940 1318.140 ;
        RECT 30.460 1269.260 30.720 1269.520 ;
        RECT 33.680 1269.260 33.940 1269.520 ;
        RECT 30.460 1221.320 30.720 1221.580 ;
        RECT 33.680 1221.320 33.940 1221.580 ;
        RECT 30.460 1172.700 30.720 1172.960 ;
        RECT 33.680 1172.700 33.940 1172.960 ;
        RECT 30.460 1124.760 30.720 1125.020 ;
        RECT 33.680 1124.760 33.940 1125.020 ;
        RECT 30.460 1076.140 30.720 1076.400 ;
        RECT 33.680 1076.140 33.940 1076.400 ;
        RECT 30.460 1028.200 30.720 1028.460 ;
        RECT 33.680 1028.200 33.940 1028.460 ;
        RECT 30.460 979.580 30.720 979.840 ;
        RECT 33.680 979.580 33.940 979.840 ;
        RECT 30.460 931.640 30.720 931.900 ;
        RECT 33.680 931.640 33.940 931.900 ;
        RECT 30.460 883.020 30.720 883.280 ;
        RECT 33.680 883.020 33.940 883.280 ;
        RECT 30.460 835.080 30.720 835.340 ;
        RECT 33.680 835.080 33.940 835.340 ;
        RECT 30.460 786.460 30.720 786.720 ;
        RECT 33.680 786.460 33.940 786.720 ;
        RECT 30.460 738.180 30.720 738.440 ;
        RECT 33.680 738.180 33.940 738.440 ;
        RECT 30.460 689.560 30.720 689.820 ;
        RECT 33.680 689.560 33.940 689.820 ;
        RECT 30.460 641.620 30.720 641.880 ;
        RECT 33.680 641.620 33.940 641.880 ;
        RECT 30.460 593.000 30.720 593.260 ;
        RECT 33.680 593.000 33.940 593.260 ;
        RECT 30.460 545.060 30.720 545.320 ;
        RECT 33.680 545.060 33.940 545.320 ;
        RECT 30.460 496.440 30.720 496.700 ;
        RECT 33.680 496.440 33.940 496.700 ;
        RECT 30.460 448.500 30.720 448.760 ;
        RECT 33.680 448.500 33.940 448.760 ;
        RECT 30.460 399.880 30.720 400.140 ;
        RECT 33.680 399.880 33.940 400.140 ;
        RECT 30.460 351.940 30.720 352.200 ;
        RECT 33.680 351.940 33.940 352.200 ;
        RECT 30.460 303.320 30.720 303.580 ;
        RECT 33.680 303.320 33.940 303.580 ;
        RECT 30.460 255.380 30.720 255.640 ;
        RECT 33.680 255.380 33.940 255.640 ;
        RECT 30.460 206.760 30.720 207.020 ;
        RECT 33.680 206.760 33.940 207.020 ;
        RECT 30.460 158.820 30.720 159.080 ;
        RECT 33.680 158.820 33.940 159.080 ;
        RECT 30.460 110.200 30.720 110.460 ;
        RECT 33.680 110.200 33.940 110.460 ;
        RECT 30.460 62.260 30.720 62.520 ;
        RECT 33.680 62.260 33.940 62.520 ;
        RECT 33.680 19.420 33.940 19.680 ;
        RECT 478.500 19.420 478.760 19.680 ;
      LAYER met2 ;
        RECT 33.670 3050.295 33.950 3050.665 ;
        RECT 33.740 3007.970 33.880 3050.295 ;
        RECT 32.300 3007.650 32.560 3007.970 ;
        RECT 33.680 3007.650 33.940 3007.970 ;
        RECT 32.360 2959.690 32.500 3007.650 ;
        RECT 32.300 2959.370 32.560 2959.690 ;
        RECT 33.680 2959.370 33.940 2959.690 ;
        RECT 33.740 2911.410 33.880 2959.370 ;
        RECT 31.840 2911.090 32.100 2911.410 ;
        RECT 33.680 2911.090 33.940 2911.410 ;
        RECT 31.900 2862.450 32.040 2911.090 ;
        RECT 31.840 2862.130 32.100 2862.450 ;
        RECT 34.140 2862.130 34.400 2862.450 ;
        RECT 34.200 2816.210 34.340 2862.130 ;
        RECT 34.140 2815.890 34.400 2816.210 ;
        RECT 32.300 2815.210 32.560 2815.530 ;
        RECT 32.360 2767.250 32.500 2815.210 ;
        RECT 32.300 2766.930 32.560 2767.250 ;
        RECT 33.680 2766.930 33.940 2767.250 ;
        RECT 33.740 2718.485 33.880 2766.930 ;
        RECT 32.290 2718.115 32.570 2718.485 ;
        RECT 33.670 2718.115 33.950 2718.485 ;
        RECT 32.360 2670.690 32.500 2718.115 ;
        RECT 32.300 2670.370 32.560 2670.690 ;
        RECT 33.680 2670.370 33.940 2670.690 ;
        RECT 33.740 2621.925 33.880 2670.370 ;
        RECT 32.290 2621.555 32.570 2621.925 ;
        RECT 33.670 2621.555 33.950 2621.925 ;
        RECT 32.360 2574.130 32.500 2621.555 ;
        RECT 32.300 2573.810 32.560 2574.130 ;
        RECT 33.680 2573.810 33.940 2574.130 ;
        RECT 33.740 2525.365 33.880 2573.810 ;
        RECT 32.290 2524.995 32.570 2525.365 ;
        RECT 33.670 2524.995 33.950 2525.365 ;
        RECT 32.360 2477.570 32.500 2524.995 ;
        RECT 32.300 2477.250 32.560 2477.570 ;
        RECT 33.680 2477.250 33.940 2477.570 ;
        RECT 33.740 2428.805 33.880 2477.250 ;
        RECT 32.290 2428.435 32.570 2428.805 ;
        RECT 33.670 2428.435 33.950 2428.805 ;
        RECT 32.360 2380.670 32.500 2428.435 ;
        RECT 32.300 2380.350 32.560 2380.670 ;
        RECT 33.680 2380.350 33.940 2380.670 ;
        RECT 33.740 2332.245 33.880 2380.350 ;
        RECT 32.290 2331.875 32.570 2332.245 ;
        RECT 33.670 2331.875 33.950 2332.245 ;
        RECT 32.360 2284.110 32.500 2331.875 ;
        RECT 32.300 2283.790 32.560 2284.110 ;
        RECT 33.680 2283.790 33.940 2284.110 ;
        RECT 33.740 2235.685 33.880 2283.790 ;
        RECT 32.290 2235.315 32.570 2235.685 ;
        RECT 33.670 2235.315 33.950 2235.685 ;
        RECT 32.360 2187.550 32.500 2235.315 ;
        RECT 32.300 2187.230 32.560 2187.550 ;
        RECT 33.680 2187.230 33.940 2187.550 ;
        RECT 33.740 2042.565 33.880 2187.230 ;
        RECT 32.290 2042.195 32.570 2042.565 ;
        RECT 33.670 2042.195 33.950 2042.565 ;
        RECT 32.360 1994.430 32.500 2042.195 ;
        RECT 32.300 1994.110 32.560 1994.430 ;
        RECT 33.680 1994.110 33.940 1994.430 ;
        RECT 33.740 1945.810 33.880 1994.110 ;
        RECT 32.300 1945.490 32.560 1945.810 ;
        RECT 33.680 1945.490 33.940 1945.810 ;
        RECT 32.360 1897.870 32.500 1945.490 ;
        RECT 32.300 1897.550 32.560 1897.870 ;
        RECT 33.680 1897.550 33.940 1897.870 ;
        RECT 33.740 1849.250 33.880 1897.550 ;
        RECT 32.300 1848.930 32.560 1849.250 ;
        RECT 33.680 1848.930 33.940 1849.250 ;
        RECT 32.360 1801.310 32.500 1848.930 ;
        RECT 32.300 1800.990 32.560 1801.310 ;
        RECT 33.680 1800.990 33.940 1801.310 ;
        RECT 33.740 1752.690 33.880 1800.990 ;
        RECT 32.300 1752.370 32.560 1752.690 ;
        RECT 33.680 1752.370 33.940 1752.690 ;
        RECT 32.360 1704.750 32.500 1752.370 ;
        RECT 32.300 1704.430 32.560 1704.750 ;
        RECT 33.680 1704.430 33.940 1704.750 ;
        RECT 33.740 1656.130 33.880 1704.430 ;
        RECT 31.840 1655.810 32.100 1656.130 ;
        RECT 33.680 1655.810 33.940 1656.130 ;
        RECT 31.900 1608.190 32.040 1655.810 ;
        RECT 31.840 1607.870 32.100 1608.190 ;
        RECT 33.680 1607.870 33.940 1608.190 ;
        RECT 33.740 1559.230 33.880 1607.870 ;
        RECT 30.460 1558.910 30.720 1559.230 ;
        RECT 33.680 1558.910 33.940 1559.230 ;
        RECT 30.520 1511.290 30.660 1558.910 ;
        RECT 30.460 1510.970 30.720 1511.290 ;
        RECT 33.680 1510.970 33.940 1511.290 ;
        RECT 33.740 1462.670 33.880 1510.970 ;
        RECT 30.460 1462.350 30.720 1462.670 ;
        RECT 33.680 1462.350 33.940 1462.670 ;
        RECT 30.520 1414.730 30.660 1462.350 ;
        RECT 30.460 1414.410 30.720 1414.730 ;
        RECT 33.680 1414.410 33.940 1414.730 ;
        RECT 33.740 1366.110 33.880 1414.410 ;
        RECT 30.460 1365.790 30.720 1366.110 ;
        RECT 33.680 1365.790 33.940 1366.110 ;
        RECT 30.520 1318.170 30.660 1365.790 ;
        RECT 30.460 1317.850 30.720 1318.170 ;
        RECT 33.680 1317.850 33.940 1318.170 ;
        RECT 33.740 1269.550 33.880 1317.850 ;
        RECT 30.460 1269.230 30.720 1269.550 ;
        RECT 33.680 1269.230 33.940 1269.550 ;
        RECT 30.520 1221.610 30.660 1269.230 ;
        RECT 30.460 1221.290 30.720 1221.610 ;
        RECT 33.680 1221.290 33.940 1221.610 ;
        RECT 33.740 1172.990 33.880 1221.290 ;
        RECT 30.460 1172.670 30.720 1172.990 ;
        RECT 33.680 1172.670 33.940 1172.990 ;
        RECT 30.520 1125.050 30.660 1172.670 ;
        RECT 30.460 1124.730 30.720 1125.050 ;
        RECT 33.680 1124.730 33.940 1125.050 ;
        RECT 33.740 1076.430 33.880 1124.730 ;
        RECT 30.460 1076.110 30.720 1076.430 ;
        RECT 33.680 1076.110 33.940 1076.430 ;
        RECT 30.520 1028.490 30.660 1076.110 ;
        RECT 30.460 1028.170 30.720 1028.490 ;
        RECT 33.680 1028.170 33.940 1028.490 ;
        RECT 33.740 979.870 33.880 1028.170 ;
        RECT 30.460 979.550 30.720 979.870 ;
        RECT 33.680 979.550 33.940 979.870 ;
        RECT 30.520 931.930 30.660 979.550 ;
        RECT 30.460 931.610 30.720 931.930 ;
        RECT 33.680 931.610 33.940 931.930 ;
        RECT 33.740 883.310 33.880 931.610 ;
        RECT 30.460 882.990 30.720 883.310 ;
        RECT 33.680 882.990 33.940 883.310 ;
        RECT 30.520 835.370 30.660 882.990 ;
        RECT 30.460 835.050 30.720 835.370 ;
        RECT 33.680 835.050 33.940 835.370 ;
        RECT 33.740 786.750 33.880 835.050 ;
        RECT 30.460 786.430 30.720 786.750 ;
        RECT 33.680 786.430 33.940 786.750 ;
        RECT 30.520 738.470 30.660 786.430 ;
        RECT 30.460 738.150 30.720 738.470 ;
        RECT 33.680 738.150 33.940 738.470 ;
        RECT 33.740 689.850 33.880 738.150 ;
        RECT 30.460 689.530 30.720 689.850 ;
        RECT 33.680 689.530 33.940 689.850 ;
        RECT 30.520 641.910 30.660 689.530 ;
        RECT 30.460 641.590 30.720 641.910 ;
        RECT 33.680 641.590 33.940 641.910 ;
        RECT 33.740 593.290 33.880 641.590 ;
        RECT 30.460 592.970 30.720 593.290 ;
        RECT 33.680 592.970 33.940 593.290 ;
        RECT 30.520 545.350 30.660 592.970 ;
        RECT 30.460 545.030 30.720 545.350 ;
        RECT 33.680 545.030 33.940 545.350 ;
        RECT 33.740 496.730 33.880 545.030 ;
        RECT 30.460 496.410 30.720 496.730 ;
        RECT 33.680 496.410 33.940 496.730 ;
        RECT 30.520 448.790 30.660 496.410 ;
        RECT 30.460 448.470 30.720 448.790 ;
        RECT 33.680 448.470 33.940 448.790 ;
        RECT 33.740 400.170 33.880 448.470 ;
        RECT 30.460 399.850 30.720 400.170 ;
        RECT 33.680 399.850 33.940 400.170 ;
        RECT 30.520 352.230 30.660 399.850 ;
        RECT 30.460 351.910 30.720 352.230 ;
        RECT 33.680 351.910 33.940 352.230 ;
        RECT 33.740 303.610 33.880 351.910 ;
        RECT 30.460 303.290 30.720 303.610 ;
        RECT 33.680 303.290 33.940 303.610 ;
        RECT 30.520 255.670 30.660 303.290 ;
        RECT 30.460 255.350 30.720 255.670 ;
        RECT 33.680 255.350 33.940 255.670 ;
        RECT 33.740 207.050 33.880 255.350 ;
        RECT 30.460 206.730 30.720 207.050 ;
        RECT 33.680 206.730 33.940 207.050 ;
        RECT 30.520 159.110 30.660 206.730 ;
        RECT 30.460 158.790 30.720 159.110 ;
        RECT 33.680 158.790 33.940 159.110 ;
        RECT 33.740 110.490 33.880 158.790 ;
        RECT 30.460 110.170 30.720 110.490 ;
        RECT 33.680 110.170 33.940 110.490 ;
        RECT 30.520 62.550 30.660 110.170 ;
        RECT 30.460 62.230 30.720 62.550 ;
        RECT 33.680 62.230 33.940 62.550 ;
        RECT 33.740 19.710 33.880 62.230 ;
        RECT 33.680 19.390 33.940 19.710 ;
        RECT 478.500 19.390 478.760 19.710 ;
        RECT 478.560 2.400 478.700 19.390 ;
        RECT 478.350 -4.800 478.910 2.400 ;
      LAYER via2 ;
        RECT 33.670 3050.340 33.950 3050.620 ;
        RECT 32.290 2718.160 32.570 2718.440 ;
        RECT 33.670 2718.160 33.950 2718.440 ;
        RECT 32.290 2621.600 32.570 2621.880 ;
        RECT 33.670 2621.600 33.950 2621.880 ;
        RECT 32.290 2525.040 32.570 2525.320 ;
        RECT 33.670 2525.040 33.950 2525.320 ;
        RECT 32.290 2428.480 32.570 2428.760 ;
        RECT 33.670 2428.480 33.950 2428.760 ;
        RECT 32.290 2331.920 32.570 2332.200 ;
        RECT 33.670 2331.920 33.950 2332.200 ;
        RECT 32.290 2235.360 32.570 2235.640 ;
        RECT 33.670 2235.360 33.950 2235.640 ;
        RECT 32.290 2042.240 32.570 2042.520 ;
        RECT 33.670 2042.240 33.950 2042.520 ;
      LAYER met3 ;
        RECT 33.645 3050.630 33.975 3050.645 ;
        RECT 35.000 3050.630 39.000 3050.760 ;
        RECT 33.645 3050.330 39.000 3050.630 ;
        RECT 33.645 3050.315 33.975 3050.330 ;
        RECT 35.000 3050.160 39.000 3050.330 ;
        RECT 32.265 2718.450 32.595 2718.465 ;
        RECT 33.645 2718.450 33.975 2718.465 ;
        RECT 32.265 2718.150 33.975 2718.450 ;
        RECT 32.265 2718.135 32.595 2718.150 ;
        RECT 33.645 2718.135 33.975 2718.150 ;
        RECT 32.265 2621.890 32.595 2621.905 ;
        RECT 33.645 2621.890 33.975 2621.905 ;
        RECT 32.265 2621.590 33.975 2621.890 ;
        RECT 32.265 2621.575 32.595 2621.590 ;
        RECT 33.645 2621.575 33.975 2621.590 ;
        RECT 32.265 2525.330 32.595 2525.345 ;
        RECT 33.645 2525.330 33.975 2525.345 ;
        RECT 32.265 2525.030 33.975 2525.330 ;
        RECT 32.265 2525.015 32.595 2525.030 ;
        RECT 33.645 2525.015 33.975 2525.030 ;
        RECT 32.265 2428.770 32.595 2428.785 ;
        RECT 33.645 2428.770 33.975 2428.785 ;
        RECT 32.265 2428.470 33.975 2428.770 ;
        RECT 32.265 2428.455 32.595 2428.470 ;
        RECT 33.645 2428.455 33.975 2428.470 ;
        RECT 32.265 2332.210 32.595 2332.225 ;
        RECT 33.645 2332.210 33.975 2332.225 ;
        RECT 32.265 2331.910 33.975 2332.210 ;
        RECT 32.265 2331.895 32.595 2331.910 ;
        RECT 33.645 2331.895 33.975 2331.910 ;
        RECT 32.265 2235.650 32.595 2235.665 ;
        RECT 33.645 2235.650 33.975 2235.665 ;
        RECT 32.265 2235.350 33.975 2235.650 ;
        RECT 32.265 2235.335 32.595 2235.350 ;
        RECT 33.645 2235.335 33.975 2235.350 ;
        RECT 32.265 2042.530 32.595 2042.545 ;
        RECT 33.645 2042.530 33.975 2042.545 ;
        RECT 32.265 2042.230 33.975 2042.530 ;
        RECT 32.265 2042.215 32.595 2042.230 ;
        RECT 33.645 2042.215 33.975 2042.230 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 33.265 3091.365 33.435 3105.475 ;
        RECT 32.805 3043.085 32.975 3090.855 ;
        RECT 33.725 2861.865 33.895 2864.415 ;
      LAYER mcon ;
        RECT 33.265 3105.305 33.435 3105.475 ;
        RECT 32.805 3090.685 32.975 3090.855 ;
        RECT 33.725 2864.245 33.895 2864.415 ;
      LAYER met1 ;
        RECT 33.650 3139.800 33.970 3139.860 ;
        RECT 34.570 3139.800 34.890 3139.860 ;
        RECT 33.650 3139.660 34.890 3139.800 ;
        RECT 33.650 3139.600 33.970 3139.660 ;
        RECT 34.570 3139.600 34.890 3139.660 ;
        RECT 33.205 3105.460 33.495 3105.505 ;
        RECT 33.650 3105.460 33.970 3105.520 ;
        RECT 33.205 3105.320 33.970 3105.460 ;
        RECT 33.205 3105.275 33.495 3105.320 ;
        RECT 33.650 3105.260 33.970 3105.320 ;
        RECT 33.190 3091.520 33.510 3091.580 ;
        RECT 32.995 3091.380 33.510 3091.520 ;
        RECT 33.190 3091.320 33.510 3091.380 ;
        RECT 32.745 3090.840 33.035 3090.885 ;
        RECT 33.190 3090.840 33.510 3090.900 ;
        RECT 32.745 3090.700 33.510 3090.840 ;
        RECT 32.745 3090.655 33.035 3090.700 ;
        RECT 33.190 3090.640 33.510 3090.700 ;
        RECT 32.730 3043.240 33.050 3043.300 ;
        RECT 32.535 3043.100 33.050 3043.240 ;
        RECT 32.730 3043.040 33.050 3043.100 ;
        RECT 32.730 3008.900 33.050 3008.960 ;
        RECT 34.570 3008.900 34.890 3008.960 ;
        RECT 32.730 3008.760 34.890 3008.900 ;
        RECT 32.730 3008.700 33.050 3008.760 ;
        RECT 34.570 3008.700 34.890 3008.760 ;
        RECT 32.730 3008.220 33.050 3008.280 ;
        RECT 34.570 3008.220 34.890 3008.280 ;
        RECT 32.730 3008.080 34.890 3008.220 ;
        RECT 32.730 3008.020 33.050 3008.080 ;
        RECT 34.570 3008.020 34.890 3008.080 ;
        RECT 32.730 2960.420 33.050 2960.680 ;
        RECT 32.820 2960.000 32.960 2960.420 ;
        RECT 32.730 2959.740 33.050 2960.000 ;
        RECT 32.730 2912.000 33.050 2912.060 ;
        RECT 34.570 2912.000 34.890 2912.060 ;
        RECT 32.730 2911.860 34.890 2912.000 ;
        RECT 32.730 2911.800 33.050 2911.860 ;
        RECT 34.570 2911.800 34.890 2911.860 ;
        RECT 33.650 2864.400 33.970 2864.460 ;
        RECT 33.455 2864.260 33.970 2864.400 ;
        RECT 33.650 2864.200 33.970 2864.260 ;
        RECT 33.650 2862.020 33.970 2862.080 ;
        RECT 33.455 2861.880 33.970 2862.020 ;
        RECT 33.650 2861.820 33.970 2861.880 ;
        RECT 31.810 2815.100 32.130 2815.160 ;
        RECT 34.570 2815.100 34.890 2815.160 ;
        RECT 31.810 2814.960 34.890 2815.100 ;
        RECT 31.810 2814.900 32.130 2814.960 ;
        RECT 34.570 2814.900 34.890 2814.960 ;
        RECT 31.810 2767.500 32.130 2767.560 ;
        RECT 31.810 2767.360 34.340 2767.500 ;
        RECT 31.810 2767.300 32.130 2767.360 ;
        RECT 34.200 2767.220 34.340 2767.360 ;
        RECT 34.110 2766.960 34.430 2767.220 ;
        RECT 32.270 2766.480 32.590 2766.540 ;
        RECT 34.110 2766.480 34.430 2766.540 ;
        RECT 32.270 2766.340 34.430 2766.480 ;
        RECT 32.270 2766.280 32.590 2766.340 ;
        RECT 34.110 2766.280 34.430 2766.340 ;
        RECT 32.270 2719.220 32.590 2719.280 ;
        RECT 34.570 2719.220 34.890 2719.280 ;
        RECT 32.270 2719.080 34.890 2719.220 ;
        RECT 32.270 2719.020 32.590 2719.080 ;
        RECT 34.570 2719.020 34.890 2719.080 ;
        RECT 31.810 2718.540 32.130 2718.600 ;
        RECT 34.570 2718.540 34.890 2718.600 ;
        RECT 31.810 2718.400 34.890 2718.540 ;
        RECT 31.810 2718.340 32.130 2718.400 ;
        RECT 34.570 2718.340 34.890 2718.400 ;
        RECT 31.810 2670.940 32.130 2671.000 ;
        RECT 31.810 2670.800 34.340 2670.940 ;
        RECT 31.810 2670.740 32.130 2670.800 ;
        RECT 34.200 2670.660 34.340 2670.800 ;
        RECT 34.110 2670.400 34.430 2670.660 ;
        RECT 32.270 2669.920 32.590 2669.980 ;
        RECT 34.110 2669.920 34.430 2669.980 ;
        RECT 32.270 2669.780 34.430 2669.920 ;
        RECT 32.270 2669.720 32.590 2669.780 ;
        RECT 34.110 2669.720 34.430 2669.780 ;
        RECT 32.270 2622.320 32.590 2622.380 ;
        RECT 34.570 2622.320 34.890 2622.380 ;
        RECT 32.270 2622.180 34.890 2622.320 ;
        RECT 32.270 2622.120 32.590 2622.180 ;
        RECT 34.570 2622.120 34.890 2622.180 ;
        RECT 33.650 2574.720 33.970 2574.780 ;
        RECT 33.650 2574.580 34.340 2574.720 ;
        RECT 33.650 2574.520 33.970 2574.580 ;
        RECT 34.200 2574.100 34.340 2574.580 ;
        RECT 34.110 2573.840 34.430 2574.100 ;
        RECT 32.270 2573.360 32.590 2573.420 ;
        RECT 34.110 2573.360 34.430 2573.420 ;
        RECT 32.270 2573.220 34.430 2573.360 ;
        RECT 32.270 2573.160 32.590 2573.220 ;
        RECT 34.110 2573.160 34.430 2573.220 ;
        RECT 32.270 2525.760 32.590 2525.820 ;
        RECT 34.570 2525.760 34.890 2525.820 ;
        RECT 32.270 2525.620 34.890 2525.760 ;
        RECT 32.270 2525.560 32.590 2525.620 ;
        RECT 34.570 2525.560 34.890 2525.620 ;
        RECT 33.650 2478.160 33.970 2478.220 ;
        RECT 33.650 2478.020 34.340 2478.160 ;
        RECT 33.650 2477.960 33.970 2478.020 ;
        RECT 34.200 2477.540 34.340 2478.020 ;
        RECT 34.110 2477.280 34.430 2477.540 ;
        RECT 32.270 2476.800 32.590 2476.860 ;
        RECT 34.110 2476.800 34.430 2476.860 ;
        RECT 32.270 2476.660 34.430 2476.800 ;
        RECT 32.270 2476.600 32.590 2476.660 ;
        RECT 34.110 2476.600 34.430 2476.660 ;
        RECT 32.270 2429.200 32.590 2429.260 ;
        RECT 34.570 2429.200 34.890 2429.260 ;
        RECT 32.270 2429.060 34.890 2429.200 ;
        RECT 32.270 2429.000 32.590 2429.060 ;
        RECT 34.570 2429.000 34.890 2429.060 ;
        RECT 33.650 2381.260 33.970 2381.320 ;
        RECT 33.650 2381.120 34.340 2381.260 ;
        RECT 33.650 2381.060 33.970 2381.120 ;
        RECT 34.200 2380.640 34.340 2381.120 ;
        RECT 34.110 2380.380 34.430 2380.640 ;
        RECT 33.650 2284.700 33.970 2284.760 ;
        RECT 33.650 2284.560 34.340 2284.700 ;
        RECT 33.650 2284.500 33.970 2284.560 ;
        RECT 34.200 2284.080 34.340 2284.560 ;
        RECT 34.110 2283.820 34.430 2284.080 ;
        RECT 33.650 2188.140 33.970 2188.200 ;
        RECT 33.650 2188.000 34.340 2188.140 ;
        RECT 33.650 2187.940 33.970 2188.000 ;
        RECT 34.200 2187.520 34.340 2188.000 ;
        RECT 34.110 2187.260 34.430 2187.520 ;
        RECT 34.110 1945.520 34.430 1945.780 ;
        RECT 31.810 1945.380 32.130 1945.440 ;
        RECT 34.200 1945.380 34.340 1945.520 ;
        RECT 31.810 1945.240 34.340 1945.380 ;
        RECT 31.810 1945.180 32.130 1945.240 ;
        RECT 31.810 1898.120 32.130 1898.180 ;
        RECT 31.810 1897.980 34.340 1898.120 ;
        RECT 31.810 1897.920 32.130 1897.980 ;
        RECT 34.200 1897.840 34.340 1897.980 ;
        RECT 34.110 1897.580 34.430 1897.840 ;
        RECT 34.110 1848.960 34.430 1849.220 ;
        RECT 31.810 1848.820 32.130 1848.880 ;
        RECT 34.200 1848.820 34.340 1848.960 ;
        RECT 31.810 1848.680 34.340 1848.820 ;
        RECT 31.810 1848.620 32.130 1848.680 ;
        RECT 31.810 1801.560 32.130 1801.620 ;
        RECT 31.810 1801.420 34.340 1801.560 ;
        RECT 31.810 1801.360 32.130 1801.420 ;
        RECT 34.200 1801.280 34.340 1801.420 ;
        RECT 34.110 1801.020 34.430 1801.280 ;
        RECT 34.110 1752.400 34.430 1752.660 ;
        RECT 31.810 1752.260 32.130 1752.320 ;
        RECT 34.200 1752.260 34.340 1752.400 ;
        RECT 31.810 1752.120 34.340 1752.260 ;
        RECT 31.810 1752.060 32.130 1752.120 ;
        RECT 31.810 1705.000 32.130 1705.060 ;
        RECT 31.810 1704.860 34.340 1705.000 ;
        RECT 31.810 1704.800 32.130 1704.860 ;
        RECT 34.200 1704.720 34.340 1704.860 ;
        RECT 34.110 1704.460 34.430 1704.720 ;
        RECT 34.110 1655.840 34.430 1656.100 ;
        RECT 30.430 1655.700 30.750 1655.760 ;
        RECT 34.200 1655.700 34.340 1655.840 ;
        RECT 30.430 1655.560 34.340 1655.700 ;
        RECT 30.430 1655.500 30.750 1655.560 ;
        RECT 30.430 1608.440 30.750 1608.500 ;
        RECT 30.430 1608.300 34.340 1608.440 ;
        RECT 30.430 1608.240 30.750 1608.300 ;
        RECT 34.200 1608.160 34.340 1608.300 ;
        RECT 34.110 1607.900 34.430 1608.160 ;
        RECT 34.110 1558.940 34.430 1559.200 ;
        RECT 31.810 1558.800 32.130 1558.860 ;
        RECT 34.200 1558.800 34.340 1558.940 ;
        RECT 31.810 1558.660 34.340 1558.800 ;
        RECT 31.810 1558.600 32.130 1558.660 ;
        RECT 31.810 1513.920 32.130 1513.980 ;
        RECT 31.810 1513.780 34.340 1513.920 ;
        RECT 31.810 1513.720 32.130 1513.780 ;
        RECT 34.200 1511.260 34.340 1513.780 ;
        RECT 34.110 1511.000 34.430 1511.260 ;
        RECT 34.110 1462.380 34.430 1462.640 ;
        RECT 29.970 1462.240 30.290 1462.300 ;
        RECT 34.200 1462.240 34.340 1462.380 ;
        RECT 29.970 1462.100 34.340 1462.240 ;
        RECT 29.970 1462.040 30.290 1462.100 ;
        RECT 29.970 1414.980 30.290 1415.040 ;
        RECT 29.970 1414.840 34.340 1414.980 ;
        RECT 29.970 1414.780 30.290 1414.840 ;
        RECT 34.200 1414.700 34.340 1414.840 ;
        RECT 34.110 1414.440 34.430 1414.700 ;
        RECT 34.110 1365.820 34.430 1366.080 ;
        RECT 29.970 1365.680 30.290 1365.740 ;
        RECT 34.200 1365.680 34.340 1365.820 ;
        RECT 29.970 1365.540 34.340 1365.680 ;
        RECT 29.970 1365.480 30.290 1365.540 ;
        RECT 29.970 1318.420 30.290 1318.480 ;
        RECT 29.970 1318.280 34.340 1318.420 ;
        RECT 29.970 1318.220 30.290 1318.280 ;
        RECT 34.200 1318.140 34.340 1318.280 ;
        RECT 34.110 1317.880 34.430 1318.140 ;
        RECT 34.110 1269.260 34.430 1269.520 ;
        RECT 29.970 1269.120 30.290 1269.180 ;
        RECT 34.200 1269.120 34.340 1269.260 ;
        RECT 29.970 1268.980 34.340 1269.120 ;
        RECT 29.970 1268.920 30.290 1268.980 ;
        RECT 29.970 1221.860 30.290 1221.920 ;
        RECT 29.970 1221.720 34.340 1221.860 ;
        RECT 29.970 1221.660 30.290 1221.720 ;
        RECT 34.200 1221.580 34.340 1221.720 ;
        RECT 34.110 1221.320 34.430 1221.580 ;
        RECT 34.110 1172.700 34.430 1172.960 ;
        RECT 29.970 1172.560 30.290 1172.620 ;
        RECT 34.200 1172.560 34.340 1172.700 ;
        RECT 29.970 1172.420 34.340 1172.560 ;
        RECT 29.970 1172.360 30.290 1172.420 ;
        RECT 29.970 1125.300 30.290 1125.360 ;
        RECT 29.970 1125.160 34.340 1125.300 ;
        RECT 29.970 1125.100 30.290 1125.160 ;
        RECT 34.200 1125.020 34.340 1125.160 ;
        RECT 34.110 1124.760 34.430 1125.020 ;
        RECT 34.110 1076.140 34.430 1076.400 ;
        RECT 29.970 1076.000 30.290 1076.060 ;
        RECT 34.200 1076.000 34.340 1076.140 ;
        RECT 29.970 1075.860 34.340 1076.000 ;
        RECT 29.970 1075.800 30.290 1075.860 ;
        RECT 29.970 1028.740 30.290 1028.800 ;
        RECT 29.970 1028.600 34.340 1028.740 ;
        RECT 29.970 1028.540 30.290 1028.600 ;
        RECT 34.200 1028.460 34.340 1028.600 ;
        RECT 34.110 1028.200 34.430 1028.460 ;
        RECT 34.110 979.580 34.430 979.840 ;
        RECT 29.970 979.440 30.290 979.500 ;
        RECT 34.200 979.440 34.340 979.580 ;
        RECT 29.970 979.300 34.340 979.440 ;
        RECT 29.970 979.240 30.290 979.300 ;
        RECT 29.970 932.180 30.290 932.240 ;
        RECT 29.970 932.040 34.340 932.180 ;
        RECT 29.970 931.980 30.290 932.040 ;
        RECT 34.200 931.900 34.340 932.040 ;
        RECT 34.110 931.640 34.430 931.900 ;
        RECT 34.110 883.020 34.430 883.280 ;
        RECT 29.970 882.880 30.290 882.940 ;
        RECT 34.200 882.880 34.340 883.020 ;
        RECT 29.970 882.740 34.340 882.880 ;
        RECT 29.970 882.680 30.290 882.740 ;
        RECT 29.970 835.620 30.290 835.680 ;
        RECT 29.970 835.480 34.340 835.620 ;
        RECT 29.970 835.420 30.290 835.480 ;
        RECT 34.200 835.340 34.340 835.480 ;
        RECT 34.110 835.080 34.430 835.340 ;
        RECT 34.110 786.460 34.430 786.720 ;
        RECT 29.970 786.320 30.290 786.380 ;
        RECT 34.200 786.320 34.340 786.460 ;
        RECT 29.970 786.180 34.340 786.320 ;
        RECT 29.970 786.120 30.290 786.180 ;
        RECT 29.970 738.720 30.290 738.780 ;
        RECT 29.970 738.580 34.340 738.720 ;
        RECT 29.970 738.520 30.290 738.580 ;
        RECT 34.200 738.440 34.340 738.580 ;
        RECT 34.110 738.180 34.430 738.440 ;
        RECT 34.110 689.560 34.430 689.820 ;
        RECT 29.970 689.420 30.290 689.480 ;
        RECT 34.200 689.420 34.340 689.560 ;
        RECT 29.970 689.280 34.340 689.420 ;
        RECT 29.970 689.220 30.290 689.280 ;
        RECT 29.970 642.160 30.290 642.220 ;
        RECT 29.970 642.020 34.340 642.160 ;
        RECT 29.970 641.960 30.290 642.020 ;
        RECT 34.200 641.880 34.340 642.020 ;
        RECT 34.110 641.620 34.430 641.880 ;
        RECT 34.110 593.000 34.430 593.260 ;
        RECT 29.970 592.860 30.290 592.920 ;
        RECT 34.200 592.860 34.340 593.000 ;
        RECT 29.970 592.720 34.340 592.860 ;
        RECT 29.970 592.660 30.290 592.720 ;
        RECT 29.970 545.600 30.290 545.660 ;
        RECT 29.970 545.460 34.340 545.600 ;
        RECT 29.970 545.400 30.290 545.460 ;
        RECT 34.200 545.320 34.340 545.460 ;
        RECT 34.110 545.060 34.430 545.320 ;
        RECT 34.110 496.440 34.430 496.700 ;
        RECT 29.970 496.300 30.290 496.360 ;
        RECT 34.200 496.300 34.340 496.440 ;
        RECT 29.970 496.160 34.340 496.300 ;
        RECT 29.970 496.100 30.290 496.160 ;
        RECT 29.970 449.040 30.290 449.100 ;
        RECT 29.970 448.900 34.340 449.040 ;
        RECT 29.970 448.840 30.290 448.900 ;
        RECT 34.200 448.760 34.340 448.900 ;
        RECT 34.110 448.500 34.430 448.760 ;
        RECT 34.110 399.880 34.430 400.140 ;
        RECT 29.970 399.740 30.290 399.800 ;
        RECT 34.200 399.740 34.340 399.880 ;
        RECT 29.970 399.600 34.340 399.740 ;
        RECT 29.970 399.540 30.290 399.600 ;
        RECT 29.970 352.480 30.290 352.540 ;
        RECT 29.970 352.340 34.340 352.480 ;
        RECT 29.970 352.280 30.290 352.340 ;
        RECT 34.200 352.200 34.340 352.340 ;
        RECT 34.110 351.940 34.430 352.200 ;
        RECT 34.110 303.320 34.430 303.580 ;
        RECT 29.970 303.180 30.290 303.240 ;
        RECT 34.200 303.180 34.340 303.320 ;
        RECT 29.970 303.040 34.340 303.180 ;
        RECT 29.970 302.980 30.290 303.040 ;
        RECT 29.970 255.920 30.290 255.980 ;
        RECT 29.970 255.780 34.340 255.920 ;
        RECT 29.970 255.720 30.290 255.780 ;
        RECT 34.200 255.640 34.340 255.780 ;
        RECT 34.110 255.380 34.430 255.640 ;
        RECT 34.110 206.760 34.430 207.020 ;
        RECT 29.970 206.620 30.290 206.680 ;
        RECT 34.200 206.620 34.340 206.760 ;
        RECT 29.970 206.480 34.340 206.620 ;
        RECT 29.970 206.420 30.290 206.480 ;
        RECT 29.970 159.360 30.290 159.420 ;
        RECT 29.970 159.220 34.340 159.360 ;
        RECT 29.970 159.160 30.290 159.220 ;
        RECT 34.200 159.080 34.340 159.220 ;
        RECT 34.110 158.820 34.430 159.080 ;
        RECT 34.110 110.200 34.430 110.460 ;
        RECT 29.970 110.060 30.290 110.120 ;
        RECT 34.200 110.060 34.340 110.200 ;
        RECT 29.970 109.920 34.340 110.060 ;
        RECT 29.970 109.860 30.290 109.920 ;
        RECT 29.970 62.800 30.290 62.860 ;
        RECT 29.970 62.660 34.340 62.800 ;
        RECT 29.970 62.600 30.290 62.660 ;
        RECT 34.200 62.520 34.340 62.660 ;
        RECT 34.110 62.260 34.430 62.520 ;
      LAYER via ;
        RECT 33.680 3139.600 33.940 3139.860 ;
        RECT 34.600 3139.600 34.860 3139.860 ;
        RECT 33.680 3105.260 33.940 3105.520 ;
        RECT 33.220 3091.320 33.480 3091.580 ;
        RECT 33.220 3090.640 33.480 3090.900 ;
        RECT 32.760 3043.040 33.020 3043.300 ;
        RECT 32.760 3008.700 33.020 3008.960 ;
        RECT 34.600 3008.700 34.860 3008.960 ;
        RECT 32.760 3008.020 33.020 3008.280 ;
        RECT 34.600 3008.020 34.860 3008.280 ;
        RECT 32.760 2960.420 33.020 2960.680 ;
        RECT 32.760 2959.740 33.020 2960.000 ;
        RECT 32.760 2911.800 33.020 2912.060 ;
        RECT 34.600 2911.800 34.860 2912.060 ;
        RECT 33.680 2864.200 33.940 2864.460 ;
        RECT 33.680 2861.820 33.940 2862.080 ;
        RECT 31.840 2814.900 32.100 2815.160 ;
        RECT 34.600 2814.900 34.860 2815.160 ;
        RECT 31.840 2767.300 32.100 2767.560 ;
        RECT 34.140 2766.960 34.400 2767.220 ;
        RECT 32.300 2766.280 32.560 2766.540 ;
        RECT 34.140 2766.280 34.400 2766.540 ;
        RECT 32.300 2719.020 32.560 2719.280 ;
        RECT 34.600 2719.020 34.860 2719.280 ;
        RECT 31.840 2718.340 32.100 2718.600 ;
        RECT 34.600 2718.340 34.860 2718.600 ;
        RECT 31.840 2670.740 32.100 2671.000 ;
        RECT 34.140 2670.400 34.400 2670.660 ;
        RECT 32.300 2669.720 32.560 2669.980 ;
        RECT 34.140 2669.720 34.400 2669.980 ;
        RECT 32.300 2622.120 32.560 2622.380 ;
        RECT 34.600 2622.120 34.860 2622.380 ;
        RECT 33.680 2574.520 33.940 2574.780 ;
        RECT 34.140 2573.840 34.400 2574.100 ;
        RECT 32.300 2573.160 32.560 2573.420 ;
        RECT 34.140 2573.160 34.400 2573.420 ;
        RECT 32.300 2525.560 32.560 2525.820 ;
        RECT 34.600 2525.560 34.860 2525.820 ;
        RECT 33.680 2477.960 33.940 2478.220 ;
        RECT 34.140 2477.280 34.400 2477.540 ;
        RECT 32.300 2476.600 32.560 2476.860 ;
        RECT 34.140 2476.600 34.400 2476.860 ;
        RECT 32.300 2429.000 32.560 2429.260 ;
        RECT 34.600 2429.000 34.860 2429.260 ;
        RECT 33.680 2381.060 33.940 2381.320 ;
        RECT 34.140 2380.380 34.400 2380.640 ;
        RECT 33.680 2284.500 33.940 2284.760 ;
        RECT 34.140 2283.820 34.400 2284.080 ;
        RECT 33.680 2187.940 33.940 2188.200 ;
        RECT 34.140 2187.260 34.400 2187.520 ;
        RECT 34.140 1945.520 34.400 1945.780 ;
        RECT 31.840 1945.180 32.100 1945.440 ;
        RECT 31.840 1897.920 32.100 1898.180 ;
        RECT 34.140 1897.580 34.400 1897.840 ;
        RECT 34.140 1848.960 34.400 1849.220 ;
        RECT 31.840 1848.620 32.100 1848.880 ;
        RECT 31.840 1801.360 32.100 1801.620 ;
        RECT 34.140 1801.020 34.400 1801.280 ;
        RECT 34.140 1752.400 34.400 1752.660 ;
        RECT 31.840 1752.060 32.100 1752.320 ;
        RECT 31.840 1704.800 32.100 1705.060 ;
        RECT 34.140 1704.460 34.400 1704.720 ;
        RECT 34.140 1655.840 34.400 1656.100 ;
        RECT 30.460 1655.500 30.720 1655.760 ;
        RECT 30.460 1608.240 30.720 1608.500 ;
        RECT 34.140 1607.900 34.400 1608.160 ;
        RECT 34.140 1558.940 34.400 1559.200 ;
        RECT 31.840 1558.600 32.100 1558.860 ;
        RECT 31.840 1513.720 32.100 1513.980 ;
        RECT 34.140 1511.000 34.400 1511.260 ;
        RECT 34.140 1462.380 34.400 1462.640 ;
        RECT 30.000 1462.040 30.260 1462.300 ;
        RECT 30.000 1414.780 30.260 1415.040 ;
        RECT 34.140 1414.440 34.400 1414.700 ;
        RECT 34.140 1365.820 34.400 1366.080 ;
        RECT 30.000 1365.480 30.260 1365.740 ;
        RECT 30.000 1318.220 30.260 1318.480 ;
        RECT 34.140 1317.880 34.400 1318.140 ;
        RECT 34.140 1269.260 34.400 1269.520 ;
        RECT 30.000 1268.920 30.260 1269.180 ;
        RECT 30.000 1221.660 30.260 1221.920 ;
        RECT 34.140 1221.320 34.400 1221.580 ;
        RECT 34.140 1172.700 34.400 1172.960 ;
        RECT 30.000 1172.360 30.260 1172.620 ;
        RECT 30.000 1125.100 30.260 1125.360 ;
        RECT 34.140 1124.760 34.400 1125.020 ;
        RECT 34.140 1076.140 34.400 1076.400 ;
        RECT 30.000 1075.800 30.260 1076.060 ;
        RECT 30.000 1028.540 30.260 1028.800 ;
        RECT 34.140 1028.200 34.400 1028.460 ;
        RECT 34.140 979.580 34.400 979.840 ;
        RECT 30.000 979.240 30.260 979.500 ;
        RECT 30.000 931.980 30.260 932.240 ;
        RECT 34.140 931.640 34.400 931.900 ;
        RECT 34.140 883.020 34.400 883.280 ;
        RECT 30.000 882.680 30.260 882.940 ;
        RECT 30.000 835.420 30.260 835.680 ;
        RECT 34.140 835.080 34.400 835.340 ;
        RECT 34.140 786.460 34.400 786.720 ;
        RECT 30.000 786.120 30.260 786.380 ;
        RECT 30.000 738.520 30.260 738.780 ;
        RECT 34.140 738.180 34.400 738.440 ;
        RECT 34.140 689.560 34.400 689.820 ;
        RECT 30.000 689.220 30.260 689.480 ;
        RECT 30.000 641.960 30.260 642.220 ;
        RECT 34.140 641.620 34.400 641.880 ;
        RECT 34.140 593.000 34.400 593.260 ;
        RECT 30.000 592.660 30.260 592.920 ;
        RECT 30.000 545.400 30.260 545.660 ;
        RECT 34.140 545.060 34.400 545.320 ;
        RECT 34.140 496.440 34.400 496.700 ;
        RECT 30.000 496.100 30.260 496.360 ;
        RECT 30.000 448.840 30.260 449.100 ;
        RECT 34.140 448.500 34.400 448.760 ;
        RECT 34.140 399.880 34.400 400.140 ;
        RECT 30.000 399.540 30.260 399.800 ;
        RECT 30.000 352.280 30.260 352.540 ;
        RECT 34.140 351.940 34.400 352.200 ;
        RECT 34.140 303.320 34.400 303.580 ;
        RECT 30.000 302.980 30.260 303.240 ;
        RECT 30.000 255.720 30.260 255.980 ;
        RECT 34.140 255.380 34.400 255.640 ;
        RECT 34.140 206.760 34.400 207.020 ;
        RECT 30.000 206.420 30.260 206.680 ;
        RECT 30.000 159.160 30.260 159.420 ;
        RECT 34.140 158.820 34.400 159.080 ;
        RECT 34.140 110.200 34.400 110.460 ;
        RECT 30.000 109.860 30.260 110.120 ;
        RECT 30.000 62.600 30.260 62.860 ;
        RECT 34.140 62.260 34.400 62.520 ;
      LAYER met2 ;
        RECT 34.590 3157.395 34.870 3157.765 ;
        RECT 34.660 3139.890 34.800 3157.395 ;
        RECT 33.680 3139.570 33.940 3139.890 ;
        RECT 34.600 3139.570 34.860 3139.890 ;
        RECT 33.740 3105.550 33.880 3139.570 ;
        RECT 33.680 3105.230 33.940 3105.550 ;
        RECT 33.220 3091.290 33.480 3091.610 ;
        RECT 33.280 3090.930 33.420 3091.290 ;
        RECT 33.220 3090.610 33.480 3090.930 ;
        RECT 32.760 3043.010 33.020 3043.330 ;
        RECT 32.820 3008.990 32.960 3043.010 ;
        RECT 32.760 3008.670 33.020 3008.990 ;
        RECT 34.600 3008.670 34.860 3008.990 ;
        RECT 34.660 3008.310 34.800 3008.670 ;
        RECT 32.760 3007.990 33.020 3008.310 ;
        RECT 34.600 3007.990 34.860 3008.310 ;
        RECT 32.820 2960.710 32.960 3007.990 ;
        RECT 32.760 2960.390 33.020 2960.710 ;
        RECT 32.760 2959.710 33.020 2960.030 ;
        RECT 32.820 2912.090 32.960 2959.710 ;
        RECT 32.760 2911.770 33.020 2912.090 ;
        RECT 34.600 2911.770 34.860 2912.090 ;
        RECT 34.660 2910.810 34.800 2911.770 ;
        RECT 33.740 2910.670 34.800 2910.810 ;
        RECT 33.740 2864.490 33.880 2910.670 ;
        RECT 33.680 2864.170 33.940 2864.490 ;
        RECT 33.680 2861.790 33.940 2862.110 ;
        RECT 33.740 2815.610 33.880 2861.790 ;
        RECT 33.740 2815.470 34.800 2815.610 ;
        RECT 34.660 2815.190 34.800 2815.470 ;
        RECT 31.840 2814.870 32.100 2815.190 ;
        RECT 34.600 2814.870 34.860 2815.190 ;
        RECT 31.900 2767.590 32.040 2814.870 ;
        RECT 31.840 2767.270 32.100 2767.590 ;
        RECT 34.140 2766.930 34.400 2767.250 ;
        RECT 34.200 2766.570 34.340 2766.930 ;
        RECT 32.300 2766.250 32.560 2766.570 ;
        RECT 34.140 2766.250 34.400 2766.570 ;
        RECT 32.360 2719.310 32.500 2766.250 ;
        RECT 32.300 2718.990 32.560 2719.310 ;
        RECT 34.600 2718.990 34.860 2719.310 ;
        RECT 34.660 2718.630 34.800 2718.990 ;
        RECT 31.840 2718.310 32.100 2718.630 ;
        RECT 34.600 2718.310 34.860 2718.630 ;
        RECT 31.900 2671.030 32.040 2718.310 ;
        RECT 31.840 2670.710 32.100 2671.030 ;
        RECT 34.140 2670.370 34.400 2670.690 ;
        RECT 34.200 2670.010 34.340 2670.370 ;
        RECT 32.300 2669.690 32.560 2670.010 ;
        RECT 34.140 2669.690 34.400 2670.010 ;
        RECT 32.360 2622.410 32.500 2669.690 ;
        RECT 32.300 2622.090 32.560 2622.410 ;
        RECT 34.600 2622.090 34.860 2622.410 ;
        RECT 34.660 2621.130 34.800 2622.090 ;
        RECT 33.740 2620.990 34.800 2621.130 ;
        RECT 33.740 2574.810 33.880 2620.990 ;
        RECT 33.680 2574.490 33.940 2574.810 ;
        RECT 34.140 2573.810 34.400 2574.130 ;
        RECT 34.200 2573.450 34.340 2573.810 ;
        RECT 32.300 2573.130 32.560 2573.450 ;
        RECT 34.140 2573.130 34.400 2573.450 ;
        RECT 32.360 2525.850 32.500 2573.130 ;
        RECT 32.300 2525.530 32.560 2525.850 ;
        RECT 34.600 2525.530 34.860 2525.850 ;
        RECT 34.660 2524.570 34.800 2525.530 ;
        RECT 33.740 2524.430 34.800 2524.570 ;
        RECT 33.740 2478.250 33.880 2524.430 ;
        RECT 33.680 2477.930 33.940 2478.250 ;
        RECT 34.140 2477.250 34.400 2477.570 ;
        RECT 34.200 2476.890 34.340 2477.250 ;
        RECT 32.300 2476.570 32.560 2476.890 ;
        RECT 34.140 2476.570 34.400 2476.890 ;
        RECT 32.360 2429.290 32.500 2476.570 ;
        RECT 32.300 2428.970 32.560 2429.290 ;
        RECT 34.600 2428.970 34.860 2429.290 ;
        RECT 34.660 2428.010 34.800 2428.970 ;
        RECT 33.740 2427.870 34.800 2428.010 ;
        RECT 33.740 2381.350 33.880 2427.870 ;
        RECT 33.680 2381.030 33.940 2381.350 ;
        RECT 34.140 2380.350 34.400 2380.670 ;
        RECT 34.200 2331.450 34.340 2380.350 ;
        RECT 33.740 2331.310 34.340 2331.450 ;
        RECT 33.740 2284.790 33.880 2331.310 ;
        RECT 33.680 2284.470 33.940 2284.790 ;
        RECT 34.140 2283.790 34.400 2284.110 ;
        RECT 34.200 2234.890 34.340 2283.790 ;
        RECT 33.740 2234.750 34.340 2234.890 ;
        RECT 33.740 2188.230 33.880 2234.750 ;
        RECT 33.680 2187.910 33.940 2188.230 ;
        RECT 34.140 2187.230 34.400 2187.550 ;
        RECT 34.200 1945.810 34.340 2187.230 ;
        RECT 34.140 1945.490 34.400 1945.810 ;
        RECT 31.840 1945.150 32.100 1945.470 ;
        RECT 31.900 1898.210 32.040 1945.150 ;
        RECT 31.840 1897.890 32.100 1898.210 ;
        RECT 34.140 1897.550 34.400 1897.870 ;
        RECT 34.200 1849.250 34.340 1897.550 ;
        RECT 34.140 1848.930 34.400 1849.250 ;
        RECT 31.840 1848.590 32.100 1848.910 ;
        RECT 31.900 1801.650 32.040 1848.590 ;
        RECT 31.840 1801.330 32.100 1801.650 ;
        RECT 34.140 1800.990 34.400 1801.310 ;
        RECT 34.200 1752.690 34.340 1800.990 ;
        RECT 34.140 1752.370 34.400 1752.690 ;
        RECT 31.840 1752.030 32.100 1752.350 ;
        RECT 31.900 1705.090 32.040 1752.030 ;
        RECT 31.840 1704.770 32.100 1705.090 ;
        RECT 34.140 1704.430 34.400 1704.750 ;
        RECT 34.200 1656.130 34.340 1704.430 ;
        RECT 34.140 1655.810 34.400 1656.130 ;
        RECT 30.460 1655.470 30.720 1655.790 ;
        RECT 30.520 1608.530 30.660 1655.470 ;
        RECT 30.460 1608.210 30.720 1608.530 ;
        RECT 34.140 1607.870 34.400 1608.190 ;
        RECT 34.200 1559.230 34.340 1607.870 ;
        RECT 34.140 1558.910 34.400 1559.230 ;
        RECT 31.840 1558.570 32.100 1558.890 ;
        RECT 31.900 1514.010 32.040 1558.570 ;
        RECT 31.840 1513.690 32.100 1514.010 ;
        RECT 34.140 1510.970 34.400 1511.290 ;
        RECT 34.200 1462.670 34.340 1510.970 ;
        RECT 34.140 1462.350 34.400 1462.670 ;
        RECT 30.000 1462.010 30.260 1462.330 ;
        RECT 30.060 1415.070 30.200 1462.010 ;
        RECT 30.000 1414.750 30.260 1415.070 ;
        RECT 34.140 1414.410 34.400 1414.730 ;
        RECT 34.200 1366.110 34.340 1414.410 ;
        RECT 34.140 1365.790 34.400 1366.110 ;
        RECT 30.000 1365.450 30.260 1365.770 ;
        RECT 30.060 1318.510 30.200 1365.450 ;
        RECT 30.000 1318.190 30.260 1318.510 ;
        RECT 34.140 1317.850 34.400 1318.170 ;
        RECT 34.200 1269.550 34.340 1317.850 ;
        RECT 34.140 1269.230 34.400 1269.550 ;
        RECT 30.000 1268.890 30.260 1269.210 ;
        RECT 30.060 1221.950 30.200 1268.890 ;
        RECT 30.000 1221.630 30.260 1221.950 ;
        RECT 34.140 1221.290 34.400 1221.610 ;
        RECT 34.200 1172.990 34.340 1221.290 ;
        RECT 34.140 1172.670 34.400 1172.990 ;
        RECT 30.000 1172.330 30.260 1172.650 ;
        RECT 30.060 1125.390 30.200 1172.330 ;
        RECT 30.000 1125.070 30.260 1125.390 ;
        RECT 34.140 1124.730 34.400 1125.050 ;
        RECT 34.200 1076.430 34.340 1124.730 ;
        RECT 34.140 1076.110 34.400 1076.430 ;
        RECT 30.000 1075.770 30.260 1076.090 ;
        RECT 30.060 1028.830 30.200 1075.770 ;
        RECT 30.000 1028.510 30.260 1028.830 ;
        RECT 34.140 1028.170 34.400 1028.490 ;
        RECT 34.200 979.870 34.340 1028.170 ;
        RECT 34.140 979.550 34.400 979.870 ;
        RECT 30.000 979.210 30.260 979.530 ;
        RECT 30.060 932.270 30.200 979.210 ;
        RECT 30.000 931.950 30.260 932.270 ;
        RECT 34.140 931.610 34.400 931.930 ;
        RECT 34.200 883.310 34.340 931.610 ;
        RECT 34.140 882.990 34.400 883.310 ;
        RECT 30.000 882.650 30.260 882.970 ;
        RECT 30.060 835.710 30.200 882.650 ;
        RECT 30.000 835.390 30.260 835.710 ;
        RECT 34.140 835.050 34.400 835.370 ;
        RECT 34.200 786.750 34.340 835.050 ;
        RECT 34.140 786.430 34.400 786.750 ;
        RECT 30.000 786.090 30.260 786.410 ;
        RECT 30.060 738.810 30.200 786.090 ;
        RECT 30.000 738.490 30.260 738.810 ;
        RECT 34.140 738.150 34.400 738.470 ;
        RECT 34.200 689.850 34.340 738.150 ;
        RECT 34.140 689.530 34.400 689.850 ;
        RECT 30.000 689.190 30.260 689.510 ;
        RECT 30.060 642.250 30.200 689.190 ;
        RECT 30.000 641.930 30.260 642.250 ;
        RECT 34.140 641.590 34.400 641.910 ;
        RECT 34.200 593.290 34.340 641.590 ;
        RECT 34.140 592.970 34.400 593.290 ;
        RECT 30.000 592.630 30.260 592.950 ;
        RECT 30.060 545.690 30.200 592.630 ;
        RECT 30.000 545.370 30.260 545.690 ;
        RECT 34.140 545.030 34.400 545.350 ;
        RECT 34.200 496.730 34.340 545.030 ;
        RECT 34.140 496.410 34.400 496.730 ;
        RECT 30.000 496.070 30.260 496.390 ;
        RECT 30.060 449.130 30.200 496.070 ;
        RECT 30.000 448.810 30.260 449.130 ;
        RECT 34.140 448.470 34.400 448.790 ;
        RECT 34.200 400.170 34.340 448.470 ;
        RECT 34.140 399.850 34.400 400.170 ;
        RECT 30.000 399.510 30.260 399.830 ;
        RECT 30.060 352.570 30.200 399.510 ;
        RECT 30.000 352.250 30.260 352.570 ;
        RECT 34.140 351.910 34.400 352.230 ;
        RECT 34.200 303.610 34.340 351.910 ;
        RECT 34.140 303.290 34.400 303.610 ;
        RECT 30.000 302.950 30.260 303.270 ;
        RECT 30.060 256.010 30.200 302.950 ;
        RECT 30.000 255.690 30.260 256.010 ;
        RECT 34.140 255.350 34.400 255.670 ;
        RECT 34.200 207.050 34.340 255.350 ;
        RECT 34.140 206.730 34.400 207.050 ;
        RECT 30.000 206.390 30.260 206.710 ;
        RECT 30.060 159.450 30.200 206.390 ;
        RECT 30.000 159.130 30.260 159.450 ;
        RECT 34.140 158.790 34.400 159.110 ;
        RECT 34.200 110.490 34.340 158.790 ;
        RECT 34.140 110.170 34.400 110.490 ;
        RECT 30.000 109.830 30.260 110.150 ;
        RECT 30.060 62.890 30.200 109.830 ;
        RECT 30.000 62.570 30.260 62.890 ;
        RECT 34.140 62.230 34.400 62.550 ;
        RECT 34.200 19.565 34.340 62.230 ;
        RECT 34.130 19.195 34.410 19.565 ;
        RECT 496.430 19.195 496.710 19.565 ;
        RECT 496.500 2.400 496.640 19.195 ;
        RECT 496.290 -4.800 496.850 2.400 ;
      LAYER via2 ;
        RECT 34.590 3157.440 34.870 3157.720 ;
        RECT 34.130 19.240 34.410 19.520 ;
        RECT 496.430 19.240 496.710 19.520 ;
      LAYER met3 ;
        RECT 35.000 3160.320 39.000 3160.920 ;
        RECT 34.565 3157.730 34.895 3157.745 ;
        RECT 35.270 3157.730 35.570 3160.320 ;
        RECT 34.565 3157.430 35.570 3157.730 ;
        RECT 34.565 3157.415 34.895 3157.430 ;
        RECT 34.105 19.530 34.435 19.545 ;
        RECT 496.405 19.530 496.735 19.545 ;
        RECT 34.105 19.230 496.735 19.530 ;
        RECT 34.105 19.215 34.435 19.230 ;
        RECT 496.405 19.215 496.735 19.230 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2501.110 3442.995 2501.390 3443.365 ;
        RECT 2501.180 3435.000 2501.320 3442.995 ;
        RECT 2501.150 3431.000 2501.430 3435.000 ;
        RECT 513.910 19.195 514.190 19.565 ;
        RECT 513.980 2.400 514.120 19.195 ;
        RECT 513.770 -4.800 514.330 2.400 ;
      LAYER via2 ;
        RECT 2501.110 3443.040 2501.390 3443.320 ;
        RECT 513.910 19.240 514.190 19.520 ;
      LAYER met3 ;
        RECT 2501.085 3443.330 2501.415 3443.345 ;
        RECT 2822.830 3443.330 2823.210 3443.340 ;
        RECT 2501.085 3443.030 2823.210 3443.330 ;
        RECT 2501.085 3443.015 2501.415 3443.030 ;
        RECT 2822.830 3443.020 2823.210 3443.030 ;
        RECT 513.885 19.530 514.215 19.545 ;
        RECT 2822.830 19.530 2823.210 19.540 ;
        RECT 513.885 19.230 2823.210 19.530 ;
        RECT 513.885 19.215 514.215 19.230 ;
        RECT 2822.830 19.220 2823.210 19.230 ;
      LAYER via3 ;
        RECT 2822.860 3443.020 2823.180 3443.340 ;
        RECT 2822.860 19.220 2823.180 19.540 ;
      LAYER met4 ;
        RECT 2822.855 3443.015 2823.185 3443.345 ;
        RECT 2822.870 19.545 2823.170 3443.015 ;
        RECT 2822.855 19.215 2823.185 19.545 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 531.830 29.820 532.150 29.880 ;
        RECT 2892.090 29.820 2892.410 29.880 ;
        RECT 531.830 29.680 2892.410 29.820 ;
        RECT 531.830 29.620 532.150 29.680 ;
        RECT 2892.090 29.620 2892.410 29.680 ;
      LAYER via ;
        RECT 531.860 29.620 532.120 29.880 ;
        RECT 2892.120 29.620 2892.380 29.880 ;
      LAYER met2 ;
        RECT 2892.110 2939.795 2892.390 2940.165 ;
        RECT 2892.180 29.910 2892.320 2939.795 ;
        RECT 531.860 29.590 532.120 29.910 ;
        RECT 2892.120 29.590 2892.380 29.910 ;
        RECT 531.920 2.400 532.060 29.590 ;
        RECT 531.710 -4.800 532.270 2.400 ;
      LAYER via2 ;
        RECT 2892.110 2939.840 2892.390 2940.120 ;
      LAYER met3 ;
        RECT 2881.000 2940.680 2885.000 2941.280 ;
        RECT 2884.510 2940.130 2884.810 2940.680 ;
        RECT 2892.085 2940.130 2892.415 2940.145 ;
        RECT 2884.510 2939.830 2892.415 2940.130 ;
        RECT 2892.085 2939.815 2892.415 2939.830 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2611.050 3443.675 2611.330 3444.045 ;
        RECT 2611.120 3435.000 2611.260 3443.675 ;
        RECT 2611.090 3431.000 2611.370 3435.000 ;
        RECT 549.790 37.555 550.070 37.925 ;
        RECT 549.860 2.400 550.000 37.555 ;
        RECT 549.650 -4.800 550.210 2.400 ;
      LAYER via2 ;
        RECT 2611.050 3443.720 2611.330 3444.000 ;
        RECT 549.790 37.600 550.070 37.880 ;
      LAYER met3 ;
        RECT 2611.025 3444.010 2611.355 3444.025 ;
        RECT 2830.190 3444.010 2830.570 3444.020 ;
        RECT 2611.025 3443.710 2830.570 3444.010 ;
        RECT 2611.025 3443.695 2611.355 3443.710 ;
        RECT 2830.190 3443.700 2830.570 3443.710 ;
        RECT 549.765 37.890 550.095 37.905 ;
        RECT 2830.190 37.890 2830.570 37.900 ;
        RECT 549.765 37.590 2830.570 37.890 ;
        RECT 549.765 37.575 550.095 37.590 ;
        RECT 2830.190 37.580 2830.570 37.590 ;
      LAYER via3 ;
        RECT 2830.220 3443.700 2830.540 3444.020 ;
        RECT 2830.220 37.580 2830.540 37.900 ;
      LAYER met4 ;
        RECT 2830.215 3443.695 2830.545 3444.025 ;
        RECT 2830.230 37.905 2830.530 3443.695 ;
        RECT 2830.215 37.575 2830.545 37.905 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2720.530 3444.355 2720.810 3444.725 ;
        RECT 2720.600 3435.000 2720.740 3444.355 ;
        RECT 2720.570 3431.000 2720.850 3435.000 ;
        RECT 567.730 38.235 568.010 38.605 ;
        RECT 567.800 2.400 567.940 38.235 ;
        RECT 567.590 -4.800 568.150 2.400 ;
      LAYER via2 ;
        RECT 2720.530 3444.400 2720.810 3444.680 ;
        RECT 567.730 38.280 568.010 38.560 ;
      LAYER met3 ;
        RECT 2720.505 3444.690 2720.835 3444.705 ;
        RECT 2823.750 3444.690 2824.130 3444.700 ;
        RECT 2720.505 3444.390 2824.130 3444.690 ;
        RECT 2720.505 3444.375 2720.835 3444.390 ;
        RECT 2823.750 3444.380 2824.130 3444.390 ;
        RECT 567.705 38.570 568.035 38.585 ;
        RECT 2823.750 38.570 2824.130 38.580 ;
        RECT 567.705 38.270 2824.130 38.570 ;
        RECT 567.705 38.255 568.035 38.270 ;
        RECT 2823.750 38.260 2824.130 38.270 ;
      LAYER via3 ;
        RECT 2823.780 3444.380 2824.100 3444.700 ;
        RECT 2823.780 38.260 2824.100 38.580 ;
      LAYER met4 ;
        RECT 2823.775 3444.375 2824.105 3444.705 ;
        RECT 2823.790 38.585 2824.090 3444.375 ;
        RECT 2823.775 38.255 2824.105 38.585 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2829.550 3431.690 2829.830 3431.805 ;
        RECT 2830.050 3431.690 2830.330 3435.000 ;
        RECT 2829.550 3431.550 2830.330 3431.690 ;
        RECT 2829.550 3431.435 2829.830 3431.550 ;
        RECT 2830.050 3431.000 2830.330 3431.550 ;
        RECT 585.670 15.795 585.950 16.165 ;
        RECT 585.740 2.400 585.880 15.795 ;
        RECT 585.530 -4.800 586.090 2.400 ;
      LAYER via2 ;
        RECT 2829.550 3431.480 2829.830 3431.760 ;
        RECT 585.670 15.840 585.950 16.120 ;
      LAYER met3 ;
        RECT 2829.525 3431.780 2829.855 3431.785 ;
        RECT 2829.270 3431.770 2829.855 3431.780 ;
        RECT 2829.070 3431.470 2829.855 3431.770 ;
        RECT 2829.270 3431.460 2829.855 3431.470 ;
        RECT 2829.525 3431.455 2829.855 3431.460 ;
        RECT 585.645 16.130 585.975 16.145 ;
        RECT 2829.270 16.130 2829.650 16.140 ;
        RECT 585.645 15.830 2829.650 16.130 ;
        RECT 585.645 15.815 585.975 15.830 ;
        RECT 2829.270 15.820 2829.650 15.830 ;
      LAYER via3 ;
        RECT 2829.300 3431.460 2829.620 3431.780 ;
        RECT 2829.300 15.820 2829.620 16.140 ;
      LAYER met4 ;
        RECT 2829.295 3431.455 2829.625 3431.785 ;
        RECT 2829.310 16.145 2829.610 3431.455 ;
        RECT 2829.295 15.815 2829.625 16.145 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 23.990 59.880 24.310 60.140 ;
        RECT 24.080 59.120 24.220 59.880 ;
        RECT 23.990 58.860 24.310 59.120 ;
        RECT 91.610 17.580 91.930 17.640 ;
        RECT 32.820 17.440 91.930 17.580 ;
        RECT 23.990 17.240 24.310 17.300 ;
        RECT 32.820 17.240 32.960 17.440 ;
        RECT 91.610 17.380 91.930 17.440 ;
        RECT 23.990 17.100 32.960 17.240 ;
        RECT 23.990 17.040 24.310 17.100 ;
      LAYER via ;
        RECT 24.020 59.880 24.280 60.140 ;
        RECT 24.020 58.860 24.280 59.120 ;
        RECT 24.020 17.040 24.280 17.300 ;
        RECT 91.640 17.380 91.900 17.640 ;
      LAYER met2 ;
        RECT 24.010 1953.115 24.290 1953.485 ;
        RECT 24.080 60.170 24.220 1953.115 ;
        RECT 24.020 59.850 24.280 60.170 ;
        RECT 24.020 58.830 24.280 59.150 ;
        RECT 24.080 17.330 24.220 58.830 ;
        RECT 91.640 17.350 91.900 17.670 ;
        RECT 24.020 17.010 24.280 17.330 ;
        RECT 91.700 2.400 91.840 17.350 ;
        RECT 91.490 -4.800 92.050 2.400 ;
      LAYER via2 ;
        RECT 24.010 1953.160 24.290 1953.440 ;
      LAYER met3 ;
        RECT 23.985 1953.450 24.315 1953.465 ;
        RECT 35.000 1953.450 39.000 1953.920 ;
        RECT 23.985 1953.320 39.000 1953.450 ;
        RECT 23.985 1953.150 35.570 1953.320 ;
        RECT 23.985 1953.135 24.315 1953.150 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2891.650 3049.955 2891.930 3050.325 ;
        RECT 2891.720 20.245 2891.860 3049.955 ;
        RECT 603.150 19.875 603.430 20.245 ;
        RECT 2891.650 19.875 2891.930 20.245 ;
        RECT 603.220 2.400 603.360 19.875 ;
        RECT 603.010 -4.800 603.570 2.400 ;
      LAYER via2 ;
        RECT 2891.650 3050.000 2891.930 3050.280 ;
        RECT 603.150 19.920 603.430 20.200 ;
        RECT 2891.650 19.920 2891.930 20.200 ;
      LAYER met3 ;
        RECT 2881.000 3050.290 2885.000 3050.760 ;
        RECT 2891.625 3050.290 2891.955 3050.305 ;
        RECT 2881.000 3050.160 2891.955 3050.290 ;
        RECT 2884.510 3049.990 2891.955 3050.160 ;
        RECT 2891.625 3049.975 2891.955 3049.990 ;
        RECT 603.125 20.210 603.455 20.225 ;
        RECT 2891.625 20.210 2891.955 20.225 ;
        RECT 603.125 19.910 2891.955 20.210 ;
        RECT 603.125 19.895 603.455 19.910 ;
        RECT 2891.625 19.895 2891.955 19.910 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 621.070 17.580 621.390 17.640 ;
        RECT 2891.170 17.580 2891.490 17.640 ;
        RECT 621.070 17.440 2891.490 17.580 ;
        RECT 621.070 17.380 621.390 17.440 ;
        RECT 2891.170 17.380 2891.490 17.440 ;
      LAYER via ;
        RECT 621.100 17.380 621.360 17.640 ;
        RECT 2891.200 17.380 2891.460 17.640 ;
      LAYER met2 ;
        RECT 2891.190 3160.115 2891.470 3160.485 ;
        RECT 2891.260 17.670 2891.400 3160.115 ;
        RECT 621.100 17.350 621.360 17.670 ;
        RECT 2891.200 17.350 2891.460 17.670 ;
        RECT 621.160 2.400 621.300 17.350 ;
        RECT 620.950 -4.800 621.510 2.400 ;
      LAYER via2 ;
        RECT 2891.190 3160.160 2891.470 3160.440 ;
      LAYER met3 ;
        RECT 2881.000 3160.450 2885.000 3160.920 ;
        RECT 2891.165 3160.450 2891.495 3160.465 ;
        RECT 2881.000 3160.320 2891.495 3160.450 ;
        RECT 2884.510 3160.150 2891.495 3160.320 ;
        RECT 2891.165 3160.135 2891.495 3160.150 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2893.490 2499.835 2893.770 2500.205 ;
        RECT 2893.560 17.525 2893.700 2499.835 ;
        RECT 115.550 17.155 115.830 17.525 ;
        RECT 2893.490 17.155 2893.770 17.525 ;
        RECT 115.620 2.400 115.760 17.155 ;
        RECT 115.410 -4.800 115.970 2.400 ;
      LAYER via2 ;
        RECT 2893.490 2499.880 2893.770 2500.160 ;
        RECT 115.550 17.200 115.830 17.480 ;
        RECT 2893.490 17.200 2893.770 17.480 ;
      LAYER met3 ;
        RECT 2881.000 2502.080 2885.000 2502.680 ;
        RECT 2884.510 2500.170 2884.810 2502.080 ;
        RECT 2893.465 2500.170 2893.795 2500.185 ;
        RECT 2884.510 2499.870 2893.795 2500.170 ;
        RECT 2893.465 2499.855 2893.795 2499.870 ;
        RECT 115.525 17.490 115.855 17.505 ;
        RECT 2893.465 17.490 2893.795 17.505 ;
        RECT 115.525 17.190 2893.795 17.490 ;
        RECT 115.525 17.175 115.855 17.190 ;
        RECT 2893.465 17.175 2893.795 17.190 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 46.145 18.445 46.315 20.315 ;
      LAYER mcon ;
        RECT 46.145 20.145 46.315 20.315 ;
      LAYER met1 ;
        RECT 35.030 20.300 35.350 20.360 ;
        RECT 46.085 20.300 46.375 20.345 ;
        RECT 35.030 20.160 46.375 20.300 ;
        RECT 35.030 20.100 35.350 20.160 ;
        RECT 46.085 20.115 46.375 20.160 ;
        RECT 46.085 18.600 46.375 18.645 ;
        RECT 139.450 18.600 139.770 18.660 ;
        RECT 46.085 18.460 139.770 18.600 ;
        RECT 46.085 18.415 46.375 18.460 ;
        RECT 139.450 18.400 139.770 18.460 ;
      LAYER via ;
        RECT 35.060 20.100 35.320 20.360 ;
        RECT 139.480 18.400 139.740 18.660 ;
      LAYER met2 ;
        RECT 35.050 2062.595 35.330 2062.965 ;
        RECT 35.120 20.390 35.260 2062.595 ;
        RECT 35.060 20.070 35.320 20.390 ;
        RECT 139.480 18.370 139.740 18.690 ;
        RECT 139.540 2.400 139.680 18.370 ;
        RECT 139.330 -4.800 139.890 2.400 ;
      LAYER via2 ;
        RECT 35.050 2062.640 35.330 2062.920 ;
      LAYER met3 ;
        RECT 35.000 2063.480 39.000 2064.080 ;
        RECT 35.270 2062.945 35.570 2063.480 ;
        RECT 35.025 2062.630 35.570 2062.945 ;
        RECT 35.025 2062.615 35.355 2062.630 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2655.710 35.000 2655.990 39.000 ;
        RECT 2655.740 27.045 2655.880 35.000 ;
        RECT 157.410 26.675 157.690 27.045 ;
        RECT 2655.670 26.675 2655.950 27.045 ;
        RECT 157.480 2.400 157.620 26.675 ;
        RECT 157.270 -4.800 157.830 2.400 ;
      LAYER via2 ;
        RECT 157.410 26.720 157.690 27.000 ;
        RECT 2655.670 26.720 2655.950 27.000 ;
      LAYER met3 ;
        RECT 157.385 27.010 157.715 27.025 ;
        RECT 2655.645 27.010 2655.975 27.025 ;
        RECT 157.385 26.710 2655.975 27.010 ;
        RECT 157.385 26.695 157.715 26.710 ;
        RECT 2655.645 26.695 2655.975 26.710 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2879.745 2427.345 2879.915 2463.215 ;
        RECT 2880.665 2089.045 2880.835 2142.595 ;
        RECT 2879.745 1896.945 2879.915 1950.495 ;
        RECT 2880.665 1829.285 2880.835 1883.515 ;
        RECT 2879.745 1796.645 2879.915 1806.335 ;
        RECT 2880.205 1659.285 2880.375 1690.395 ;
        RECT 2880.665 1578.025 2880.835 1597.575 ;
        RECT 2880.665 1124.465 2880.835 1125.315 ;
        RECT 2881.125 1125.145 2881.295 1184.135 ;
        RECT 2880.205 987.105 2880.375 1015.495 ;
        RECT 2880.205 873.885 2880.375 934.575 ;
        RECT 2880.205 789.225 2880.375 851.275 ;
        RECT 2880.665 627.725 2880.835 638.435 ;
        RECT 2879.745 521.985 2879.915 592.195 ;
        RECT 2881.585 592.025 2881.755 627.895 ;
        RECT 2880.665 406.725 2880.835 453.135 ;
        RECT 2880.665 83.385 2880.835 107.695 ;
      LAYER mcon ;
        RECT 2879.745 2463.045 2879.915 2463.215 ;
        RECT 2880.665 2142.425 2880.835 2142.595 ;
        RECT 2879.745 1950.325 2879.915 1950.495 ;
        RECT 2880.665 1883.345 2880.835 1883.515 ;
        RECT 2879.745 1806.165 2879.915 1806.335 ;
        RECT 2880.205 1690.225 2880.375 1690.395 ;
        RECT 2880.665 1597.405 2880.835 1597.575 ;
        RECT 2881.125 1183.965 2881.295 1184.135 ;
        RECT 2880.665 1125.145 2880.835 1125.315 ;
        RECT 2880.205 1015.325 2880.375 1015.495 ;
        RECT 2880.205 934.405 2880.375 934.575 ;
        RECT 2880.205 851.105 2880.375 851.275 ;
        RECT 2880.665 638.265 2880.835 638.435 ;
        RECT 2881.585 627.725 2881.755 627.895 ;
        RECT 2879.745 592.025 2879.915 592.195 ;
        RECT 2880.665 452.965 2880.835 453.135 ;
        RECT 2880.665 107.525 2880.835 107.695 ;
      LAYER met1 ;
        RECT 2879.670 2599.880 2879.990 2599.940 ;
        RECT 2881.510 2599.880 2881.830 2599.940 ;
        RECT 2879.670 2599.740 2881.830 2599.880 ;
        RECT 2879.670 2599.680 2879.990 2599.740 ;
        RECT 2881.510 2599.680 2881.830 2599.740 ;
        RECT 2879.685 2463.200 2879.975 2463.245 ;
        RECT 2880.130 2463.200 2880.450 2463.260 ;
        RECT 2879.685 2463.060 2880.450 2463.200 ;
        RECT 2879.685 2463.015 2879.975 2463.060 ;
        RECT 2880.130 2463.000 2880.450 2463.060 ;
        RECT 2879.670 2427.500 2879.990 2427.560 ;
        RECT 2879.475 2427.360 2879.990 2427.500 ;
        RECT 2879.670 2427.300 2879.990 2427.360 ;
        RECT 2879.670 2332.640 2879.990 2332.700 ;
        RECT 2879.670 2332.500 2880.820 2332.640 ;
        RECT 2879.670 2332.440 2879.990 2332.500 ;
        RECT 2880.680 2331.340 2880.820 2332.500 ;
        RECT 2880.590 2331.080 2880.910 2331.340 ;
        RECT 2880.130 2235.540 2880.450 2235.800 ;
        RECT 2880.220 2235.400 2880.360 2235.540 ;
        RECT 2880.590 2235.400 2880.910 2235.460 ;
        RECT 2880.220 2235.260 2880.910 2235.400 ;
        RECT 2880.590 2235.200 2880.910 2235.260 ;
        RECT 2880.130 2142.580 2880.450 2142.640 ;
        RECT 2880.605 2142.580 2880.895 2142.625 ;
        RECT 2880.130 2142.440 2880.895 2142.580 ;
        RECT 2880.130 2142.380 2880.450 2142.440 ;
        RECT 2880.605 2142.395 2880.895 2142.440 ;
        RECT 2880.590 2089.200 2880.910 2089.260 ;
        RECT 2880.395 2089.060 2880.910 2089.200 ;
        RECT 2880.590 2089.000 2880.910 2089.060 ;
        RECT 2879.670 1985.160 2879.990 1985.220 ;
        RECT 2880.590 1985.160 2880.910 1985.220 ;
        RECT 2879.670 1985.020 2880.910 1985.160 ;
        RECT 2879.670 1984.960 2879.990 1985.020 ;
        RECT 2880.590 1984.960 2880.910 1985.020 ;
        RECT 2879.670 1950.480 2879.990 1950.540 ;
        RECT 2879.475 1950.340 2879.990 1950.480 ;
        RECT 2879.670 1950.280 2879.990 1950.340 ;
        RECT 2879.685 1897.100 2879.975 1897.145 ;
        RECT 2880.590 1897.100 2880.910 1897.160 ;
        RECT 2879.685 1896.960 2880.910 1897.100 ;
        RECT 2879.685 1896.915 2879.975 1896.960 ;
        RECT 2880.590 1896.900 2880.910 1896.960 ;
        RECT 2880.590 1883.500 2880.910 1883.560 ;
        RECT 2880.395 1883.360 2880.910 1883.500 ;
        RECT 2880.590 1883.300 2880.910 1883.360 ;
        RECT 2879.670 1829.440 2879.990 1829.500 ;
        RECT 2880.605 1829.440 2880.895 1829.485 ;
        RECT 2879.670 1829.300 2880.895 1829.440 ;
        RECT 2879.670 1829.240 2879.990 1829.300 ;
        RECT 2880.605 1829.255 2880.895 1829.300 ;
        RECT 2879.670 1806.320 2879.990 1806.380 ;
        RECT 2879.475 1806.180 2879.990 1806.320 ;
        RECT 2879.670 1806.120 2879.990 1806.180 ;
        RECT 2879.670 1796.800 2879.990 1796.860 ;
        RECT 2879.475 1796.660 2879.990 1796.800 ;
        RECT 2879.670 1796.600 2879.990 1796.660 ;
        RECT 2879.670 1690.380 2879.990 1690.440 ;
        RECT 2880.145 1690.380 2880.435 1690.425 ;
        RECT 2879.670 1690.240 2880.435 1690.380 ;
        RECT 2879.670 1690.180 2879.990 1690.240 ;
        RECT 2880.145 1690.195 2880.435 1690.240 ;
        RECT 2879.670 1659.440 2879.990 1659.500 ;
        RECT 2880.145 1659.440 2880.435 1659.485 ;
        RECT 2879.670 1659.300 2880.435 1659.440 ;
        RECT 2879.670 1659.240 2879.990 1659.300 ;
        RECT 2880.145 1659.255 2880.435 1659.300 ;
        RECT 2879.670 1597.560 2879.990 1597.620 ;
        RECT 2880.605 1597.560 2880.895 1597.605 ;
        RECT 2879.670 1597.420 2880.895 1597.560 ;
        RECT 2879.670 1597.360 2879.990 1597.420 ;
        RECT 2880.605 1597.375 2880.895 1597.420 ;
        RECT 2879.670 1578.180 2879.990 1578.240 ;
        RECT 2880.605 1578.180 2880.895 1578.225 ;
        RECT 2879.670 1578.040 2880.895 1578.180 ;
        RECT 2879.670 1577.980 2879.990 1578.040 ;
        RECT 2880.605 1577.995 2880.895 1578.040 ;
        RECT 2879.670 1442.520 2879.990 1442.580 ;
        RECT 2880.590 1442.520 2880.910 1442.580 ;
        RECT 2879.670 1442.380 2880.910 1442.520 ;
        RECT 2879.670 1442.320 2879.990 1442.380 ;
        RECT 2880.590 1442.320 2880.910 1442.380 ;
        RECT 2879.670 1314.680 2879.990 1314.740 ;
        RECT 2881.050 1314.680 2881.370 1314.740 ;
        RECT 2879.670 1314.540 2881.370 1314.680 ;
        RECT 2879.670 1314.480 2879.990 1314.540 ;
        RECT 2881.050 1314.480 2881.370 1314.540 ;
        RECT 2881.050 1184.120 2881.370 1184.180 ;
        RECT 2880.855 1183.980 2881.370 1184.120 ;
        RECT 2881.050 1183.920 2881.370 1183.980 ;
        RECT 2880.605 1125.300 2880.895 1125.345 ;
        RECT 2881.065 1125.300 2881.355 1125.345 ;
        RECT 2880.605 1125.160 2881.355 1125.300 ;
        RECT 2880.605 1125.115 2880.895 1125.160 ;
        RECT 2881.065 1125.115 2881.355 1125.160 ;
        RECT 2880.590 1124.620 2880.910 1124.680 ;
        RECT 2880.395 1124.480 2880.910 1124.620 ;
        RECT 2880.590 1124.420 2880.910 1124.480 ;
        RECT 2880.130 1015.480 2880.450 1015.540 ;
        RECT 2879.935 1015.340 2880.450 1015.480 ;
        RECT 2880.130 1015.280 2880.450 1015.340 ;
        RECT 2880.145 987.260 2880.435 987.305 ;
        RECT 2880.145 987.120 2880.820 987.260 ;
        RECT 2880.145 987.075 2880.435 987.120 ;
        RECT 2880.680 986.980 2880.820 987.120 ;
        RECT 2880.590 986.720 2880.910 986.980 ;
        RECT 2879.670 934.560 2879.990 934.620 ;
        RECT 2880.145 934.560 2880.435 934.605 ;
        RECT 2879.670 934.420 2880.435 934.560 ;
        RECT 2879.670 934.360 2879.990 934.420 ;
        RECT 2880.145 934.375 2880.435 934.420 ;
        RECT 2879.670 874.040 2879.990 874.100 ;
        RECT 2880.145 874.040 2880.435 874.085 ;
        RECT 2879.670 873.900 2880.435 874.040 ;
        RECT 2879.670 873.840 2879.990 873.900 ;
        RECT 2880.145 873.855 2880.435 873.900 ;
        RECT 2879.670 851.260 2879.990 851.320 ;
        RECT 2880.145 851.260 2880.435 851.305 ;
        RECT 2879.670 851.120 2880.435 851.260 ;
        RECT 2879.670 851.060 2879.990 851.120 ;
        RECT 2880.145 851.075 2880.435 851.120 ;
        RECT 2880.145 789.380 2880.435 789.425 ;
        RECT 2880.590 789.380 2880.910 789.440 ;
        RECT 2880.145 789.240 2880.910 789.380 ;
        RECT 2880.145 789.195 2880.435 789.240 ;
        RECT 2880.590 789.180 2880.910 789.240 ;
        RECT 2879.670 699.620 2879.990 699.680 ;
        RECT 2880.590 699.620 2880.910 699.680 ;
        RECT 2879.670 699.480 2880.910 699.620 ;
        RECT 2879.670 699.420 2879.990 699.480 ;
        RECT 2880.590 699.420 2880.910 699.480 ;
        RECT 2879.670 638.420 2879.990 638.480 ;
        RECT 2880.605 638.420 2880.895 638.465 ;
        RECT 2879.670 638.280 2880.895 638.420 ;
        RECT 2879.670 638.220 2879.990 638.280 ;
        RECT 2880.605 638.235 2880.895 638.280 ;
        RECT 2880.605 627.880 2880.895 627.925 ;
        RECT 2881.525 627.880 2881.815 627.925 ;
        RECT 2880.605 627.740 2881.815 627.880 ;
        RECT 2880.605 627.695 2880.895 627.740 ;
        RECT 2881.525 627.695 2881.815 627.740 ;
        RECT 2879.685 592.180 2879.975 592.225 ;
        RECT 2881.525 592.180 2881.815 592.225 ;
        RECT 2879.685 592.040 2881.815 592.180 ;
        RECT 2879.685 591.995 2879.975 592.040 ;
        RECT 2881.525 591.995 2881.815 592.040 ;
        RECT 2879.670 522.140 2879.990 522.200 ;
        RECT 2879.475 522.000 2879.990 522.140 ;
        RECT 2879.670 521.940 2879.990 522.000 ;
        RECT 2879.670 453.120 2879.990 453.180 ;
        RECT 2880.605 453.120 2880.895 453.165 ;
        RECT 2879.670 452.980 2880.895 453.120 ;
        RECT 2879.670 452.920 2879.990 452.980 ;
        RECT 2880.605 452.935 2880.895 452.980 ;
        RECT 2880.590 406.880 2880.910 406.940 ;
        RECT 2880.395 406.740 2880.910 406.880 ;
        RECT 2880.590 406.680 2880.910 406.740 ;
        RECT 2880.590 307.940 2880.910 308.000 ;
        RECT 2881.970 307.940 2882.290 308.000 ;
        RECT 2880.590 307.800 2882.290 307.940 ;
        RECT 2880.590 307.740 2880.910 307.800 ;
        RECT 2881.970 307.740 2882.290 307.800 ;
        RECT 2880.590 169.220 2880.910 169.280 ;
        RECT 2881.970 169.220 2882.290 169.280 ;
        RECT 2880.590 169.080 2882.290 169.220 ;
        RECT 2880.590 169.020 2880.910 169.080 ;
        RECT 2881.970 169.020 2882.290 169.080 ;
        RECT 2880.590 107.680 2880.910 107.740 ;
        RECT 2880.395 107.540 2880.910 107.680 ;
        RECT 2880.590 107.480 2880.910 107.540 ;
        RECT 2879.670 83.540 2879.990 83.600 ;
        RECT 2880.605 83.540 2880.895 83.585 ;
        RECT 2879.670 83.400 2880.895 83.540 ;
        RECT 2879.670 83.340 2879.990 83.400 ;
        RECT 2880.605 83.355 2880.895 83.400 ;
      LAYER via ;
        RECT 2879.700 2599.680 2879.960 2599.940 ;
        RECT 2881.540 2599.680 2881.800 2599.940 ;
        RECT 2880.160 2463.000 2880.420 2463.260 ;
        RECT 2879.700 2427.300 2879.960 2427.560 ;
        RECT 2879.700 2332.440 2879.960 2332.700 ;
        RECT 2880.620 2331.080 2880.880 2331.340 ;
        RECT 2880.160 2235.540 2880.420 2235.800 ;
        RECT 2880.620 2235.200 2880.880 2235.460 ;
        RECT 2880.160 2142.380 2880.420 2142.640 ;
        RECT 2880.620 2089.000 2880.880 2089.260 ;
        RECT 2879.700 1984.960 2879.960 1985.220 ;
        RECT 2880.620 1984.960 2880.880 1985.220 ;
        RECT 2879.700 1950.280 2879.960 1950.540 ;
        RECT 2880.620 1896.900 2880.880 1897.160 ;
        RECT 2880.620 1883.300 2880.880 1883.560 ;
        RECT 2879.700 1829.240 2879.960 1829.500 ;
        RECT 2879.700 1806.120 2879.960 1806.380 ;
        RECT 2879.700 1796.600 2879.960 1796.860 ;
        RECT 2879.700 1690.180 2879.960 1690.440 ;
        RECT 2879.700 1659.240 2879.960 1659.500 ;
        RECT 2879.700 1597.360 2879.960 1597.620 ;
        RECT 2879.700 1577.980 2879.960 1578.240 ;
        RECT 2879.700 1442.320 2879.960 1442.580 ;
        RECT 2880.620 1442.320 2880.880 1442.580 ;
        RECT 2879.700 1314.480 2879.960 1314.740 ;
        RECT 2881.080 1314.480 2881.340 1314.740 ;
        RECT 2881.080 1183.920 2881.340 1184.180 ;
        RECT 2880.620 1124.420 2880.880 1124.680 ;
        RECT 2880.160 1015.280 2880.420 1015.540 ;
        RECT 2880.620 986.720 2880.880 986.980 ;
        RECT 2879.700 934.360 2879.960 934.620 ;
        RECT 2879.700 873.840 2879.960 874.100 ;
        RECT 2879.700 851.060 2879.960 851.320 ;
        RECT 2880.620 789.180 2880.880 789.440 ;
        RECT 2879.700 699.420 2879.960 699.680 ;
        RECT 2880.620 699.420 2880.880 699.680 ;
        RECT 2879.700 638.220 2879.960 638.480 ;
        RECT 2879.700 521.940 2879.960 522.200 ;
        RECT 2879.700 452.920 2879.960 453.180 ;
        RECT 2880.620 406.680 2880.880 406.940 ;
        RECT 2880.620 307.740 2880.880 308.000 ;
        RECT 2882.000 307.740 2882.260 308.000 ;
        RECT 2880.620 169.020 2880.880 169.280 ;
        RECT 2882.000 169.020 2882.260 169.280 ;
        RECT 2880.620 107.480 2880.880 107.740 ;
        RECT 2879.700 83.340 2879.960 83.600 ;
      LAYER met2 ;
        RECT 2881.530 2608.635 2881.810 2609.005 ;
        RECT 2881.600 2599.970 2881.740 2608.635 ;
        RECT 2879.700 2599.650 2879.960 2599.970 ;
        RECT 2881.540 2599.650 2881.800 2599.970 ;
        RECT 2879.760 2591.210 2879.900 2599.650 ;
        RECT 2877.920 2591.070 2879.900 2591.210 ;
        RECT 2877.920 2574.210 2878.060 2591.070 ;
        RECT 2877.920 2574.070 2878.520 2574.210 ;
        RECT 2878.380 2551.090 2878.520 2574.070 ;
        RECT 2878.380 2550.950 2880.360 2551.090 ;
        RECT 2880.220 2515.730 2880.360 2550.950 ;
        RECT 2878.380 2515.590 2880.360 2515.730 ;
        RECT 2878.380 2476.970 2878.520 2515.590 ;
        RECT 2878.380 2476.830 2880.360 2476.970 ;
        RECT 2880.220 2463.290 2880.360 2476.830 ;
        RECT 2880.160 2462.970 2880.420 2463.290 ;
        RECT 2879.700 2427.270 2879.960 2427.590 ;
        RECT 2879.760 2381.090 2879.900 2427.270 ;
        RECT 2878.380 2380.950 2879.900 2381.090 ;
        RECT 2878.380 2380.410 2878.520 2380.950 ;
        RECT 2878.380 2380.270 2879.440 2380.410 ;
        RECT 2879.300 2342.330 2879.440 2380.270 ;
        RECT 2879.300 2342.190 2879.900 2342.330 ;
        RECT 2879.760 2332.730 2879.900 2342.190 ;
        RECT 2879.700 2332.410 2879.960 2332.730 ;
        RECT 2880.620 2331.050 2880.880 2331.370 ;
        RECT 2880.680 2318.530 2880.820 2331.050 ;
        RECT 2880.220 2318.390 2880.820 2318.530 ;
        RECT 2880.220 2235.830 2880.360 2318.390 ;
        RECT 2880.160 2235.510 2880.420 2235.830 ;
        RECT 2880.620 2235.170 2880.880 2235.490 ;
        RECT 2880.680 2187.290 2880.820 2235.170 ;
        RECT 2880.220 2187.150 2880.820 2187.290 ;
        RECT 2880.220 2142.670 2880.360 2187.150 ;
        RECT 2880.160 2142.350 2880.420 2142.670 ;
        RECT 2880.620 2088.970 2880.880 2089.290 ;
        RECT 2880.680 1985.250 2880.820 2088.970 ;
        RECT 2879.700 1984.930 2879.960 1985.250 ;
        RECT 2880.620 1984.930 2880.880 1985.250 ;
        RECT 2879.760 1950.570 2879.900 1984.930 ;
        RECT 2879.700 1950.250 2879.960 1950.570 ;
        RECT 2880.620 1896.870 2880.880 1897.190 ;
        RECT 2880.680 1883.590 2880.820 1896.870 ;
        RECT 2880.620 1883.270 2880.880 1883.590 ;
        RECT 2879.700 1829.210 2879.960 1829.530 ;
        RECT 2879.760 1806.410 2879.900 1829.210 ;
        RECT 2879.700 1806.090 2879.960 1806.410 ;
        RECT 2879.700 1796.570 2879.960 1796.890 ;
        RECT 2879.760 1795.610 2879.900 1796.570 ;
        RECT 2878.380 1795.470 2879.900 1795.610 ;
        RECT 2878.380 1762.970 2878.520 1795.470 ;
        RECT 2878.380 1762.830 2880.820 1762.970 ;
        RECT 2880.680 1735.090 2880.820 1762.830 ;
        RECT 2879.760 1734.950 2880.820 1735.090 ;
        RECT 2879.760 1690.470 2879.900 1734.950 ;
        RECT 2879.700 1690.150 2879.960 1690.470 ;
        RECT 2879.700 1659.210 2879.960 1659.530 ;
        RECT 2879.760 1641.250 2879.900 1659.210 ;
        RECT 2877.920 1641.110 2879.900 1641.250 ;
        RECT 2877.920 1639.210 2878.060 1641.110 ;
        RECT 2877.920 1639.070 2878.520 1639.210 ;
        RECT 2878.380 1597.730 2878.520 1639.070 ;
        RECT 2878.380 1597.650 2879.900 1597.730 ;
        RECT 2878.380 1597.590 2879.960 1597.650 ;
        RECT 2879.700 1597.330 2879.960 1597.590 ;
        RECT 2879.700 1578.010 2879.960 1578.270 ;
        RECT 2879.300 1577.950 2879.960 1578.010 ;
        RECT 2879.300 1577.870 2879.900 1577.950 ;
        RECT 2879.300 1563.050 2879.440 1577.870 ;
        RECT 2878.380 1562.910 2879.440 1563.050 ;
        RECT 2878.380 1461.730 2878.520 1562.910 ;
        RECT 2878.380 1461.590 2878.980 1461.730 ;
        RECT 2878.840 1443.370 2878.980 1461.590 ;
        RECT 2878.840 1443.230 2879.900 1443.370 ;
        RECT 2879.760 1442.610 2879.900 1443.230 ;
        RECT 2879.700 1442.290 2879.960 1442.610 ;
        RECT 2880.620 1442.290 2880.880 1442.610 ;
        RECT 2880.680 1431.810 2880.820 1442.290 ;
        RECT 2877.920 1431.670 2880.820 1431.810 ;
        RECT 2877.920 1399.170 2878.060 1431.670 ;
        RECT 2877.460 1399.030 2878.060 1399.170 ;
        RECT 2877.460 1397.810 2877.600 1399.030 ;
        RECT 2877.000 1397.670 2877.600 1397.810 ;
        RECT 2877.000 1367.210 2877.140 1397.670 ;
        RECT 2877.000 1367.070 2877.600 1367.210 ;
        RECT 2877.460 1365.850 2877.600 1367.070 ;
        RECT 2877.000 1365.710 2877.600 1365.850 ;
        RECT 2877.000 1348.850 2877.140 1365.710 ;
        RECT 2877.000 1348.710 2877.600 1348.850 ;
        RECT 2877.460 1314.850 2877.600 1348.710 ;
        RECT 2877.460 1314.770 2879.900 1314.850 ;
        RECT 2877.460 1314.710 2879.960 1314.770 ;
        RECT 2879.700 1314.450 2879.960 1314.710 ;
        RECT 2881.080 1314.450 2881.340 1314.770 ;
        RECT 2881.140 1184.210 2881.280 1314.450 ;
        RECT 2881.080 1183.890 2881.340 1184.210 ;
        RECT 2880.620 1124.390 2880.880 1124.710 ;
        RECT 2880.680 1087.050 2880.820 1124.390 ;
        RECT 2880.220 1086.910 2880.820 1087.050 ;
        RECT 2880.220 1015.570 2880.360 1086.910 ;
        RECT 2880.160 1015.250 2880.420 1015.570 ;
        RECT 2880.620 986.690 2880.880 987.010 ;
        RECT 2880.680 963.290 2880.820 986.690 ;
        RECT 2880.220 963.150 2880.820 963.290 ;
        RECT 2880.220 961.250 2880.360 963.150 ;
        RECT 2879.300 961.110 2880.360 961.250 ;
        RECT 2879.300 934.730 2879.440 961.110 ;
        RECT 2879.300 934.650 2879.900 934.730 ;
        RECT 2879.300 934.590 2879.960 934.650 ;
        RECT 2879.700 934.330 2879.960 934.590 ;
        RECT 2879.700 873.810 2879.960 874.130 ;
        RECT 2879.760 873.530 2879.900 873.810 ;
        RECT 2879.300 873.390 2879.900 873.530 ;
        RECT 2879.300 851.770 2879.440 873.390 ;
        RECT 2879.300 851.630 2879.900 851.770 ;
        RECT 2879.760 851.350 2879.900 851.630 ;
        RECT 2879.700 851.030 2879.960 851.350 ;
        RECT 2880.620 789.150 2880.880 789.470 ;
        RECT 2880.680 699.710 2880.820 789.150 ;
        RECT 2879.700 699.390 2879.960 699.710 ;
        RECT 2880.620 699.390 2880.880 699.710 ;
        RECT 2879.760 686.530 2879.900 699.390 ;
        RECT 2878.380 686.390 2879.900 686.530 ;
        RECT 2878.380 638.930 2878.520 686.390 ;
        RECT 2878.380 638.790 2879.900 638.930 ;
        RECT 2879.760 638.510 2879.900 638.790 ;
        RECT 2879.700 638.190 2879.960 638.510 ;
        RECT 2879.700 521.970 2879.960 522.230 ;
        RECT 2878.380 521.910 2879.960 521.970 ;
        RECT 2878.380 521.830 2879.900 521.910 ;
        RECT 2878.380 461.450 2878.520 521.830 ;
        RECT 2878.380 461.310 2879.900 461.450 ;
        RECT 2879.760 453.210 2879.900 461.310 ;
        RECT 2879.700 452.890 2879.960 453.210 ;
        RECT 2880.620 406.650 2880.880 406.970 ;
        RECT 2880.680 308.030 2880.820 406.650 ;
        RECT 2880.620 307.710 2880.880 308.030 ;
        RECT 2882.000 307.710 2882.260 308.030 ;
        RECT 2882.060 169.310 2882.200 307.710 ;
        RECT 2880.620 168.990 2880.880 169.310 ;
        RECT 2882.000 168.990 2882.260 169.310 ;
        RECT 2880.680 107.770 2880.820 168.990 ;
        RECT 2880.620 107.450 2880.880 107.770 ;
        RECT 2879.700 83.370 2879.960 83.630 ;
        RECT 2877.460 83.310 2879.960 83.370 ;
        RECT 2877.460 83.230 2879.900 83.310 ;
        RECT 2877.460 75.890 2877.600 83.230 ;
        RECT 2877.000 75.750 2877.600 75.890 ;
        RECT 2877.000 74.530 2877.140 75.750 ;
        RECT 2877.000 74.390 2877.600 74.530 ;
        RECT 2877.460 58.890 2877.600 74.390 ;
        RECT 2877.460 58.750 2878.060 58.890 ;
        RECT 2877.920 18.885 2878.060 58.750 ;
        RECT 174.890 18.515 175.170 18.885 ;
        RECT 2877.850 18.515 2878.130 18.885 ;
        RECT 174.960 2.400 175.100 18.515 ;
        RECT 174.750 -4.800 175.310 2.400 ;
      LAYER via2 ;
        RECT 2881.530 2608.680 2881.810 2608.960 ;
        RECT 174.890 18.560 175.170 18.840 ;
        RECT 2877.850 18.560 2878.130 18.840 ;
      LAYER met3 ;
        RECT 2881.000 2611.560 2885.000 2612.160 ;
        RECT 2881.750 2608.985 2882.050 2611.560 ;
        RECT 2881.505 2608.670 2882.050 2608.985 ;
        RECT 2881.505 2608.655 2881.835 2608.670 ;
        RECT 174.865 18.850 175.195 18.865 ;
        RECT 2877.825 18.850 2878.155 18.865 ;
        RECT 174.865 18.550 2878.155 18.850 ;
        RECT 174.865 18.535 175.195 18.550 ;
        RECT 2877.825 18.535 2878.155 18.550 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 23.530 14.860 23.850 14.920 ;
        RECT 192.810 14.860 193.130 14.920 ;
        RECT 23.530 14.720 193.130 14.860 ;
        RECT 23.530 14.660 23.850 14.720 ;
        RECT 192.810 14.660 193.130 14.720 ;
      LAYER via ;
        RECT 23.560 14.660 23.820 14.920 ;
        RECT 192.840 14.660 193.100 14.920 ;
      LAYER met2 ;
        RECT 24.470 2170.035 24.750 2170.405 ;
        RECT 24.540 59.570 24.680 2170.035 ;
        RECT 23.620 59.430 24.680 59.570 ;
        RECT 23.620 14.950 23.760 59.430 ;
        RECT 23.560 14.630 23.820 14.950 ;
        RECT 192.840 14.630 193.100 14.950 ;
        RECT 192.900 2.400 193.040 14.630 ;
        RECT 192.690 -4.800 193.250 2.400 ;
      LAYER via2 ;
        RECT 24.470 2170.080 24.750 2170.360 ;
      LAYER met3 ;
        RECT 35.000 2172.960 39.000 2173.560 ;
        RECT 24.445 2170.370 24.775 2170.385 ;
        RECT 35.270 2170.370 35.570 2172.960 ;
        RECT 24.445 2170.070 35.570 2170.370 ;
        RECT 24.445 2170.055 24.775 2170.070 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2706.770 35.000 2707.050 39.000 ;
        RECT 2706.800 26.365 2706.940 35.000 ;
        RECT 210.770 25.995 211.050 26.365 ;
        RECT 2706.730 25.995 2707.010 26.365 ;
        RECT 210.840 2.400 210.980 25.995 ;
        RECT 210.630 -4.800 211.190 2.400 ;
      LAYER via2 ;
        RECT 210.770 26.040 211.050 26.320 ;
        RECT 2706.730 26.040 2707.010 26.320 ;
      LAYER met3 ;
        RECT 210.745 26.330 211.075 26.345 ;
        RECT 2706.705 26.330 2707.035 26.345 ;
        RECT 210.745 26.030 2707.035 26.330 ;
        RECT 210.745 26.015 211.075 26.030 ;
        RECT 2706.705 26.015 2707.035 26.030 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 24.450 15.880 24.770 15.940 ;
        RECT 228.690 15.880 229.010 15.940 ;
        RECT 24.450 15.740 229.010 15.880 ;
        RECT 24.450 15.680 24.770 15.740 ;
        RECT 228.690 15.680 229.010 15.740 ;
      LAYER via ;
        RECT 24.480 15.680 24.740 15.940 ;
        RECT 228.720 15.680 228.980 15.940 ;
      LAYER met2 ;
        RECT 24.930 2279.515 25.210 2279.885 ;
        RECT 25.000 58.890 25.140 2279.515 ;
        RECT 24.540 58.750 25.140 58.890 ;
        RECT 24.540 15.970 24.680 58.750 ;
        RECT 24.480 15.650 24.740 15.970 ;
        RECT 228.720 15.650 228.980 15.970 ;
        RECT 228.780 2.400 228.920 15.650 ;
        RECT 228.570 -4.800 229.130 2.400 ;
      LAYER via2 ;
        RECT 24.930 2279.560 25.210 2279.840 ;
      LAYER met3 ;
        RECT 35.000 2282.440 39.000 2283.040 ;
        RECT 24.905 2279.850 25.235 2279.865 ;
        RECT 35.270 2279.850 35.570 2282.440 ;
        RECT 24.905 2279.550 35.570 2279.850 ;
        RECT 24.905 2279.535 25.235 2279.550 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 50.210 20.300 50.530 20.360 ;
        RECT 467.430 20.300 467.750 20.360 ;
        RECT 50.210 20.160 467.750 20.300 ;
        RECT 50.210 20.100 50.530 20.160 ;
        RECT 467.430 20.100 467.750 20.160 ;
      LAYER via ;
        RECT 50.240 20.100 50.500 20.360 ;
        RECT 467.460 20.100 467.720 20.360 ;
      LAYER met2 ;
        RECT 467.490 35.000 467.770 39.000 ;
        RECT 467.520 20.390 467.660 35.000 ;
        RECT 50.240 20.070 50.500 20.390 ;
        RECT 467.460 20.070 467.720 20.390 ;
        RECT 50.300 2.400 50.440 20.070 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 252.610 15.540 252.930 15.600 ;
        RECT 976.190 15.540 976.510 15.600 ;
        RECT 252.610 15.400 976.510 15.540 ;
        RECT 252.610 15.340 252.930 15.400 ;
        RECT 976.190 15.340 976.510 15.400 ;
      LAYER via ;
        RECT 252.640 15.340 252.900 15.600 ;
        RECT 976.220 15.340 976.480 15.600 ;
      LAYER met2 ;
        RECT 976.250 35.000 976.530 39.000 ;
        RECT 976.280 15.630 976.420 35.000 ;
        RECT 252.640 15.310 252.900 15.630 ;
        RECT 976.220 15.310 976.480 15.630 ;
        RECT 252.700 2.400 252.840 15.310 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 270.090 21.660 270.410 21.720 ;
        RECT 1027.250 21.660 1027.570 21.720 ;
        RECT 270.090 21.520 1027.570 21.660 ;
        RECT 270.090 21.460 270.410 21.520 ;
        RECT 1027.250 21.460 1027.570 21.520 ;
      LAYER via ;
        RECT 270.120 21.460 270.380 21.720 ;
        RECT 1027.280 21.460 1027.540 21.720 ;
      LAYER met2 ;
        RECT 1027.310 35.000 1027.590 39.000 ;
        RECT 1027.340 21.750 1027.480 35.000 ;
        RECT 270.120 21.430 270.380 21.750 ;
        RECT 1027.280 21.430 1027.540 21.750 ;
        RECT 270.180 2.400 270.320 21.430 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 288.030 22.000 288.350 22.060 ;
        RECT 1077.850 22.000 1078.170 22.060 ;
        RECT 288.030 21.860 1078.170 22.000 ;
        RECT 288.030 21.800 288.350 21.860 ;
        RECT 1077.850 21.800 1078.170 21.860 ;
      LAYER via ;
        RECT 288.060 21.800 288.320 22.060 ;
        RECT 1077.880 21.800 1078.140 22.060 ;
      LAYER met2 ;
        RECT 1077.910 35.000 1078.190 39.000 ;
        RECT 1077.940 22.090 1078.080 35.000 ;
        RECT 288.060 21.770 288.320 22.090 ;
        RECT 1077.880 21.770 1078.140 22.090 ;
        RECT 288.120 2.400 288.260 21.770 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 305.970 15.880 306.290 15.940 ;
        RECT 1128.910 15.880 1129.230 15.940 ;
        RECT 305.970 15.740 1129.230 15.880 ;
        RECT 305.970 15.680 306.290 15.740 ;
        RECT 1128.910 15.680 1129.230 15.740 ;
      LAYER via ;
        RECT 306.000 15.680 306.260 15.940 ;
        RECT 1128.940 15.680 1129.200 15.940 ;
      LAYER met2 ;
        RECT 1128.970 35.000 1129.250 39.000 ;
        RECT 1129.000 15.970 1129.140 35.000 ;
        RECT 306.000 15.650 306.260 15.970 ;
        RECT 1128.940 15.650 1129.200 15.970 ;
        RECT 306.060 2.400 306.200 15.650 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 323.910 22.340 324.230 22.400 ;
        RECT 1179.970 22.340 1180.290 22.400 ;
        RECT 323.910 22.200 1180.290 22.340 ;
        RECT 323.910 22.140 324.230 22.200 ;
        RECT 1179.970 22.140 1180.290 22.200 ;
      LAYER via ;
        RECT 323.940 22.140 324.200 22.400 ;
        RECT 1180.000 22.140 1180.260 22.400 ;
      LAYER met2 ;
        RECT 1180.030 35.000 1180.310 39.000 ;
        RECT 1180.060 22.430 1180.200 35.000 ;
        RECT 323.940 22.110 324.200 22.430 ;
        RECT 1180.000 22.110 1180.260 22.430 ;
        RECT 324.000 2.400 324.140 22.110 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 341.390 22.680 341.710 22.740 ;
        RECT 1230.570 22.680 1230.890 22.740 ;
        RECT 341.390 22.540 1230.890 22.680 ;
        RECT 341.390 22.480 341.710 22.540 ;
        RECT 1230.570 22.480 1230.890 22.540 ;
      LAYER via ;
        RECT 341.420 22.480 341.680 22.740 ;
        RECT 1230.600 22.480 1230.860 22.740 ;
      LAYER met2 ;
        RECT 1230.630 35.000 1230.910 39.000 ;
        RECT 1230.660 22.770 1230.800 35.000 ;
        RECT 341.420 22.450 341.680 22.770 ;
        RECT 1230.600 22.450 1230.860 22.770 ;
        RECT 341.480 2.400 341.620 22.450 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 359.330 16.220 359.650 16.280 ;
        RECT 1281.630 16.220 1281.950 16.280 ;
        RECT 359.330 16.080 1281.950 16.220 ;
        RECT 359.330 16.020 359.650 16.080 ;
        RECT 1281.630 16.020 1281.950 16.080 ;
      LAYER via ;
        RECT 359.360 16.020 359.620 16.280 ;
        RECT 1281.660 16.020 1281.920 16.280 ;
      LAYER met2 ;
        RECT 1281.690 35.000 1281.970 39.000 ;
        RECT 1281.720 16.310 1281.860 35.000 ;
        RECT 359.360 15.990 359.620 16.310 ;
        RECT 1281.660 15.990 1281.920 16.310 ;
        RECT 359.420 2.400 359.560 15.990 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 377.270 23.020 377.590 23.080 ;
        RECT 1332.690 23.020 1333.010 23.080 ;
        RECT 377.270 22.880 1333.010 23.020 ;
        RECT 377.270 22.820 377.590 22.880 ;
        RECT 1332.690 22.820 1333.010 22.880 ;
      LAYER via ;
        RECT 377.300 22.820 377.560 23.080 ;
        RECT 1332.720 22.820 1332.980 23.080 ;
      LAYER met2 ;
        RECT 1332.750 35.000 1333.030 39.000 ;
        RECT 1332.780 23.110 1332.920 35.000 ;
        RECT 377.300 22.790 377.560 23.110 ;
        RECT 1332.720 22.790 1332.980 23.110 ;
        RECT 377.360 2.400 377.500 22.790 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 395.210 16.560 395.530 16.620 ;
        RECT 1383.290 16.560 1383.610 16.620 ;
        RECT 395.210 16.420 1383.610 16.560 ;
        RECT 395.210 16.360 395.530 16.420 ;
        RECT 1383.290 16.360 1383.610 16.420 ;
      LAYER via ;
        RECT 395.240 16.360 395.500 16.620 ;
        RECT 1383.320 16.360 1383.580 16.620 ;
      LAYER met2 ;
        RECT 1383.350 35.000 1383.630 39.000 ;
        RECT 1383.380 16.650 1383.520 35.000 ;
        RECT 395.240 16.330 395.500 16.650 ;
        RECT 1383.320 16.330 1383.580 16.650 ;
        RECT 395.300 2.400 395.440 16.330 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 413.150 23.360 413.470 23.420 ;
        RECT 1434.350 23.360 1434.670 23.420 ;
        RECT 413.150 23.220 1434.670 23.360 ;
        RECT 413.150 23.160 413.470 23.220 ;
        RECT 1434.350 23.160 1434.670 23.220 ;
      LAYER via ;
        RECT 413.180 23.160 413.440 23.420 ;
        RECT 1434.380 23.160 1434.640 23.420 ;
      LAYER met2 ;
        RECT 1434.410 35.000 1434.690 39.000 ;
        RECT 1434.440 23.450 1434.580 35.000 ;
        RECT 413.180 23.130 413.440 23.450 ;
        RECT 1434.380 23.130 1434.640 23.450 ;
        RECT 413.240 2.400 413.380 23.130 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 74.130 19.280 74.450 19.340 ;
        RECT 518.030 19.280 518.350 19.340 ;
        RECT 74.130 19.140 518.350 19.280 ;
        RECT 74.130 19.080 74.450 19.140 ;
        RECT 518.030 19.080 518.350 19.140 ;
      LAYER via ;
        RECT 74.160 19.080 74.420 19.340 ;
        RECT 518.060 19.080 518.320 19.340 ;
      LAYER met2 ;
        RECT 518.090 35.000 518.370 39.000 ;
        RECT 518.120 19.370 518.260 35.000 ;
        RECT 74.160 19.050 74.420 19.370 ;
        RECT 518.060 19.050 518.320 19.370 ;
        RECT 74.220 2.400 74.360 19.050 ;
        RECT 74.010 -4.800 74.570 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 430.630 16.900 430.950 16.960 ;
        RECT 1485.410 16.900 1485.730 16.960 ;
        RECT 430.630 16.760 1485.730 16.900 ;
        RECT 430.630 16.700 430.950 16.760 ;
        RECT 1485.410 16.700 1485.730 16.760 ;
      LAYER via ;
        RECT 430.660 16.700 430.920 16.960 ;
        RECT 1485.440 16.700 1485.700 16.960 ;
      LAYER met2 ;
        RECT 1485.470 35.000 1485.750 39.000 ;
        RECT 1485.500 16.990 1485.640 35.000 ;
        RECT 430.660 16.670 430.920 16.990 ;
        RECT 1485.440 16.670 1485.700 16.990 ;
        RECT 430.720 2.400 430.860 16.670 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 448.570 23.700 448.890 23.760 ;
        RECT 1536.010 23.700 1536.330 23.760 ;
        RECT 448.570 23.560 1536.330 23.700 ;
        RECT 448.570 23.500 448.890 23.560 ;
        RECT 1536.010 23.500 1536.330 23.560 ;
      LAYER via ;
        RECT 448.600 23.500 448.860 23.760 ;
        RECT 1536.040 23.500 1536.300 23.760 ;
      LAYER met2 ;
        RECT 1536.070 35.000 1536.350 39.000 ;
        RECT 1536.100 23.790 1536.240 35.000 ;
        RECT 448.600 23.470 448.860 23.790 ;
        RECT 1536.040 23.470 1536.300 23.790 ;
        RECT 448.660 2.400 448.800 23.470 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 466.510 20.640 466.830 20.700 ;
        RECT 1587.070 20.640 1587.390 20.700 ;
        RECT 466.510 20.500 1587.390 20.640 ;
        RECT 466.510 20.440 466.830 20.500 ;
        RECT 1587.070 20.440 1587.390 20.500 ;
      LAYER via ;
        RECT 466.540 20.440 466.800 20.700 ;
        RECT 1587.100 20.440 1587.360 20.700 ;
      LAYER met2 ;
        RECT 1587.130 35.000 1587.410 39.000 ;
        RECT 1587.160 20.730 1587.300 35.000 ;
        RECT 466.540 20.410 466.800 20.730 ;
        RECT 1587.100 20.410 1587.360 20.730 ;
        RECT 466.600 2.400 466.740 20.410 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 484.450 27.440 484.770 27.500 ;
        RECT 1637.670 27.440 1637.990 27.500 ;
        RECT 484.450 27.300 1637.990 27.440 ;
        RECT 484.450 27.240 484.770 27.300 ;
        RECT 1637.670 27.240 1637.990 27.300 ;
      LAYER via ;
        RECT 484.480 27.240 484.740 27.500 ;
        RECT 1637.700 27.240 1637.960 27.500 ;
      LAYER met2 ;
        RECT 1637.730 35.000 1638.010 39.000 ;
        RECT 1637.760 27.530 1637.900 35.000 ;
        RECT 484.480 27.210 484.740 27.530 ;
        RECT 1637.700 27.210 1637.960 27.530 ;
        RECT 484.540 2.400 484.680 27.210 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 502.390 20.300 502.710 20.360 ;
        RECT 1688.730 20.300 1689.050 20.360 ;
        RECT 502.390 20.160 1689.050 20.300 ;
        RECT 502.390 20.100 502.710 20.160 ;
        RECT 1688.730 20.100 1689.050 20.160 ;
      LAYER via ;
        RECT 502.420 20.100 502.680 20.360 ;
        RECT 1688.760 20.100 1689.020 20.360 ;
      LAYER met2 ;
        RECT 1688.790 35.000 1689.070 39.000 ;
        RECT 1688.820 20.390 1688.960 35.000 ;
        RECT 502.420 20.070 502.680 20.390 ;
        RECT 1688.760 20.070 1689.020 20.390 ;
        RECT 502.480 2.400 502.620 20.070 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 519.870 27.100 520.190 27.160 ;
        RECT 1739.790 27.100 1740.110 27.160 ;
        RECT 519.870 26.960 1740.110 27.100 ;
        RECT 519.870 26.900 520.190 26.960 ;
        RECT 1739.790 26.900 1740.110 26.960 ;
      LAYER via ;
        RECT 519.900 26.900 520.160 27.160 ;
        RECT 1739.820 26.900 1740.080 27.160 ;
      LAYER met2 ;
        RECT 1739.850 35.000 1740.130 39.000 ;
        RECT 1739.880 27.190 1740.020 35.000 ;
        RECT 519.900 26.870 520.160 27.190 ;
        RECT 1739.820 26.870 1740.080 27.190 ;
        RECT 519.960 2.400 520.100 26.870 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 537.810 19.960 538.130 20.020 ;
        RECT 1790.390 19.960 1790.710 20.020 ;
        RECT 537.810 19.820 1790.710 19.960 ;
        RECT 537.810 19.760 538.130 19.820 ;
        RECT 1790.390 19.760 1790.710 19.820 ;
      LAYER via ;
        RECT 537.840 19.760 538.100 20.020 ;
        RECT 1790.420 19.760 1790.680 20.020 ;
      LAYER met2 ;
        RECT 1790.450 35.000 1790.730 39.000 ;
        RECT 1790.480 20.050 1790.620 35.000 ;
        RECT 537.840 19.730 538.100 20.050 ;
        RECT 1790.420 19.730 1790.680 20.050 ;
        RECT 537.900 2.400 538.040 19.730 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 555.750 26.760 556.070 26.820 ;
        RECT 1841.450 26.760 1841.770 26.820 ;
        RECT 555.750 26.620 1841.770 26.760 ;
        RECT 555.750 26.560 556.070 26.620 ;
        RECT 1841.450 26.560 1841.770 26.620 ;
      LAYER via ;
        RECT 555.780 26.560 556.040 26.820 ;
        RECT 1841.480 26.560 1841.740 26.820 ;
      LAYER met2 ;
        RECT 1841.510 35.000 1841.790 39.000 ;
        RECT 1841.540 26.850 1841.680 35.000 ;
        RECT 555.780 26.530 556.040 26.850 ;
        RECT 1841.480 26.530 1841.740 26.850 ;
        RECT 555.840 2.400 555.980 26.530 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 573.690 19.620 574.010 19.680 ;
        RECT 1892.510 19.620 1892.830 19.680 ;
        RECT 573.690 19.480 1892.830 19.620 ;
        RECT 573.690 19.420 574.010 19.480 ;
        RECT 1892.510 19.420 1892.830 19.480 ;
      LAYER via ;
        RECT 573.720 19.420 573.980 19.680 ;
        RECT 1892.540 19.420 1892.800 19.680 ;
      LAYER met2 ;
        RECT 1892.570 35.000 1892.850 39.000 ;
        RECT 1892.600 19.710 1892.740 35.000 ;
        RECT 573.720 19.390 573.980 19.710 ;
        RECT 1892.540 19.390 1892.800 19.710 ;
        RECT 573.780 2.400 573.920 19.390 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 591.170 26.420 591.490 26.480 ;
        RECT 1943.110 26.420 1943.430 26.480 ;
        RECT 591.170 26.280 1943.430 26.420 ;
        RECT 591.170 26.220 591.490 26.280 ;
        RECT 1943.110 26.220 1943.430 26.280 ;
      LAYER via ;
        RECT 591.200 26.220 591.460 26.480 ;
        RECT 1943.140 26.220 1943.400 26.480 ;
      LAYER met2 ;
        RECT 1943.170 35.000 1943.450 39.000 ;
        RECT 1943.200 26.510 1943.340 35.000 ;
        RECT 591.200 26.190 591.460 26.510 ;
        RECT 1943.140 26.190 1943.400 26.510 ;
        RECT 591.260 2.400 591.400 26.190 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 97.590 26.080 97.910 26.140 ;
        RECT 569.090 26.080 569.410 26.140 ;
        RECT 97.590 25.940 569.410 26.080 ;
        RECT 97.590 25.880 97.910 25.940 ;
        RECT 569.090 25.880 569.410 25.940 ;
      LAYER via ;
        RECT 97.620 25.880 97.880 26.140 ;
        RECT 569.120 25.880 569.380 26.140 ;
      LAYER met2 ;
        RECT 569.150 35.000 569.430 39.000 ;
        RECT 569.180 26.170 569.320 35.000 ;
        RECT 97.620 25.850 97.880 26.170 ;
        RECT 569.120 25.850 569.380 26.170 ;
        RECT 97.680 2.400 97.820 25.850 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 609.110 19.280 609.430 19.340 ;
        RECT 1994.170 19.280 1994.490 19.340 ;
        RECT 609.110 19.140 1994.490 19.280 ;
        RECT 609.110 19.080 609.430 19.140 ;
        RECT 1994.170 19.080 1994.490 19.140 ;
      LAYER via ;
        RECT 609.140 19.080 609.400 19.340 ;
        RECT 1994.200 19.080 1994.460 19.340 ;
      LAYER met2 ;
        RECT 1994.230 35.000 1994.510 39.000 ;
        RECT 1994.260 19.370 1994.400 35.000 ;
        RECT 609.140 19.050 609.400 19.370 ;
        RECT 1994.200 19.050 1994.460 19.370 ;
        RECT 609.200 2.400 609.340 19.050 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 627.050 26.080 627.370 26.140 ;
        RECT 2045.230 26.080 2045.550 26.140 ;
        RECT 627.050 25.940 2045.550 26.080 ;
        RECT 627.050 25.880 627.370 25.940 ;
        RECT 2045.230 25.880 2045.550 25.940 ;
      LAYER via ;
        RECT 627.080 25.880 627.340 26.140 ;
        RECT 2045.260 25.880 2045.520 26.140 ;
      LAYER met2 ;
        RECT 2045.290 35.000 2045.570 39.000 ;
        RECT 2045.320 26.170 2045.460 35.000 ;
        RECT 627.080 25.850 627.340 26.170 ;
        RECT 2045.260 25.850 2045.520 26.170 ;
        RECT 627.140 2.400 627.280 25.850 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 17.580 121.830 17.640 ;
        RECT 620.150 17.580 620.470 17.640 ;
        RECT 121.510 17.440 620.470 17.580 ;
        RECT 121.510 17.380 121.830 17.440 ;
        RECT 620.150 17.380 620.470 17.440 ;
      LAYER via ;
        RECT 121.540 17.380 121.800 17.640 ;
        RECT 620.180 17.380 620.440 17.640 ;
      LAYER met2 ;
        RECT 620.210 35.000 620.490 39.000 ;
        RECT 620.240 17.670 620.380 35.000 ;
        RECT 121.540 17.350 121.800 17.670 ;
        RECT 620.180 17.350 620.440 17.670 ;
        RECT 121.600 2.400 121.740 17.350 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 145.430 14.180 145.750 14.240 ;
        RECT 670.750 14.180 671.070 14.240 ;
        RECT 145.430 14.040 671.070 14.180 ;
        RECT 145.430 13.980 145.750 14.040 ;
        RECT 670.750 13.980 671.070 14.040 ;
      LAYER via ;
        RECT 145.460 13.980 145.720 14.240 ;
        RECT 670.780 13.980 671.040 14.240 ;
      LAYER met2 ;
        RECT 670.810 35.000 671.090 39.000 ;
        RECT 670.840 14.270 670.980 35.000 ;
        RECT 145.460 13.950 145.720 14.270 ;
        RECT 670.780 13.950 671.040 14.270 ;
        RECT 145.520 2.400 145.660 13.950 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 163.370 14.520 163.690 14.580 ;
        RECT 721.810 14.520 722.130 14.580 ;
        RECT 163.370 14.380 722.130 14.520 ;
        RECT 163.370 14.320 163.690 14.380 ;
        RECT 721.810 14.320 722.130 14.380 ;
      LAYER via ;
        RECT 163.400 14.320 163.660 14.580 ;
        RECT 721.840 14.320 722.100 14.580 ;
      LAYER met2 ;
        RECT 721.870 35.000 722.150 39.000 ;
        RECT 721.900 14.610 722.040 35.000 ;
        RECT 163.400 14.290 163.660 14.610 ;
        RECT 721.840 14.290 722.100 14.610 ;
        RECT 163.460 2.400 163.600 14.290 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 180.850 20.980 181.170 21.040 ;
        RECT 772.870 20.980 773.190 21.040 ;
        RECT 180.850 20.840 773.190 20.980 ;
        RECT 180.850 20.780 181.170 20.840 ;
        RECT 772.870 20.780 773.190 20.840 ;
      LAYER via ;
        RECT 180.880 20.780 181.140 21.040 ;
        RECT 772.900 20.780 773.160 21.040 ;
      LAYER met2 ;
        RECT 772.930 35.000 773.210 39.000 ;
        RECT 772.960 21.070 773.100 35.000 ;
        RECT 180.880 20.750 181.140 21.070 ;
        RECT 772.900 20.750 773.160 21.070 ;
        RECT 180.940 2.400 181.080 20.750 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 198.790 14.860 199.110 14.920 ;
        RECT 823.470 14.860 823.790 14.920 ;
        RECT 198.790 14.720 823.790 14.860 ;
        RECT 198.790 14.660 199.110 14.720 ;
        RECT 823.470 14.660 823.790 14.720 ;
      LAYER via ;
        RECT 198.820 14.660 199.080 14.920 ;
        RECT 823.500 14.660 823.760 14.920 ;
      LAYER met2 ;
        RECT 823.530 35.000 823.810 39.000 ;
        RECT 823.560 14.950 823.700 35.000 ;
        RECT 198.820 14.630 199.080 14.950 ;
        RECT 823.500 14.630 823.760 14.950 ;
        RECT 198.880 2.400 199.020 14.630 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 216.730 21.320 217.050 21.380 ;
        RECT 874.530 21.320 874.850 21.380 ;
        RECT 216.730 21.180 874.850 21.320 ;
        RECT 216.730 21.120 217.050 21.180 ;
        RECT 874.530 21.120 874.850 21.180 ;
      LAYER via ;
        RECT 216.760 21.120 217.020 21.380 ;
        RECT 874.560 21.120 874.820 21.380 ;
      LAYER met2 ;
        RECT 874.590 35.000 874.870 39.000 ;
        RECT 874.620 21.410 874.760 35.000 ;
        RECT 216.760 21.090 217.020 21.410 ;
        RECT 874.560 21.090 874.820 21.410 ;
        RECT 216.820 2.400 216.960 21.090 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 234.670 15.880 234.990 15.940 ;
        RECT 234.670 15.740 247.320 15.880 ;
        RECT 234.670 15.680 234.990 15.740 ;
        RECT 247.180 15.200 247.320 15.740 ;
        RECT 925.130 15.200 925.450 15.260 ;
        RECT 247.180 15.060 925.450 15.200 ;
        RECT 925.130 15.000 925.450 15.060 ;
      LAYER via ;
        RECT 234.700 15.680 234.960 15.940 ;
        RECT 925.160 15.000 925.420 15.260 ;
      LAYER met2 ;
        RECT 925.190 35.000 925.470 39.000 ;
        RECT 234.700 15.650 234.960 15.970 ;
        RECT 234.760 2.400 234.900 15.650 ;
        RECT 925.220 15.290 925.360 35.000 ;
        RECT 925.160 14.970 925.420 15.290 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2880.205 3173.985 2880.375 3239.095 ;
        RECT 2880.205 2987.665 2880.375 3011.975 ;
        RECT 2879.745 2773.805 2879.915 2821.915 ;
        RECT 2880.205 2428.025 2880.375 2439.075 ;
        RECT 2880.205 1897.965 2880.375 1921.935 ;
        RECT 2880.205 1832.345 2880.375 1859.715 ;
        RECT 2880.205 1794.945 2880.375 1797.495 ;
        RECT 2879.745 1737.145 2879.915 1763.495 ;
        RECT 2880.205 1580.235 2880.375 1596.215 ;
        RECT 2879.745 1580.065 2880.375 1580.235 ;
        RECT 2879.745 1578.705 2879.915 1580.065 ;
        RECT 2880.665 824.585 2880.835 878.475 ;
        RECT 2880.205 701.505 2880.375 726.495 ;
        RECT 2880.665 554.625 2880.835 579.275 ;
        RECT 2880.205 141.525 2880.375 165.495 ;
      LAYER mcon ;
        RECT 2880.205 3238.925 2880.375 3239.095 ;
        RECT 2880.205 3011.805 2880.375 3011.975 ;
        RECT 2879.745 2821.745 2879.915 2821.915 ;
        RECT 2880.205 2438.905 2880.375 2439.075 ;
        RECT 2880.205 1921.765 2880.375 1921.935 ;
        RECT 2880.205 1859.545 2880.375 1859.715 ;
        RECT 2880.205 1797.325 2880.375 1797.495 ;
        RECT 2879.745 1763.325 2879.915 1763.495 ;
        RECT 2880.205 1596.045 2880.375 1596.215 ;
        RECT 2880.665 878.305 2880.835 878.475 ;
        RECT 2880.205 726.325 2880.375 726.495 ;
        RECT 2880.665 579.105 2880.835 579.275 ;
        RECT 2880.205 165.325 2880.375 165.495 ;
      LAYER met1 ;
        RECT 2879.670 3264.580 2879.990 3264.640 ;
        RECT 2881.510 3264.580 2881.830 3264.640 ;
        RECT 2879.670 3264.440 2881.830 3264.580 ;
        RECT 2879.670 3264.380 2879.990 3264.440 ;
        RECT 2881.510 3264.380 2881.830 3264.440 ;
        RECT 2879.670 3239.080 2879.990 3239.140 ;
        RECT 2880.145 3239.080 2880.435 3239.125 ;
        RECT 2879.670 3238.940 2880.435 3239.080 ;
        RECT 2879.670 3238.880 2879.990 3238.940 ;
        RECT 2880.145 3238.895 2880.435 3238.940 ;
        RECT 2880.130 3174.140 2880.450 3174.200 ;
        RECT 2879.935 3174.000 2880.450 3174.140 ;
        RECT 2880.130 3173.940 2880.450 3174.000 ;
        RECT 2879.670 3011.960 2879.990 3012.020 ;
        RECT 2880.145 3011.960 2880.435 3012.005 ;
        RECT 2879.670 3011.820 2880.435 3011.960 ;
        RECT 2879.670 3011.760 2879.990 3011.820 ;
        RECT 2880.145 3011.775 2880.435 3011.820 ;
        RECT 2880.130 2987.820 2880.450 2987.880 ;
        RECT 2879.935 2987.680 2880.450 2987.820 ;
        RECT 2880.130 2987.620 2880.450 2987.680 ;
        RECT 2879.670 2835.980 2879.990 2836.240 ;
        RECT 2879.760 2835.560 2879.900 2835.980 ;
        RECT 2879.670 2835.300 2879.990 2835.560 ;
        RECT 2879.670 2821.900 2879.990 2821.960 ;
        RECT 2879.475 2821.760 2879.990 2821.900 ;
        RECT 2879.670 2821.700 2879.990 2821.760 ;
        RECT 2879.685 2773.960 2879.975 2774.005 ;
        RECT 2880.130 2773.960 2880.450 2774.020 ;
        RECT 2879.685 2773.820 2880.450 2773.960 ;
        RECT 2879.685 2773.775 2879.975 2773.820 ;
        RECT 2880.130 2773.760 2880.450 2773.820 ;
        RECT 2879.670 2684.200 2879.990 2684.260 ;
        RECT 2880.130 2684.200 2880.450 2684.260 ;
        RECT 2879.670 2684.060 2880.450 2684.200 ;
        RECT 2879.670 2684.000 2879.990 2684.060 ;
        RECT 2880.130 2684.000 2880.450 2684.060 ;
        RECT 2880.130 2573.700 2880.450 2573.760 ;
        RECT 2881.050 2573.700 2881.370 2573.760 ;
        RECT 2880.130 2573.560 2881.370 2573.700 ;
        RECT 2880.130 2573.500 2880.450 2573.560 ;
        RECT 2881.050 2573.500 2881.370 2573.560 ;
        RECT 2879.670 2526.780 2879.990 2526.840 ;
        RECT 2881.050 2526.780 2881.370 2526.840 ;
        RECT 2879.670 2526.640 2881.370 2526.780 ;
        RECT 2879.670 2526.580 2879.990 2526.640 ;
        RECT 2881.050 2526.580 2881.370 2526.640 ;
        RECT 2879.670 2439.060 2879.990 2439.120 ;
        RECT 2880.145 2439.060 2880.435 2439.105 ;
        RECT 2879.670 2438.920 2880.435 2439.060 ;
        RECT 2879.670 2438.860 2879.990 2438.920 ;
        RECT 2880.145 2438.875 2880.435 2438.920 ;
        RECT 2879.670 2428.180 2879.990 2428.240 ;
        RECT 2880.145 2428.180 2880.435 2428.225 ;
        RECT 2879.670 2428.040 2880.435 2428.180 ;
        RECT 2879.670 2427.980 2879.990 2428.040 ;
        RECT 2880.145 2427.995 2880.435 2428.040 ;
        RECT 2879.670 1921.920 2879.990 1921.980 ;
        RECT 2880.145 1921.920 2880.435 1921.965 ;
        RECT 2879.670 1921.780 2880.435 1921.920 ;
        RECT 2879.670 1921.720 2879.990 1921.780 ;
        RECT 2880.145 1921.735 2880.435 1921.780 ;
        RECT 2880.145 1898.120 2880.435 1898.165 ;
        RECT 2879.760 1897.980 2880.435 1898.120 ;
        RECT 2879.760 1897.440 2879.900 1897.980 ;
        RECT 2880.145 1897.935 2880.435 1897.980 ;
        RECT 2880.130 1897.440 2880.450 1897.500 ;
        RECT 2879.760 1897.300 2880.450 1897.440 ;
        RECT 2880.130 1897.240 2880.450 1897.300 ;
        RECT 2880.130 1859.700 2880.450 1859.760 ;
        RECT 2879.935 1859.560 2880.450 1859.700 ;
        RECT 2880.130 1859.500 2880.450 1859.560 ;
        RECT 2879.670 1832.500 2879.990 1832.560 ;
        RECT 2880.145 1832.500 2880.435 1832.545 ;
        RECT 2879.670 1832.360 2880.435 1832.500 ;
        RECT 2879.670 1832.300 2879.990 1832.360 ;
        RECT 2880.145 1832.315 2880.435 1832.360 ;
        RECT 2879.670 1797.480 2879.990 1797.540 ;
        RECT 2880.145 1797.480 2880.435 1797.525 ;
        RECT 2879.670 1797.340 2880.435 1797.480 ;
        RECT 2879.670 1797.280 2879.990 1797.340 ;
        RECT 2880.145 1797.295 2880.435 1797.340 ;
        RECT 2879.670 1795.100 2879.990 1795.160 ;
        RECT 2880.145 1795.100 2880.435 1795.145 ;
        RECT 2879.670 1794.960 2880.435 1795.100 ;
        RECT 2879.670 1794.900 2879.990 1794.960 ;
        RECT 2880.145 1794.915 2880.435 1794.960 ;
        RECT 2879.670 1763.480 2879.990 1763.540 ;
        RECT 2879.475 1763.340 2879.990 1763.480 ;
        RECT 2879.670 1763.280 2879.990 1763.340 ;
        RECT 2879.670 1737.300 2879.990 1737.360 ;
        RECT 2879.475 1737.160 2879.990 1737.300 ;
        RECT 2879.670 1737.100 2879.990 1737.160 ;
        RECT 2879.670 1596.200 2879.990 1596.260 ;
        RECT 2880.145 1596.200 2880.435 1596.245 ;
        RECT 2879.670 1596.060 2880.435 1596.200 ;
        RECT 2879.670 1596.000 2879.990 1596.060 ;
        RECT 2880.145 1596.015 2880.435 1596.060 ;
        RECT 2879.670 1578.860 2879.990 1578.920 ;
        RECT 2879.475 1578.720 2879.990 1578.860 ;
        RECT 2879.670 1578.660 2879.990 1578.720 ;
        RECT 2879.670 1432.120 2879.990 1432.380 ;
        RECT 2879.760 1431.360 2879.900 1432.120 ;
        RECT 2879.670 1431.100 2879.990 1431.360 ;
        RECT 2879.670 1394.580 2879.990 1394.640 ;
        RECT 2880.590 1394.580 2880.910 1394.640 ;
        RECT 2879.670 1394.440 2880.910 1394.580 ;
        RECT 2879.670 1394.380 2879.990 1394.440 ;
        RECT 2880.590 1394.380 2880.910 1394.440 ;
        RECT 2879.670 878.460 2879.990 878.520 ;
        RECT 2880.605 878.460 2880.895 878.505 ;
        RECT 2879.670 878.320 2880.895 878.460 ;
        RECT 2879.670 878.260 2879.990 878.320 ;
        RECT 2880.605 878.275 2880.895 878.320 ;
        RECT 2879.670 824.740 2879.990 824.800 ;
        RECT 2880.605 824.740 2880.895 824.785 ;
        RECT 2879.670 824.600 2880.895 824.740 ;
        RECT 2879.670 824.540 2879.990 824.600 ;
        RECT 2880.605 824.555 2880.895 824.600 ;
        RECT 2879.670 726.480 2879.990 726.540 ;
        RECT 2880.145 726.480 2880.435 726.525 ;
        RECT 2879.670 726.340 2880.435 726.480 ;
        RECT 2879.670 726.280 2879.990 726.340 ;
        RECT 2880.145 726.295 2880.435 726.340 ;
        RECT 2879.670 701.660 2879.990 701.720 ;
        RECT 2880.145 701.660 2880.435 701.705 ;
        RECT 2879.670 701.520 2880.435 701.660 ;
        RECT 2879.670 701.460 2879.990 701.520 ;
        RECT 2880.145 701.475 2880.435 701.520 ;
        RECT 2880.130 579.400 2880.450 579.660 ;
        RECT 2880.220 579.260 2880.360 579.400 ;
        RECT 2880.605 579.260 2880.895 579.305 ;
        RECT 2880.220 579.120 2880.895 579.260 ;
        RECT 2880.605 579.075 2880.895 579.120 ;
        RECT 2879.670 554.780 2879.990 554.840 ;
        RECT 2880.605 554.780 2880.895 554.825 ;
        RECT 2879.670 554.640 2880.895 554.780 ;
        RECT 2879.670 554.580 2879.990 554.640 ;
        RECT 2880.605 554.595 2880.895 554.640 ;
        RECT 2879.670 231.920 2879.990 232.180 ;
        RECT 2879.760 231.100 2879.900 231.920 ;
        RECT 2880.130 231.100 2880.450 231.160 ;
        RECT 2879.760 230.960 2880.450 231.100 ;
        RECT 2880.130 230.900 2880.450 230.960 ;
        RECT 2879.670 165.480 2879.990 165.540 ;
        RECT 2880.145 165.480 2880.435 165.525 ;
        RECT 2879.670 165.340 2880.435 165.480 ;
        RECT 2879.670 165.280 2879.990 165.340 ;
        RECT 2880.145 165.295 2880.435 165.340 ;
        RECT 2879.670 141.680 2879.990 141.740 ;
        RECT 2880.145 141.680 2880.435 141.725 ;
        RECT 2879.670 141.540 2880.435 141.680 ;
        RECT 2879.670 141.480 2879.990 141.540 ;
        RECT 2880.145 141.495 2880.435 141.540 ;
        RECT 2875.530 37.640 2875.850 37.700 ;
        RECT 2879.670 37.640 2879.990 37.700 ;
        RECT 2875.530 37.500 2879.990 37.640 ;
        RECT 2875.530 37.440 2875.850 37.500 ;
        RECT 2879.670 37.440 2879.990 37.500 ;
      LAYER via ;
        RECT 2879.700 3264.380 2879.960 3264.640 ;
        RECT 2881.540 3264.380 2881.800 3264.640 ;
        RECT 2879.700 3238.880 2879.960 3239.140 ;
        RECT 2880.160 3173.940 2880.420 3174.200 ;
        RECT 2879.700 3011.760 2879.960 3012.020 ;
        RECT 2880.160 2987.620 2880.420 2987.880 ;
        RECT 2879.700 2835.980 2879.960 2836.240 ;
        RECT 2879.700 2835.300 2879.960 2835.560 ;
        RECT 2879.700 2821.700 2879.960 2821.960 ;
        RECT 2880.160 2773.760 2880.420 2774.020 ;
        RECT 2879.700 2684.000 2879.960 2684.260 ;
        RECT 2880.160 2684.000 2880.420 2684.260 ;
        RECT 2880.160 2573.500 2880.420 2573.760 ;
        RECT 2881.080 2573.500 2881.340 2573.760 ;
        RECT 2879.700 2526.580 2879.960 2526.840 ;
        RECT 2881.080 2526.580 2881.340 2526.840 ;
        RECT 2879.700 2438.860 2879.960 2439.120 ;
        RECT 2879.700 2427.980 2879.960 2428.240 ;
        RECT 2879.700 1921.720 2879.960 1921.980 ;
        RECT 2880.160 1897.240 2880.420 1897.500 ;
        RECT 2880.160 1859.500 2880.420 1859.760 ;
        RECT 2879.700 1832.300 2879.960 1832.560 ;
        RECT 2879.700 1797.280 2879.960 1797.540 ;
        RECT 2879.700 1794.900 2879.960 1795.160 ;
        RECT 2879.700 1763.280 2879.960 1763.540 ;
        RECT 2879.700 1737.100 2879.960 1737.360 ;
        RECT 2879.700 1596.000 2879.960 1596.260 ;
        RECT 2879.700 1578.660 2879.960 1578.920 ;
        RECT 2879.700 1432.120 2879.960 1432.380 ;
        RECT 2879.700 1431.100 2879.960 1431.360 ;
        RECT 2879.700 1394.380 2879.960 1394.640 ;
        RECT 2880.620 1394.380 2880.880 1394.640 ;
        RECT 2879.700 878.260 2879.960 878.520 ;
        RECT 2879.700 824.540 2879.960 824.800 ;
        RECT 2879.700 726.280 2879.960 726.540 ;
        RECT 2879.700 701.460 2879.960 701.720 ;
        RECT 2880.160 579.400 2880.420 579.660 ;
        RECT 2879.700 554.580 2879.960 554.840 ;
        RECT 2879.700 231.920 2879.960 232.180 ;
        RECT 2880.160 230.900 2880.420 231.160 ;
        RECT 2879.700 165.280 2879.960 165.540 ;
        RECT 2879.700 141.480 2879.960 141.740 ;
        RECT 2875.560 37.440 2875.820 37.700 ;
        RECT 2879.700 37.440 2879.960 37.700 ;
      LAYER met2 ;
        RECT 2881.530 3266.875 2881.810 3267.245 ;
        RECT 2881.600 3264.670 2881.740 3266.875 ;
        RECT 2879.700 3264.580 2879.960 3264.670 ;
        RECT 2879.300 3264.440 2879.960 3264.580 ;
        RECT 2879.300 3239.250 2879.440 3264.440 ;
        RECT 2879.700 3264.350 2879.960 3264.440 ;
        RECT 2881.540 3264.350 2881.800 3264.670 ;
        RECT 2879.300 3239.170 2879.900 3239.250 ;
        RECT 2879.300 3239.110 2879.960 3239.170 ;
        RECT 2879.700 3238.850 2879.960 3239.110 ;
        RECT 2880.160 3173.910 2880.420 3174.230 ;
        RECT 2880.220 3152.890 2880.360 3173.910 ;
        RECT 2879.760 3152.750 2880.360 3152.890 ;
        RECT 2879.760 3108.690 2879.900 3152.750 ;
        RECT 2879.300 3108.550 2879.900 3108.690 ;
        RECT 2879.300 3042.730 2879.440 3108.550 ;
        RECT 2878.840 3042.590 2879.440 3042.730 ;
        RECT 2878.840 3035.930 2878.980 3042.590 ;
        RECT 2878.840 3035.790 2879.440 3035.930 ;
        RECT 2879.300 3034.570 2879.440 3035.790 ;
        RECT 2879.300 3034.430 2879.900 3034.570 ;
        RECT 2879.760 3012.050 2879.900 3034.430 ;
        RECT 2879.700 3011.730 2879.960 3012.050 ;
        RECT 2880.160 2987.590 2880.420 2987.910 ;
        RECT 2880.220 2884.970 2880.360 2987.590 ;
        RECT 2879.760 2884.830 2880.360 2884.970 ;
        RECT 2879.760 2836.270 2879.900 2884.830 ;
        RECT 2879.700 2835.950 2879.960 2836.270 ;
        RECT 2879.700 2835.270 2879.960 2835.590 ;
        RECT 2879.760 2821.990 2879.900 2835.270 ;
        RECT 2879.700 2821.670 2879.960 2821.990 ;
        RECT 2880.160 2773.730 2880.420 2774.050 ;
        RECT 2880.220 2755.770 2880.360 2773.730 ;
        RECT 2879.760 2755.630 2880.360 2755.770 ;
        RECT 2879.760 2731.970 2879.900 2755.630 ;
        RECT 2879.760 2731.830 2880.360 2731.970 ;
        RECT 2880.220 2684.290 2880.360 2731.830 ;
        RECT 2879.700 2683.970 2879.960 2684.290 ;
        RECT 2880.160 2683.970 2880.420 2684.290 ;
        RECT 2879.760 2642.890 2879.900 2683.970 ;
        RECT 2879.760 2642.750 2880.360 2642.890 ;
        RECT 2880.220 2573.790 2880.360 2642.750 ;
        RECT 2880.160 2573.470 2880.420 2573.790 ;
        RECT 2881.080 2573.470 2881.340 2573.790 ;
        RECT 2881.140 2526.870 2881.280 2573.470 ;
        RECT 2879.700 2526.780 2879.960 2526.870 ;
        RECT 2879.300 2526.640 2879.960 2526.780 ;
        RECT 2879.300 2517.090 2879.440 2526.640 ;
        RECT 2879.700 2526.550 2879.960 2526.640 ;
        RECT 2881.080 2526.550 2881.340 2526.870 ;
        RECT 2877.920 2516.950 2879.440 2517.090 ;
        RECT 2877.920 2476.290 2878.060 2516.950 ;
        RECT 2877.920 2476.150 2879.900 2476.290 ;
        RECT 2879.760 2439.150 2879.900 2476.150 ;
        RECT 2879.700 2438.830 2879.960 2439.150 ;
        RECT 2879.700 2428.010 2879.960 2428.270 ;
        RECT 2878.840 2427.950 2879.960 2428.010 ;
        RECT 2878.840 2427.870 2879.900 2427.950 ;
        RECT 2878.840 2415.090 2878.980 2427.870 ;
        RECT 2877.920 2414.950 2878.980 2415.090 ;
        RECT 2877.920 2379.730 2878.060 2414.950 ;
        RECT 2877.920 2379.590 2878.520 2379.730 ;
        RECT 2878.380 2283.850 2878.520 2379.590 ;
        RECT 2876.080 2283.710 2878.520 2283.850 ;
        RECT 2876.080 2222.650 2876.220 2283.710 ;
        RECT 2876.080 2222.510 2877.140 2222.650 ;
        RECT 2877.000 2221.970 2877.140 2222.510 ;
        RECT 2877.000 2221.830 2878.060 2221.970 ;
        RECT 2877.920 2197.490 2878.060 2221.830 ;
        RECT 2877.920 2197.350 2878.980 2197.490 ;
        RECT 2878.840 2186.610 2878.980 2197.350 ;
        RECT 2878.380 2186.470 2878.980 2186.610 ;
        RECT 2878.380 2141.730 2878.520 2186.470 ;
        RECT 2877.460 2141.590 2878.520 2141.730 ;
        RECT 2877.460 2136.970 2877.600 2141.590 ;
        RECT 2877.460 2136.830 2878.060 2136.970 ;
        RECT 2877.920 2077.130 2878.060 2136.830 ;
        RECT 2877.920 2076.990 2878.520 2077.130 ;
        RECT 2878.380 2045.850 2878.520 2076.990 ;
        RECT 2877.000 2045.710 2878.520 2045.850 ;
        RECT 2877.000 1980.570 2877.140 2045.710 ;
        RECT 2877.000 1980.430 2877.600 1980.570 ;
        RECT 2877.460 1950.650 2877.600 1980.430 ;
        RECT 2877.460 1950.510 2878.520 1950.650 ;
        RECT 2878.380 1946.570 2878.520 1950.510 ;
        RECT 2877.920 1946.430 2878.520 1946.570 ;
        RECT 2877.920 1943.170 2878.060 1946.430 ;
        RECT 2877.920 1943.030 2878.520 1943.170 ;
        RECT 2878.380 1942.490 2878.520 1943.030 ;
        RECT 2878.380 1942.350 2879.900 1942.490 ;
        RECT 2879.760 1922.010 2879.900 1942.350 ;
        RECT 2879.700 1921.690 2879.960 1922.010 ;
        RECT 2880.160 1897.210 2880.420 1897.530 ;
        RECT 2880.220 1859.790 2880.360 1897.210 ;
        RECT 2880.160 1859.470 2880.420 1859.790 ;
        RECT 2879.700 1832.330 2879.960 1832.590 ;
        RECT 2879.300 1832.270 2879.960 1832.330 ;
        RECT 2879.300 1832.190 2879.900 1832.270 ;
        RECT 2879.300 1805.130 2879.440 1832.190 ;
        RECT 2879.300 1804.990 2879.900 1805.130 ;
        RECT 2879.760 1797.570 2879.900 1804.990 ;
        RECT 2879.700 1797.250 2879.960 1797.570 ;
        RECT 2879.700 1794.870 2879.960 1795.190 ;
        RECT 2879.760 1794.250 2879.900 1794.870 ;
        RECT 2879.300 1794.110 2879.900 1794.250 ;
        RECT 2879.300 1763.650 2879.440 1794.110 ;
        RECT 2879.300 1763.570 2879.900 1763.650 ;
        RECT 2879.300 1763.510 2879.960 1763.570 ;
        RECT 2879.700 1763.250 2879.960 1763.510 ;
        RECT 2879.700 1737.130 2879.960 1737.390 ;
        RECT 2877.920 1737.070 2879.960 1737.130 ;
        RECT 2877.920 1736.990 2879.900 1737.070 ;
        RECT 2877.920 1663.690 2878.060 1736.990 ;
        RECT 2876.540 1663.550 2878.060 1663.690 ;
        RECT 2876.540 1637.850 2876.680 1663.550 ;
        RECT 2876.540 1637.710 2878.060 1637.850 ;
        RECT 2877.920 1597.050 2878.060 1637.710 ;
        RECT 2877.920 1596.910 2879.900 1597.050 ;
        RECT 2879.760 1596.290 2879.900 1596.910 ;
        RECT 2879.700 1595.970 2879.960 1596.290 ;
        RECT 2879.700 1578.690 2879.960 1578.950 ;
        RECT 2877.920 1578.630 2879.960 1578.690 ;
        RECT 2877.920 1578.550 2879.900 1578.630 ;
        RECT 2877.920 1462.410 2878.060 1578.550 ;
        RECT 2877.460 1462.270 2878.060 1462.410 ;
        RECT 2877.460 1442.010 2877.600 1462.270 ;
        RECT 2877.460 1441.870 2879.900 1442.010 ;
        RECT 2879.760 1432.410 2879.900 1441.870 ;
        RECT 2879.700 1432.090 2879.960 1432.410 ;
        RECT 2879.700 1431.070 2879.960 1431.390 ;
        RECT 2879.760 1394.670 2879.900 1431.070 ;
        RECT 2879.700 1394.350 2879.960 1394.670 ;
        RECT 2880.620 1394.350 2880.880 1394.670 ;
        RECT 2878.380 1265.750 2880.360 1265.890 ;
        RECT 2878.380 1245.660 2878.520 1265.750 ;
        RECT 2880.220 1265.210 2880.360 1265.750 ;
        RECT 2880.680 1265.210 2880.820 1394.350 ;
        RECT 2880.220 1265.070 2880.820 1265.210 ;
        RECT 2877.000 1245.520 2878.520 1245.660 ;
        RECT 2877.000 1233.250 2877.140 1245.520 ;
        RECT 2876.540 1233.110 2877.140 1233.250 ;
        RECT 2876.540 1148.930 2876.680 1233.110 ;
        RECT 2876.540 1148.790 2878.060 1148.930 ;
        RECT 2877.920 1088.410 2878.060 1148.790 ;
        RECT 2875.160 1088.270 2878.060 1088.410 ;
        RECT 2875.160 1011.570 2875.300 1088.270 ;
        RECT 2875.160 1011.430 2876.680 1011.570 ;
        RECT 2876.540 976.890 2876.680 1011.430 ;
        RECT 2874.240 976.750 2876.680 976.890 ;
        RECT 2874.240 882.370 2874.380 976.750 ;
        RECT 2874.240 882.230 2878.980 882.370 ;
        RECT 2878.840 878.460 2878.980 882.230 ;
        RECT 2879.700 878.460 2879.960 878.550 ;
        RECT 2878.840 878.320 2879.960 878.460 ;
        RECT 2879.700 878.230 2879.960 878.320 ;
        RECT 2879.700 824.740 2879.960 824.830 ;
        RECT 2878.840 824.600 2879.960 824.740 ;
        RECT 2878.840 817.770 2878.980 824.600 ;
        RECT 2879.700 824.510 2879.960 824.600 ;
        RECT 2877.000 817.630 2878.980 817.770 ;
        RECT 2877.000 726.480 2877.140 817.630 ;
        RECT 2879.700 726.480 2879.960 726.570 ;
        RECT 2877.000 726.340 2879.960 726.480 ;
        RECT 2879.700 726.250 2879.960 726.340 ;
        RECT 2879.700 701.660 2879.960 701.750 ;
        RECT 2877.920 701.520 2879.960 701.660 ;
        RECT 2877.920 644.370 2878.060 701.520 ;
        RECT 2879.700 701.430 2879.960 701.520 ;
        RECT 2877.000 644.230 2878.060 644.370 ;
        RECT 2877.000 640.460 2877.140 644.230 ;
        RECT 2877.000 640.320 2878.060 640.460 ;
        RECT 2877.920 624.650 2878.060 640.320 ;
        RECT 2877.920 624.510 2880.360 624.650 ;
        RECT 2880.220 579.690 2880.360 624.510 ;
        RECT 2880.160 579.370 2880.420 579.690 ;
        RECT 2879.700 554.550 2879.960 554.870 ;
        RECT 2879.760 531.490 2879.900 554.550 ;
        RECT 2877.000 531.350 2879.900 531.490 ;
        RECT 2877.000 483.210 2877.140 531.350 ;
        RECT 2877.000 483.070 2878.060 483.210 ;
        RECT 2877.920 445.130 2878.060 483.070 ;
        RECT 2877.920 444.990 2878.520 445.130 ;
        RECT 2878.380 407.050 2878.520 444.990 ;
        RECT 2877.920 406.910 2878.520 407.050 ;
        RECT 2877.920 396.850 2878.060 406.910 ;
        RECT 2877.920 396.710 2878.980 396.850 ;
        RECT 2878.840 292.810 2878.980 396.710 ;
        RECT 2878.840 292.670 2879.440 292.810 ;
        RECT 2879.300 266.290 2879.440 292.670 ;
        RECT 2879.300 266.150 2880.360 266.290 ;
        RECT 2880.220 263.570 2880.360 266.150 ;
        RECT 2878.840 263.430 2880.360 263.570 ;
        RECT 2878.840 261.530 2878.980 263.430 ;
        RECT 2877.920 261.390 2878.980 261.530 ;
        RECT 2877.920 260.170 2878.060 261.390 ;
        RECT 2877.460 260.030 2878.060 260.170 ;
        RECT 2877.460 232.970 2877.600 260.030 ;
        RECT 2877.460 232.830 2879.900 232.970 ;
        RECT 2879.760 232.210 2879.900 232.830 ;
        RECT 2879.700 231.890 2879.960 232.210 ;
        RECT 2880.160 230.870 2880.420 231.190 ;
        RECT 2880.220 207.130 2880.360 230.870 ;
        RECT 2878.380 206.990 2880.360 207.130 ;
        RECT 2878.380 197.610 2878.520 206.990 ;
        RECT 2878.380 197.470 2880.360 197.610 ;
        RECT 2880.220 167.010 2880.360 197.470 ;
        RECT 2879.760 166.870 2880.360 167.010 ;
        RECT 2879.760 165.570 2879.900 166.870 ;
        RECT 2879.700 165.250 2879.960 165.570 ;
        RECT 2879.700 141.450 2879.960 141.770 ;
        RECT 2879.760 106.490 2879.900 141.450 ;
        RECT 2879.760 106.350 2880.360 106.490 ;
        RECT 2880.220 102.410 2880.360 106.350 ;
        RECT 2877.000 102.270 2880.360 102.410 ;
        RECT 2877.000 76.570 2877.140 102.270 ;
        RECT 2875.620 76.430 2877.140 76.570 ;
        RECT 2875.620 37.730 2875.760 76.430 ;
        RECT 2875.560 37.410 2875.820 37.730 ;
        RECT 2879.700 37.410 2879.960 37.730 ;
        RECT 2879.760 16.845 2879.900 37.410 ;
        RECT 56.210 16.475 56.490 16.845 ;
        RECT 2879.690 16.475 2879.970 16.845 ;
        RECT 56.280 2.400 56.420 16.475 ;
        RECT 56.070 -4.800 56.630 2.400 ;
      LAYER via2 ;
        RECT 2881.530 3266.920 2881.810 3267.200 ;
        RECT 56.210 16.520 56.490 16.800 ;
        RECT 2879.690 16.520 2879.970 16.800 ;
      LAYER met3 ;
        RECT 2881.000 3269.800 2885.000 3270.400 ;
        RECT 2881.750 3267.225 2882.050 3269.800 ;
        RECT 2881.505 3266.910 2882.050 3267.225 ;
        RECT 2881.505 3266.895 2881.835 3266.910 ;
        RECT 56.185 16.810 56.515 16.825 ;
        RECT 2879.665 16.810 2879.995 16.825 ;
        RECT 56.185 16.510 2879.995 16.810 ;
        RECT 56.185 16.495 56.515 16.510 ;
        RECT 2879.665 16.495 2879.995 16.510 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 44.305 18.955 44.475 19.295 ;
        RECT 44.305 18.785 45.395 18.955 ;
      LAYER mcon ;
        RECT 44.305 19.125 44.475 19.295 ;
        RECT 45.225 18.785 45.395 18.955 ;
      LAYER met1 ;
        RECT 26.750 19.280 27.070 19.340 ;
        RECT 44.245 19.280 44.535 19.325 ;
        RECT 26.750 19.140 44.535 19.280 ;
        RECT 26.750 19.080 27.070 19.140 ;
        RECT 44.245 19.095 44.535 19.140 ;
        RECT 45.165 18.940 45.455 18.985 ;
        RECT 80.110 18.940 80.430 19.000 ;
        RECT 45.165 18.800 80.430 18.940 ;
        RECT 45.165 18.755 45.455 18.800 ;
        RECT 80.110 18.740 80.430 18.800 ;
      LAYER via ;
        RECT 26.780 19.080 27.040 19.340 ;
        RECT 80.140 18.740 80.400 19.000 ;
      LAYER met2 ;
        RECT 26.770 3266.875 27.050 3267.245 ;
        RECT 26.840 19.370 26.980 3266.875 ;
        RECT 26.780 19.050 27.040 19.370 ;
        RECT 80.140 18.710 80.400 19.030 ;
        RECT 80.200 2.400 80.340 18.710 ;
        RECT 79.990 -4.800 80.550 2.400 ;
      LAYER via2 ;
        RECT 26.770 3266.920 27.050 3267.200 ;
      LAYER met3 ;
        RECT 35.000 3269.800 39.000 3270.400 ;
        RECT 26.745 3267.210 27.075 3267.225 ;
        RECT 35.270 3267.210 35.570 3269.800 ;
        RECT 26.745 3266.910 35.570 3267.210 ;
        RECT 26.745 3266.895 27.075 3266.910 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2879.745 2589.865 2879.915 2611.455 ;
        RECT 2879.745 2547.365 2879.915 2573.715 ;
        RECT 2880.205 1980.245 2880.375 2028.015 ;
        RECT 2879.745 1639.905 2879.915 1673.055 ;
        RECT 2879.745 1595.365 2879.915 1609.815 ;
        RECT 2880.665 1077.545 2880.835 1088.255 ;
        RECT 2880.205 955.485 2880.375 963.815 ;
        RECT 2881.125 862.665 2881.295 886.295 ;
        RECT 2880.665 766.105 2880.835 790.075 ;
        RECT 2881.125 724.285 2881.295 729.895 ;
        RECT 2880.205 588.625 2880.375 612.935 ;
        RECT 2880.665 175.865 2880.835 218.195 ;
      LAYER mcon ;
        RECT 2879.745 2611.285 2879.915 2611.455 ;
        RECT 2879.745 2573.545 2879.915 2573.715 ;
        RECT 2880.205 2027.845 2880.375 2028.015 ;
        RECT 2879.745 1672.885 2879.915 1673.055 ;
        RECT 2879.745 1609.645 2879.915 1609.815 ;
        RECT 2880.665 1088.085 2880.835 1088.255 ;
        RECT 2880.205 963.645 2880.375 963.815 ;
        RECT 2881.125 886.125 2881.295 886.295 ;
        RECT 2880.665 789.905 2880.835 790.075 ;
        RECT 2881.125 729.725 2881.295 729.895 ;
        RECT 2880.205 612.765 2880.375 612.935 ;
        RECT 2880.665 218.025 2880.835 218.195 ;
      LAYER met1 ;
        RECT 2879.670 3374.740 2879.990 3374.800 ;
        RECT 2881.510 3374.740 2881.830 3374.800 ;
        RECT 2879.670 3374.600 2881.830 3374.740 ;
        RECT 2879.670 3374.540 2879.990 3374.600 ;
        RECT 2881.510 3374.540 2881.830 3374.600 ;
        RECT 2879.670 2611.440 2879.990 2611.500 ;
        RECT 2879.475 2611.300 2879.990 2611.440 ;
        RECT 2879.670 2611.240 2879.990 2611.300 ;
        RECT 2879.670 2590.020 2879.990 2590.080 ;
        RECT 2879.475 2589.880 2879.990 2590.020 ;
        RECT 2879.670 2589.820 2879.990 2589.880 ;
        RECT 2879.670 2573.700 2879.990 2573.760 ;
        RECT 2879.475 2573.560 2879.990 2573.700 ;
        RECT 2879.670 2573.500 2879.990 2573.560 ;
        RECT 2879.670 2547.520 2879.990 2547.580 ;
        RECT 2879.475 2547.380 2879.990 2547.520 ;
        RECT 2879.670 2547.320 2879.990 2547.380 ;
        RECT 2879.670 2428.860 2879.990 2428.920 ;
        RECT 2880.130 2428.860 2880.450 2428.920 ;
        RECT 2879.670 2428.720 2880.450 2428.860 ;
        RECT 2879.670 2428.660 2879.990 2428.720 ;
        RECT 2880.130 2428.660 2880.450 2428.720 ;
        RECT 2880.130 2332.300 2880.450 2332.360 ;
        RECT 2879.760 2332.160 2880.450 2332.300 ;
        RECT 2879.760 2331.340 2879.900 2332.160 ;
        RECT 2880.130 2332.100 2880.450 2332.160 ;
        RECT 2879.670 2331.080 2879.990 2331.340 ;
        RECT 2879.670 2138.300 2879.990 2138.560 ;
        RECT 2879.760 2137.880 2879.900 2138.300 ;
        RECT 2879.670 2137.620 2879.990 2137.880 ;
        RECT 2879.670 2028.000 2879.990 2028.060 ;
        RECT 2880.145 2028.000 2880.435 2028.045 ;
        RECT 2879.670 2027.860 2880.435 2028.000 ;
        RECT 2879.670 2027.800 2879.990 2027.860 ;
        RECT 2880.145 2027.815 2880.435 2027.860 ;
        RECT 2880.130 1980.400 2880.450 1980.460 ;
        RECT 2879.935 1980.260 2880.450 1980.400 ;
        RECT 2880.130 1980.200 2880.450 1980.260 ;
        RECT 2879.670 1673.040 2879.990 1673.100 ;
        RECT 2879.475 1672.900 2879.990 1673.040 ;
        RECT 2879.670 1672.840 2879.990 1672.900 ;
        RECT 2879.670 1640.060 2879.990 1640.120 ;
        RECT 2879.475 1639.920 2879.990 1640.060 ;
        RECT 2879.670 1639.860 2879.990 1639.920 ;
        RECT 2879.670 1609.800 2879.990 1609.860 ;
        RECT 2879.475 1609.660 2879.990 1609.800 ;
        RECT 2879.670 1609.600 2879.990 1609.660 ;
        RECT 2879.670 1595.520 2879.990 1595.580 ;
        RECT 2879.475 1595.380 2879.990 1595.520 ;
        RECT 2879.670 1595.320 2879.990 1595.380 ;
        RECT 2879.670 1266.200 2879.990 1266.460 ;
        RECT 2879.760 1265.440 2879.900 1266.200 ;
        RECT 2879.670 1265.180 2879.990 1265.440 ;
        RECT 2879.670 1088.240 2879.990 1088.300 ;
        RECT 2880.605 1088.240 2880.895 1088.285 ;
        RECT 2879.670 1088.100 2880.895 1088.240 ;
        RECT 2879.670 1088.040 2879.990 1088.100 ;
        RECT 2880.605 1088.055 2880.895 1088.100 ;
        RECT 2879.670 1077.700 2879.990 1077.760 ;
        RECT 2880.605 1077.700 2880.895 1077.745 ;
        RECT 2879.670 1077.560 2880.895 1077.700 ;
        RECT 2879.670 1077.500 2879.990 1077.560 ;
        RECT 2880.605 1077.515 2880.895 1077.560 ;
        RECT 2880.130 963.800 2880.450 963.860 ;
        RECT 2879.935 963.660 2880.450 963.800 ;
        RECT 2880.130 963.600 2880.450 963.660 ;
        RECT 2880.130 955.640 2880.450 955.700 ;
        RECT 2879.935 955.500 2880.450 955.640 ;
        RECT 2880.130 955.440 2880.450 955.500 ;
        RECT 2879.670 886.280 2879.990 886.340 ;
        RECT 2881.065 886.280 2881.355 886.325 ;
        RECT 2879.670 886.140 2881.355 886.280 ;
        RECT 2879.670 886.080 2879.990 886.140 ;
        RECT 2881.065 886.095 2881.355 886.140 ;
        RECT 2880.590 862.820 2880.910 862.880 ;
        RECT 2881.065 862.820 2881.355 862.865 ;
        RECT 2880.590 862.680 2881.355 862.820 ;
        RECT 2880.590 862.620 2880.910 862.680 ;
        RECT 2881.065 862.635 2881.355 862.680 ;
        RECT 2879.670 850.580 2879.990 850.640 ;
        RECT 2880.590 850.580 2880.910 850.640 ;
        RECT 2879.670 850.440 2880.910 850.580 ;
        RECT 2879.670 850.380 2879.990 850.440 ;
        RECT 2880.590 850.380 2880.910 850.440 ;
        RECT 2880.590 790.060 2880.910 790.120 ;
        RECT 2880.395 789.920 2880.910 790.060 ;
        RECT 2880.590 789.860 2880.910 789.920 ;
        RECT 2879.670 766.260 2879.990 766.320 ;
        RECT 2880.605 766.260 2880.895 766.305 ;
        RECT 2879.670 766.120 2880.895 766.260 ;
        RECT 2879.670 766.060 2879.990 766.120 ;
        RECT 2880.605 766.075 2880.895 766.120 ;
        RECT 2879.670 729.880 2879.990 729.940 ;
        RECT 2881.065 729.880 2881.355 729.925 ;
        RECT 2879.670 729.740 2881.355 729.880 ;
        RECT 2879.670 729.680 2879.990 729.740 ;
        RECT 2881.065 729.695 2881.355 729.740 ;
        RECT 2879.670 724.440 2879.990 724.500 ;
        RECT 2881.065 724.440 2881.355 724.485 ;
        RECT 2879.670 724.300 2881.355 724.440 ;
        RECT 2879.670 724.240 2879.990 724.300 ;
        RECT 2881.065 724.255 2881.355 724.300 ;
        RECT 2879.670 612.920 2879.990 612.980 ;
        RECT 2880.145 612.920 2880.435 612.965 ;
        RECT 2879.670 612.780 2880.435 612.920 ;
        RECT 2879.670 612.720 2879.990 612.780 ;
        RECT 2880.145 612.735 2880.435 612.780 ;
        RECT 2879.670 588.780 2879.990 588.840 ;
        RECT 2880.145 588.780 2880.435 588.825 ;
        RECT 2879.670 588.640 2880.435 588.780 ;
        RECT 2879.670 588.580 2879.990 588.640 ;
        RECT 2880.145 588.595 2880.435 588.640 ;
        RECT 2879.670 263.880 2879.990 264.140 ;
        RECT 2879.760 263.120 2879.900 263.880 ;
        RECT 2879.670 262.860 2879.990 263.120 ;
        RECT 2879.670 218.180 2879.990 218.240 ;
        RECT 2880.605 218.180 2880.895 218.225 ;
        RECT 2879.670 218.040 2880.895 218.180 ;
        RECT 2879.670 217.980 2879.990 218.040 ;
        RECT 2880.605 217.995 2880.895 218.040 ;
        RECT 2879.670 176.020 2879.990 176.080 ;
        RECT 2880.605 176.020 2880.895 176.065 ;
        RECT 2879.670 175.880 2880.895 176.020 ;
        RECT 2879.670 175.820 2879.990 175.880 ;
        RECT 2880.605 175.835 2880.895 175.880 ;
        RECT 2875.070 37.300 2875.390 37.360 ;
        RECT 2877.370 37.300 2877.690 37.360 ;
        RECT 2875.070 37.160 2877.690 37.300 ;
        RECT 2875.070 37.100 2875.390 37.160 ;
        RECT 2877.370 37.100 2877.690 37.160 ;
      LAYER via ;
        RECT 2879.700 3374.540 2879.960 3374.800 ;
        RECT 2881.540 3374.540 2881.800 3374.800 ;
        RECT 2879.700 2611.240 2879.960 2611.500 ;
        RECT 2879.700 2589.820 2879.960 2590.080 ;
        RECT 2879.700 2573.500 2879.960 2573.760 ;
        RECT 2879.700 2547.320 2879.960 2547.580 ;
        RECT 2879.700 2428.660 2879.960 2428.920 ;
        RECT 2880.160 2428.660 2880.420 2428.920 ;
        RECT 2880.160 2332.100 2880.420 2332.360 ;
        RECT 2879.700 2331.080 2879.960 2331.340 ;
        RECT 2879.700 2138.300 2879.960 2138.560 ;
        RECT 2879.700 2137.620 2879.960 2137.880 ;
        RECT 2879.700 2027.800 2879.960 2028.060 ;
        RECT 2880.160 1980.200 2880.420 1980.460 ;
        RECT 2879.700 1672.840 2879.960 1673.100 ;
        RECT 2879.700 1639.860 2879.960 1640.120 ;
        RECT 2879.700 1609.600 2879.960 1609.860 ;
        RECT 2879.700 1595.320 2879.960 1595.580 ;
        RECT 2879.700 1266.200 2879.960 1266.460 ;
        RECT 2879.700 1265.180 2879.960 1265.440 ;
        RECT 2879.700 1088.040 2879.960 1088.300 ;
        RECT 2879.700 1077.500 2879.960 1077.760 ;
        RECT 2880.160 963.600 2880.420 963.860 ;
        RECT 2880.160 955.440 2880.420 955.700 ;
        RECT 2879.700 886.080 2879.960 886.340 ;
        RECT 2880.620 862.620 2880.880 862.880 ;
        RECT 2879.700 850.380 2879.960 850.640 ;
        RECT 2880.620 850.380 2880.880 850.640 ;
        RECT 2880.620 789.860 2880.880 790.120 ;
        RECT 2879.700 766.060 2879.960 766.320 ;
        RECT 2879.700 729.680 2879.960 729.940 ;
        RECT 2879.700 724.240 2879.960 724.500 ;
        RECT 2879.700 612.720 2879.960 612.980 ;
        RECT 2879.700 588.580 2879.960 588.840 ;
        RECT 2879.700 263.880 2879.960 264.140 ;
        RECT 2879.700 262.860 2879.960 263.120 ;
        RECT 2879.700 217.980 2879.960 218.240 ;
        RECT 2879.700 175.820 2879.960 176.080 ;
        RECT 2875.100 37.100 2875.360 37.360 ;
        RECT 2877.400 37.100 2877.660 37.360 ;
      LAYER met2 ;
        RECT 2881.530 3376.355 2881.810 3376.725 ;
        RECT 2881.600 3374.830 2881.740 3376.355 ;
        RECT 2879.700 3374.570 2879.960 3374.830 ;
        RECT 2879.300 3374.510 2879.960 3374.570 ;
        RECT 2881.540 3374.510 2881.800 3374.830 ;
        RECT 2879.300 3374.430 2879.900 3374.510 ;
        RECT 2879.300 3346.690 2879.440 3374.430 ;
        RECT 2878.840 3346.550 2879.440 3346.690 ;
        RECT 2878.840 3263.050 2878.980 3346.550 ;
        RECT 2877.920 3262.910 2878.980 3263.050 ;
        RECT 2877.920 3261.690 2878.060 3262.910 ;
        RECT 2876.540 3261.550 2878.060 3261.690 ;
        RECT 2876.540 3236.530 2876.680 3261.550 ;
        RECT 2876.540 3236.390 2878.060 3236.530 ;
        RECT 2877.920 3221.570 2878.060 3236.390 ;
        RECT 2877.920 3221.430 2878.980 3221.570 ;
        RECT 2878.840 3126.370 2878.980 3221.430 ;
        RECT 2877.920 3126.230 2878.980 3126.370 ;
        RECT 2877.920 3115.490 2878.060 3126.230 ;
        RECT 2876.540 3115.350 2878.060 3115.490 ;
        RECT 2876.540 3042.730 2876.680 3115.350 ;
        RECT 2876.540 3042.590 2878.520 3042.730 ;
        RECT 2878.380 3011.450 2878.520 3042.590 ;
        RECT 2878.380 3011.310 2878.980 3011.450 ;
        RECT 2878.840 2958.410 2878.980 3011.310 ;
        RECT 2877.920 2958.270 2878.980 2958.410 ;
        RECT 2877.920 2908.090 2878.060 2958.270 ;
        RECT 2877.460 2907.950 2878.060 2908.090 ;
        RECT 2877.460 2814.930 2877.600 2907.950 ;
        RECT 2877.460 2814.790 2878.980 2814.930 ;
        RECT 2878.840 2780.250 2878.980 2814.790 ;
        RECT 2877.460 2780.110 2878.980 2780.250 ;
        RECT 2877.460 2718.370 2877.600 2780.110 ;
        RECT 2877.460 2718.230 2878.060 2718.370 ;
        RECT 2877.920 2704.770 2878.060 2718.230 ;
        RECT 2877.920 2704.630 2878.520 2704.770 ;
        RECT 2878.380 2611.610 2878.520 2704.630 ;
        RECT 2878.380 2611.530 2879.900 2611.610 ;
        RECT 2878.380 2611.470 2879.960 2611.530 ;
        RECT 2879.700 2611.210 2879.960 2611.470 ;
        RECT 2879.700 2589.850 2879.960 2590.110 ;
        RECT 2879.300 2589.790 2879.960 2589.850 ;
        RECT 2879.300 2589.710 2879.900 2589.790 ;
        RECT 2879.300 2573.700 2879.440 2589.710 ;
        RECT 2879.700 2573.700 2879.960 2573.790 ;
        RECT 2879.300 2573.560 2879.960 2573.700 ;
        RECT 2879.700 2573.470 2879.960 2573.560 ;
        RECT 2879.700 2547.290 2879.960 2547.610 ;
        RECT 2879.760 2547.010 2879.900 2547.290 ;
        RECT 2877.460 2546.870 2879.900 2547.010 ;
        RECT 2877.460 2525.250 2877.600 2546.870 ;
        RECT 2877.000 2525.110 2877.600 2525.250 ;
        RECT 2877.000 2523.890 2877.140 2525.110 ;
        RECT 2877.000 2523.750 2877.600 2523.890 ;
        RECT 2877.460 2475.610 2877.600 2523.750 ;
        RECT 2877.460 2475.470 2878.060 2475.610 ;
        RECT 2877.920 2434.810 2878.060 2475.470 ;
        RECT 2877.920 2434.670 2879.900 2434.810 ;
        RECT 2879.760 2428.950 2879.900 2434.670 ;
        RECT 2879.700 2428.630 2879.960 2428.950 ;
        RECT 2880.160 2428.630 2880.420 2428.950 ;
        RECT 2880.220 2332.390 2880.360 2428.630 ;
        RECT 2880.160 2332.070 2880.420 2332.390 ;
        RECT 2879.300 2331.370 2879.900 2331.450 ;
        RECT 2879.300 2331.310 2879.960 2331.370 ;
        RECT 2879.300 2318.530 2879.440 2331.310 ;
        RECT 2879.700 2331.050 2879.960 2331.310 ;
        RECT 2878.840 2318.390 2879.440 2318.530 ;
        RECT 2878.840 2246.450 2878.980 2318.390 ;
        RECT 2878.840 2246.310 2879.900 2246.450 ;
        RECT 2879.760 2234.890 2879.900 2246.310 ;
        RECT 2878.840 2234.750 2879.900 2234.890 ;
        RECT 2878.840 2211.090 2878.980 2234.750 ;
        RECT 2878.840 2210.950 2879.440 2211.090 ;
        RECT 2879.300 2166.210 2879.440 2210.950 ;
        RECT 2879.300 2166.070 2879.900 2166.210 ;
        RECT 2879.760 2138.590 2879.900 2166.070 ;
        RECT 2879.700 2138.270 2879.960 2138.590 ;
        RECT 2879.700 2137.590 2879.960 2137.910 ;
        RECT 2879.760 2118.610 2879.900 2137.590 ;
        RECT 2878.840 2118.470 2879.900 2118.610 ;
        RECT 2878.840 2114.530 2878.980 2118.470 ;
        RECT 2878.840 2114.390 2879.440 2114.530 ;
        RECT 2879.300 2028.000 2879.440 2114.390 ;
        RECT 2879.700 2028.000 2879.960 2028.090 ;
        RECT 2879.300 2027.860 2879.960 2028.000 ;
        RECT 2879.700 2027.770 2879.960 2027.860 ;
        RECT 2880.160 1980.170 2880.420 1980.490 ;
        RECT 2880.220 1921.410 2880.360 1980.170 ;
        RECT 2877.000 1921.270 2880.360 1921.410 ;
        RECT 2877.000 1895.570 2877.140 1921.270 ;
        RECT 2877.000 1895.430 2878.980 1895.570 ;
        RECT 2878.840 1860.890 2878.980 1895.430 ;
        RECT 2878.840 1860.750 2879.900 1860.890 ;
        RECT 2879.760 1847.970 2879.900 1860.750 ;
        RECT 2877.460 1847.830 2879.900 1847.970 ;
        RECT 2877.460 1800.370 2877.600 1847.830 ;
        RECT 2876.540 1800.230 2877.600 1800.370 ;
        RECT 2876.540 1782.010 2876.680 1800.230 ;
        RECT 2876.540 1781.870 2877.140 1782.010 ;
        RECT 2877.000 1751.410 2877.140 1781.870 ;
        RECT 2877.000 1751.270 2878.520 1751.410 ;
        RECT 2878.380 1750.050 2878.520 1751.270 ;
        RECT 2878.380 1749.910 2880.360 1750.050 ;
        RECT 2880.220 1736.450 2880.360 1749.910 ;
        RECT 2879.300 1736.310 2880.360 1736.450 ;
        RECT 2879.300 1735.770 2879.440 1736.310 ;
        RECT 2878.380 1735.630 2879.440 1735.770 ;
        RECT 2878.380 1684.090 2878.520 1735.630 ;
        RECT 2878.380 1683.950 2878.980 1684.090 ;
        RECT 2878.840 1683.410 2878.980 1683.950 ;
        RECT 2878.840 1683.270 2879.900 1683.410 ;
        RECT 2879.760 1673.130 2879.900 1683.270 ;
        RECT 2879.700 1672.810 2879.960 1673.130 ;
        RECT 2879.700 1639.830 2879.960 1640.150 ;
        RECT 2879.760 1609.890 2879.900 1639.830 ;
        RECT 2879.700 1609.570 2879.960 1609.890 ;
        RECT 2879.700 1595.290 2879.960 1595.610 ;
        RECT 2879.760 1595.010 2879.900 1595.290 ;
        RECT 2877.460 1594.870 2879.900 1595.010 ;
        RECT 2877.460 1483.490 2877.600 1594.870 ;
        RECT 2876.080 1483.350 2877.600 1483.490 ;
        RECT 2876.080 1439.970 2876.220 1483.350 ;
        RECT 2876.080 1439.830 2878.060 1439.970 ;
        RECT 2877.920 1438.610 2878.060 1439.830 ;
        RECT 2877.460 1438.470 2878.060 1438.610 ;
        RECT 2877.460 1399.850 2877.600 1438.470 ;
        RECT 2876.080 1399.710 2877.600 1399.850 ;
        RECT 2876.080 1307.370 2876.220 1399.710 ;
        RECT 2876.080 1307.230 2877.600 1307.370 ;
        RECT 2877.460 1266.570 2877.600 1307.230 ;
        RECT 2877.460 1266.490 2879.900 1266.570 ;
        RECT 2877.460 1266.430 2879.960 1266.490 ;
        RECT 2879.700 1266.170 2879.960 1266.430 ;
        RECT 2879.700 1265.210 2879.960 1265.470 ;
        RECT 2879.300 1265.150 2879.960 1265.210 ;
        RECT 2879.300 1265.070 2879.900 1265.150 ;
        RECT 2879.300 1233.250 2879.440 1265.070 ;
        RECT 2878.840 1233.110 2879.440 1233.250 ;
        RECT 2878.840 1172.730 2878.980 1233.110 ;
        RECT 2878.380 1172.590 2878.980 1172.730 ;
        RECT 2878.380 1088.240 2878.520 1172.590 ;
        RECT 2879.700 1088.240 2879.960 1088.330 ;
        RECT 2878.380 1088.100 2879.960 1088.240 ;
        RECT 2879.700 1088.010 2879.960 1088.100 ;
        RECT 2879.700 1077.470 2879.960 1077.790 ;
        RECT 2879.760 1061.210 2879.900 1077.470 ;
        RECT 2878.840 1061.070 2879.900 1061.210 ;
        RECT 2878.840 1014.800 2878.980 1061.070 ;
        RECT 2878.840 1014.660 2880.360 1014.800 ;
        RECT 2880.220 963.890 2880.360 1014.660 ;
        RECT 2880.160 963.570 2880.420 963.890 ;
        RECT 2880.160 955.410 2880.420 955.730 ;
        RECT 2880.220 931.330 2880.360 955.410 ;
        RECT 2878.380 931.190 2880.360 931.330 ;
        RECT 2878.380 886.450 2878.520 931.190 ;
        RECT 2878.380 886.370 2879.900 886.450 ;
        RECT 2878.380 886.310 2879.960 886.370 ;
        RECT 2879.700 886.050 2879.960 886.310 ;
        RECT 2880.620 862.590 2880.880 862.910 ;
        RECT 2880.680 850.670 2880.820 862.590 ;
        RECT 2879.700 850.350 2879.960 850.670 ;
        RECT 2880.620 850.350 2880.880 850.670 ;
        RECT 2879.760 849.050 2879.900 850.350 ;
        RECT 2878.380 848.910 2879.900 849.050 ;
        RECT 2878.380 830.010 2878.520 848.910 ;
        RECT 2878.380 829.870 2880.820 830.010 ;
        RECT 2880.680 790.150 2880.820 829.870 ;
        RECT 2880.620 789.830 2880.880 790.150 ;
        RECT 2879.700 766.090 2879.960 766.350 ;
        RECT 2879.300 766.030 2879.960 766.090 ;
        RECT 2879.300 765.950 2879.900 766.030 ;
        RECT 2879.300 730.730 2879.440 765.950 ;
        RECT 2879.300 730.590 2879.900 730.730 ;
        RECT 2879.760 729.970 2879.900 730.590 ;
        RECT 2879.700 729.650 2879.960 729.970 ;
        RECT 2873.780 724.530 2879.900 724.610 ;
        RECT 2873.780 724.470 2879.960 724.530 ;
        RECT 2873.780 679.730 2873.920 724.470 ;
        RECT 2879.700 724.210 2879.960 724.470 ;
        RECT 2877.000 680.950 2877.600 681.090 ;
        RECT 2877.000 679.730 2877.140 680.950 ;
        RECT 2873.780 679.590 2877.140 679.730 ;
        RECT 2877.460 645.050 2877.600 680.950 ;
        RECT 2876.080 644.910 2877.600 645.050 ;
        RECT 2876.080 639.780 2876.220 644.910 ;
        RECT 2876.080 639.640 2877.600 639.780 ;
        RECT 2877.460 627.370 2877.600 639.640 ;
        RECT 2877.000 627.230 2877.600 627.370 ;
        RECT 2877.000 620.740 2877.140 627.230 ;
        RECT 2877.000 620.600 2879.900 620.740 ;
        RECT 2879.760 613.010 2879.900 620.600 ;
        RECT 2879.700 612.690 2879.960 613.010 ;
        RECT 2879.700 588.610 2879.960 588.870 ;
        RECT 2879.300 588.550 2879.960 588.610 ;
        RECT 2879.300 588.470 2879.900 588.550 ;
        RECT 2879.300 579.770 2879.440 588.470 ;
        RECT 2878.840 579.630 2879.440 579.770 ;
        RECT 2878.840 570.930 2878.980 579.630 ;
        RECT 2878.840 570.790 2880.360 570.930 ;
        RECT 2880.220 555.290 2880.360 570.790 ;
        RECT 2875.620 555.150 2880.360 555.290 ;
        RECT 2875.620 507.010 2875.760 555.150 ;
        RECT 2875.160 506.870 2875.760 507.010 ;
        RECT 2875.160 460.090 2875.300 506.870 ;
        RECT 2875.160 459.950 2876.680 460.090 ;
        RECT 2876.540 421.330 2876.680 459.950 ;
        RECT 2876.080 421.190 2876.680 421.330 ;
        RECT 2876.080 310.490 2876.220 421.190 ;
        RECT 2876.080 310.350 2876.680 310.490 ;
        RECT 2876.540 262.210 2876.680 310.350 ;
        RECT 2877.920 264.790 2879.900 264.930 ;
        RECT 2877.920 262.210 2878.060 264.790 ;
        RECT 2879.760 264.170 2879.900 264.790 ;
        RECT 2879.700 263.850 2879.960 264.170 ;
        RECT 2879.700 262.830 2879.960 263.150 ;
        RECT 2876.540 262.070 2878.060 262.210 ;
        RECT 2879.760 257.450 2879.900 262.830 ;
        RECT 2879.760 257.310 2880.360 257.450 ;
        RECT 2877.460 232.150 2879.440 232.290 ;
        RECT 2877.460 218.690 2877.600 232.150 ;
        RECT 2879.300 231.610 2879.440 232.150 ;
        RECT 2880.220 231.610 2880.360 257.310 ;
        RECT 2879.300 231.470 2880.360 231.610 ;
        RECT 2877.460 218.550 2879.900 218.690 ;
        RECT 2879.760 218.270 2879.900 218.550 ;
        RECT 2879.700 217.950 2879.960 218.270 ;
        RECT 2879.700 175.790 2879.960 176.110 ;
        RECT 2879.760 175.170 2879.900 175.790 ;
        RECT 2878.840 175.030 2879.900 175.170 ;
        RECT 2878.840 107.850 2878.980 175.030 ;
        RECT 2877.000 107.710 2878.980 107.850 ;
        RECT 2877.000 107.170 2877.140 107.710 ;
        RECT 2876.540 107.030 2877.140 107.170 ;
        RECT 2876.540 82.690 2876.680 107.030 ;
        RECT 2875.160 82.550 2876.680 82.690 ;
        RECT 2875.160 37.390 2875.300 82.550 ;
        RECT 2875.100 37.070 2875.360 37.390 ;
        RECT 2877.400 37.070 2877.660 37.390 ;
        RECT 2877.460 18.205 2877.600 37.070 ;
        RECT 103.590 17.835 103.870 18.205 ;
        RECT 2877.390 17.835 2877.670 18.205 ;
        RECT 103.660 2.400 103.800 17.835 ;
        RECT 103.450 -4.800 104.010 2.400 ;
      LAYER via2 ;
        RECT 2881.530 3376.400 2881.810 3376.680 ;
        RECT 103.590 17.880 103.870 18.160 ;
        RECT 2877.390 17.880 2877.670 18.160 ;
      LAYER met3 ;
        RECT 2881.000 3379.280 2885.000 3379.880 ;
        RECT 2881.750 3376.705 2882.050 3379.280 ;
        RECT 2881.505 3376.390 2882.050 3376.705 ;
        RECT 2881.505 3376.375 2881.835 3376.390 ;
        RECT 103.565 18.170 103.895 18.185 ;
        RECT 2877.365 18.170 2877.695 18.185 ;
        RECT 103.565 17.870 2877.695 18.170 ;
        RECT 103.565 17.855 103.895 17.870 ;
        RECT 2877.365 17.855 2877.695 17.870 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2808.430 35.000 2808.710 39.000 ;
        RECT 2808.460 25.005 2808.600 35.000 ;
        RECT 127.510 24.635 127.790 25.005 ;
        RECT 2808.390 24.635 2808.670 25.005 ;
        RECT 127.580 2.400 127.720 24.635 ;
        RECT 127.370 -4.800 127.930 2.400 ;
      LAYER via2 ;
        RECT 127.510 24.680 127.790 24.960 ;
        RECT 2808.390 24.680 2808.670 24.960 ;
      LAYER met3 ;
        RECT 127.485 24.970 127.815 24.985 ;
        RECT 2808.365 24.970 2808.695 24.985 ;
        RECT 127.485 24.670 2808.695 24.970 ;
        RECT 127.485 24.655 127.815 24.670 ;
        RECT 2808.365 24.655 2808.695 24.670 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2859.490 35.000 2859.770 39.000 ;
        RECT 2859.520 24.325 2859.660 35.000 ;
        RECT 26.310 23.955 26.590 24.325 ;
        RECT 2859.450 23.955 2859.730 24.325 ;
        RECT 26.380 2.400 26.520 23.955 ;
        RECT 26.170 -4.800 26.730 2.400 ;
      LAYER via2 ;
        RECT 26.310 24.000 26.590 24.280 ;
        RECT 2859.450 24.000 2859.730 24.280 ;
      LAYER met3 ;
        RECT 26.285 24.290 26.615 24.305 ;
        RECT 2859.425 24.290 2859.755 24.305 ;
        RECT 26.285 23.990 2859.755 24.290 ;
        RECT 26.285 23.975 26.615 23.990 ;
        RECT 2859.425 23.975 2859.755 23.990 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 27.210 17.580 27.530 17.640 ;
        RECT 32.270 17.580 32.590 17.640 ;
        RECT 27.210 17.440 32.590 17.580 ;
        RECT 27.210 17.380 27.530 17.440 ;
        RECT 32.270 17.380 32.590 17.440 ;
      LAYER via ;
        RECT 27.240 17.380 27.500 17.640 ;
        RECT 32.300 17.380 32.560 17.640 ;
      LAYER met2 ;
        RECT 27.230 3376.355 27.510 3376.725 ;
        RECT 27.300 17.670 27.440 3376.355 ;
        RECT 27.240 17.350 27.500 17.670 ;
        RECT 32.300 17.350 32.560 17.670 ;
        RECT 32.360 2.400 32.500 17.350 ;
        RECT 32.150 -4.800 32.710 2.400 ;
      LAYER via2 ;
        RECT 27.230 3376.400 27.510 3376.680 ;
      LAYER met3 ;
        RECT 35.000 3379.280 39.000 3379.880 ;
        RECT 27.205 3376.690 27.535 3376.705 ;
        RECT 35.270 3376.690 35.570 3379.280 ;
        RECT 27.205 3376.390 35.570 3376.690 ;
        RECT 27.205 3376.375 27.535 3376.390 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -14.580 -9.220 -11.580 3528.900 ;
        RECT 2931.200 -9.220 2934.200 3528.900 ;
      LAYER via4 ;
        RECT -13.670 3527.610 -12.490 3528.790 ;
        RECT -13.670 3526.010 -12.490 3527.190 ;
        RECT -13.670 -7.510 -12.490 -6.330 ;
        RECT -13.670 -9.110 -12.490 -7.930 ;
        RECT 2932.110 3527.610 2933.290 3528.790 ;
        RECT 2932.110 3526.010 2933.290 3527.190 ;
        RECT 2932.110 -7.510 2933.290 -6.330 ;
        RECT 2932.110 -9.110 2933.290 -7.930 ;
      LAYER met5 ;
        RECT -14.580 3528.900 -11.580 3528.910 ;
        RECT 2931.200 3528.900 2934.200 3528.910 ;
        RECT -14.580 3525.900 2934.200 3528.900 ;
        RECT -14.580 3525.890 -11.580 3525.900 ;
        RECT 2931.200 3525.890 2934.200 3525.900 ;
        RECT -14.580 -6.220 -11.580 -6.210 ;
        RECT 2931.200 -6.220 2934.200 -6.210 ;
        RECT -14.580 -9.220 2934.200 -6.220 ;
        RECT -14.580 -9.230 -11.580 -9.220 ;
        RECT 2931.200 -9.230 2934.200 -9.220 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.180 -13.820 -16.180 3533.500 ;
        RECT 2935.800 -13.820 2938.800 3533.500 ;
      LAYER via4 ;
        RECT -18.270 3532.210 -17.090 3533.390 ;
        RECT -18.270 3530.610 -17.090 3531.790 ;
        RECT -18.270 -12.110 -17.090 -10.930 ;
        RECT -18.270 -13.710 -17.090 -12.530 ;
        RECT 2936.710 3532.210 2937.890 3533.390 ;
        RECT 2936.710 3530.610 2937.890 3531.790 ;
        RECT 2936.710 -12.110 2937.890 -10.930 ;
        RECT 2936.710 -13.710 2937.890 -12.530 ;
      LAYER met5 ;
        RECT -19.180 3533.500 -16.180 3533.510 ;
        RECT 2935.800 3533.500 2938.800 3533.510 ;
        RECT -19.180 3530.500 2938.800 3533.500 ;
        RECT -19.180 3530.490 -16.180 3530.500 ;
        RECT 2935.800 3530.490 2938.800 3530.500 ;
        RECT -19.180 -10.820 -16.180 -10.810 ;
        RECT 2935.800 -10.820 2938.800 -10.810 ;
        RECT -19.180 -13.820 2938.800 -10.820 ;
        RECT -19.180 -13.830 -16.180 -13.820 ;
        RECT 2935.800 -13.830 2938.800 -13.820 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -23.780 -18.420 -20.780 3538.100 ;
        RECT 2940.400 -18.420 2943.400 3538.100 ;
      LAYER via4 ;
        RECT -22.870 3536.810 -21.690 3537.990 ;
        RECT -22.870 3535.210 -21.690 3536.390 ;
        RECT -22.870 -16.710 -21.690 -15.530 ;
        RECT -22.870 -18.310 -21.690 -17.130 ;
        RECT 2941.310 3536.810 2942.490 3537.990 ;
        RECT 2941.310 3535.210 2942.490 3536.390 ;
        RECT 2941.310 -16.710 2942.490 -15.530 ;
        RECT 2941.310 -18.310 2942.490 -17.130 ;
      LAYER met5 ;
        RECT -23.780 3538.100 -20.780 3538.110 ;
        RECT 2940.400 3538.100 2943.400 3538.110 ;
        RECT -23.780 3535.100 2943.400 3538.100 ;
        RECT -23.780 3535.090 -20.780 3535.100 ;
        RECT 2940.400 3535.090 2943.400 3535.100 ;
        RECT -23.780 -15.420 -20.780 -15.410 ;
        RECT 2940.400 -15.420 2943.400 -15.410 ;
        RECT -23.780 -18.420 2943.400 -15.420 ;
        RECT -23.780 -18.430 -20.780 -18.420 ;
        RECT 2940.400 -18.430 2943.400 -18.420 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -28.380 -23.020 -25.380 3542.700 ;
        RECT 2945.000 -23.020 2948.000 3542.700 ;
      LAYER via4 ;
        RECT -27.470 3541.410 -26.290 3542.590 ;
        RECT -27.470 3539.810 -26.290 3540.990 ;
        RECT -27.470 -21.310 -26.290 -20.130 ;
        RECT -27.470 -22.910 -26.290 -21.730 ;
        RECT 2945.910 3541.410 2947.090 3542.590 ;
        RECT 2945.910 3539.810 2947.090 3540.990 ;
        RECT 2945.910 -21.310 2947.090 -20.130 ;
        RECT 2945.910 -22.910 2947.090 -21.730 ;
      LAYER met5 ;
        RECT -28.380 3542.700 -25.380 3542.710 ;
        RECT 2945.000 3542.700 2948.000 3542.710 ;
        RECT -28.380 3539.700 2948.000 3542.700 ;
        RECT -28.380 3539.690 -25.380 3539.700 ;
        RECT 2945.000 3539.690 2948.000 3539.700 ;
        RECT -28.380 -20.020 -25.380 -20.010 ;
        RECT 2945.000 -20.020 2948.000 -20.010 ;
        RECT -28.380 -23.020 2948.000 -20.020 ;
        RECT -28.380 -23.030 -25.380 -23.020 ;
        RECT 2945.000 -23.030 2948.000 -23.020 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -32.980 -27.620 -29.980 3547.300 ;
        RECT 2949.600 -27.620 2952.600 3547.300 ;
      LAYER via4 ;
        RECT -32.070 3546.010 -30.890 3547.190 ;
        RECT -32.070 3544.410 -30.890 3545.590 ;
        RECT -32.070 -25.910 -30.890 -24.730 ;
        RECT -32.070 -27.510 -30.890 -26.330 ;
        RECT 2950.510 3546.010 2951.690 3547.190 ;
        RECT 2950.510 3544.410 2951.690 3545.590 ;
        RECT 2950.510 -25.910 2951.690 -24.730 ;
        RECT 2950.510 -27.510 2951.690 -26.330 ;
      LAYER met5 ;
        RECT -32.980 3547.300 -29.980 3547.310 ;
        RECT 2949.600 3547.300 2952.600 3547.310 ;
        RECT -32.980 3544.300 2952.600 3547.300 ;
        RECT -32.980 3544.290 -29.980 3544.300 ;
        RECT 2949.600 3544.290 2952.600 3544.300 ;
        RECT -32.980 -24.620 -29.980 -24.610 ;
        RECT 2949.600 -24.620 2952.600 -24.610 ;
        RECT -32.980 -27.620 2952.600 -24.620 ;
        RECT -32.980 -27.630 -29.980 -27.620 ;
        RECT 2949.600 -27.630 2952.600 -27.620 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -37.580 -32.220 -34.580 3551.900 ;
        RECT 2954.200 -32.220 2957.200 3551.900 ;
      LAYER via4 ;
        RECT -36.670 3550.610 -35.490 3551.790 ;
        RECT -36.670 3549.010 -35.490 3550.190 ;
        RECT -36.670 -30.510 -35.490 -29.330 ;
        RECT -36.670 -32.110 -35.490 -30.930 ;
        RECT 2955.110 3550.610 2956.290 3551.790 ;
        RECT 2955.110 3549.010 2956.290 3550.190 ;
        RECT 2955.110 -30.510 2956.290 -29.330 ;
        RECT 2955.110 -32.110 2956.290 -30.930 ;
      LAYER met5 ;
        RECT -37.580 3551.900 -34.580 3551.910 ;
        RECT 2954.200 3551.900 2957.200 3551.910 ;
        RECT -37.580 3548.900 2957.200 3551.900 ;
        RECT -37.580 3548.890 -34.580 3548.900 ;
        RECT 2954.200 3548.890 2957.200 3548.900 ;
        RECT -37.580 -29.220 -34.580 -29.210 ;
        RECT 2954.200 -29.220 2957.200 -29.210 ;
        RECT -37.580 -32.220 2957.200 -29.220 ;
        RECT -37.580 -32.230 -34.580 -32.220 ;
        RECT 2954.200 -32.230 2957.200 -32.220 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -42.180 -36.820 -39.180 3556.500 ;
        RECT 2958.800 -36.820 2961.800 3556.500 ;
      LAYER via4 ;
        RECT -41.270 3555.210 -40.090 3556.390 ;
        RECT -41.270 3553.610 -40.090 3554.790 ;
        RECT -41.270 -35.110 -40.090 -33.930 ;
        RECT -41.270 -36.710 -40.090 -35.530 ;
        RECT 2959.710 3555.210 2960.890 3556.390 ;
        RECT 2959.710 3553.610 2960.890 3554.790 ;
        RECT 2959.710 -35.110 2960.890 -33.930 ;
        RECT 2959.710 -36.710 2960.890 -35.530 ;
      LAYER met5 ;
        RECT -42.180 3556.500 -39.180 3556.510 ;
        RECT 2958.800 3556.500 2961.800 3556.510 ;
        RECT -42.180 3553.500 2961.800 3556.500 ;
        RECT -42.180 3553.490 -39.180 3553.500 ;
        RECT 2958.800 3553.490 2961.800 3553.500 ;
        RECT -42.180 -33.820 -39.180 -33.810 ;
        RECT 2958.800 -33.820 2961.800 -33.810 ;
        RECT -42.180 -36.820 2961.800 -33.820 ;
        RECT -42.180 -36.830 -39.180 -36.820 ;
        RECT 2958.800 -36.830 2961.800 -36.820 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 40.520 45.795 2879.180 3424.205 ;
      LAYER met1 ;
        RECT 40.520 39.460 2879.180 3424.360 ;
      LAYER met2 ;
        RECT 49.350 3430.720 89.550 3431.000 ;
        RECT 90.390 3430.720 199.030 3431.000 ;
        RECT 199.870 3430.720 308.510 3431.000 ;
        RECT 309.350 3430.720 417.990 3431.000 ;
        RECT 418.830 3430.720 527.930 3431.000 ;
        RECT 528.770 3430.720 637.410 3431.000 ;
        RECT 638.250 3430.720 746.890 3431.000 ;
        RECT 747.730 3430.720 856.830 3431.000 ;
        RECT 857.670 3430.720 966.310 3431.000 ;
        RECT 967.150 3430.720 1075.790 3431.000 ;
        RECT 1076.630 3430.720 1185.730 3431.000 ;
        RECT 1186.570 3430.720 1295.210 3431.000 ;
        RECT 1296.050 3430.720 1404.690 3431.000 ;
        RECT 1405.530 3430.720 1514.630 3431.000 ;
        RECT 1515.470 3430.720 1624.110 3431.000 ;
        RECT 1624.950 3430.720 1733.590 3431.000 ;
        RECT 1734.430 3430.720 1843.070 3431.000 ;
        RECT 1843.910 3430.720 1953.010 3431.000 ;
        RECT 1953.850 3430.720 2062.490 3431.000 ;
        RECT 2063.330 3430.720 2171.970 3431.000 ;
        RECT 2172.810 3430.720 2281.910 3431.000 ;
        RECT 2282.750 3430.720 2391.390 3431.000 ;
        RECT 2392.230 3430.720 2500.870 3431.000 ;
        RECT 2501.710 3430.720 2610.810 3431.000 ;
        RECT 2611.650 3430.720 2720.290 3431.000 ;
        RECT 2721.130 3430.720 2829.770 3431.000 ;
        RECT 2830.610 3430.720 2870.810 3431.000 ;
        RECT 49.350 39.280 2870.810 3430.720 ;
        RECT 49.350 39.000 60.110 39.280 ;
        RECT 60.950 39.000 110.710 39.280 ;
        RECT 111.550 39.000 161.770 39.280 ;
        RECT 162.610 39.000 212.370 39.280 ;
        RECT 213.210 39.000 263.430 39.280 ;
        RECT 264.270 39.000 314.490 39.280 ;
        RECT 315.330 39.000 365.090 39.280 ;
        RECT 365.930 39.000 416.150 39.280 ;
        RECT 416.990 39.000 467.210 39.280 ;
        RECT 468.050 39.000 517.810 39.280 ;
        RECT 518.650 39.000 568.870 39.280 ;
        RECT 569.710 39.000 619.930 39.280 ;
        RECT 620.770 39.000 670.530 39.280 ;
        RECT 671.370 39.000 721.590 39.280 ;
        RECT 722.430 39.000 772.650 39.280 ;
        RECT 773.490 39.000 823.250 39.280 ;
        RECT 824.090 39.000 874.310 39.280 ;
        RECT 875.150 39.000 924.910 39.280 ;
        RECT 925.750 39.000 975.970 39.280 ;
        RECT 976.810 39.000 1027.030 39.280 ;
        RECT 1027.870 39.000 1077.630 39.280 ;
        RECT 1078.470 39.000 1128.690 39.280 ;
        RECT 1129.530 39.000 1179.750 39.280 ;
        RECT 1180.590 39.000 1230.350 39.280 ;
        RECT 1231.190 39.000 1281.410 39.280 ;
        RECT 1282.250 39.000 1332.470 39.280 ;
        RECT 1333.310 39.000 1383.070 39.280 ;
        RECT 1383.910 39.000 1434.130 39.280 ;
        RECT 1434.970 39.000 1485.190 39.280 ;
        RECT 1486.030 39.000 1535.790 39.280 ;
        RECT 1536.630 39.000 1586.850 39.280 ;
        RECT 1587.690 39.000 1637.450 39.280 ;
        RECT 1638.290 39.000 1688.510 39.280 ;
        RECT 1689.350 39.000 1739.570 39.280 ;
        RECT 1740.410 39.000 1790.170 39.280 ;
        RECT 1791.010 39.000 1841.230 39.280 ;
        RECT 1842.070 39.000 1892.290 39.280 ;
        RECT 1893.130 39.000 1942.890 39.280 ;
        RECT 1943.730 39.000 1993.950 39.280 ;
        RECT 1994.790 39.000 2045.010 39.280 ;
        RECT 2045.850 39.000 2095.610 39.280 ;
        RECT 2096.450 39.000 2146.670 39.280 ;
        RECT 2147.510 39.000 2197.730 39.280 ;
        RECT 2198.570 39.000 2248.330 39.280 ;
        RECT 2249.170 39.000 2299.390 39.280 ;
        RECT 2300.230 39.000 2349.990 39.280 ;
        RECT 2350.830 39.000 2401.050 39.280 ;
        RECT 2401.890 39.000 2452.110 39.280 ;
        RECT 2452.950 39.000 2502.710 39.280 ;
        RECT 2503.550 39.000 2553.770 39.280 ;
        RECT 2554.610 39.000 2604.830 39.280 ;
        RECT 2605.670 39.000 2655.430 39.280 ;
        RECT 2656.270 39.000 2706.490 39.280 ;
        RECT 2707.330 39.000 2757.550 39.280 ;
        RECT 2758.390 39.000 2808.150 39.280 ;
        RECT 2808.990 39.000 2859.210 39.280 ;
        RECT 2860.050 39.000 2870.810 39.280 ;
      LAYER met3 ;
        RECT 39.000 3380.280 2881.000 3430.745 ;
        RECT 39.400 3378.880 2880.600 3380.280 ;
        RECT 39.000 3270.800 2881.000 3378.880 ;
        RECT 39.400 3269.400 2880.600 3270.800 ;
        RECT 39.000 3161.320 2881.000 3269.400 ;
        RECT 39.400 3159.920 2880.600 3161.320 ;
        RECT 39.000 3051.160 2881.000 3159.920 ;
        RECT 39.400 3049.760 2880.600 3051.160 ;
        RECT 39.000 2941.680 2881.000 3049.760 ;
        RECT 39.400 2940.280 2880.600 2941.680 ;
        RECT 39.000 2832.200 2881.000 2940.280 ;
        RECT 39.400 2830.800 2880.600 2832.200 ;
        RECT 39.000 2722.040 2881.000 2830.800 ;
        RECT 39.400 2720.640 2880.600 2722.040 ;
        RECT 39.000 2612.560 2881.000 2720.640 ;
        RECT 39.400 2611.160 2880.600 2612.560 ;
        RECT 39.000 2503.080 2881.000 2611.160 ;
        RECT 39.400 2501.680 2880.600 2503.080 ;
        RECT 39.000 2393.600 2881.000 2501.680 ;
        RECT 39.400 2392.200 2880.600 2393.600 ;
        RECT 39.000 2283.440 2881.000 2392.200 ;
        RECT 39.400 2282.040 2880.600 2283.440 ;
        RECT 39.000 2173.960 2881.000 2282.040 ;
        RECT 39.400 2172.560 2880.600 2173.960 ;
        RECT 39.000 2064.480 2881.000 2172.560 ;
        RECT 39.400 2063.080 2880.600 2064.480 ;
        RECT 39.000 1954.320 2881.000 2063.080 ;
        RECT 39.400 1952.920 2880.600 1954.320 ;
        RECT 39.000 1844.840 2881.000 1952.920 ;
        RECT 39.400 1843.440 2880.600 1844.840 ;
        RECT 39.000 1735.360 2881.000 1843.440 ;
        RECT 39.400 1733.960 2880.600 1735.360 ;
        RECT 39.000 1625.880 2881.000 1733.960 ;
        RECT 39.400 1624.480 2880.600 1625.880 ;
        RECT 39.000 1515.720 2881.000 1624.480 ;
        RECT 39.400 1514.320 2880.600 1515.720 ;
        RECT 39.000 1406.240 2881.000 1514.320 ;
        RECT 39.400 1404.840 2880.600 1406.240 ;
        RECT 39.000 1296.760 2881.000 1404.840 ;
        RECT 39.400 1295.360 2880.600 1296.760 ;
        RECT 39.000 1186.600 2881.000 1295.360 ;
        RECT 39.400 1185.200 2880.600 1186.600 ;
        RECT 39.000 1077.120 2881.000 1185.200 ;
        RECT 39.400 1075.720 2880.600 1077.120 ;
        RECT 39.000 967.640 2881.000 1075.720 ;
        RECT 39.400 966.240 2880.600 967.640 ;
        RECT 39.000 858.160 2881.000 966.240 ;
        RECT 39.400 856.760 2880.600 858.160 ;
        RECT 39.000 748.000 2881.000 856.760 ;
        RECT 39.400 746.600 2880.600 748.000 ;
        RECT 39.000 638.520 2881.000 746.600 ;
        RECT 39.400 637.120 2880.600 638.520 ;
        RECT 39.000 529.040 2881.000 637.120 ;
        RECT 39.400 527.640 2880.600 529.040 ;
        RECT 39.000 418.880 2881.000 527.640 ;
        RECT 39.400 417.480 2880.600 418.880 ;
        RECT 39.000 309.400 2881.000 417.480 ;
        RECT 39.400 308.000 2880.600 309.400 ;
        RECT 39.000 199.920 2881.000 308.000 ;
        RECT 39.400 198.520 2880.600 199.920 ;
        RECT 39.000 90.440 2881.000 198.520 ;
        RECT 39.400 89.040 2880.600 90.440 ;
        RECT 39.000 45.715 2881.000 89.040 ;
      LAYER met4 ;
        RECT 56.040 45.640 123.500 3424.360 ;
      LAYER met4 ;
        RECT 123.500 35.000 126.500 3435.000 ;
      LAYER met4 ;
        RECT 126.500 45.640 313.500 3424.360 ;
      LAYER met4 ;
        RECT 313.500 35.000 316.500 3435.000 ;
      LAYER met4 ;
        RECT 316.500 45.640 503.500 3424.360 ;
      LAYER met4 ;
        RECT 503.500 35.000 506.500 3435.000 ;
      LAYER met4 ;
        RECT 506.500 45.640 693.500 3424.360 ;
      LAYER met4 ;
        RECT 693.500 35.000 696.500 3435.000 ;
      LAYER met4 ;
        RECT 696.500 45.640 883.500 3424.360 ;
      LAYER met4 ;
        RECT 883.500 35.000 886.500 3435.000 ;
      LAYER met4 ;
        RECT 886.500 45.640 1073.500 3424.360 ;
      LAYER met4 ;
        RECT 1073.500 35.000 1076.500 3435.000 ;
      LAYER met4 ;
        RECT 1076.500 45.640 1263.500 3424.360 ;
      LAYER met4 ;
        RECT 1263.500 35.000 1266.500 3435.000 ;
      LAYER met4 ;
        RECT 1266.500 45.640 1453.500 3424.360 ;
      LAYER met4 ;
        RECT 1453.500 35.000 1456.500 3435.000 ;
      LAYER met4 ;
        RECT 1456.500 45.640 1643.500 3424.360 ;
      LAYER met4 ;
        RECT 1643.500 35.000 1646.500 3435.000 ;
      LAYER met4 ;
        RECT 1646.500 45.640 1833.500 3424.360 ;
      LAYER met4 ;
        RECT 1833.500 35.000 1836.500 3435.000 ;
      LAYER met4 ;
        RECT 1836.500 45.640 2023.500 3424.360 ;
      LAYER met4 ;
        RECT 2023.500 35.000 2026.500 3435.000 ;
      LAYER met4 ;
        RECT 2026.500 45.640 2213.500 3424.360 ;
      LAYER met4 ;
        RECT 2213.500 35.000 2216.500 3435.000 ;
      LAYER met4 ;
        RECT 2216.500 45.640 2403.500 3424.360 ;
      LAYER met4 ;
        RECT 2403.500 35.000 2406.500 3435.000 ;
      LAYER met4 ;
        RECT 2406.500 45.640 2593.500 3424.360 ;
      LAYER met4 ;
        RECT 2593.500 35.000 2596.500 3435.000 ;
      LAYER met4 ;
        RECT 2596.500 45.640 2783.500 3424.360 ;
      LAYER met4 ;
        RECT 2783.500 35.000 2786.500 3435.000 ;
      LAYER met4 ;
        RECT 2786.500 45.640 2822.440 3424.360 ;
      LAYER met5 ;
        RECT 40.520 138.080 2879.180 3394.755 ;
      LAYER met5 ;
        RECT 40.520 99.785 2879.180 101.385 ;
        RECT 40.520 61.490 2879.180 63.090 ;
  END
END user_project_wrapper
END LIBRARY


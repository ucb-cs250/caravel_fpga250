magic
tech sky130A
magscale 1 2
timestamp 1607933928
<< locali >>
rect 11713 679711 11747 679813
rect 16589 679711 16623 679813
rect 31033 679711 31067 679813
rect 35909 679711 35943 679813
rect 50353 679711 50387 679813
rect 55229 679711 55263 679813
rect 69673 679711 69707 679813
rect 74549 679711 74583 679813
rect 88993 679711 89027 679813
rect 93869 679711 93903 679813
rect 108313 679711 108347 679813
rect 113189 679711 113223 679813
rect 127633 679711 127667 679813
rect 132509 679711 132543 679813
rect 146953 679711 146987 679813
rect 151829 679711 151863 679813
rect 166273 679711 166307 679813
rect 171149 679711 171183 679813
rect 185593 679711 185627 679813
rect 190469 679711 190503 679813
rect 204913 679711 204947 679813
rect 207029 679167 207063 680289
rect 209789 679711 209823 679813
rect 216597 679779 216631 680357
rect 222059 679813 222151 679847
rect 222117 679779 222151 679813
rect 231961 679779 231995 680357
rect 222209 679575 222243 679677
rect 231777 679575 231811 679745
rect 364809 679575 364843 680289
rect 370237 679575 370271 680289
rect 380081 679575 380115 680357
rect 394525 680255 394559 680357
rect 394709 679575 394743 680357
rect 403173 679575 403207 680357
rect 412649 680051 412683 680221
rect 412741 679575 412775 680357
rect 418629 679575 418663 680357
rect 428013 679983 428047 680357
rect 428197 679575 428231 680357
rect 434729 679847 434763 679949
rect 437765 679575 437799 680357
rect 443561 679167 443595 680357
rect 444297 679847 444331 680085
rect 451289 679983 451323 680221
rect 451381 679575 451415 680357
rect 457177 679575 457211 680357
rect 461593 679983 461627 680221
rect 466561 679575 466595 680357
rect 469597 680119 469631 680221
rect 474749 680051 474783 680357
rect 481039 680289 481131 680323
rect 478003 680153 478153 680187
rect 481097 679983 481131 680289
rect 481189 679575 481223 680289
rect 485697 679915 485731 680085
rect 485639 679881 485731 679915
rect 485789 679575 485823 680289
rect 489745 679983 489779 680289
rect 490481 679847 490515 680221
rect 494069 679983 494103 680357
rect 495449 679575 495483 680357
rect 500233 679847 500267 680221
rect 502257 679235 502291 680357
rect 505937 679575 505971 680357
rect 506489 679915 506523 680085
rect 509801 679779 509835 680221
rect 515413 679575 515447 680357
rect 516333 679779 516367 680085
rect 519553 679847 519587 680153
rect 522129 679303 522163 680357
rect 524429 679575 524463 680357
rect 529029 679779 529063 680085
rect 529121 679847 529155 680153
rect 529213 679915 529247 680085
rect 533997 679779 534031 680221
rect 534365 679575 534399 680357
rect 538873 679915 538907 680221
rect 543749 679779 543783 680357
rect 544025 679575 544059 680357
rect 546877 679915 546911 680221
rect 553409 679779 553443 680221
rect 553501 679847 553535 680289
rect 554881 679167 554915 680289
rect 557733 680119 557767 680425
rect 559205 679983 559239 680289
rect 560769 679167 560803 680289
rect 561597 679915 561631 680289
rect 561781 679847 561815 680289
rect 561873 679303 561907 680289
rect 562517 679235 562551 680289
rect 569969 654075 570003 659209
rect 1869 633471 1903 642617
rect 1961 639319 1995 648057
rect 1685 600559 1719 601069
rect 1777 599743 1811 601953
rect 1869 597023 1903 602361
rect 1961 599879 1995 602089
rect 1869 566627 1903 580465
rect 1961 566559 1995 580193
rect 1869 566525 1995 566559
rect 1685 563431 1719 564417
rect 1777 563159 1811 565505
rect 1869 561119 1903 566525
rect 1961 547723 1995 563737
rect 569969 551055 570003 552041
rect 1685 526983 1719 527085
rect 1685 526167 1719 526473
rect 1777 522495 1811 527153
rect 1869 522359 1903 527697
rect 1961 510663 1995 529193
rect 569969 528887 570003 530961
rect 570061 528751 570095 531097
rect 569969 518483 570003 522597
rect 570061 521067 570095 522461
rect 1501 502231 1535 507161
rect 1593 501823 1627 507297
rect 1777 504883 1811 506073
rect 1869 504475 1903 509881
rect 1685 493391 1719 502265
rect 1777 497539 1811 504101
rect 1961 497539 1995 510017
rect 569969 503047 570003 505121
rect 570061 503183 570095 504169
rect 1685 464967 1719 483701
rect 1777 464355 1811 472073
rect 1869 467619 1903 474045
rect 1685 464321 1811 464355
rect 1409 447967 1443 449905
rect 1593 449055 1627 450721
rect 1593 448511 1627 448749
rect 1685 448715 1719 464321
rect 1961 462383 1995 474657
rect 569877 468537 569969 468571
rect 569877 461431 569911 468537
rect 569969 461703 570003 466565
rect 570061 465511 570095 467041
rect 570153 466871 570187 468265
rect 570245 466599 570279 467585
rect 570061 463607 570095 465205
rect 570153 462791 570187 465341
rect 570337 463879 570371 465477
rect 569877 461397 569969 461431
rect 1777 447831 1811 450041
rect 1777 441439 1811 442289
rect 1869 440963 1903 449157
rect 1961 439195 1995 454597
rect 570061 436815 570095 441609
rect 1961 425731 1995 434197
rect 569969 418183 570003 432497
rect 1961 407303 1995 414953
rect 1869 393975 1903 405569
rect 1961 393499 1995 405637
rect 569969 402271 570003 418013
rect 569969 393771 570003 399517
rect 569877 393737 570003 393771
rect 1409 381191 1443 387073
rect 1593 379151 1627 381429
rect 1685 379015 1719 380681
rect 1777 376771 1811 387345
rect 1869 380715 1903 387209
rect 1961 381463 1995 387073
rect 569877 382687 569911 393737
rect 569969 389895 570003 393669
rect 570061 392343 570095 396797
rect 570153 389079 570187 393805
rect 570245 388535 570279 394961
rect 570337 390031 570371 393125
rect 569969 376703 570003 382789
rect 570061 376567 570095 381837
rect 1409 358071 1443 369257
rect 1685 367795 1719 370481
rect 1777 358343 1811 370209
rect 1685 358309 1811 358343
rect 1685 345831 1719 358309
rect 1593 345797 1719 345831
rect 1409 333455 1443 334169
rect 1501 331891 1535 336005
rect 1225 304147 1259 312137
rect 1317 311831 1351 315129
rect 1501 312715 1535 326485
rect 1593 326383 1627 345797
rect 1685 329783 1719 345729
rect 1777 345695 1811 358241
rect 1869 358139 1903 370345
rect 1869 352971 1903 353209
rect 1777 335971 1811 340697
rect 1869 336039 1903 340833
rect 1961 340255 1995 370617
rect 569877 369393 569969 369427
rect 569877 358071 569911 369393
rect 569969 358139 570003 368305
rect 570061 358275 570095 359533
rect 569877 358037 570095 358071
rect 569877 357629 569969 357663
rect 569877 344879 569911 357629
rect 569969 353651 570003 353957
rect 569969 348959 570003 352597
rect 570061 352495 570095 358037
rect 570153 347735 570187 369733
rect 570245 357663 570279 376669
rect 570337 358071 570371 359873
rect 570245 348007 570279 352461
rect 570429 352359 570463 367761
rect 570521 353719 570555 359125
rect 569877 344845 569969 344879
rect 1777 335937 1903 335971
rect 1777 332027 1811 334033
rect 1409 312171 1443 312273
rect 1133 294491 1167 298061
rect 1225 293131 1259 303365
rect 1317 298095 1351 304521
rect 1409 304011 1443 312001
rect 1501 308431 1535 312409
rect 1593 311695 1627 318937
rect 1685 311559 1719 313905
rect 1777 312035 1811 331857
rect 1869 326519 1903 335937
rect 1961 329171 1995 338045
rect 569969 331279 570003 342193
rect 1869 313939 1903 326349
rect 569877 321011 569911 329545
rect 569969 321147 570003 331041
rect 570061 325023 570095 329681
rect 570153 321147 570187 330497
rect 570245 325703 570279 329409
rect 570337 327063 570371 329273
rect 569877 320977 570061 321011
rect 569877 320841 569969 320875
rect 1961 315027 1995 319141
rect 569877 315979 569911 320841
rect 570245 320807 570279 325533
rect 570061 320773 570279 320807
rect 569969 317951 570003 320705
rect 569877 315945 569969 315979
rect 570061 315911 570095 320773
rect 569877 315877 570095 315911
rect 1869 309655 1903 312545
rect 1961 309859 1995 312681
rect 1501 308397 1627 308431
rect 1317 292179 1351 296021
rect 1501 294627 1535 304385
rect 1593 296055 1627 308397
rect 1685 301495 1719 305609
rect 1777 303263 1811 305473
rect 1869 296259 1903 305337
rect 1317 284631 1351 287113
rect 1409 284767 1443 293369
rect 1501 287147 1535 294457
rect 1593 287079 1627 292145
rect 1501 287045 1627 287079
rect 1501 284359 1535 287045
rect 1409 283475 1443 283917
rect 1593 283271 1627 286977
rect 1685 283339 1719 295817
rect 1777 283407 1811 296089
rect 1869 283951 1903 295953
rect 1685 283305 1811 283339
rect 1685 270215 1719 273921
rect 1777 269807 1811 283305
rect 581 251855 615 266577
rect 1869 266543 1903 283441
rect 1961 269399 1995 306629
rect 569877 304351 569911 315877
rect 570003 315809 570095 315843
rect 569969 306187 570003 315605
rect 570061 309111 570095 315809
rect 570153 305031 570187 320705
rect 570245 315503 570279 320705
rect 570337 314755 570371 321113
rect 570521 309247 570555 314721
rect 569877 304317 570187 304351
rect 569877 304249 569969 304283
rect 569877 292791 569911 304249
rect 569969 300883 570003 301869
rect 570061 300271 570095 302889
rect 569969 298571 570003 300033
rect 570061 296599 570095 300101
rect 570153 296191 570187 304317
rect 570245 302923 570279 309145
rect 570245 298435 570279 302753
rect 570337 300407 570371 303841
rect 570429 301903 570463 306969
rect 569877 292757 569969 292791
rect 570153 292655 570187 296021
rect 569877 292621 570187 292655
rect 569877 285651 569911 292621
rect 569969 288303 570003 292553
rect 570153 289799 570187 291941
rect 569877 285617 569969 285651
rect 569969 285379 570003 285481
rect 569877 285345 570003 285379
rect 569877 274023 569911 285345
rect 569969 283747 570003 285141
rect 570061 283679 570095 289765
rect 570245 288167 570279 295137
rect 570337 291975 570371 296565
rect 570429 292451 570463 301121
rect 570521 296123 570555 304929
rect 569969 283645 570095 283679
rect 569969 274227 570003 283645
rect 570061 274295 570095 283577
rect 570153 274363 570187 285345
rect 570245 283611 570279 285617
rect 570061 274261 570187 274295
rect 569969 274193 570095 274227
rect 569877 273989 569969 274023
rect 570061 273955 570095 274193
rect 569877 273921 570095 273955
rect 1777 266509 1903 266543
rect 1777 264163 1811 266509
rect 857 251855 891 261545
rect 1133 242063 1167 261477
rect 1777 251855 1811 261477
rect 1501 238323 1535 250257
rect 305 199495 339 221017
rect 673 193987 707 201841
rect 857 199495 891 221697
rect 1501 221527 1535 238153
rect 1593 222615 1627 242097
rect 1685 237983 1719 242233
rect 1777 228395 1811 242165
rect 1869 242131 1903 266441
rect 1961 250155 1995 264673
rect 569877 245735 569911 273921
rect 569969 271575 570003 273037
rect 570061 269807 570095 273853
rect 570153 270487 570187 274261
rect 570245 270351 570279 283441
rect 570337 283407 570371 284937
rect 570337 270079 570371 274329
rect 570429 269943 570463 288133
rect 570521 283543 570555 289629
rect 570521 271031 570555 277253
rect 570613 272527 570647 284801
rect 570705 272935 570739 274465
rect 569969 259879 570003 267257
rect 569969 246007 570003 254745
rect 570061 250495 570095 266373
rect 1961 242947 1995 243049
rect 1869 222683 1903 241961
rect 1777 222649 1903 222683
rect 1317 212891 1351 221493
rect 1041 200923 1075 204901
rect 949 200889 1075 200923
rect 949 199427 983 200889
rect 857 199393 983 199427
rect 857 196231 891 199393
rect 1041 198883 1075 200821
rect 1133 197931 1167 207757
rect 949 195959 983 197625
rect 1133 194735 1167 197761
rect 1225 195075 1259 207689
rect 1317 197999 1351 209933
rect 1409 198067 1443 216801
rect 1593 207791 1627 219929
rect 1501 200855 1535 204697
rect 1317 197965 1443 197999
rect 1317 195823 1351 197897
rect 1409 193987 1443 197965
rect 1501 195211 1535 200685
rect 1593 198203 1627 198713
rect 213 165903 247 174573
rect 305 171003 339 182801
rect 489 170323 523 179197
rect 1225 176647 1259 188921
rect 1317 176511 1351 189193
rect 1409 176375 1443 189737
rect 1501 188547 1535 189601
rect 1501 176783 1535 188377
rect 1593 175967 1627 198033
rect 1685 197523 1719 221493
rect 1777 221323 1811 222649
rect 1777 217719 1811 218297
rect 1777 205751 1811 217413
rect 1869 205819 1903 222581
rect 1961 221527 1995 242505
rect 569877 230231 569911 245361
rect 569969 241111 570003 245701
rect 570061 243559 570095 246653
rect 570153 241179 570187 265897
rect 570245 259607 570279 263993
rect 570245 246551 570279 250937
rect 570245 243695 570279 245973
rect 570153 241145 570279 241179
rect 569969 241077 570187 241111
rect 569877 230197 569969 230231
rect 569877 229653 569969 229687
rect 1777 205717 1903 205751
rect 1685 182903 1719 195653
rect 1777 195279 1811 205649
rect 1869 200719 1903 205717
rect 1869 196095 1903 198169
rect 1961 198067 1995 221357
rect 569877 205003 569911 229653
rect 569969 205207 570003 228701
rect 570061 227035 570095 236045
rect 570153 229891 570187 241077
rect 570245 229755 570279 241145
rect 570337 228735 570371 247265
rect 570521 245395 570555 250597
rect 570061 205479 570095 226865
rect 570429 225879 570463 239445
rect 570521 229279 570555 233665
rect 570245 225845 570463 225879
rect 569877 204969 570095 205003
rect 569969 202623 570003 204901
rect 570061 204799 570095 204969
rect 570061 203167 570095 203677
rect 570153 203031 570187 214557
rect 570245 205547 570279 225845
rect 570337 214659 570371 225777
rect 570245 205513 570371 205547
rect 570245 204459 570279 205445
rect 570337 203575 570371 205513
rect 1961 196367 1995 197625
rect 1777 195245 1995 195279
rect 1777 179095 1811 195177
rect 1869 186507 1903 195109
rect 305 145639 339 167773
rect 397 146999 431 153833
rect 673 146183 707 153901
rect 765 146999 799 159613
rect 857 159307 891 166889
rect 949 154819 983 167637
rect 1041 159171 1075 167365
rect 949 150127 983 154037
rect 1133 153867 1167 166141
rect 1225 153935 1259 167637
rect 1317 159443 1351 167229
rect 1409 165495 1443 166413
rect 1501 163659 1535 175593
rect 1685 173043 1719 176953
rect 1777 176239 1811 178381
rect 1869 176171 1903 179605
rect 1961 179231 1995 195245
rect 1961 176239 1995 177633
rect 569969 177463 570003 192457
rect 570061 188411 570095 192185
rect 569877 177293 569969 177327
rect 1777 176137 1903 176171
rect 1409 163625 1535 163659
rect 1409 159375 1443 163625
rect 1501 159511 1535 163557
rect 1593 163455 1627 167977
rect 1133 153833 1351 153867
rect 581 141627 615 142953
rect 305 130271 339 138941
rect 489 129455 523 130373
rect 581 109327 615 130577
rect 673 126259 707 132073
rect 765 130407 799 141185
rect 857 140743 891 146285
rect 949 142851 983 146965
rect 1041 141151 1075 150229
rect 1225 146999 1259 153765
rect 1317 146319 1351 153833
rect 857 140709 983 140743
rect 673 117419 707 126021
rect 765 117487 799 130237
rect 857 126123 891 140641
rect 949 139111 983 140709
rect 1133 138907 1167 145673
rect 949 134623 983 138737
rect 949 134589 1075 134623
rect 949 128367 983 134521
rect 1041 126667 1075 134589
rect 949 117419 983 126225
rect 1041 119595 1075 126497
rect 673 117385 891 117419
rect 673 109191 707 109429
rect 765 108783 799 109701
rect 857 107695 891 117385
rect 1041 115243 1075 117453
rect 949 108919 983 115073
rect 1041 108103 1075 110993
rect 1133 96067 1167 138669
rect 1225 108375 1259 134453
rect 1317 107219 1351 146149
rect 1409 141423 1443 159205
rect 1501 150263 1535 156349
rect 1501 141491 1535 150093
rect 1593 148767 1627 163285
rect 1685 159647 1719 167229
rect 1777 159579 1811 176137
rect 1869 163591 1903 176069
rect 1961 163523 1995 169065
rect 1869 163489 1995 163523
rect 569877 163523 569911 177293
rect 570061 176851 570095 180421
rect 570153 179843 570187 193885
rect 569969 163727 570003 174913
rect 569877 163489 569969 163523
rect 1685 148699 1719 159477
rect 1593 148665 1719 148699
rect 1593 145979 1627 148665
rect 1409 141389 1627 141423
rect 1409 138771 1443 141253
rect 949 86139 983 92021
rect 1041 90423 1075 94673
rect 1133 91647 1167 93993
rect 1225 91783 1259 93585
rect 1317 93551 1351 98277
rect 1317 91511 1351 93381
rect 1409 91375 1443 138601
rect 1501 137955 1535 141321
rect 1501 126259 1535 134589
rect 1593 131155 1627 141389
rect 1685 134623 1719 148597
rect 1777 146387 1811 159409
rect 1869 159239 1903 163489
rect 1869 146931 1903 159069
rect 1961 146999 1995 163421
rect 569877 158729 569969 158763
rect 569877 158015 569911 158729
rect 569877 157981 569969 158015
rect 569969 149311 570003 157845
rect 1869 146897 1995 146931
rect 1777 140743 1811 146217
rect 1869 143123 1903 145877
rect 1777 138975 1811 139961
rect 1777 138295 1811 138805
rect 1685 134589 1811 134623
rect 1593 129183 1627 130849
rect 1593 126531 1627 128877
rect 1501 116467 1535 126089
rect 1501 108511 1535 115209
rect 1593 108647 1627 126361
rect 1685 124899 1719 134521
rect 1777 134419 1811 134589
rect 1777 124763 1811 133433
rect 1869 133331 1903 142953
rect 1961 131155 1995 146897
rect 569969 134555 570003 148325
rect 570061 134215 570095 169065
rect 570153 161959 570187 178041
rect 570245 178007 570279 191913
rect 570337 178075 570371 192049
rect 570429 191539 570463 192729
rect 570245 177973 570371 178007
rect 570245 162027 570279 175185
rect 570153 161925 570279 161959
rect 570153 147679 570187 157981
rect 570245 153459 570279 161925
rect 570337 158763 570371 177973
rect 570429 162231 570463 171921
rect 570521 169099 570555 177429
rect 570337 155703 570371 157369
rect 570337 155669 570463 155703
rect 570337 153935 570371 155601
rect 570429 153391 570463 155669
rect 570521 155023 570555 157641
rect 570245 153357 570463 153391
rect 570245 147951 570279 153357
rect 570337 133127 570371 148461
rect 570521 146999 570555 149549
rect 1869 131121 1995 131155
rect 1869 124967 1903 131121
rect 1961 124967 1995 131053
rect 1685 108103 1719 124729
rect 1777 102595 1811 119561
rect 949 82127 983 84745
rect 1041 83623 1075 87601
rect 1133 70431 1167 84609
rect 1225 80699 1259 88757
rect 1317 80767 1351 83793
rect 765 64651 799 66725
rect 857 57919 891 66589
rect 949 63155 983 67201
rect 1041 62883 1075 67473
rect 1133 62271 1167 65433
rect 1225 62747 1259 69581
rect 1225 55879 1259 57069
rect 1317 52751 1351 70261
rect 1409 69479 1443 90389
rect 1501 87635 1535 93517
rect 1501 80835 1535 87329
rect 1409 63019 1443 69309
rect 1501 66963 1535 80665
rect 1593 72335 1627 96033
rect 1685 87363 1719 98277
rect 1777 91239 1811 98413
rect 1869 96271 1903 117793
rect 1961 107083 1995 117997
rect 1869 93279 1903 94741
rect 1685 80971 1719 86309
rect 1593 66283 1627 71961
rect 1685 69615 1719 80801
rect 1777 72403 1811 86173
rect 1869 72471 1903 93109
rect 1961 88791 1995 98141
rect 1777 72369 1903 72403
rect 1685 66351 1719 69445
rect 1501 66249 1627 66283
rect 1409 55199 1443 56729
rect 1501 52615 1535 66249
rect 1593 64243 1627 65433
rect 1685 64787 1719 65841
rect 1593 64209 1719 64243
rect 29 35003 63 50405
rect 1041 37043 1075 50337
rect 1593 45543 1627 62713
rect 1409 43095 1443 45509
rect 1685 43571 1719 64209
rect 1777 47651 1811 72301
rect 1869 65467 1903 72369
rect 1961 66487 1995 86377
rect 569877 76313 569969 76347
rect 1869 50439 1903 64753
rect 1961 47719 1995 66317
rect 569877 58871 569911 76313
rect 569969 56967 570003 75905
rect 570061 53771 570095 77265
rect 570153 56695 570187 76721
rect 570245 75939 570279 76585
rect 570337 75871 570371 76177
rect 570245 75837 570371 75871
rect 570245 59959 570279 75837
rect 570337 72471 570371 74817
rect 570429 73015 570463 73593
rect 570337 60775 570371 68017
rect 570521 66147 570555 73389
rect 570429 58735 570463 64957
rect 570521 56627 570555 65977
rect 1869 47685 1995 47719
rect 1593 43537 1719 43571
rect 1593 42823 1627 43537
rect 121 16983 155 24225
rect 581 15487 615 24021
rect 673 22083 707 33541
rect 1041 29563 1075 35377
rect 1133 29631 1167 39457
rect 949 23783 983 28849
rect 1225 27319 1259 35513
rect 1133 27285 1259 27319
rect 489 323 523 8653
rect 581 1751 615 10353
rect 673 10115 707 16541
rect 765 12087 799 18445
rect 765 3723 799 10421
rect 857 10319 891 17085
rect 949 7531 983 20009
rect 1041 18615 1075 27081
rect 1041 14603 1075 17901
rect 1133 15215 1167 27285
rect 1225 15351 1259 27217
rect 1317 21199 1351 35649
rect 1409 29019 1443 39321
rect 1409 22219 1443 28305
rect 1501 27115 1535 29461
rect 1317 21165 1443 21199
rect 1133 14535 1167 14773
rect 1041 14501 1167 14535
rect 1041 13379 1075 14501
rect 1041 1683 1075 10353
rect 1133 1343 1167 14433
rect 1225 3315 1259 13481
rect 1317 12359 1351 16405
rect 1409 12767 1443 21165
rect 1501 16099 1535 21573
rect 1593 18411 1627 29665
rect 1501 14671 1535 15929
rect 1409 12733 1535 12767
rect 1317 1547 1351 11849
rect 1409 10523 1443 12325
rect 1409 1071 1443 10353
rect 1501 391 1535 12733
rect 1593 10455 1627 18241
rect 1685 17119 1719 43469
rect 1777 39219 1811 47481
rect 1869 43435 1903 47685
rect 1961 43503 1995 47617
rect 1869 43401 1995 43435
rect 1869 29699 1903 39321
rect 1961 29903 1995 43401
rect 569877 42313 569969 42347
rect 1777 29665 1903 29699
rect 1777 20043 1811 29665
rect 1869 20111 1903 29597
rect 1777 20009 1903 20043
rect 1685 10387 1719 16949
rect 1777 12359 1811 19941
rect 1593 1207 1627 10285
rect 1685 1139 1719 10217
rect 1777 51 1811 12189
rect 1869 3723 1903 20009
rect 1961 18887 1995 29733
rect 1961 9435 1995 18717
rect 569877 18139 569911 42313
rect 569969 39695 570003 40953
rect 570061 39423 570095 41633
rect 570153 39899 570187 41089
rect 569969 23103 570003 27897
rect 569877 18105 570003 18139
rect 1961 1615 1995 8721
rect 569969 8143 570003 18105
rect 570061 14739 570095 25721
rect 570153 23239 570187 39729
rect 570245 27931 570279 42177
rect 570337 39763 570371 41769
rect 570429 40035 570463 40409
rect 570521 39083 570555 43265
rect 570613 34799 570647 40273
rect 570245 23783 570279 26469
rect 570153 17663 570187 23069
rect 570337 7871 570371 31025
rect 570429 24191 570463 25517
rect 124321 3043 124355 3077
rect 125609 3077 126839 3111
rect 177991 3077 179187 3111
rect 125609 3043 125643 3077
rect 124321 3009 125827 3043
rect 125609 2771 125643 3009
rect 122665 2737 125643 2771
rect 106289 1989 112855 2023
rect 3525 1853 6135 1887
rect 3525 1479 3559 1853
rect 5089 1785 5491 1819
rect 3709 1683 3743 1717
rect 3709 1649 4169 1683
rect 5089 1547 5123 1785
rect 5457 1683 5491 1785
rect 5549 1683 5583 1785
rect 5273 1615 5307 1649
rect 5273 1581 5583 1615
rect 3467 1445 3559 1479
rect 5181 1411 5215 1513
rect 5399 1445 5457 1479
rect 5123 1241 5273 1275
rect 5215 1173 5365 1207
rect 5273 731 5307 1037
rect 5549 867 5583 1581
rect 5641 1411 5675 1785
rect 5549 833 5641 867
rect 5365 663 5399 697
rect 5123 629 5399 663
rect 4721 561 5181 595
rect 4721 459 4755 561
rect 6101 527 6135 1853
rect 87153 1853 92983 1887
rect 10149 1479 10183 1649
rect 10149 1445 10609 1479
rect 6929 1207 6963 1445
rect 7297 663 7331 1377
rect 10425 1139 10459 1241
rect 10517 1139 10551 1377
rect 11161 1275 11195 1581
rect 11069 1207 11103 1241
rect 11253 1207 11287 1581
rect 12909 1343 12943 1445
rect 12909 1309 13185 1343
rect 11069 1173 11287 1207
rect 25145 1207 25179 1649
rect 25789 867 25823 1649
rect 25973 1003 26007 1377
rect 26249 1343 26283 1717
rect 26985 1683 27019 1785
rect 27077 1411 27111 1649
rect 25881 867 25915 969
rect 19383 765 19441 799
rect 5089 459 5123 493
rect 5089 425 5457 459
rect 5549 425 5859 459
rect 5549 391 5583 425
rect 5825 391 5859 425
rect 5399 357 5583 391
rect 5273 51 5307 289
rect 5733 255 5767 357
rect 5675 221 5767 255
rect 6009 255 6043 493
rect 9689 323 9723 561
rect 10241 323 10275 425
rect 10425 391 10459 561
rect 10241 289 10643 323
rect 5399 153 5549 187
rect 9781 119 9815 289
rect 5491 85 5641 119
rect 10517 119 10551 221
rect 10609 119 10643 289
rect 6009 51 6043 85
rect 5273 17 6043 51
rect 13185 51 13219 697
rect 14289 391 14323 561
rect 14473 51 14507 357
rect 26801 323 26835 1377
rect 28273 1275 28307 1513
rect 34345 1139 34379 1309
rect 28181 187 28215 833
rect 34989 323 35023 1717
rect 35081 1411 35115 1649
rect 35265 1547 35299 1785
rect 35357 1003 35391 1717
rect 34989 289 35265 323
rect 38025 187 38059 1649
rect 38301 867 38335 969
rect 38393 867 38427 1105
rect 38117 187 38151 765
rect 38669 255 38703 357
rect 39037 323 39071 1377
rect 39129 1343 39163 1649
rect 39221 1377 39405 1411
rect 39221 1207 39255 1377
rect 39497 799 39531 1241
rect 39589 663 39623 1785
rect 39313 391 39347 629
rect 39221 119 39255 357
rect 39681 187 39715 1785
rect 48697 1785 48973 1819
rect 48697 1751 48731 1785
rect 48789 1717 49065 1751
rect 50847 1717 50997 1751
rect 42441 867 42475 1581
rect 42901 799 42935 1581
rect 48789 1547 48823 1717
rect 56793 1683 56827 1785
rect 48973 1649 49191 1683
rect 48973 1615 49007 1649
rect 49065 1547 49099 1581
rect 48915 1513 49099 1547
rect 48881 1275 48915 1377
rect 49065 1207 49099 1445
rect 49157 1411 49191 1649
rect 49157 799 49191 1173
rect 49709 663 49743 765
rect 49249 323 49283 561
rect 39773 187 39807 289
rect 39865 119 39899 289
rect 49801 187 49835 629
rect 53297 255 53331 1377
rect 55781 935 55815 1649
rect 56609 1547 56643 1649
rect 56609 1513 56701 1547
rect 58081 1513 58265 1547
rect 58081 1343 58115 1513
rect 55781 901 56885 935
rect 39221 85 39899 119
rect 55321 119 55355 765
rect 57989 187 58023 901
rect 58173 255 58207 1445
rect 60749 1445 60933 1479
rect 59093 323 59127 1309
rect 58265 187 58299 221
rect 57989 153 58299 187
rect 60749 187 60783 1445
rect 62129 1343 62163 1445
rect 61301 935 61335 1309
rect 63233 1275 63267 1649
rect 63325 1343 63359 1649
rect 65441 1411 65475 1785
rect 65533 1479 65567 1785
rect 74641 1717 78723 1751
rect 71789 1649 71881 1683
rect 66821 1581 67131 1615
rect 66821 1547 66855 1581
rect 66729 1513 66855 1547
rect 66729 1479 66763 1513
rect 65625 1411 65659 1445
rect 65441 1377 65659 1411
rect 63417 1275 63451 1309
rect 63233 1241 63451 1275
rect 66821 1207 66855 1445
rect 67005 1343 67039 1513
rect 67097 1343 67131 1581
rect 71789 1411 71823 1649
rect 72525 1377 72927 1411
rect 63325 935 63359 1173
rect 63509 1139 63543 1173
rect 63509 1105 63819 1139
rect 63785 867 63819 1105
rect 67373 1037 68937 1071
rect 64981 867 65015 901
rect 63543 833 63635 867
rect 60841 187 60875 289
rect 63601 255 63635 833
rect 63785 833 65015 867
rect 63509 187 63543 221
rect 63693 187 63727 833
rect 67373 255 67407 1037
rect 68845 969 69523 1003
rect 68845 935 68879 969
rect 69489 935 69523 969
rect 67315 221 67407 255
rect 63509 153 63727 187
rect 69397 187 69431 901
rect 70593 119 70627 901
rect 72525 187 72559 1377
rect 72893 1343 72927 1377
rect 72801 1139 72835 1309
rect 73019 1173 73169 1207
rect 72801 1105 73111 1139
rect 73077 1071 73111 1105
rect 72985 935 73019 1037
rect 72835 833 73111 867
rect 73077 323 73111 833
rect 73169 697 73387 731
rect 73169 663 73203 697
rect 72985 255 73019 289
rect 72985 221 73111 255
rect 73077 187 73111 221
rect 73261 187 73295 629
rect 73353 527 73387 697
rect 74641 459 74675 1717
rect 76205 1513 76423 1547
rect 74825 1343 74859 1377
rect 74825 1309 75009 1343
rect 76205 1207 76239 1513
rect 76389 1479 76423 1513
rect 78689 1479 78723 1717
rect 87153 1683 87187 1853
rect 92949 1751 92983 1853
rect 101413 1853 106139 1887
rect 92949 1717 93351 1751
rect 82645 1649 87187 1683
rect 82645 1479 82679 1649
rect 83933 1581 87095 1615
rect 82863 1513 83473 1547
rect 81541 1445 81943 1479
rect 83231 1445 83381 1479
rect 76297 1207 76331 1445
rect 78815 1377 81449 1411
rect 81541 1343 81575 1445
rect 75469 969 76055 1003
rect 75469 935 75503 969
rect 75561 663 75595 901
rect 76021 867 76055 969
rect 75929 663 75963 833
rect 76573 799 76607 901
rect 76757 867 76791 1309
rect 78689 1309 81575 1343
rect 78689 1275 78723 1309
rect 78965 799 78999 1105
rect 75837 595 75871 629
rect 76665 595 76699 765
rect 75837 561 76699 595
rect 73537 425 74675 459
rect 73537 255 73571 425
rect 73939 357 74365 391
rect 73077 153 73295 187
rect 73445 187 73479 221
rect 73721 187 73755 221
rect 76573 187 76607 357
rect 73445 153 73755 187
rect 72617 119 72651 153
rect 70593 85 72651 119
rect 76481 119 76515 153
rect 76665 119 76699 357
rect 76481 85 76699 119
rect 81725 51 81759 1377
rect 81909 119 81943 1445
rect 82737 1139 82771 1445
rect 83231 1309 83381 1343
rect 83105 1275 83139 1309
rect 83105 1241 83415 1275
rect 82863 1173 83013 1207
rect 83013 1105 83289 1139
rect 82829 663 82863 969
rect 82921 731 82955 901
rect 83013 799 83047 1105
rect 83105 731 83139 901
rect 83381 867 83415 1241
rect 83565 1071 83599 1309
rect 83473 1037 83599 1071
rect 83473 1003 83507 1037
rect 83565 731 83599 969
rect 82921 697 83139 731
rect 83197 697 83599 731
rect 83197 663 83231 697
rect 82277 595 82311 629
rect 82829 629 83231 663
rect 82737 595 82771 629
rect 82277 561 82771 595
rect 83933 187 83967 1581
rect 85957 1513 86451 1547
rect 83415 153 83967 187
rect 84025 1445 85807 1479
rect 84025 119 84059 1445
rect 84117 867 84151 1377
rect 81909 85 84059 119
rect 84209 51 84243 1377
rect 85773 1343 85807 1445
rect 85957 1411 85991 1513
rect 85773 1309 85991 1343
rect 85957 1275 85991 1309
rect 86049 1275 86083 1377
rect 84577 1241 85715 1275
rect 85957 1241 86083 1275
rect 84577 187 84611 1241
rect 84853 867 84887 1173
rect 81725 17 84243 51
rect 84393 51 84427 153
rect 85681 119 85715 1241
rect 85773 731 85807 1173
rect 86417 867 86451 1513
rect 87061 1343 87095 1581
rect 87429 1581 93259 1615
rect 87429 1411 87463 1581
rect 87521 1411 87555 1513
rect 87613 1513 93167 1547
rect 87613 1343 87647 1513
rect 87705 1275 87739 1445
rect 87429 1241 87739 1275
rect 87797 1445 92765 1479
rect 85865 799 85899 833
rect 87429 799 87463 1241
rect 87797 867 87831 1445
rect 91879 1377 92431 1411
rect 92615 1377 93041 1411
rect 92397 1343 92431 1377
rect 87889 1309 92063 1343
rect 93133 1343 93167 1513
rect 87889 1207 87923 1309
rect 90925 1241 91787 1275
rect 85865 765 87463 799
rect 85773 697 87647 731
rect 87613 255 87647 697
rect 87613 221 87831 255
rect 87797 187 87831 221
rect 89637 119 89671 357
rect 85681 85 89671 119
rect 90925 51 90959 1241
rect 91753 1207 91787 1241
rect 91845 1207 91879 1241
rect 91845 1173 91971 1207
rect 91661 731 91695 1173
rect 91937 1071 91971 1173
rect 92029 1139 92063 1309
rect 92155 1173 93167 1207
rect 92029 1105 92305 1139
rect 92029 1037 92247 1071
rect 91845 1003 91879 1037
rect 92029 1003 92063 1037
rect 91845 969 92063 1003
rect 92213 1003 92247 1037
rect 92673 1003 92707 1105
rect 92213 969 92523 1003
rect 92673 969 93075 1003
rect 92489 935 92523 969
rect 92489 901 92983 935
rect 92949 799 92983 901
rect 92615 765 92799 799
rect 91569 187 91603 697
rect 92155 629 92489 663
rect 92765 391 92799 765
rect 93041 391 93075 969
rect 93133 799 93167 1173
rect 93225 1139 93259 1581
rect 93317 1207 93351 1717
rect 101413 1547 101447 1853
rect 106105 1819 106139 1853
rect 93409 1513 96755 1547
rect 101505 1717 102459 1751
rect 93409 1139 93443 1513
rect 96721 1411 96755 1513
rect 101505 1479 101539 1717
rect 102425 1683 102459 1717
rect 101597 1649 102275 1683
rect 102425 1649 103839 1683
rect 101597 1479 101631 1649
rect 102241 1615 102275 1649
rect 101689 1581 102183 1615
rect 102241 1581 103747 1615
rect 101689 1411 101723 1581
rect 102149 1411 102183 1581
rect 102333 1411 102367 1445
rect 96721 1377 101723 1411
rect 101781 1377 102057 1411
rect 102149 1377 102367 1411
rect 101781 1343 101815 1377
rect 102425 1343 102459 1513
rect 93317 1105 93443 1139
rect 96629 1309 101815 1343
rect 101907 1309 102091 1343
rect 102275 1309 102459 1343
rect 102517 1513 103437 1547
rect 93317 595 93351 1105
rect 96629 1071 96663 1309
rect 102057 1275 102091 1309
rect 93409 1037 96663 1071
rect 97457 1241 100401 1275
rect 100711 1241 100769 1275
rect 102149 1241 102425 1275
rect 93409 867 93443 1037
rect 96353 901 97365 935
rect 96353 867 96387 901
rect 97457 867 97491 1241
rect 102149 1207 102183 1241
rect 97031 833 97491 867
rect 97549 1173 102183 1207
rect 93961 799 93995 833
rect 96445 799 96479 833
rect 97549 799 97583 1173
rect 93961 765 96479 799
rect 96537 765 97583 799
rect 97641 1105 100987 1139
rect 96537 595 96571 765
rect 93317 561 93409 595
rect 94179 561 96571 595
rect 97365 527 97399 697
rect 93259 493 94329 527
rect 94421 493 96847 527
rect 92765 357 92857 391
rect 93041 357 94329 391
rect 92673 323 92707 357
rect 94421 323 94455 493
rect 92673 289 94455 323
rect 95709 323 95743 425
rect 95801 425 96721 459
rect 95801 391 95835 425
rect 96813 391 96847 493
rect 97457 459 97491 697
rect 97215 425 97491 459
rect 97641 391 97675 1105
rect 100953 1071 100987 1105
rect 100861 799 100895 1037
rect 102517 1003 102551 1513
rect 102701 1377 103655 1411
rect 102701 1275 102735 1377
rect 102793 1309 103471 1343
rect 101873 969 102551 1003
rect 101873 935 101907 969
rect 102793 935 102827 1309
rect 103287 1241 103379 1275
rect 100619 765 100803 799
rect 101045 799 101079 901
rect 101137 901 101321 935
rect 102333 901 102827 935
rect 101137 867 101171 901
rect 101229 799 101263 833
rect 101045 765 101263 799
rect 102149 765 102241 799
rect 100769 731 100803 765
rect 102149 731 102183 765
rect 96813 357 97675 391
rect 97733 697 98503 731
rect 97733 323 97767 697
rect 95709 289 97767 323
rect 97825 629 98319 663
rect 97825 255 97859 629
rect 98285 595 98319 629
rect 92581 221 97859 255
rect 92581 187 92615 221
rect 91661 153 92615 187
rect 91477 119 91511 153
rect 91661 119 91695 153
rect 91477 85 91695 119
rect 84393 17 90959 51
rect 92121 51 92155 85
rect 92489 51 92523 85
rect 92121 17 92523 51
rect 98193 51 98227 561
rect 98469 323 98503 697
rect 100125 391 100159 697
rect 100493 595 100527 697
rect 100309 561 100527 595
rect 100769 697 102183 731
rect 102333 731 102367 901
rect 102885 799 102919 901
rect 102517 765 102919 799
rect 100309 527 100343 561
rect 100677 527 100711 697
rect 102241 629 102459 663
rect 102241 459 102275 629
rect 102425 595 102459 629
rect 102333 527 102367 561
rect 102517 527 102551 765
rect 103345 731 103379 1241
rect 103437 799 103471 1309
rect 103529 867 103563 1105
rect 103621 1071 103655 1377
rect 103713 1139 103747 1581
rect 103805 1547 103839 1649
rect 104357 1139 104391 1513
rect 104541 1207 104575 1513
rect 106013 1411 106047 1785
rect 105921 1139 105955 1377
rect 106289 1207 106323 1989
rect 108405 1921 112027 1955
rect 108405 1887 108439 1921
rect 111993 1887 112027 1921
rect 106381 1853 108439 1887
rect 110061 1853 111935 1887
rect 111993 1853 112487 1887
rect 103805 1105 104081 1139
rect 104357 1105 104909 1139
rect 103805 1071 103839 1105
rect 103621 1037 103839 1071
rect 106381 867 106415 1853
rect 106875 1785 110003 1819
rect 106841 1717 107025 1751
rect 106841 1479 106875 1717
rect 109969 1411 110003 1785
rect 110061 867 110095 1853
rect 111901 1819 111935 1853
rect 106599 833 107301 867
rect 107577 833 109175 867
rect 109359 833 110095 867
rect 110153 1785 111751 1819
rect 107577 799 107611 833
rect 109141 799 109175 833
rect 110153 799 110187 1785
rect 103437 765 107611 799
rect 109141 765 110187 799
rect 110245 1649 110555 1683
rect 109049 731 109083 765
rect 110245 731 110279 1649
rect 110521 1615 110555 1649
rect 111073 1649 111567 1683
rect 110521 1581 111015 1615
rect 102643 697 103287 731
rect 103345 697 109083 731
rect 109141 697 110279 731
rect 103253 595 103287 697
rect 109141 663 109175 697
rect 103345 629 109175 663
rect 103345 595 103379 629
rect 102333 493 102551 527
rect 102609 561 103161 595
rect 103253 561 103379 595
rect 100953 425 102275 459
rect 100953 391 100987 425
rect 102609 391 102643 561
rect 100125 357 100987 391
rect 101045 357 102643 391
rect 101045 323 101079 357
rect 98469 289 101079 323
rect 106841 289 107025 323
rect 106841 255 106875 289
rect 110705 119 110739 1445
rect 110797 867 110831 1445
rect 110889 595 110923 833
rect 110981 595 111015 1581
rect 111073 1479 111107 1649
rect 111165 799 111199 1377
rect 111257 1275 111291 1581
rect 111073 731 111107 765
rect 111349 731 111383 1377
rect 111441 1139 111475 1581
rect 111533 1411 111567 1649
rect 111625 1479 111659 1717
rect 111717 1547 111751 1785
rect 111809 1785 111935 1819
rect 112453 1819 112487 1853
rect 112453 1785 112671 1819
rect 111809 1615 111843 1785
rect 111901 1581 112361 1615
rect 111901 1547 111935 1581
rect 111717 1513 111935 1547
rect 111993 1513 112303 1547
rect 111993 1479 112027 1513
rect 111625 1445 112027 1479
rect 111809 1309 112119 1343
rect 111809 1275 111843 1309
rect 112085 1207 112119 1309
rect 111993 1139 112027 1173
rect 111441 1105 112027 1139
rect 111843 1037 112085 1071
rect 112269 867 112303 1513
rect 111843 833 111935 867
rect 112269 833 112545 867
rect 111901 799 111935 833
rect 112637 799 112671 1785
rect 112821 1547 112855 1989
rect 115857 1921 116351 1955
rect 115155 1581 115339 1615
rect 112821 1513 115247 1547
rect 114845 867 114879 1445
rect 114937 1275 114971 1445
rect 114753 799 114787 833
rect 115029 799 115063 1241
rect 115213 1071 115247 1513
rect 115305 1411 115339 1581
rect 115857 1139 115891 1921
rect 116317 1887 116351 1921
rect 115949 1853 116259 1887
rect 116317 1853 122423 1887
rect 115949 1071 115983 1853
rect 116225 1819 116259 1853
rect 116317 1785 122331 1819
rect 116133 1343 116167 1785
rect 116317 1479 116351 1785
rect 116225 1445 116351 1479
rect 116409 1717 121561 1751
rect 116225 1411 116259 1445
rect 116317 1343 116351 1377
rect 116133 1309 116351 1343
rect 116409 1139 116443 1717
rect 121411 1649 121503 1683
rect 116133 1105 116443 1139
rect 116133 1071 116167 1105
rect 116501 1071 116535 1581
rect 116593 1207 116627 1581
rect 116961 1513 120123 1547
rect 116685 1207 116719 1241
rect 116685 1173 116869 1207
rect 115213 1037 115983 1071
rect 116041 1037 116167 1071
rect 116041 935 116075 1037
rect 111751 765 111843 799
rect 111901 765 111993 799
rect 112637 765 112913 799
rect 114753 765 115063 799
rect 115213 901 116075 935
rect 111073 697 111383 731
rect 111809 731 111843 765
rect 115213 731 115247 901
rect 116133 867 116167 969
rect 116409 935 116443 1037
rect 116409 901 116685 935
rect 116961 867 116995 1513
rect 120089 1479 120123 1513
rect 120089 1445 120583 1479
rect 117053 1377 120457 1411
rect 117053 935 117087 1377
rect 119445 1241 119663 1275
rect 119445 1207 119479 1241
rect 119261 1139 119295 1173
rect 119537 1139 119571 1173
rect 119261 1105 119571 1139
rect 119629 1139 119663 1241
rect 120549 1207 120583 1445
rect 120951 1377 121319 1411
rect 121009 1309 121227 1343
rect 121009 1275 121043 1309
rect 120549 1173 121043 1207
rect 119629 1105 120859 1139
rect 116133 833 116995 867
rect 111809 697 115247 731
rect 111441 629 111717 663
rect 112211 629 113223 663
rect 111441 595 111475 629
rect 112027 493 112177 527
rect 111843 425 112269 459
rect 111809 357 112395 391
rect 111809 187 111843 357
rect 112027 289 112303 323
rect 112269 255 112303 289
rect 112361 187 112395 357
rect 111901 119 111935 153
rect 112453 119 112487 561
rect 110705 85 111935 119
rect 111993 85 112487 119
rect 111993 51 112027 85
rect 98193 17 112027 51
rect 113189 51 113223 629
rect 120181 51 120215 969
rect 120733 187 120767 765
rect 120825 255 120859 1105
rect 121009 323 121043 1173
rect 121101 391 121135 1241
rect 121193 867 121227 1309
rect 121285 1071 121319 1377
rect 121469 1003 121503 1649
rect 121929 1003 121963 1377
rect 122113 1275 122147 1445
rect 122297 1411 122331 1785
rect 122389 1207 122423 1853
rect 122665 1479 122699 2737
rect 125793 2567 125827 3009
rect 124873 2533 125919 2567
rect 124413 1649 124689 1683
rect 122021 1173 122423 1207
rect 121377 935 121411 969
rect 121377 901 121503 935
rect 121193 833 121377 867
rect 121469 799 121503 901
rect 121285 731 121319 765
rect 121285 697 121595 731
rect 121561 663 121595 697
rect 121469 459 121503 629
rect 121837 527 121871 969
rect 122021 595 122055 1173
rect 123677 1105 123895 1139
rect 123033 1003 123067 1037
rect 123677 1003 123711 1105
rect 123033 969 123711 1003
rect 123861 1003 123895 1105
rect 123861 969 124045 1003
rect 124229 969 124321 1003
rect 122389 935 122423 969
rect 122389 901 122665 935
rect 124229 867 124263 969
rect 122113 833 124263 867
rect 122113 663 122147 833
rect 124413 595 124447 1649
rect 124873 799 124907 2533
rect 125793 2227 125827 2533
rect 125241 2193 125827 2227
rect 125241 1207 125275 2193
rect 125885 2159 125919 2533
rect 126805 2363 126839 3077
rect 142169 2465 147447 2499
rect 142169 2431 142203 2465
rect 132509 2397 142203 2431
rect 147413 2431 147447 2465
rect 147413 2397 156187 2431
rect 132509 2363 132543 2397
rect 126805 2329 132543 2363
rect 156153 2363 156187 2397
rect 156153 2329 160235 2363
rect 160201 2295 160235 2329
rect 156153 2261 157475 2295
rect 129749 2193 129967 2227
rect 129749 2159 129783 2193
rect 125885 2125 129783 2159
rect 129933 2159 129967 2193
rect 129933 2125 139167 2159
rect 128093 2057 129783 2091
rect 125333 1921 126379 1955
rect 125333 1615 125367 1921
rect 126345 1887 126379 1921
rect 125425 1853 126287 1887
rect 126345 1853 127575 1887
rect 125425 1275 125459 1853
rect 125609 1683 125643 1785
rect 125701 1615 125735 1785
rect 126253 1683 126287 1853
rect 125885 1649 126195 1683
rect 126253 1649 127483 1683
rect 125885 1479 125919 1649
rect 125517 1275 125551 1445
rect 125609 1207 125643 1445
rect 125241 1173 125643 1207
rect 125977 1207 126011 1581
rect 126069 1275 126103 1581
rect 126161 1411 126195 1649
rect 127449 1615 127483 1649
rect 127357 1479 127391 1581
rect 127541 1547 127575 1853
rect 128093 1751 128127 2057
rect 129749 2023 129783 2057
rect 139133 2023 139167 2125
rect 147873 2125 154531 2159
rect 129749 1989 134567 2023
rect 139133 1989 143767 2023
rect 134533 1955 134567 1989
rect 128185 1921 134475 1955
rect 134533 1921 138891 1955
rect 128185 1683 128219 1921
rect 134441 1887 134475 1921
rect 128461 1853 134383 1887
rect 134441 1853 138799 1887
rect 128461 1819 128495 1853
rect 134349 1819 134383 1853
rect 130301 1785 130485 1819
rect 134441 1785 134625 1819
rect 130301 1751 130335 1785
rect 128093 1649 128219 1683
rect 128093 1615 128127 1649
rect 128185 1547 128219 1581
rect 127541 1513 128219 1547
rect 127357 1445 128093 1479
rect 128277 1411 128311 1717
rect 128369 1717 129231 1751
rect 128369 1479 128403 1717
rect 128645 1479 128679 1649
rect 129197 1547 129231 1717
rect 129381 1717 129565 1751
rect 134257 1751 134291 1785
rect 134441 1751 134475 1785
rect 138765 1751 138799 1853
rect 138857 1819 138891 1921
rect 139133 1921 141835 1955
rect 139133 1819 139167 1921
rect 138857 1785 139167 1819
rect 140605 1785 141743 1819
rect 134257 1717 134383 1751
rect 134717 1717 138615 1751
rect 138765 1717 140513 1751
rect 129381 1683 129415 1717
rect 134349 1683 134383 1717
rect 134349 1649 134625 1683
rect 129197 1513 132819 1547
rect 129323 1445 129749 1479
rect 131773 1445 132727 1479
rect 126161 1377 128311 1411
rect 128737 1343 128771 1445
rect 131773 1411 131807 1445
rect 128001 1309 128185 1343
rect 128001 1275 128035 1309
rect 128127 1241 128829 1275
rect 128921 1207 128955 1309
rect 125977 1173 128955 1207
rect 129013 1309 129415 1343
rect 129013 1139 129047 1309
rect 129381 1275 129415 1309
rect 125977 1105 129047 1139
rect 129197 1139 129231 1241
rect 131957 1139 131991 1309
rect 129197 1105 131991 1139
rect 125977 1003 126011 1105
rect 132601 1071 132635 1377
rect 132693 1343 132727 1445
rect 132785 1411 132819 1513
rect 132877 1513 134291 1547
rect 132877 1343 132911 1513
rect 134257 1479 134291 1513
rect 132693 1309 132911 1343
rect 134257 1445 134567 1479
rect 134165 1139 134199 1445
rect 134441 1275 134475 1377
rect 134533 1343 134567 1445
rect 134717 1411 134751 1717
rect 138581 1683 138615 1717
rect 140605 1683 140639 1785
rect 141709 1751 141743 1785
rect 141801 1751 141835 1921
rect 143733 1819 143767 1989
rect 144837 1921 146895 1955
rect 143733 1785 144687 1819
rect 141801 1717 144595 1751
rect 141617 1683 141651 1717
rect 135119 1649 137293 1683
rect 140363 1649 140639 1683
rect 140915 1649 141099 1683
rect 141617 1649 143215 1683
rect 136591 1581 137017 1615
rect 138489 1547 138523 1649
rect 141065 1615 141099 1649
rect 143181 1615 143215 1649
rect 141341 1581 143123 1615
rect 143181 1581 144503 1615
rect 134809 1513 135027 1547
rect 136683 1513 136833 1547
rect 138489 1513 141191 1547
rect 134809 1343 134843 1513
rect 134993 1479 135027 1513
rect 134993 1445 141099 1479
rect 134533 1309 134843 1343
rect 134901 1377 135913 1411
rect 138707 1377 141007 1411
rect 134901 1275 134935 1377
rect 135453 1309 139535 1343
rect 134751 1241 134935 1275
rect 134165 1105 134901 1139
rect 125551 969 126011 1003
rect 128921 1037 131899 1071
rect 132601 1037 134843 1071
rect 128921 1003 128955 1037
rect 129473 969 131773 1003
rect 124505 765 124907 799
rect 125241 901 129105 935
rect 124505 663 124539 765
rect 125241 731 125275 901
rect 124597 697 125275 731
rect 122021 561 124447 595
rect 124597 527 124631 697
rect 121837 493 124631 527
rect 124689 459 124723 629
rect 121469 425 124723 459
rect 129289 391 129323 901
rect 121101 357 129323 391
rect 129473 323 129507 969
rect 121009 289 129507 323
rect 129565 255 129599 901
rect 131865 799 131899 1037
rect 132785 969 134751 1003
rect 132785 799 132819 969
rect 131865 765 132819 799
rect 134625 731 134659 901
rect 134717 799 134751 969
rect 134809 935 134843 1037
rect 135361 935 135395 1241
rect 135269 867 135303 901
rect 135453 867 135487 1309
rect 139501 1275 139535 1309
rect 140789 1309 140915 1343
rect 140789 1275 140823 1309
rect 135269 833 135487 867
rect 135545 799 135579 1241
rect 136097 1241 139443 1275
rect 139501 1241 140823 1275
rect 140881 1275 140915 1309
rect 136097 935 136131 1241
rect 139409 1207 139443 1241
rect 139501 1173 139593 1207
rect 139317 1139 139351 1173
rect 139501 1139 139535 1173
rect 139317 1105 139535 1139
rect 139685 1105 140697 1139
rect 134717 765 135579 799
rect 136189 731 136223 901
rect 134625 697 136223 731
rect 139685 595 139719 1105
rect 140087 1037 140605 1071
rect 140421 969 140639 1003
rect 140731 969 140881 1003
rect 140421 935 140455 969
rect 140513 663 140547 901
rect 140605 731 140639 969
rect 140973 799 141007 1377
rect 141065 867 141099 1445
rect 141157 935 141191 1513
rect 141249 867 141283 1377
rect 141065 833 141283 867
rect 141341 799 141375 1581
rect 143089 1547 143123 1581
rect 142479 1513 142997 1547
rect 143089 1513 143859 1547
rect 144135 1513 144377 1547
rect 143089 1445 143767 1479
rect 143089 1411 143123 1445
rect 143181 1377 143641 1411
rect 142445 1241 142905 1275
rect 142261 1071 142295 1105
rect 142445 1071 142479 1241
rect 142261 1037 142479 1071
rect 143181 935 143215 1377
rect 143733 1071 143767 1445
rect 143825 1411 143859 1513
rect 144043 1445 144285 1479
rect 144469 1411 144503 1581
rect 144561 1547 144595 1717
rect 144653 1615 144687 1785
rect 144837 1751 144871 1921
rect 146861 1887 146895 1921
rect 144929 1853 146803 1887
rect 146861 1853 147263 1887
rect 144653 1581 144837 1615
rect 144929 1547 144963 1853
rect 144561 1513 144963 1547
rect 145021 1785 146711 1819
rect 145021 1479 145055 1785
rect 145297 1649 146619 1683
rect 145147 1513 145205 1547
rect 145297 1411 145331 1649
rect 146585 1547 146619 1649
rect 146677 1615 146711 1785
rect 146769 1751 146803 1853
rect 147229 1819 147263 1853
rect 146895 1785 147137 1819
rect 147873 1819 147907 2125
rect 147965 2057 154347 2091
rect 147965 1819 147999 2057
rect 148333 1989 151679 2023
rect 148057 1751 148091 1785
rect 146769 1717 148091 1751
rect 148333 1615 148367 1989
rect 148425 1921 151587 1955
rect 148425 1751 148459 1921
rect 149161 1853 150391 1887
rect 149161 1819 149195 1853
rect 150357 1819 150391 1853
rect 146677 1581 148367 1615
rect 148517 1547 148551 1785
rect 149253 1785 150207 1819
rect 149069 1751 149103 1785
rect 149253 1751 149287 1785
rect 148885 1717 148977 1751
rect 149069 1717 149287 1751
rect 149713 1717 150081 1751
rect 148885 1615 148919 1717
rect 148977 1649 149195 1683
rect 148977 1547 149011 1649
rect 149161 1615 149195 1649
rect 145573 1513 145791 1547
rect 146585 1513 148459 1547
rect 148517 1513 149011 1547
rect 145573 1479 145607 1513
rect 143825 1377 144043 1411
rect 144009 1139 144043 1377
rect 144469 1377 145331 1411
rect 144101 1343 144135 1377
rect 144101 1309 145055 1343
rect 145021 1275 145055 1309
rect 145665 1275 145699 1445
rect 145021 1241 145699 1275
rect 145757 1207 145791 1513
rect 147413 1411 147447 1445
rect 147413 1377 147781 1411
rect 148425 1343 148459 1513
rect 149069 1479 149103 1581
rect 149529 1479 149563 1581
rect 149069 1445 149345 1479
rect 149621 1411 149655 1581
rect 148827 1377 149655 1411
rect 149713 1343 149747 1717
rect 150173 1411 150207 1785
rect 151093 1785 151403 1819
rect 150265 1547 150299 1785
rect 150449 1615 150483 1717
rect 150265 1513 150575 1547
rect 150541 1479 150575 1513
rect 150173 1377 150299 1411
rect 148425 1309 149747 1343
rect 145757 1173 148275 1207
rect 149563 1173 149897 1207
rect 144009 1105 147815 1139
rect 147781 1071 147815 1105
rect 143733 1037 146343 1071
rect 145607 969 145791 1003
rect 145757 935 145791 969
rect 146309 935 146343 1037
rect 147965 1071 147999 1105
rect 148241 1071 148275 1173
rect 149345 1105 149713 1139
rect 149345 1071 149379 1105
rect 147965 1037 148149 1071
rect 148241 1037 148977 1071
rect 147413 935 147447 1037
rect 149437 935 149471 1037
rect 150081 935 150115 1105
rect 142353 867 142387 901
rect 143273 867 143307 901
rect 142353 833 143307 867
rect 147321 867 147355 901
rect 150173 867 150207 901
rect 147321 833 150207 867
rect 150265 867 150299 1377
rect 150449 1275 150483 1445
rect 151093 1275 151127 1785
rect 151369 1751 151403 1785
rect 151185 1003 151219 1581
rect 151277 1275 151311 1717
rect 151461 1547 151495 1785
rect 151553 1751 151587 1921
rect 151645 1819 151679 1989
rect 152197 1853 153427 1887
rect 151737 1785 152139 1819
rect 151737 1751 151771 1785
rect 152105 1751 152139 1785
rect 151553 1717 151771 1751
rect 152013 1683 152047 1717
rect 152197 1683 152231 1853
rect 153393 1819 153427 1853
rect 152013 1649 152231 1683
rect 152289 1615 152323 1785
rect 151369 1071 151403 1377
rect 151461 1139 151495 1377
rect 151553 1139 151587 1581
rect 151645 1071 151679 1581
rect 151737 1581 152047 1615
rect 151737 1275 151771 1581
rect 151921 1411 151955 1513
rect 152013 1479 152047 1581
rect 152381 1547 152415 1785
rect 152139 1513 152415 1547
rect 152473 1649 152783 1683
rect 152473 1479 152507 1649
rect 152749 1615 152783 1649
rect 152013 1445 152507 1479
rect 152657 1479 152691 1581
rect 153301 1547 153335 1785
rect 154221 1683 154255 1785
rect 154313 1751 154347 2057
rect 154497 1819 154531 2125
rect 156153 1819 156187 2261
rect 157441 2159 157475 2261
rect 157809 2261 159591 2295
rect 160201 2261 161799 2295
rect 157809 2159 157843 2261
rect 159557 2227 159591 2261
rect 159557 2193 161247 2227
rect 157441 2125 157843 2159
rect 161213 2023 161247 2193
rect 161213 1989 161707 2023
rect 156245 1921 161431 1955
rect 154313 1717 155359 1751
rect 154221 1649 155267 1683
rect 153577 1547 153611 1581
rect 153577 1513 153761 1547
rect 153209 1479 153243 1513
rect 153209 1445 153887 1479
rect 153853 1411 153887 1445
rect 151921 1377 152691 1411
rect 151829 1241 152565 1275
rect 151369 1037 151679 1071
rect 151829 1003 151863 1241
rect 152657 1207 152691 1377
rect 152749 1275 152783 1377
rect 153853 1377 155083 1411
rect 152473 1173 152691 1207
rect 151185 969 151863 1003
rect 152013 935 152047 969
rect 152289 935 152323 969
rect 152013 901 152323 935
rect 152473 935 152507 1173
rect 152841 1139 152875 1377
rect 152933 1309 153151 1343
rect 152933 935 152967 1309
rect 152565 901 152967 935
rect 152565 867 152599 901
rect 150265 833 152599 867
rect 140973 765 141375 799
rect 144929 765 150207 799
rect 152047 765 152323 799
rect 144929 731 144963 765
rect 140605 697 144963 731
rect 145021 697 149931 731
rect 145021 663 145055 697
rect 140513 629 145055 663
rect 120825 221 129599 255
rect 129657 561 139719 595
rect 129657 187 129691 561
rect 135395 425 144837 459
rect 120733 153 129691 187
rect 149713 187 149747 629
rect 149897 595 149931 697
rect 150081 527 150115 629
rect 150173 595 150207 765
rect 152289 731 152323 765
rect 153025 731 153059 1241
rect 150449 697 151679 731
rect 152381 697 153059 731
rect 150449 663 150483 697
rect 151645 663 151679 697
rect 152381 663 152415 697
rect 150299 629 150483 663
rect 151369 629 151587 663
rect 151645 629 152415 663
rect 151369 595 151403 629
rect 150173 561 150449 595
rect 151461 527 151495 561
rect 150081 493 151495 527
rect 151553 459 151587 629
rect 153117 595 153151 1309
rect 153301 1309 153703 1343
rect 153301 1275 153335 1309
rect 153669 1275 153703 1309
rect 155049 1275 155083 1377
rect 153393 1241 153577 1275
rect 153669 1241 154531 1275
rect 154623 1241 154899 1275
rect 153393 1207 153427 1241
rect 153209 1173 153427 1207
rect 153485 1173 153795 1207
rect 153209 799 153243 1173
rect 153485 1139 153519 1173
rect 153427 1105 153519 1139
rect 153761 1139 153795 1173
rect 154037 1173 154439 1207
rect 154037 1139 154071 1173
rect 153335 833 153979 867
rect 153945 799 153979 833
rect 153393 663 153427 765
rect 153853 731 153887 765
rect 154129 731 154163 1105
rect 154313 799 154347 1105
rect 154405 799 154439 1173
rect 154497 1139 154531 1241
rect 154497 1105 154807 1139
rect 153853 697 154163 731
rect 154531 629 154589 663
rect 153117 561 153979 595
rect 151461 425 151587 459
rect 151461 323 151495 425
rect 151645 357 153301 391
rect 153485 357 153853 391
rect 151645 323 151679 357
rect 151461 289 151679 323
rect 153485 255 153519 357
rect 151311 221 151829 255
rect 152013 221 153519 255
rect 152013 187 152047 221
rect 149713 153 152047 187
rect 153945 119 153979 561
rect 154589 187 154623 357
rect 154681 255 154715 697
rect 154773 323 154807 1105
rect 154865 595 154899 1241
rect 155233 935 155267 1649
rect 155325 799 155359 1717
rect 156245 799 156279 1921
rect 156889 1853 157843 1887
rect 156337 1547 156371 1717
rect 156521 1547 156555 1785
rect 156889 1547 156923 1853
rect 157291 1785 157751 1819
rect 156981 1717 157441 1751
rect 156981 1615 157015 1717
rect 157717 1683 157751 1785
rect 157809 1751 157843 1853
rect 157901 1853 161339 1887
rect 157901 1683 157935 1853
rect 157257 1649 157567 1683
rect 157717 1649 157935 1683
rect 158729 1785 161155 1819
rect 156521 1275 156555 1377
rect 155325 765 156279 799
rect 156613 731 156647 1377
rect 157165 1343 157199 1513
rect 156797 1309 157199 1343
rect 156797 731 156831 1309
rect 156889 901 157165 935
rect 156889 799 156923 901
rect 157165 663 157199 697
rect 156739 629 157199 663
rect 157257 595 157291 1649
rect 157533 1615 157567 1649
rect 158729 1615 158763 1785
rect 157533 1581 157625 1615
rect 158821 1717 160511 1751
rect 157349 1275 157383 1513
rect 157441 1275 157475 1581
rect 157935 1513 158487 1547
rect 158453 1275 158487 1513
rect 157441 1241 158269 1275
rect 158453 1241 158729 1275
rect 158821 1207 158855 1717
rect 160477 1683 160511 1717
rect 159005 1547 159039 1649
rect 159097 1649 160051 1683
rect 159097 1343 159131 1649
rect 159315 1581 159683 1615
rect 157809 1173 158855 1207
rect 158913 1309 159131 1343
rect 157441 867 157475 1105
rect 157809 799 157843 1173
rect 157993 663 158027 765
rect 157659 629 158027 663
rect 154865 561 157291 595
rect 158269 595 158303 1105
rect 158913 1071 158947 1309
rect 158361 1037 158947 1071
rect 158361 935 158395 1037
rect 159005 663 159039 1241
rect 159189 595 159223 1513
rect 159557 1003 159591 1241
rect 159649 1071 159683 1581
rect 160017 1275 160051 1649
rect 160845 1649 161029 1683
rect 160385 1547 160419 1649
rect 160845 1615 160879 1649
rect 161121 1615 161155 1785
rect 160017 1241 160143 1275
rect 160109 1207 160143 1241
rect 160109 1173 160971 1207
rect 159649 1037 160051 1071
rect 159557 969 159867 1003
rect 158269 561 159223 595
rect 156521 459 156555 493
rect 156981 459 157015 493
rect 156521 425 157015 459
rect 159281 391 159315 629
rect 157199 357 159315 391
rect 159649 323 159683 901
rect 154773 289 159683 323
rect 159741 255 159775 629
rect 154681 221 159775 255
rect 159833 187 159867 969
rect 160017 731 160051 1037
rect 160937 935 160971 1173
rect 160937 901 161213 935
rect 160845 867 160879 901
rect 161305 867 161339 1853
rect 161397 1071 161431 1921
rect 161673 1751 161707 1989
rect 161765 1275 161799 2261
rect 161857 2057 170171 2091
rect 161489 1139 161523 1241
rect 161857 1139 161891 2057
rect 170137 2023 170171 2057
rect 170137 1989 170539 2023
rect 161949 1921 162167 1955
rect 161949 1411 161983 1921
rect 162133 1887 162167 1921
rect 162133 1853 170263 1887
rect 164065 1785 169803 1819
rect 164065 1479 164099 1785
rect 169309 1717 169677 1751
rect 164617 1649 169217 1683
rect 164617 1479 164651 1649
rect 169309 1615 169343 1717
rect 164985 1581 169343 1615
rect 162041 1445 163087 1479
rect 161489 1105 161891 1139
rect 162041 1071 162075 1445
rect 163053 1411 163087 1445
rect 164157 1411 164191 1445
rect 161397 1037 162075 1071
rect 162133 935 162167 1377
rect 163053 1377 164191 1411
rect 164709 1445 164927 1479
rect 164525 1411 164559 1445
rect 164709 1411 164743 1445
rect 164893 1411 164927 1445
rect 164525 1377 164743 1411
rect 160845 833 160971 867
rect 160603 765 160787 799
rect 154589 153 159867 187
rect 159925 187 159959 697
rect 160661 459 160695 697
rect 160753 595 160787 765
rect 160937 595 160971 833
rect 161397 901 162167 935
rect 162409 935 162443 1241
rect 162593 969 162811 1003
rect 161029 663 161063 833
rect 161155 765 161213 799
rect 161397 595 161431 901
rect 162501 867 162535 901
rect 160753 561 160879 595
rect 160937 561 161431 595
rect 161489 833 162535 867
rect 160845 527 160879 561
rect 161489 527 161523 833
rect 162593 799 162627 969
rect 160845 493 161523 527
rect 161581 765 162627 799
rect 161581 459 161615 765
rect 162225 697 162443 731
rect 162225 663 162259 697
rect 160661 425 161615 459
rect 162317 187 162351 629
rect 162409 255 162443 697
rect 162685 255 162719 901
rect 162409 221 162719 255
rect 162777 187 162811 969
rect 162961 527 162995 1377
rect 164801 1343 164835 1377
rect 163605 1309 164835 1343
rect 163605 1275 163639 1309
rect 164985 1207 165019 1581
rect 169769 1547 169803 1785
rect 170045 1683 170079 1785
rect 170229 1751 170263 1853
rect 170505 1751 170539 1989
rect 173909 1921 178359 1955
rect 173909 1751 173943 1921
rect 170505 1717 173943 1751
rect 174185 1853 178267 1887
rect 174185 1751 174219 1853
rect 175599 1785 175875 1819
rect 174277 1717 175381 1751
rect 174277 1683 174311 1717
rect 170045 1649 174311 1683
rect 169217 1513 169803 1547
rect 170137 1581 172103 1615
rect 169217 1411 169251 1513
rect 170137 1479 170171 1581
rect 169343 1445 169619 1479
rect 170137 1445 170263 1479
rect 169585 1411 169619 1445
rect 166767 1377 167227 1411
rect 169217 1377 169493 1411
rect 169585 1377 170171 1411
rect 163053 1173 165019 1207
rect 163053 935 163087 1173
rect 165905 1105 167009 1139
rect 164375 901 164559 935
rect 163145 799 163179 901
rect 164525 867 164559 901
rect 165905 867 165939 1105
rect 163087 765 163179 799
rect 166089 663 166123 765
rect 166181 697 166399 731
rect 163053 595 163087 629
rect 166181 595 166215 697
rect 163053 561 166215 595
rect 162961 493 163179 527
rect 159925 153 162351 187
rect 162409 153 162903 187
rect 162409 119 162443 153
rect 153945 85 162443 119
rect 113189 17 120215 51
rect 162777 51 162811 153
rect 162869 119 162903 153
rect 163145 119 163179 493
rect 166273 459 166307 629
rect 166365 527 166399 697
rect 167193 663 167227 1377
rect 167285 1241 170045 1275
rect 167101 595 167135 629
rect 167285 595 167319 1241
rect 170137 1207 170171 1377
rect 168941 1173 169711 1207
rect 168941 1139 168975 1173
rect 169677 1139 169711 1173
rect 169861 1173 170171 1207
rect 168941 697 169125 731
rect 168941 663 168975 697
rect 167101 561 167319 595
rect 169585 595 169619 1105
rect 169861 663 169895 1173
rect 170229 867 170263 1445
rect 169953 833 170263 867
rect 170321 1445 171609 1479
rect 169953 731 169987 833
rect 170321 799 170355 1445
rect 172069 1343 172103 1581
rect 173541 1581 174219 1615
rect 173541 1479 173575 1581
rect 174185 1479 174219 1581
rect 175749 1547 175783 1717
rect 175841 1547 175875 1785
rect 175933 1785 178175 1819
rect 175933 1479 175967 1785
rect 174185 1445 175967 1479
rect 173449 1411 173483 1445
rect 173725 1411 173759 1445
rect 176577 1411 176611 1513
rect 173449 1377 173759 1411
rect 173817 1377 176059 1411
rect 173817 1343 173851 1377
rect 172069 1309 173851 1343
rect 175783 1309 175933 1343
rect 176025 1275 176059 1377
rect 176761 1445 177715 1479
rect 176485 1343 176519 1377
rect 176761 1343 176795 1445
rect 176485 1309 176795 1343
rect 176853 1275 176887 1377
rect 176025 1241 176887 1275
rect 176945 1377 177589 1411
rect 176945 1275 176979 1377
rect 177681 1275 177715 1445
rect 177773 1275 177807 1717
rect 177865 1649 178083 1683
rect 177865 1615 177899 1649
rect 177957 1411 177991 1581
rect 178049 1479 178083 1649
rect 178141 1547 178175 1785
rect 178233 1615 178267 1853
rect 178325 1819 178359 1921
rect 178325 1785 179095 1819
rect 178601 1717 178877 1751
rect 178601 1683 178635 1717
rect 178233 1581 178785 1615
rect 178141 1513 178727 1547
rect 178693 1411 178727 1513
rect 178969 1479 179003 1581
rect 177773 1241 177865 1275
rect 175841 1207 175875 1241
rect 175841 1173 178267 1207
rect 170045 765 170355 799
rect 170413 833 173943 867
rect 170045 731 170079 765
rect 170413 731 170447 833
rect 170137 697 170447 731
rect 173909 731 173943 833
rect 176669 833 178175 867
rect 173909 697 176577 731
rect 170137 663 170171 697
rect 169861 629 170171 663
rect 170229 595 170263 629
rect 169585 561 170263 595
rect 170321 527 170355 629
rect 175657 629 176209 663
rect 175657 595 175691 629
rect 176669 595 176703 833
rect 177037 765 178083 799
rect 177037 663 177071 765
rect 177347 697 177623 731
rect 177589 663 177623 697
rect 178049 663 178083 765
rect 178141 731 178175 833
rect 178233 799 178267 1173
rect 179061 867 179095 1785
rect 179153 1479 179187 3077
rect 262965 3077 268393 3111
rect 231501 2261 232547 2295
rect 179245 2057 191883 2091
rect 179245 1683 179279 2057
rect 191849 2023 191883 2057
rect 191849 1989 197403 2023
rect 179797 1853 180843 1887
rect 179371 1037 179613 1071
rect 179279 969 179429 1003
rect 179371 901 179521 935
rect 179705 867 179739 1717
rect 179061 833 179739 867
rect 179797 799 179831 1853
rect 180441 1785 180659 1819
rect 180441 1751 180475 1785
rect 179889 1479 179923 1513
rect 179889 1445 180441 1479
rect 178233 765 179831 799
rect 179889 731 179923 1377
rect 180073 1207 180107 1377
rect 180533 1207 180567 1717
rect 180625 1207 180659 1785
rect 180809 1479 180843 1853
rect 183569 1853 190043 1887
rect 183569 1819 183603 1853
rect 184063 1581 189583 1615
rect 189549 1547 189583 1581
rect 184029 1513 184121 1547
rect 178141 697 179923 731
rect 179981 833 180073 867
rect 176427 561 176703 595
rect 166365 493 170355 527
rect 170413 493 175841 527
rect 170413 459 170447 493
rect 175933 459 175967 561
rect 176243 493 176485 527
rect 177405 459 177439 629
rect 179981 459 180015 833
rect 166273 425 170447 459
rect 170505 425 171275 459
rect 170505 323 170539 425
rect 162869 85 163179 119
rect 164157 289 170539 323
rect 171241 323 171275 425
rect 175841 425 175967 459
rect 176025 425 176427 459
rect 177405 425 180015 459
rect 171241 289 175323 323
rect 164157 51 164191 289
rect 175289 187 175323 289
rect 175841 255 175875 425
rect 176025 391 176059 425
rect 176393 391 176427 425
rect 175967 357 176059 391
rect 176301 323 176335 357
rect 180165 323 180199 1173
rect 176301 289 180199 323
rect 180257 255 180291 833
rect 180717 731 180751 1445
rect 182557 1071 182591 1445
rect 183845 1139 183879 1173
rect 184029 1139 184063 1513
rect 183845 1105 184063 1139
rect 189457 1071 189491 1513
rect 189733 1445 189951 1479
rect 189733 1275 189767 1445
rect 189825 1275 189859 1377
rect 189917 1343 189951 1445
rect 190009 1411 190043 1853
rect 190101 1853 191423 1887
rect 190101 1343 190135 1853
rect 191021 1785 191331 1819
rect 191021 1751 191055 1785
rect 191297 1751 191331 1785
rect 190285 1683 190319 1717
rect 190469 1717 191055 1751
rect 190469 1683 190503 1717
rect 190285 1649 190503 1683
rect 190377 1581 190837 1615
rect 190377 1479 190411 1581
rect 190469 1513 190779 1547
rect 190469 1411 190503 1513
rect 190745 1479 190779 1513
rect 190745 1445 191113 1479
rect 190561 1343 190595 1377
rect 189917 1309 190135 1343
rect 190285 1309 190595 1343
rect 190653 1343 190687 1445
rect 190745 1377 191147 1411
rect 189825 1241 190135 1275
rect 190101 1207 190135 1241
rect 190285 1207 190319 1309
rect 190745 1275 190779 1377
rect 191113 1343 191147 1377
rect 191021 1275 191055 1309
rect 191021 1241 191147 1275
rect 190101 1173 190319 1207
rect 190929 1173 191021 1207
rect 190929 1071 190963 1173
rect 182557 1037 189123 1071
rect 189457 1037 190963 1071
rect 189089 935 189123 1037
rect 191113 935 191147 1241
rect 189089 901 191147 935
rect 183569 833 190319 867
rect 183569 731 183603 833
rect 190285 799 190319 833
rect 191205 799 191239 1717
rect 191389 1683 191423 1853
rect 191297 1649 191423 1683
rect 191481 1853 197311 1887
rect 191297 1275 191331 1649
rect 191389 1343 191423 1445
rect 183695 765 184247 799
rect 180717 697 183603 731
rect 183971 697 184063 731
rect 183511 629 183603 663
rect 183787 629 183971 663
rect 183569 595 183603 629
rect 183569 561 183845 595
rect 183695 493 183879 527
rect 183511 425 183695 459
rect 183661 391 183695 425
rect 183569 323 183603 357
rect 183845 323 183879 493
rect 183937 459 183971 629
rect 184029 527 184063 697
rect 184213 663 184247 765
rect 190469 765 191239 799
rect 190193 731 190227 765
rect 190469 731 190503 765
rect 191481 731 191515 1853
rect 196633 1785 197035 1819
rect 191665 1683 191699 1717
rect 196633 1683 196667 1785
rect 191665 1649 191883 1683
rect 196725 1717 196909 1751
rect 191849 1615 191883 1649
rect 196725 1615 196759 1717
rect 197001 1683 197035 1785
rect 191849 1581 196759 1615
rect 191665 1513 196759 1547
rect 191665 1479 191699 1513
rect 191975 1445 196633 1479
rect 191573 1207 191607 1445
rect 192125 1377 195471 1411
rect 192125 1207 192159 1377
rect 191573 1173 192159 1207
rect 194609 1309 195345 1343
rect 190193 697 190503 731
rect 190653 697 191515 731
rect 190653 663 190687 697
rect 194609 663 194643 1309
rect 184213 629 190687 663
rect 191297 629 194643 663
rect 191297 595 191331 629
rect 190561 561 191331 595
rect 190561 527 190595 561
rect 184029 493 190595 527
rect 195437 527 195471 1377
rect 196633 1207 196667 1309
rect 196725 1275 196759 1513
rect 196817 1343 196851 1649
rect 197185 1479 197219 1717
rect 197277 1547 197311 1853
rect 197369 1751 197403 1989
rect 214113 1989 222151 2023
rect 214113 1615 214147 1989
rect 216781 1921 221047 1955
rect 216781 1819 216815 1921
rect 215125 1785 216815 1819
rect 220277 1853 220771 1887
rect 220277 1819 220311 1853
rect 220737 1819 220771 1853
rect 198013 1581 200899 1615
rect 197277 1513 197921 1547
rect 198013 1479 198047 1581
rect 197185 1445 198047 1479
rect 196909 1411 196943 1445
rect 198749 1411 198783 1513
rect 196909 1377 198783 1411
rect 198841 1513 199209 1547
rect 199393 1513 200807 1547
rect 197219 1309 198565 1343
rect 196725 1241 196943 1275
rect 196633 1173 196851 1207
rect 196817 527 196851 1173
rect 196909 595 196943 1241
rect 198841 731 198875 1513
rect 199393 1479 199427 1513
rect 197001 697 198875 731
rect 198933 1445 199427 1479
rect 197001 663 197035 697
rect 197093 595 197127 629
rect 196909 561 197127 595
rect 195437 493 196207 527
rect 196817 493 198599 527
rect 183937 425 184339 459
rect 193447 425 196115 459
rect 183569 289 183753 323
rect 175841 221 180291 255
rect 183603 221 184213 255
rect 184305 187 184339 425
rect 193355 357 196023 391
rect 175289 153 183753 187
rect 195989 119 196023 357
rect 196081 187 196115 425
rect 196173 323 196207 493
rect 196541 425 198473 459
rect 196541 391 196575 425
rect 198565 391 198599 493
rect 198933 459 198967 1445
rect 199025 1377 199243 1411
rect 199025 663 199059 1377
rect 199209 1343 199243 1377
rect 199117 663 199151 1309
rect 200405 731 200439 1309
rect 200773 1139 200807 1513
rect 200865 1479 200899 1581
rect 211077 1581 211295 1615
rect 214423 1581 214515 1615
rect 211077 1547 211111 1581
rect 202889 1479 202923 1513
rect 211169 1479 211203 1513
rect 202889 1445 211203 1479
rect 211261 1479 211295 1581
rect 211261 1445 211445 1479
rect 211169 1377 211387 1411
rect 211169 1343 211203 1377
rect 202923 1309 211203 1343
rect 211261 1139 211295 1309
rect 211353 1275 211387 1377
rect 214205 1377 214423 1411
rect 214205 1343 214239 1377
rect 211353 1241 212767 1275
rect 200773 1105 211295 1139
rect 199209 697 200439 731
rect 204303 697 204545 731
rect 196943 357 198289 391
rect 198565 357 198657 391
rect 199209 323 199243 697
rect 199301 629 204453 663
rect 199301 391 199335 629
rect 208041 595 208075 765
rect 208961 765 210007 799
rect 208133 663 208167 697
rect 208409 697 208777 731
rect 208409 663 208443 697
rect 208133 629 208443 663
rect 208961 595 208995 765
rect 209973 731 210007 765
rect 209973 697 212675 731
rect 208041 561 208995 595
rect 212549 459 212583 629
rect 212641 527 212675 697
rect 212733 663 212767 1241
rect 214297 935 214331 1309
rect 214389 1275 214423 1377
rect 214481 1343 214515 1581
rect 214849 1343 214883 1581
rect 215125 1275 215159 1785
rect 220645 1649 220955 1683
rect 220645 1615 220679 1649
rect 220921 1615 220955 1649
rect 217977 1581 220369 1615
rect 220771 1581 220863 1615
rect 214389 1241 215159 1275
rect 217609 1445 217827 1479
rect 217609 1207 217643 1445
rect 217793 1411 217827 1445
rect 217977 1207 218011 1581
rect 220829 1547 220863 1581
rect 218345 1445 218655 1479
rect 218345 1411 218379 1445
rect 218621 1343 218655 1445
rect 218713 1445 218931 1479
rect 220219 1445 220369 1479
rect 218713 1411 218747 1445
rect 213745 901 214331 935
rect 214573 1173 217643 1207
rect 217793 1173 218011 1207
rect 218897 1207 218931 1445
rect 221013 1275 221047 1921
rect 222117 1615 222151 1989
rect 231501 1751 231535 2261
rect 231593 2193 232455 2227
rect 231593 1819 231627 2193
rect 231961 1853 232271 1887
rect 224049 1717 224727 1751
rect 224049 1683 224083 1717
rect 224693 1683 224727 1717
rect 224601 1615 224635 1649
rect 231685 1615 231719 1785
rect 231811 1649 231903 1683
rect 224601 1581 224969 1615
rect 225245 1581 231719 1615
rect 222025 1479 222059 1581
rect 224417 1547 224451 1581
rect 224359 1513 224451 1547
rect 225245 1479 225279 1581
rect 222025 1445 225279 1479
rect 224543 1377 225061 1411
rect 228189 1377 228591 1411
rect 228189 1343 228223 1377
rect 224325 1309 224601 1343
rect 224693 1309 225003 1343
rect 225463 1309 225831 1343
rect 221013 1241 224267 1275
rect 224233 1207 224267 1241
rect 218897 1173 223991 1207
rect 213745 799 213779 901
rect 213963 697 214297 731
rect 214573 663 214607 1173
rect 214055 629 214607 663
rect 214941 765 215343 799
rect 214941 663 214975 765
rect 215309 663 215343 765
rect 215309 629 217701 663
rect 212641 493 217609 527
rect 217793 459 217827 1173
rect 217919 1105 218195 1139
rect 218161 1071 218195 1105
rect 218161 1037 221691 1071
rect 218379 969 218529 1003
rect 218103 901 218437 935
rect 221657 731 221691 1037
rect 223865 799 223899 1105
rect 223957 1071 223991 1173
rect 224141 1139 224175 1173
rect 224325 1139 224359 1309
rect 224693 1275 224727 1309
rect 224451 1241 224727 1275
rect 224969 1275 225003 1309
rect 224141 1105 224359 1139
rect 224417 1173 225187 1207
rect 224417 1071 224451 1173
rect 225153 1139 225187 1173
rect 223957 1037 224451 1071
rect 224601 1105 225095 1139
rect 225245 1173 225647 1207
rect 224601 799 224635 1105
rect 225061 1071 225095 1105
rect 225245 1071 225279 1173
rect 225613 1139 225647 1173
rect 225797 1139 225831 1309
rect 228281 1207 228315 1309
rect 228557 1207 228591 1377
rect 228557 1173 231811 1207
rect 228373 1139 228407 1173
rect 231777 1139 231811 1173
rect 225797 1105 228407 1139
rect 225061 1037 225279 1071
rect 224969 1003 225003 1037
rect 225429 1003 225463 1037
rect 224969 969 225463 1003
rect 225521 935 225555 1105
rect 224141 765 224233 799
rect 224325 765 224635 799
rect 225061 901 225555 935
rect 224141 731 224175 765
rect 218161 697 219759 731
rect 218161 527 218195 697
rect 219725 595 219759 697
rect 221657 697 224175 731
rect 221473 663 221507 697
rect 224325 663 224359 765
rect 225061 731 225095 901
rect 231685 799 231719 1105
rect 231869 1071 231903 1649
rect 231961 1479 231995 1853
rect 232237 1819 232271 1853
rect 232237 1785 232363 1819
rect 232145 1683 232179 1785
rect 232329 1547 232363 1785
rect 232421 1751 232455 2193
rect 232513 2023 232547 2261
rect 260941 2057 261435 2091
rect 232513 1989 239355 2023
rect 232789 1921 239263 1955
rect 232605 1615 232639 1785
rect 232789 1547 232823 1921
rect 233893 1785 236745 1819
rect 232329 1513 232823 1547
rect 232237 1139 232271 1241
rect 233249 1139 233283 1445
rect 232237 1105 233283 1139
rect 233341 1071 233375 1649
rect 231869 1037 233375 1071
rect 233893 935 233927 1785
rect 233985 1615 234019 1717
rect 236561 1513 236779 1547
rect 236561 1479 236595 1513
rect 236653 1207 236687 1445
rect 236745 1207 236779 1513
rect 237941 1445 239045 1479
rect 237941 1207 237975 1445
rect 239137 1411 239171 1717
rect 239229 1479 239263 1921
rect 239321 1751 239355 1989
rect 260941 1955 260975 2057
rect 250085 1921 251223 1955
rect 250085 1751 250119 1921
rect 251189 1887 251223 1921
rect 258641 1921 260975 1955
rect 258641 1887 258675 1921
rect 251189 1853 251591 1887
rect 251557 1751 251591 1853
rect 240091 1717 241621 1751
rect 250821 1479 250855 1717
rect 239229 1445 241437 1479
rect 249809 1411 249843 1445
rect 250913 1411 250947 1717
rect 239137 1377 239447 1411
rect 249809 1377 250947 1411
rect 251833 1853 252971 1887
rect 251465 1411 251499 1717
rect 251465 1377 251591 1411
rect 238585 1309 239171 1343
rect 238033 1241 238217 1275
rect 231869 901 233927 935
rect 231869 799 231903 901
rect 238033 867 238067 1241
rect 231685 765 231903 799
rect 231961 833 238067 867
rect 231961 799 231995 833
rect 232915 765 233433 799
rect 221047 629 221507 663
rect 224417 697 224635 731
rect 224417 663 224451 697
rect 224601 663 224635 697
rect 225153 663 225187 697
rect 225521 697 231777 731
rect 224601 629 225187 663
rect 224141 595 224175 629
rect 225429 595 225463 629
rect 219725 561 222243 595
rect 224141 561 225463 595
rect 217919 493 218195 527
rect 222209 527 222243 561
rect 225521 527 225555 697
rect 231593 595 231627 629
rect 232053 595 232087 765
rect 238401 731 238435 765
rect 238585 731 238619 1309
rect 239137 1275 239171 1309
rect 238711 1241 238987 1275
rect 238953 1207 238987 1241
rect 239321 1207 239355 1241
rect 238803 1173 238895 1207
rect 238953 1173 239355 1207
rect 238861 799 238895 1173
rect 239413 1139 239447 1377
rect 251557 1275 251591 1377
rect 239229 1105 239447 1139
rect 239505 1241 239597 1275
rect 239229 1071 239263 1105
rect 239045 1003 239079 1037
rect 239321 1003 239355 1037
rect 239045 969 239355 1003
rect 239079 833 239413 867
rect 239505 799 239539 1241
rect 251465 1207 251499 1241
rect 251833 1207 251867 1853
rect 252569 1785 252787 1819
rect 252569 1751 252603 1785
rect 251465 1173 251867 1207
rect 247359 1105 247601 1139
rect 245519 1037 248337 1071
rect 241839 969 242081 1003
rect 241931 901 242173 935
rect 241747 833 242081 867
rect 238401 697 238619 731
rect 238861 765 239539 799
rect 239597 765 241897 799
rect 238769 731 238803 765
rect 239597 731 239631 765
rect 238769 697 239631 731
rect 231593 561 232087 595
rect 241529 561 247083 595
rect 222209 493 225555 527
rect 241529 527 241563 561
rect 247049 527 247083 561
rect 251189 527 251223 1173
rect 252661 663 252695 1717
rect 252603 629 252695 663
rect 252753 663 252787 1785
rect 252937 1343 252971 1853
rect 258457 1853 258675 1887
rect 258457 1819 258491 1853
rect 261401 1819 261435 2057
rect 261401 1785 262045 1819
rect 253615 1717 257169 1751
rect 258215 1717 258365 1751
rect 258273 1615 258307 1649
rect 258549 1615 258583 1785
rect 261895 1717 262321 1751
rect 262539 1717 262631 1751
rect 262597 1683 262631 1717
rect 260699 1649 261401 1683
rect 262229 1649 262539 1683
rect 262597 1649 262873 1683
rect 262229 1615 262263 1649
rect 262505 1615 262539 1649
rect 258273 1581 258583 1615
rect 260331 1581 260849 1615
rect 262505 1581 262781 1615
rect 262413 1547 262447 1581
rect 262965 1547 262999 3077
rect 290473 1921 294187 1955
rect 280169 1853 282135 1887
rect 258549 1513 260975 1547
rect 262413 1513 262999 1547
rect 258549 1479 258583 1513
rect 258365 1445 258583 1479
rect 260607 1445 260883 1479
rect 258365 1411 258399 1445
rect 258457 1343 258491 1377
rect 252937 1309 258491 1343
rect 260849 1343 260883 1445
rect 260941 1411 260975 1513
rect 261125 1445 263149 1479
rect 260941 1377 261033 1411
rect 261125 1343 261159 1445
rect 260849 1309 261159 1343
rect 259653 1173 260757 1207
rect 252753 629 259377 663
rect 259653 527 259687 1173
rect 261309 595 261343 697
rect 263241 595 263275 1785
rect 268761 1785 268945 1819
rect 268761 1751 268795 1785
rect 280169 1751 280203 1853
rect 280261 1785 281951 1819
rect 279985 1683 280019 1717
rect 280261 1683 280295 1785
rect 279985 1649 280295 1683
rect 280445 1649 280755 1683
rect 265265 1513 265667 1547
rect 265265 1479 265299 1513
rect 265633 1479 265667 1513
rect 270509 1479 270543 1581
rect 274557 1581 280353 1615
rect 273269 1513 274039 1547
rect 265483 1445 265575 1479
rect 265633 1445 268853 1479
rect 270509 1445 271429 1479
rect 265081 663 265115 1445
rect 265541 1139 265575 1445
rect 270727 1241 272349 1275
rect 265541 1105 267231 1139
rect 267197 663 267231 1105
rect 273269 731 273303 1513
rect 274005 1479 274039 1513
rect 274557 1479 274591 1581
rect 280445 1547 280479 1649
rect 280169 1513 280479 1547
rect 280169 1479 280203 1513
rect 279559 1445 280203 1479
rect 273855 1241 279985 1275
rect 280077 799 280111 1173
rect 280629 867 280663 1581
rect 279341 765 279651 799
rect 279341 731 279375 765
rect 279617 663 279651 765
rect 279893 765 280111 799
rect 280261 833 280663 867
rect 279801 663 279835 697
rect 265081 629 267105 663
rect 267197 629 267289 663
rect 279617 629 279835 663
rect 261309 561 263275 595
rect 279893 527 279927 765
rect 280261 731 280295 833
rect 279985 697 280295 731
rect 279985 663 280019 697
rect 280721 595 280755 1649
rect 281917 1479 281951 1785
rect 282101 1547 282135 1853
rect 290473 1751 290507 1921
rect 290565 1853 294095 1887
rect 289737 1615 289771 1717
rect 289737 1581 290473 1615
rect 290565 1547 290599 1853
rect 282101 1513 285873 1547
rect 289679 1513 290599 1547
rect 290749 1649 293819 1683
rect 282193 1445 285597 1479
rect 285723 1445 285965 1479
rect 289587 1445 290323 1479
rect 281825 1241 282135 1275
rect 281549 1139 281583 1173
rect 281825 1139 281859 1241
rect 282101 1207 282135 1241
rect 281549 1105 281859 1139
rect 282009 1139 282043 1173
rect 282193 1139 282227 1445
rect 282009 1105 282227 1139
rect 281457 663 281491 697
rect 281457 629 281641 663
rect 281733 595 281767 697
rect 280721 561 281767 595
rect 247049 493 247601 527
rect 251189 493 251649 527
rect 260883 493 265541 527
rect 268887 493 270417 527
rect 270543 493 270785 527
rect 279835 493 279927 527
rect 203107 425 212457 459
rect 212549 425 217827 459
rect 241655 425 251005 459
rect 251407 425 260665 459
rect 260975 425 265081 459
rect 268979 425 270325 459
rect 270635 425 279985 459
rect 280295 425 281641 459
rect 196173 289 199243 323
rect 199393 187 199427 425
rect 196081 153 199427 187
rect 251591 357 259837 391
rect 270543 357 280077 391
rect 199485 119 199519 357
rect 285137 187 285171 1377
rect 285781 731 285815 1377
rect 285505 663 285539 697
rect 286149 663 286183 833
rect 285505 629 285631 663
rect 285597 595 285631 629
rect 285597 561 285723 595
rect 285689 527 285723 561
rect 285689 493 285907 527
rect 285539 425 285781 459
rect 285873 323 285907 493
rect 287345 391 287379 1377
rect 289277 867 289311 1445
rect 290289 1207 290323 1445
rect 289277 833 289737 867
rect 287437 731 287471 833
rect 290657 731 290691 1173
rect 287437 697 290691 731
rect 290231 629 290657 663
rect 289645 595 289679 629
rect 290749 595 290783 1649
rect 293785 1615 293819 1649
rect 290841 1581 291025 1615
rect 290841 1207 290875 1581
rect 293877 1547 293911 1717
rect 290933 1513 293911 1547
rect 290933 1275 290967 1513
rect 291117 867 291151 1241
rect 289645 561 290783 595
rect 290841 833 291151 867
rect 293877 867 293911 1445
rect 294061 1207 294095 1853
rect 294153 1819 294187 1921
rect 294153 1785 295291 1819
rect 295257 1751 295291 1785
rect 297005 1785 298695 1819
rect 295165 1411 295199 1717
rect 296763 1445 296855 1479
rect 295165 1377 295383 1411
rect 295349 1207 295383 1377
rect 296821 1275 296855 1445
rect 290841 527 290875 833
rect 289829 493 290875 527
rect 293969 527 294003 1173
rect 295257 731 295291 1173
rect 296913 1003 296947 1649
rect 296855 969 296947 1003
rect 297005 663 297039 1785
rect 298385 1717 298603 1751
rect 298385 1683 298419 1717
rect 298477 1547 298511 1649
rect 298569 1615 298603 1717
rect 298661 1683 298695 1785
rect 309701 1717 315071 1751
rect 298661 1649 300041 1683
rect 298569 1581 298845 1615
rect 298695 1513 300167 1547
rect 296947 629 297039 663
rect 297281 1445 300041 1479
rect 297281 595 297315 1445
rect 297925 1207 297959 1241
rect 297925 1173 298109 1207
rect 297189 561 297315 595
rect 297465 561 297683 595
rect 297189 527 297223 561
rect 296763 493 297223 527
rect 297465 527 297499 561
rect 289829 391 289863 493
rect 289955 425 296855 459
rect 287345 357 289311 391
rect 285965 289 289185 323
rect 285781 255 285815 289
rect 285965 255 285999 289
rect 289277 255 289311 357
rect 285781 221 285999 255
rect 286057 221 289311 255
rect 296821 255 296855 425
rect 297005 255 297039 425
rect 297557 391 297591 493
rect 297649 391 297683 561
rect 300133 323 300167 1513
rect 304089 1479 304123 1649
rect 304181 1547 304215 1649
rect 304273 1479 304307 1513
rect 304089 1445 304307 1479
rect 309149 1207 309183 1445
rect 309701 1411 309735 1717
rect 314703 1649 314795 1683
rect 309425 1275 309459 1377
rect 309275 1241 309459 1275
rect 300685 1173 300777 1207
rect 309149 1173 309425 1207
rect 300685 391 300719 1173
rect 306849 867 306883 969
rect 314761 799 314795 1649
rect 315037 1275 315071 1717
rect 319361 1649 319821 1683
rect 319361 1547 319395 1649
rect 318717 1513 318993 1547
rect 318475 1445 318625 1479
rect 315037 1241 318625 1275
rect 318717 1071 318751 1513
rect 314853 1037 318751 1071
rect 314669 731 314703 765
rect 314853 731 314887 1037
rect 317521 969 318717 1003
rect 317521 799 317555 969
rect 317613 799 317647 901
rect 319453 799 319487 1513
rect 320189 1513 320499 1547
rect 320189 1479 320223 1513
rect 320465 1479 320499 1513
rect 320465 1445 320591 1479
rect 329699 1445 329791 1479
rect 320557 1411 320591 1445
rect 319637 867 319671 1377
rect 320557 1377 321879 1411
rect 319729 731 319763 1377
rect 314669 697 314887 731
rect 319361 697 319763 731
rect 319361 663 319395 697
rect 321845 527 321879 1377
rect 329757 1275 329791 1445
rect 327089 1207 327123 1241
rect 326939 1173 327123 1207
rect 335863 1241 336139 1275
rect 322949 969 323535 1003
rect 322949 527 322983 969
rect 323501 935 323535 969
rect 323409 527 323443 901
rect 327457 527 327491 1241
rect 335495 561 335737 595
rect 336013 527 336047 1173
rect 327457 493 328009 527
rect 335587 493 335771 527
rect 336105 527 336139 1241
rect 337577 527 337611 1241
rect 337945 1003 337979 1717
rect 338773 527 338807 969
rect 338865 527 338899 1241
rect 345397 1071 345431 1241
rect 342211 1037 343223 1071
rect 343189 935 343223 1037
rect 345765 1003 345799 1649
rect 348985 1207 349019 1717
rect 347363 561 347513 595
rect 318809 459 318843 493
rect 335737 459 335771 493
rect 309275 425 318625 459
rect 318809 425 323225 459
rect 337485 391 337519 493
rect 337945 391 337979 425
rect 300777 323 300811 357
rect 300133 289 300811 323
rect 322949 323 322983 357
rect 337485 357 337979 391
rect 348249 391 348283 901
rect 348525 527 348559 1173
rect 349445 935 349479 1717
rect 352665 527 352699 1037
rect 352849 527 352883 1717
rect 348341 391 348375 493
rect 323409 323 323443 357
rect 354137 323 354171 1173
rect 322949 289 323443 323
rect 351963 289 354171 323
rect 355977 323 356011 1173
rect 356161 935 356195 1173
rect 356437 799 356471 1445
rect 358093 1411 358127 1649
rect 367293 1275 367327 1377
rect 357081 1071 357115 1173
rect 357909 1071 357943 1241
rect 368397 1207 368431 1785
rect 367051 1173 367109 1207
rect 364165 1105 364383 1139
rect 364165 1071 364199 1105
rect 364257 935 364291 1037
rect 364349 935 364383 1105
rect 368489 935 368523 1377
rect 374653 1275 374687 1377
rect 374745 1207 374779 1377
rect 374837 1207 374871 1785
rect 372721 1105 372939 1139
rect 372721 1003 372755 1105
rect 372905 1003 372939 1105
rect 376033 1071 376067 1717
rect 372905 969 373089 1003
rect 378425 867 378459 1037
rect 372445 833 372813 867
rect 386429 867 386463 1241
rect 386521 1207 386555 1445
rect 388453 1411 388487 1785
rect 390419 1309 390753 1343
rect 391213 1207 391247 1445
rect 391581 1411 391615 1785
rect 390695 1105 390845 1139
rect 393605 1071 393639 1445
rect 404277 867 404311 1241
rect 386429 833 386521 867
rect 372445 799 372479 833
rect 356529 561 356747 595
rect 356529 527 356563 561
rect 356621 391 356655 493
rect 356713 391 356747 561
rect 386337 459 386371 765
rect 386429 527 386463 765
rect 395997 527 396031 765
rect 412189 731 412223 1581
rect 432245 1275 432279 1513
rect 459569 1275 459603 1445
rect 473185 1275 473219 1445
rect 500969 1275 501003 1513
rect 509525 1275 509559 1513
rect 473369 1071 473403 1241
rect 521703 1105 521761 1139
rect 493885 1071 493919 1105
rect 493885 1037 494069 1071
rect 516793 935 516827 1037
rect 528201 935 528235 1649
rect 555433 1275 555467 1445
rect 556169 1275 556203 1581
rect 560217 1343 560251 1445
rect 538229 867 538263 1105
rect 425069 527 425103 833
rect 386521 459 386555 493
rect 372663 425 372755 459
rect 386337 425 386555 459
rect 372721 391 372755 425
rect 367143 357 368615 391
rect 368581 323 368615 357
rect 372353 357 372663 391
rect 372721 357 372813 391
rect 372997 357 373181 391
rect 372353 323 372387 357
rect 372629 323 372663 357
rect 372997 323 373031 357
rect 372629 289 373031 323
rect 296821 221 297039 255
rect 372571 221 372997 255
rect 286057 187 286091 221
rect 285137 153 286091 187
rect 335403 153 335645 187
rect 347547 153 347697 187
rect 372387 153 373273 187
rect 376803 153 376953 187
rect 430773 119 430807 765
rect 430865 527 430899 833
rect 162777 17 164191 51
rect 183569 51 183603 85
rect 195989 85 199519 119
rect 335587 85 335737 119
rect 347455 85 347605 119
rect 372479 85 372721 119
rect 436109 119 436143 765
rect 463709 527 463743 765
rect 473185 527 473219 765
rect 473369 663 473403 765
rect 473495 561 473553 595
rect 481097 527 481131 833
rect 473403 493 473645 527
rect 549303 1105 549361 1139
rect 543105 867 543139 1105
rect 559481 935 559515 1105
rect 508881 527 508915 833
rect 514769 527 514803 765
rect 459603 425 459753 459
rect 473495 425 473553 459
rect 473403 357 473645 391
rect 507811 357 507869 391
rect 473495 289 473737 323
rect 473495 153 473645 187
rect 184029 51 184063 85
rect 568313 51 568347 1717
rect 183569 17 184063 51
rect 335495 17 335645 51
rect 347363 17 347697 51
<< viali >>
rect 557733 680425 557767 680459
rect 216597 680357 216631 680391
rect 207029 680289 207063 680323
rect 11713 679813 11747 679847
rect 11713 679677 11747 679711
rect 16589 679813 16623 679847
rect 16589 679677 16623 679711
rect 31033 679813 31067 679847
rect 31033 679677 31067 679711
rect 35909 679813 35943 679847
rect 35909 679677 35943 679711
rect 50353 679813 50387 679847
rect 50353 679677 50387 679711
rect 55229 679813 55263 679847
rect 55229 679677 55263 679711
rect 69673 679813 69707 679847
rect 69673 679677 69707 679711
rect 74549 679813 74583 679847
rect 74549 679677 74583 679711
rect 88993 679813 89027 679847
rect 88993 679677 89027 679711
rect 93869 679813 93903 679847
rect 93869 679677 93903 679711
rect 108313 679813 108347 679847
rect 108313 679677 108347 679711
rect 113189 679813 113223 679847
rect 113189 679677 113223 679711
rect 127633 679813 127667 679847
rect 127633 679677 127667 679711
rect 132509 679813 132543 679847
rect 132509 679677 132543 679711
rect 146953 679813 146987 679847
rect 146953 679677 146987 679711
rect 151829 679813 151863 679847
rect 151829 679677 151863 679711
rect 166273 679813 166307 679847
rect 166273 679677 166307 679711
rect 171149 679813 171183 679847
rect 171149 679677 171183 679711
rect 185593 679813 185627 679847
rect 185593 679677 185627 679711
rect 190469 679813 190503 679847
rect 190469 679677 190503 679711
rect 204913 679813 204947 679847
rect 204913 679677 204947 679711
rect 209789 679813 209823 679847
rect 231961 680357 231995 680391
rect 222025 679813 222059 679847
rect 216597 679745 216631 679779
rect 380081 680357 380115 680391
rect 222117 679745 222151 679779
rect 231777 679745 231811 679779
rect 231961 679745 231995 679779
rect 364809 680289 364843 680323
rect 209789 679677 209823 679711
rect 222209 679677 222243 679711
rect 222209 679541 222243 679575
rect 231777 679541 231811 679575
rect 364809 679541 364843 679575
rect 370237 680289 370271 680323
rect 370237 679541 370271 679575
rect 394525 680357 394559 680391
rect 394525 680221 394559 680255
rect 394709 680357 394743 680391
rect 380081 679541 380115 679575
rect 394709 679541 394743 679575
rect 403173 680357 403207 680391
rect 412741 680357 412775 680391
rect 412649 680221 412683 680255
rect 412649 680017 412683 680051
rect 403173 679541 403207 679575
rect 412741 679541 412775 679575
rect 418629 680357 418663 680391
rect 428013 680357 428047 680391
rect 428013 679949 428047 679983
rect 428197 680357 428231 680391
rect 418629 679541 418663 679575
rect 437765 680357 437799 680391
rect 434729 679949 434763 679983
rect 434729 679813 434763 679847
rect 428197 679541 428231 679575
rect 437765 679541 437799 679575
rect 443561 680357 443595 680391
rect 207029 679133 207063 679167
rect 451381 680357 451415 680391
rect 451289 680221 451323 680255
rect 444297 680085 444331 680119
rect 451289 679949 451323 679983
rect 444297 679813 444331 679847
rect 451381 679541 451415 679575
rect 457177 680357 457211 680391
rect 466561 680357 466595 680391
rect 461593 680221 461627 680255
rect 461593 679949 461627 679983
rect 457177 679541 457211 679575
rect 474749 680357 474783 680391
rect 469597 680221 469631 680255
rect 469597 680085 469631 680119
rect 494069 680357 494103 680391
rect 481005 680289 481039 680323
rect 477969 680153 478003 680187
rect 478153 680153 478187 680187
rect 474749 680017 474783 680051
rect 481097 679949 481131 679983
rect 481189 680289 481223 680323
rect 466561 679541 466595 679575
rect 485789 680289 485823 680323
rect 485697 680085 485731 680119
rect 485605 679881 485639 679915
rect 481189 679541 481223 679575
rect 489745 680289 489779 680323
rect 489745 679949 489779 679983
rect 490481 680221 490515 680255
rect 494069 679949 494103 679983
rect 495449 680357 495483 680391
rect 490481 679813 490515 679847
rect 485789 679541 485823 679575
rect 502257 680357 502291 680391
rect 500233 680221 500267 680255
rect 500233 679813 500267 679847
rect 495449 679541 495483 679575
rect 505937 680357 505971 680391
rect 515413 680357 515447 680391
rect 509801 680221 509835 680255
rect 506489 680085 506523 680119
rect 506489 679881 506523 679915
rect 509801 679745 509835 679779
rect 505937 679541 505971 679575
rect 522129 680357 522163 680391
rect 519553 680153 519587 680187
rect 516333 680085 516367 680119
rect 519553 679813 519587 679847
rect 516333 679745 516367 679779
rect 515413 679541 515447 679575
rect 524429 680357 524463 680391
rect 534365 680357 534399 680391
rect 533997 680221 534031 680255
rect 529121 680153 529155 680187
rect 529029 680085 529063 680119
rect 529213 680085 529247 680119
rect 529213 679881 529247 679915
rect 529121 679813 529155 679847
rect 529029 679745 529063 679779
rect 533997 679745 534031 679779
rect 524429 679541 524463 679575
rect 543749 680357 543783 680391
rect 538873 680221 538907 680255
rect 538873 679881 538907 679915
rect 543749 679745 543783 679779
rect 544025 680357 544059 680391
rect 534365 679541 534399 679575
rect 553501 680289 553535 680323
rect 546877 680221 546911 680255
rect 546877 679881 546911 679915
rect 553409 680221 553443 680255
rect 553501 679813 553535 679847
rect 554881 680289 554915 680323
rect 553409 679745 553443 679779
rect 544025 679541 544059 679575
rect 522129 679269 522163 679303
rect 502257 679201 502291 679235
rect 443561 679133 443595 679167
rect 557733 680085 557767 680119
rect 559205 680289 559239 680323
rect 559205 679949 559239 679983
rect 560769 680289 560803 680323
rect 554881 679133 554915 679167
rect 561597 680289 561631 680323
rect 561597 679881 561631 679915
rect 561781 680289 561815 680323
rect 561781 679813 561815 679847
rect 561873 680289 561907 680323
rect 561873 679269 561907 679303
rect 562517 680289 562551 680323
rect 562517 679201 562551 679235
rect 560769 679133 560803 679167
rect 569969 659209 570003 659243
rect 569969 654041 570003 654075
rect 1961 648057 1995 648091
rect 1869 642617 1903 642651
rect 1961 639285 1995 639319
rect 1869 633437 1903 633471
rect 1869 602361 1903 602395
rect 1777 601953 1811 601987
rect 1685 601069 1719 601103
rect 1685 600525 1719 600559
rect 1777 599709 1811 599743
rect 1961 602089 1995 602123
rect 1961 599845 1995 599879
rect 1869 596989 1903 597023
rect 1869 580465 1903 580499
rect 1869 566593 1903 566627
rect 1961 580193 1995 580227
rect 1777 565505 1811 565539
rect 1685 564417 1719 564451
rect 1685 563397 1719 563431
rect 1777 563125 1811 563159
rect 1869 561085 1903 561119
rect 1961 563737 1995 563771
rect 569969 552041 570003 552075
rect 569969 551021 570003 551055
rect 1961 547689 1995 547723
rect 570061 531097 570095 531131
rect 569969 530961 570003 530995
rect 1961 529193 1995 529227
rect 1869 527697 1903 527731
rect 1777 527153 1811 527187
rect 1685 527085 1719 527119
rect 1685 526949 1719 526983
rect 1685 526473 1719 526507
rect 1685 526133 1719 526167
rect 1777 522461 1811 522495
rect 1869 522325 1903 522359
rect 569969 528853 570003 528887
rect 570061 528717 570095 528751
rect 569969 522597 570003 522631
rect 570061 522461 570095 522495
rect 570061 521033 570095 521067
rect 569969 518449 570003 518483
rect 1961 510629 1995 510663
rect 1961 510017 1995 510051
rect 1869 509881 1903 509915
rect 1593 507297 1627 507331
rect 1501 507161 1535 507195
rect 1501 502197 1535 502231
rect 1777 506073 1811 506107
rect 1777 504849 1811 504883
rect 1869 504441 1903 504475
rect 1777 504101 1811 504135
rect 1593 501789 1627 501823
rect 1685 502265 1719 502299
rect 1777 497505 1811 497539
rect 569969 505121 570003 505155
rect 570061 504169 570095 504203
rect 570061 503149 570095 503183
rect 569969 503013 570003 503047
rect 1961 497505 1995 497539
rect 1685 493357 1719 493391
rect 1685 483701 1719 483735
rect 1961 474657 1995 474691
rect 1869 474045 1903 474079
rect 1685 464933 1719 464967
rect 1777 472073 1811 472107
rect 1869 467585 1903 467619
rect 1593 450721 1627 450755
rect 1409 449905 1443 449939
rect 1593 449021 1627 449055
rect 1593 448749 1627 448783
rect 1961 462349 1995 462383
rect 569969 468537 570003 468571
rect 570153 468265 570187 468299
rect 570061 467041 570095 467075
rect 569969 466565 570003 466599
rect 570153 466837 570187 466871
rect 570245 467585 570279 467619
rect 570245 466565 570279 466599
rect 570061 465477 570095 465511
rect 570337 465477 570371 465511
rect 570153 465341 570187 465375
rect 570061 465205 570095 465239
rect 570061 463573 570095 463607
rect 570337 463845 570371 463879
rect 570153 462757 570187 462791
rect 569969 461669 570003 461703
rect 569969 461397 570003 461431
rect 1961 454597 1995 454631
rect 1685 448681 1719 448715
rect 1777 450041 1811 450075
rect 1593 448477 1627 448511
rect 1409 447933 1443 447967
rect 1777 447797 1811 447831
rect 1869 449157 1903 449191
rect 1777 442289 1811 442323
rect 1777 441405 1811 441439
rect 1869 440929 1903 440963
rect 1961 439161 1995 439195
rect 570061 441609 570095 441643
rect 570061 436781 570095 436815
rect 1961 434197 1995 434231
rect 1961 425697 1995 425731
rect 569969 432497 570003 432531
rect 569969 418149 570003 418183
rect 569969 418013 570003 418047
rect 1961 414953 1995 414987
rect 1961 407269 1995 407303
rect 1961 405637 1995 405671
rect 1869 405569 1903 405603
rect 1869 393941 1903 393975
rect 569969 402237 570003 402271
rect 569969 399517 570003 399551
rect 1961 393465 1995 393499
rect 570061 396797 570095 396831
rect 1777 387345 1811 387379
rect 1409 387073 1443 387107
rect 1409 381157 1443 381191
rect 1593 381429 1627 381463
rect 1593 379117 1627 379151
rect 1685 380681 1719 380715
rect 1685 378981 1719 379015
rect 1869 387209 1903 387243
rect 1961 387073 1995 387107
rect 569969 393669 570003 393703
rect 570245 394961 570279 394995
rect 570061 392309 570095 392343
rect 570153 393805 570187 393839
rect 569969 389861 570003 389895
rect 570153 389045 570187 389079
rect 570337 393125 570371 393159
rect 570337 389997 570371 390031
rect 570245 388501 570279 388535
rect 569877 382653 569911 382687
rect 569969 382789 570003 382823
rect 1961 381429 1995 381463
rect 1869 380681 1903 380715
rect 1777 376737 1811 376771
rect 569969 376669 570003 376703
rect 570061 381837 570095 381871
rect 570061 376533 570095 376567
rect 570245 376669 570279 376703
rect 1961 370617 1995 370651
rect 1685 370481 1719 370515
rect 1409 369257 1443 369291
rect 1869 370345 1903 370379
rect 1685 367761 1719 367795
rect 1777 370209 1811 370243
rect 1409 358037 1443 358071
rect 1777 358241 1811 358275
rect 1501 336005 1535 336039
rect 1409 334169 1443 334203
rect 1409 333421 1443 333455
rect 1501 331857 1535 331891
rect 1501 326485 1535 326519
rect 1317 315129 1351 315163
rect 1225 312137 1259 312171
rect 1685 345729 1719 345763
rect 1869 358105 1903 358139
rect 1869 353209 1903 353243
rect 1869 352937 1903 352971
rect 1777 345661 1811 345695
rect 1869 340833 1903 340867
rect 1777 340697 1811 340731
rect 570153 369733 570187 369767
rect 569969 369393 570003 369427
rect 569969 368305 570003 368339
rect 570061 359533 570095 359567
rect 570061 358241 570095 358275
rect 569969 358105 570003 358139
rect 569969 357629 570003 357663
rect 569969 353957 570003 353991
rect 569969 353617 570003 353651
rect 569969 352597 570003 352631
rect 570061 352461 570095 352495
rect 569969 348925 570003 348959
rect 570429 367761 570463 367795
rect 570337 359873 570371 359907
rect 570337 358037 570371 358071
rect 570245 357629 570279 357663
rect 570245 352461 570279 352495
rect 570521 359125 570555 359159
rect 570521 353685 570555 353719
rect 570429 352325 570463 352359
rect 570245 347973 570279 348007
rect 570153 347701 570187 347735
rect 569969 344845 570003 344879
rect 1961 340221 1995 340255
rect 569969 342193 570003 342227
rect 1869 336005 1903 336039
rect 1961 338045 1995 338079
rect 1777 334033 1811 334067
rect 1777 331993 1811 332027
rect 1685 329749 1719 329783
rect 1777 331857 1811 331891
rect 1593 326349 1627 326383
rect 1501 312681 1535 312715
rect 1593 318937 1627 318971
rect 1501 312409 1535 312443
rect 1409 312273 1443 312307
rect 1409 312137 1443 312171
rect 1317 311797 1351 311831
rect 1409 312001 1443 312035
rect 1225 304113 1259 304147
rect 1317 304521 1351 304555
rect 1225 303365 1259 303399
rect 1133 298061 1167 298095
rect 1133 294457 1167 294491
rect 1593 311661 1627 311695
rect 1685 313905 1719 313939
rect 569969 331245 570003 331279
rect 569969 331041 570003 331075
rect 1961 329137 1995 329171
rect 569877 329545 569911 329579
rect 1869 326485 1903 326519
rect 1869 326349 1903 326383
rect 570153 330497 570187 330531
rect 570061 329681 570095 329715
rect 570061 324989 570095 325023
rect 569969 321113 570003 321147
rect 570245 329409 570279 329443
rect 570337 329273 570371 329307
rect 570337 327029 570371 327063
rect 570245 325669 570279 325703
rect 570153 321113 570187 321147
rect 570245 325533 570279 325567
rect 570061 320977 570095 321011
rect 569969 320841 570003 320875
rect 1961 319141 1995 319175
rect 570337 321113 570371 321147
rect 569969 320705 570003 320739
rect 569969 317917 570003 317951
rect 569969 315945 570003 315979
rect 1961 314993 1995 315027
rect 570153 320705 570187 320739
rect 1869 313905 1903 313939
rect 1961 312681 1995 312715
rect 1777 312001 1811 312035
rect 1869 312545 1903 312579
rect 1685 311525 1719 311559
rect 1961 309825 1995 309859
rect 1869 309621 1903 309655
rect 1409 303977 1443 304011
rect 1501 304385 1535 304419
rect 1317 298061 1351 298095
rect 1225 293097 1259 293131
rect 1317 296021 1351 296055
rect 1961 306629 1995 306663
rect 1685 305609 1719 305643
rect 1777 305473 1811 305507
rect 1777 303229 1811 303263
rect 1869 305337 1903 305371
rect 1685 301461 1719 301495
rect 1869 296225 1903 296259
rect 1593 296021 1627 296055
rect 1777 296089 1811 296123
rect 1501 294593 1535 294627
rect 1685 295817 1719 295851
rect 1501 294457 1535 294491
rect 1317 292145 1351 292179
rect 1409 293369 1443 293403
rect 1317 287113 1351 287147
rect 1501 287113 1535 287147
rect 1593 292145 1627 292179
rect 1409 284733 1443 284767
rect 1317 284597 1351 284631
rect 1501 284325 1535 284359
rect 1593 286977 1627 287011
rect 1409 283917 1443 283951
rect 1409 283441 1443 283475
rect 1869 295953 1903 295987
rect 1869 283917 1903 283951
rect 1777 283373 1811 283407
rect 1869 283441 1903 283475
rect 1593 283237 1627 283271
rect 1685 273921 1719 273955
rect 1685 270181 1719 270215
rect 1777 269773 1811 269807
rect 581 266577 615 266611
rect 569969 315809 570003 315843
rect 569969 315605 570003 315639
rect 570061 309077 570095 309111
rect 569969 306153 570003 306187
rect 570245 320705 570279 320739
rect 570245 315469 570279 315503
rect 570337 314721 570371 314755
rect 570521 314721 570555 314755
rect 570521 309213 570555 309247
rect 570153 304997 570187 305031
rect 570245 309145 570279 309179
rect 569969 304249 570003 304283
rect 570061 302889 570095 302923
rect 569969 301869 570003 301903
rect 569969 300849 570003 300883
rect 570061 300237 570095 300271
rect 570061 300101 570095 300135
rect 569969 300033 570003 300067
rect 569969 298537 570003 298571
rect 570061 296565 570095 296599
rect 570429 306969 570463 307003
rect 570245 302889 570279 302923
rect 570337 303841 570371 303875
rect 570245 302753 570279 302787
rect 570429 301869 570463 301903
rect 570521 304929 570555 304963
rect 570337 300373 570371 300407
rect 570429 301121 570463 301155
rect 570245 298401 570279 298435
rect 570153 296157 570187 296191
rect 570337 296565 570371 296599
rect 570153 296021 570187 296055
rect 569969 292757 570003 292791
rect 570245 295137 570279 295171
rect 569969 292553 570003 292587
rect 570153 291941 570187 291975
rect 569969 288269 570003 288303
rect 570061 289765 570095 289799
rect 570153 289765 570187 289799
rect 569969 285617 570003 285651
rect 569969 285481 570003 285515
rect 569969 285141 570003 285175
rect 569969 283713 570003 283747
rect 570521 296089 570555 296123
rect 570429 292417 570463 292451
rect 570337 291941 570371 291975
rect 570521 289629 570555 289663
rect 570245 288133 570279 288167
rect 570429 288133 570463 288167
rect 570245 285617 570279 285651
rect 570153 285345 570187 285379
rect 570061 283577 570095 283611
rect 570245 283577 570279 283611
rect 570337 284937 570371 284971
rect 570153 274329 570187 274363
rect 570245 283441 570279 283475
rect 569969 273989 570003 274023
rect 1961 269365 1995 269399
rect 1777 264129 1811 264163
rect 1869 266441 1903 266475
rect 581 251821 615 251855
rect 857 261545 891 261579
rect 857 251821 891 251855
rect 1133 261477 1167 261511
rect 1777 261477 1811 261511
rect 1777 251821 1811 251855
rect 1133 242029 1167 242063
rect 1501 250257 1535 250291
rect 1685 242233 1719 242267
rect 1501 238289 1535 238323
rect 1593 242097 1627 242131
rect 1501 238153 1535 238187
rect 857 221697 891 221731
rect 305 221017 339 221051
rect 305 199461 339 199495
rect 673 201841 707 201875
rect 1685 237949 1719 237983
rect 1777 242165 1811 242199
rect 1961 264673 1995 264707
rect 1961 250121 1995 250155
rect 570061 273853 570095 273887
rect 569969 273037 570003 273071
rect 569969 271541 570003 271575
rect 570153 270453 570187 270487
rect 570337 283373 570371 283407
rect 570245 270317 570279 270351
rect 570337 274329 570371 274363
rect 570337 270045 570371 270079
rect 570521 283509 570555 283543
rect 570613 284801 570647 284835
rect 570521 277253 570555 277287
rect 570705 274465 570739 274499
rect 570705 272901 570739 272935
rect 570613 272493 570647 272527
rect 570521 270997 570555 271031
rect 570429 269909 570463 269943
rect 570061 269773 570095 269807
rect 569969 267257 570003 267291
rect 569969 259845 570003 259879
rect 570061 266373 570095 266407
rect 569969 254745 570003 254779
rect 570061 250461 570095 250495
rect 570153 265897 570187 265931
rect 569969 245973 570003 246007
rect 570061 246653 570095 246687
rect 569877 245701 569911 245735
rect 569969 245701 570003 245735
rect 569877 245361 569911 245395
rect 1961 243049 1995 243083
rect 1961 242913 1995 242947
rect 1869 242097 1903 242131
rect 1961 242505 1995 242539
rect 1777 228361 1811 228395
rect 1869 241961 1903 241995
rect 1593 222581 1627 222615
rect 1317 221493 1351 221527
rect 1501 221493 1535 221527
rect 1685 221493 1719 221527
rect 1593 219929 1627 219963
rect 1317 212857 1351 212891
rect 1409 216801 1443 216835
rect 1317 209933 1351 209967
rect 1133 207757 1167 207791
rect 1041 204901 1075 204935
rect 857 199461 891 199495
rect 1041 200821 1075 200855
rect 1041 198849 1075 198883
rect 1133 197897 1167 197931
rect 1225 207689 1259 207723
rect 1133 197761 1167 197795
rect 857 196197 891 196231
rect 949 197625 983 197659
rect 949 195925 983 195959
rect 1593 207757 1627 207791
rect 1501 204697 1535 204731
rect 1501 200821 1535 200855
rect 1409 198033 1443 198067
rect 1501 200685 1535 200719
rect 1317 197897 1351 197931
rect 1317 195789 1351 195823
rect 1225 195041 1259 195075
rect 1133 194701 1167 194735
rect 673 193953 707 193987
rect 1593 198713 1627 198747
rect 1593 198169 1627 198203
rect 1501 195177 1535 195211
rect 1593 198033 1627 198067
rect 1409 193953 1443 193987
rect 1409 189737 1443 189771
rect 1317 189193 1351 189227
rect 1225 188921 1259 188955
rect 305 182801 339 182835
rect 213 174573 247 174607
rect 305 170969 339 171003
rect 489 179197 523 179231
rect 1225 176613 1259 176647
rect 1317 176477 1351 176511
rect 1501 189601 1535 189635
rect 1501 188513 1535 188547
rect 1501 188377 1535 188411
rect 1501 176749 1535 176783
rect 1409 176341 1443 176375
rect 1777 221289 1811 221323
rect 1869 222581 1903 222615
rect 1777 218297 1811 218331
rect 1777 217685 1811 217719
rect 1777 217413 1811 217447
rect 570061 243525 570095 243559
rect 570245 263993 570279 264027
rect 570245 259573 570279 259607
rect 570245 250937 570279 250971
rect 570521 250597 570555 250631
rect 570245 246517 570279 246551
rect 570337 247265 570371 247299
rect 570245 245973 570279 246007
rect 570245 243661 570279 243695
rect 570061 236045 570095 236079
rect 569969 230197 570003 230231
rect 1961 221493 1995 221527
rect 569969 229653 570003 229687
rect 1869 205785 1903 205819
rect 1961 221357 1995 221391
rect 1685 197489 1719 197523
rect 1777 205649 1811 205683
rect 1685 195653 1719 195687
rect 1869 200685 1903 200719
rect 1869 198169 1903 198203
rect 569969 228701 570003 228735
rect 570153 229857 570187 229891
rect 570245 229721 570279 229755
rect 570521 245361 570555 245395
rect 570337 228701 570371 228735
rect 570429 239445 570463 239479
rect 570061 227001 570095 227035
rect 570061 226865 570095 226899
rect 570521 233665 570555 233699
rect 570521 229245 570555 229279
rect 570061 205445 570095 205479
rect 570153 214557 570187 214591
rect 569969 205173 570003 205207
rect 569969 204901 570003 204935
rect 570061 204765 570095 204799
rect 570061 203677 570095 203711
rect 570061 203133 570095 203167
rect 570337 225777 570371 225811
rect 570337 214625 570371 214659
rect 570245 205445 570279 205479
rect 570245 204425 570279 204459
rect 570337 203541 570371 203575
rect 570153 202997 570187 203031
rect 569969 202589 570003 202623
rect 1961 198033 1995 198067
rect 1961 197625 1995 197659
rect 1961 196333 1995 196367
rect 1869 196061 1903 196095
rect 1685 182869 1719 182903
rect 1777 195177 1811 195211
rect 1869 195109 1903 195143
rect 1869 186473 1903 186507
rect 1777 179061 1811 179095
rect 1869 179605 1903 179639
rect 1777 178381 1811 178415
rect 1593 175933 1627 175967
rect 1685 176953 1719 176987
rect 489 170289 523 170323
rect 1501 175593 1535 175627
rect 213 165869 247 165903
rect 305 167773 339 167807
rect 949 167637 983 167671
rect 857 166889 891 166923
rect 765 159613 799 159647
rect 673 153901 707 153935
rect 397 153833 431 153867
rect 397 146965 431 146999
rect 857 159273 891 159307
rect 1225 167637 1259 167671
rect 1041 167365 1075 167399
rect 1041 159137 1075 159171
rect 1133 166141 1167 166175
rect 949 154785 983 154819
rect 949 154037 983 154071
rect 1317 167229 1351 167263
rect 1409 166413 1443 166447
rect 1409 165461 1443 165495
rect 1777 176205 1811 176239
rect 570153 193885 570187 193919
rect 1961 179197 1995 179231
rect 569969 192457 570003 192491
rect 1961 177633 1995 177667
rect 570061 192185 570095 192219
rect 570061 188377 570095 188411
rect 569969 177429 570003 177463
rect 570061 180421 570095 180455
rect 1961 176205 1995 176239
rect 569969 177293 570003 177327
rect 1685 173009 1719 173043
rect 1317 159409 1351 159443
rect 1593 167977 1627 168011
rect 1501 163557 1535 163591
rect 1593 163421 1627 163455
rect 1685 167229 1719 167263
rect 1501 159477 1535 159511
rect 1593 163285 1627 163319
rect 1409 159341 1443 159375
rect 1225 153901 1259 153935
rect 1409 159205 1443 159239
rect 1225 153765 1259 153799
rect 949 150093 983 150127
rect 1041 150229 1075 150263
rect 765 146965 799 146999
rect 949 146965 983 146999
rect 673 146149 707 146183
rect 857 146285 891 146319
rect 305 145605 339 145639
rect 581 142953 615 142987
rect 581 141593 615 141627
rect 765 141185 799 141219
rect 305 138941 339 138975
rect 673 132073 707 132107
rect 581 130577 615 130611
rect 305 130237 339 130271
rect 489 130373 523 130407
rect 489 129421 523 129455
rect 949 142817 983 142851
rect 1225 146965 1259 146999
rect 1317 146285 1351 146319
rect 1317 146149 1351 146183
rect 1041 141117 1075 141151
rect 1133 145673 1167 145707
rect 765 130373 799 130407
rect 857 140641 891 140675
rect 673 126225 707 126259
rect 765 130237 799 130271
rect 673 126021 707 126055
rect 949 139077 983 139111
rect 1133 138873 1167 138907
rect 949 138737 983 138771
rect 1133 138669 1167 138703
rect 949 134521 983 134555
rect 949 128333 983 128367
rect 1041 126633 1075 126667
rect 1041 126497 1075 126531
rect 857 126089 891 126123
rect 949 126225 983 126259
rect 765 117453 799 117487
rect 1041 119561 1075 119595
rect 949 117385 983 117419
rect 1041 117453 1075 117487
rect 765 109701 799 109735
rect 581 109293 615 109327
rect 673 109429 707 109463
rect 673 109157 707 109191
rect 765 108749 799 108783
rect 1041 115209 1075 115243
rect 949 115073 983 115107
rect 949 108885 983 108919
rect 1041 110993 1075 111027
rect 1041 108069 1075 108103
rect 857 107661 891 107695
rect 1225 134453 1259 134487
rect 1225 108341 1259 108375
rect 1501 156349 1535 156383
rect 1501 150229 1535 150263
rect 1501 150093 1535 150127
rect 1685 159613 1719 159647
rect 1869 176069 1903 176103
rect 1869 163557 1903 163591
rect 1961 169065 1995 169099
rect 1777 159545 1811 159579
rect 570429 192729 570463 192763
rect 570337 192049 570371 192083
rect 570153 179809 570187 179843
rect 570245 191913 570279 191947
rect 570061 176817 570095 176851
rect 570153 178041 570187 178075
rect 569969 174913 570003 174947
rect 569969 163693 570003 163727
rect 570061 169065 570095 169099
rect 569969 163489 570003 163523
rect 1593 148733 1627 148767
rect 1685 159477 1719 159511
rect 1777 159409 1811 159443
rect 1593 145945 1627 145979
rect 1685 148597 1719 148631
rect 1501 141457 1535 141491
rect 1501 141321 1535 141355
rect 1409 141253 1443 141287
rect 1409 138737 1443 138771
rect 1317 107185 1351 107219
rect 1409 138601 1443 138635
rect 1133 96033 1167 96067
rect 1317 98277 1351 98311
rect 1041 94673 1075 94707
rect 949 92021 983 92055
rect 1133 93993 1167 94027
rect 1225 93585 1259 93619
rect 1317 93517 1351 93551
rect 1225 91749 1259 91783
rect 1317 93381 1351 93415
rect 1133 91613 1167 91647
rect 1317 91477 1351 91511
rect 1501 137921 1535 137955
rect 1501 134589 1535 134623
rect 1869 159205 1903 159239
rect 1961 163421 1995 163455
rect 1869 159069 1903 159103
rect 569969 158729 570003 158763
rect 569969 157981 570003 158015
rect 569969 157845 570003 157879
rect 569969 149277 570003 149311
rect 1961 146965 1995 146999
rect 569969 148325 570003 148359
rect 1777 146353 1811 146387
rect 1777 146217 1811 146251
rect 1869 145877 1903 145911
rect 1869 143089 1903 143123
rect 1777 140709 1811 140743
rect 1869 142953 1903 142987
rect 1777 139961 1811 139995
rect 1777 138941 1811 138975
rect 1777 138805 1811 138839
rect 1777 138261 1811 138295
rect 1593 131121 1627 131155
rect 1685 134521 1719 134555
rect 1593 130849 1627 130883
rect 1593 129149 1627 129183
rect 1593 128877 1627 128911
rect 1593 126497 1627 126531
rect 1501 126225 1535 126259
rect 1593 126361 1627 126395
rect 1501 126089 1535 126123
rect 1501 116433 1535 116467
rect 1501 115209 1535 115243
rect 1777 134385 1811 134419
rect 1685 124865 1719 124899
rect 1777 133433 1811 133467
rect 1869 133297 1903 133331
rect 569969 134521 570003 134555
rect 570429 191505 570463 191539
rect 570337 178041 570371 178075
rect 570245 175185 570279 175219
rect 570245 161993 570279 162027
rect 570153 157981 570187 158015
rect 570521 177429 570555 177463
rect 570429 171921 570463 171955
rect 570521 169065 570555 169099
rect 570429 162197 570463 162231
rect 570337 158729 570371 158763
rect 570521 157641 570555 157675
rect 570337 157369 570371 157403
rect 570337 155601 570371 155635
rect 570337 153901 570371 153935
rect 570245 153425 570279 153459
rect 570521 154989 570555 155023
rect 570521 149549 570555 149583
rect 570245 147917 570279 147951
rect 570337 148461 570371 148495
rect 570153 147645 570187 147679
rect 570061 134181 570095 134215
rect 570521 146965 570555 146999
rect 570337 133093 570371 133127
rect 1869 124933 1903 124967
rect 1961 131053 1995 131087
rect 1961 124933 1995 124967
rect 1593 108613 1627 108647
rect 1685 124729 1719 124763
rect 1777 124729 1811 124763
rect 1501 108477 1535 108511
rect 1685 108069 1719 108103
rect 1777 119561 1811 119595
rect 1961 117997 1995 118031
rect 1777 102561 1811 102595
rect 1869 117793 1903 117827
rect 1777 98413 1811 98447
rect 1685 98277 1719 98311
rect 1593 96033 1627 96067
rect 1409 91341 1443 91375
rect 1501 93517 1535 93551
rect 1041 90389 1075 90423
rect 1409 90389 1443 90423
rect 1225 88757 1259 88791
rect 949 86105 983 86139
rect 1041 87601 1075 87635
rect 949 84745 983 84779
rect 1041 83589 1075 83623
rect 1133 84609 1167 84643
rect 949 82093 983 82127
rect 1317 83793 1351 83827
rect 1317 80733 1351 80767
rect 1225 80665 1259 80699
rect 1133 70397 1167 70431
rect 1317 70261 1351 70295
rect 1225 69581 1259 69615
rect 1041 67473 1075 67507
rect 949 67201 983 67235
rect 765 66725 799 66759
rect 765 64617 799 64651
rect 857 66589 891 66623
rect 949 63121 983 63155
rect 1041 62849 1075 62883
rect 1133 65433 1167 65467
rect 1225 62713 1259 62747
rect 1133 62237 1167 62271
rect 857 57885 891 57919
rect 1225 57069 1259 57103
rect 1225 55845 1259 55879
rect 1501 87601 1535 87635
rect 1501 87329 1535 87363
rect 1501 80801 1535 80835
rect 1409 69445 1443 69479
rect 1501 80665 1535 80699
rect 1409 69309 1443 69343
rect 1961 107049 1995 107083
rect 1869 96237 1903 96271
rect 1961 98141 1995 98175
rect 1869 94741 1903 94775
rect 1869 93245 1903 93279
rect 1777 91205 1811 91239
rect 1869 93109 1903 93143
rect 1685 87329 1719 87363
rect 1685 86309 1719 86343
rect 1685 80937 1719 80971
rect 1777 86173 1811 86207
rect 1593 72301 1627 72335
rect 1685 80801 1719 80835
rect 1501 66929 1535 66963
rect 1593 71961 1627 71995
rect 1961 88757 1995 88791
rect 1869 72437 1903 72471
rect 1961 86377 1995 86411
rect 1685 69581 1719 69615
rect 1777 72301 1811 72335
rect 1685 69445 1719 69479
rect 1685 66317 1719 66351
rect 1409 62985 1443 63019
rect 1409 56729 1443 56763
rect 1409 55165 1443 55199
rect 1317 52717 1351 52751
rect 1685 65841 1719 65875
rect 1593 65433 1627 65467
rect 1685 64753 1719 64787
rect 1501 52581 1535 52615
rect 1593 62713 1627 62747
rect 29 50405 63 50439
rect 1041 50337 1075 50371
rect 1409 45509 1443 45543
rect 1593 45509 1627 45543
rect 570061 77265 570095 77299
rect 1961 66453 1995 66487
rect 569969 76313 570003 76347
rect 1869 65433 1903 65467
rect 1961 66317 1995 66351
rect 1869 64753 1903 64787
rect 1869 50405 1903 50439
rect 569877 58837 569911 58871
rect 569969 75905 570003 75939
rect 569969 56933 570003 56967
rect 570153 76721 570187 76755
rect 570245 76585 570279 76619
rect 570245 75905 570279 75939
rect 570337 76177 570371 76211
rect 570337 74817 570371 74851
rect 570429 73593 570463 73627
rect 570429 72981 570463 73015
rect 570521 73389 570555 73423
rect 570337 72437 570371 72471
rect 570337 68017 570371 68051
rect 570521 66113 570555 66147
rect 570521 65977 570555 66011
rect 570337 60741 570371 60775
rect 570429 64957 570463 64991
rect 570245 59925 570279 59959
rect 570429 58701 570463 58735
rect 570153 56661 570187 56695
rect 570521 56593 570555 56627
rect 570061 53737 570095 53771
rect 1777 47617 1811 47651
rect 1409 43061 1443 43095
rect 1777 47481 1811 47515
rect 1593 42789 1627 42823
rect 1685 43469 1719 43503
rect 1041 37009 1075 37043
rect 1133 39457 1167 39491
rect 29 34969 63 35003
rect 1041 35377 1075 35411
rect 673 33541 707 33575
rect 121 24225 155 24259
rect 121 16949 155 16983
rect 581 24021 615 24055
rect 1409 39321 1443 39355
rect 1317 35649 1351 35683
rect 1133 29597 1167 29631
rect 1225 35513 1259 35547
rect 1041 29529 1075 29563
rect 949 28849 983 28883
rect 949 23749 983 23783
rect 1041 27081 1075 27115
rect 673 22049 707 22083
rect 949 20009 983 20043
rect 765 18445 799 18479
rect 581 15453 615 15487
rect 673 16541 707 16575
rect 581 10353 615 10387
rect 489 8653 523 8687
rect 765 12053 799 12087
rect 857 17085 891 17119
rect 673 10081 707 10115
rect 765 10421 799 10455
rect 857 10285 891 10319
rect 1041 18581 1075 18615
rect 1041 17901 1075 17935
rect 1225 27217 1259 27251
rect 1593 29665 1627 29699
rect 1409 28985 1443 29019
rect 1501 29461 1535 29495
rect 1409 28305 1443 28339
rect 1501 27081 1535 27115
rect 1409 22185 1443 22219
rect 1501 21573 1535 21607
rect 1225 15317 1259 15351
rect 1317 16405 1351 16439
rect 1133 15181 1167 15215
rect 1041 14569 1075 14603
rect 1133 14773 1167 14807
rect 1041 13345 1075 13379
rect 1133 14433 1167 14467
rect 949 7497 983 7531
rect 1041 10353 1075 10387
rect 765 3689 799 3723
rect 581 1717 615 1751
rect 1041 1649 1075 1683
rect 1225 13481 1259 13515
rect 1593 18377 1627 18411
rect 1501 16065 1535 16099
rect 1593 18241 1627 18275
rect 1501 15929 1535 15963
rect 1501 14637 1535 14671
rect 1317 12325 1351 12359
rect 1409 12325 1443 12359
rect 1225 3281 1259 3315
rect 1317 11849 1351 11883
rect 1409 10489 1443 10523
rect 1317 1513 1351 1547
rect 1409 10353 1443 10387
rect 1133 1309 1167 1343
rect 1409 1037 1443 1071
rect 1961 47617 1995 47651
rect 1961 43469 1995 43503
rect 1777 39185 1811 39219
rect 1869 39321 1903 39355
rect 570521 43265 570555 43299
rect 1961 29869 1995 29903
rect 569969 42313 570003 42347
rect 1961 29733 1995 29767
rect 1869 29597 1903 29631
rect 1869 20077 1903 20111
rect 1685 17085 1719 17119
rect 1777 19941 1811 19975
rect 1593 10421 1627 10455
rect 1685 16949 1719 16983
rect 1777 12325 1811 12359
rect 1685 10353 1719 10387
rect 1777 12189 1811 12223
rect 1593 10285 1627 10319
rect 1593 1173 1627 1207
rect 1685 10217 1719 10251
rect 1685 1105 1719 1139
rect 1501 357 1535 391
rect 489 289 523 323
rect 1961 18853 1995 18887
rect 1961 18717 1995 18751
rect 570245 42177 570279 42211
rect 570061 41633 570095 41667
rect 569969 40953 570003 40987
rect 569969 39661 570003 39695
rect 570153 41089 570187 41123
rect 570153 39865 570187 39899
rect 570061 39389 570095 39423
rect 570153 39729 570187 39763
rect 569969 27897 570003 27931
rect 569969 23069 570003 23103
rect 570061 25721 570095 25755
rect 1961 9401 1995 9435
rect 1869 3689 1903 3723
rect 1961 8721 1995 8755
rect 570337 41769 570371 41803
rect 570429 40409 570463 40443
rect 570429 40001 570463 40035
rect 570337 39729 570371 39763
rect 570521 39049 570555 39083
rect 570613 40273 570647 40307
rect 570613 34765 570647 34799
rect 570245 27897 570279 27931
rect 570337 31025 570371 31059
rect 570245 26469 570279 26503
rect 570245 23749 570279 23783
rect 570153 23205 570187 23239
rect 570153 23069 570187 23103
rect 570153 17629 570187 17663
rect 570061 14705 570095 14739
rect 569969 8109 570003 8143
rect 570429 25517 570463 25551
rect 570429 24157 570463 24191
rect 570337 7837 570371 7871
rect 124321 3077 124355 3111
rect 177957 3077 177991 3111
rect 1961 1581 1995 1615
rect 3709 1717 3743 1751
rect 4169 1649 4203 1683
rect 5273 1649 5307 1683
rect 5457 1649 5491 1683
rect 5549 1785 5583 1819
rect 5549 1649 5583 1683
rect 5641 1785 5675 1819
rect 5089 1513 5123 1547
rect 5181 1513 5215 1547
rect 3433 1445 3467 1479
rect 5365 1445 5399 1479
rect 5457 1445 5491 1479
rect 5181 1377 5215 1411
rect 5089 1241 5123 1275
rect 5273 1241 5307 1275
rect 5181 1173 5215 1207
rect 5365 1173 5399 1207
rect 5273 1037 5307 1071
rect 5641 1377 5675 1411
rect 5641 833 5675 867
rect 5273 697 5307 731
rect 5365 697 5399 731
rect 5089 629 5123 663
rect 5181 561 5215 595
rect 26985 1785 27019 1819
rect 26249 1717 26283 1751
rect 10149 1649 10183 1683
rect 25145 1649 25179 1683
rect 11161 1581 11195 1615
rect 6929 1445 6963 1479
rect 10609 1445 10643 1479
rect 6929 1173 6963 1207
rect 7297 1377 7331 1411
rect 10517 1377 10551 1411
rect 10425 1241 10459 1275
rect 10425 1105 10459 1139
rect 11069 1241 11103 1275
rect 11161 1241 11195 1275
rect 11253 1581 11287 1615
rect 12909 1445 12943 1479
rect 13185 1309 13219 1343
rect 25145 1173 25179 1207
rect 25789 1649 25823 1683
rect 10517 1105 10551 1139
rect 25973 1377 26007 1411
rect 35265 1785 35299 1819
rect 34989 1717 35023 1751
rect 26985 1649 27019 1683
rect 27077 1649 27111 1683
rect 26249 1309 26283 1343
rect 26801 1377 26835 1411
rect 27077 1377 27111 1411
rect 28273 1513 28307 1547
rect 25789 833 25823 867
rect 25881 969 25915 1003
rect 25973 969 26007 1003
rect 25881 833 25915 867
rect 19349 765 19383 799
rect 19441 765 19475 799
rect 7297 629 7331 663
rect 13185 697 13219 731
rect 4721 425 4755 459
rect 5089 493 5123 527
rect 6009 493 6043 527
rect 6101 493 6135 527
rect 9689 561 9723 595
rect 5457 425 5491 459
rect 5365 357 5399 391
rect 5733 357 5767 391
rect 5825 357 5859 391
rect 1777 17 1811 51
rect 5273 289 5307 323
rect 5641 221 5675 255
rect 10425 561 10459 595
rect 10241 425 10275 459
rect 10425 357 10459 391
rect 9689 289 9723 323
rect 9781 289 9815 323
rect 6009 221 6043 255
rect 5365 153 5399 187
rect 5549 153 5583 187
rect 5457 85 5491 119
rect 5641 85 5675 119
rect 6009 85 6043 119
rect 9781 85 9815 119
rect 10517 221 10551 255
rect 10517 85 10551 119
rect 10609 85 10643 119
rect 14289 561 14323 595
rect 14289 357 14323 391
rect 14473 357 14507 391
rect 13185 17 13219 51
rect 28273 1241 28307 1275
rect 34345 1309 34379 1343
rect 34345 1105 34379 1139
rect 26801 289 26835 323
rect 28181 833 28215 867
rect 35081 1649 35115 1683
rect 39589 1785 39623 1819
rect 35265 1513 35299 1547
rect 35357 1717 35391 1751
rect 35081 1377 35115 1411
rect 35357 969 35391 1003
rect 38025 1649 38059 1683
rect 35265 289 35299 323
rect 28181 153 28215 187
rect 39129 1649 39163 1683
rect 39037 1377 39071 1411
rect 38393 1105 38427 1139
rect 38301 969 38335 1003
rect 38301 833 38335 867
rect 38393 833 38427 867
rect 38025 153 38059 187
rect 38117 765 38151 799
rect 38669 357 38703 391
rect 39129 1309 39163 1343
rect 39405 1377 39439 1411
rect 39221 1173 39255 1207
rect 39497 1241 39531 1275
rect 39497 765 39531 799
rect 39313 629 39347 663
rect 39589 629 39623 663
rect 39681 1785 39715 1819
rect 39037 289 39071 323
rect 39221 357 39255 391
rect 39313 357 39347 391
rect 38669 221 38703 255
rect 38117 153 38151 187
rect 48973 1785 49007 1819
rect 56793 1785 56827 1819
rect 48697 1717 48731 1751
rect 49065 1717 49099 1751
rect 50813 1717 50847 1751
rect 50997 1717 51031 1751
rect 42441 1581 42475 1615
rect 42441 833 42475 867
rect 42901 1581 42935 1615
rect 65441 1785 65475 1819
rect 48973 1581 49007 1615
rect 49065 1581 49099 1615
rect 48789 1513 48823 1547
rect 48881 1513 48915 1547
rect 49065 1445 49099 1479
rect 48881 1377 48915 1411
rect 48881 1241 48915 1275
rect 55781 1649 55815 1683
rect 49157 1377 49191 1411
rect 53297 1377 53331 1411
rect 49065 1173 49099 1207
rect 49157 1173 49191 1207
rect 42901 765 42935 799
rect 49157 765 49191 799
rect 49709 765 49743 799
rect 49709 629 49743 663
rect 49801 629 49835 663
rect 49249 561 49283 595
rect 39681 153 39715 187
rect 39773 289 39807 323
rect 39773 153 39807 187
rect 39865 289 39899 323
rect 49249 289 49283 323
rect 56609 1649 56643 1683
rect 56793 1649 56827 1683
rect 63233 1649 63267 1683
rect 56701 1513 56735 1547
rect 58265 1513 58299 1547
rect 58081 1309 58115 1343
rect 58173 1445 58207 1479
rect 56885 901 56919 935
rect 57989 901 58023 935
rect 53297 221 53331 255
rect 55321 765 55355 799
rect 49801 153 49835 187
rect 60933 1445 60967 1479
rect 62129 1445 62163 1479
rect 59093 1309 59127 1343
rect 59093 289 59127 323
rect 58173 221 58207 255
rect 58265 221 58299 255
rect 61301 1309 61335 1343
rect 62129 1309 62163 1343
rect 63325 1649 63359 1683
rect 65533 1785 65567 1819
rect 71881 1649 71915 1683
rect 67005 1513 67039 1547
rect 65533 1445 65567 1479
rect 65625 1445 65659 1479
rect 66729 1445 66763 1479
rect 66821 1445 66855 1479
rect 63325 1309 63359 1343
rect 63417 1309 63451 1343
rect 67005 1309 67039 1343
rect 71789 1377 71823 1411
rect 67097 1309 67131 1343
rect 61301 901 61335 935
rect 63325 1173 63359 1207
rect 63509 1173 63543 1207
rect 66821 1173 66855 1207
rect 63325 901 63359 935
rect 68937 1037 68971 1071
rect 64981 901 65015 935
rect 63509 833 63543 867
rect 60749 153 60783 187
rect 60841 289 60875 323
rect 60841 153 60875 187
rect 63509 221 63543 255
rect 63601 221 63635 255
rect 63693 833 63727 867
rect 68845 901 68879 935
rect 69397 901 69431 935
rect 69489 901 69523 935
rect 70593 901 70627 935
rect 67281 221 67315 255
rect 69397 153 69431 187
rect 55321 85 55355 119
rect 72801 1309 72835 1343
rect 72893 1309 72927 1343
rect 72985 1173 73019 1207
rect 73169 1173 73203 1207
rect 72985 1037 73019 1071
rect 73077 1037 73111 1071
rect 72985 901 73019 935
rect 72801 833 72835 867
rect 73169 629 73203 663
rect 73261 629 73295 663
rect 72985 289 73019 323
rect 73077 289 73111 323
rect 73353 493 73387 527
rect 74825 1377 74859 1411
rect 75009 1309 75043 1343
rect 76205 1173 76239 1207
rect 76297 1445 76331 1479
rect 76389 1445 76423 1479
rect 82829 1513 82863 1547
rect 83473 1513 83507 1547
rect 78689 1445 78723 1479
rect 82645 1445 82679 1479
rect 82737 1445 82771 1479
rect 83197 1445 83231 1479
rect 83381 1445 83415 1479
rect 78781 1377 78815 1411
rect 81449 1377 81483 1411
rect 76297 1173 76331 1207
rect 76757 1309 76791 1343
rect 75469 901 75503 935
rect 75561 901 75595 935
rect 75929 833 75963 867
rect 76021 833 76055 867
rect 76573 901 76607 935
rect 81725 1377 81759 1411
rect 78689 1241 78723 1275
rect 76757 833 76791 867
rect 78965 1105 78999 1139
rect 76573 765 76607 799
rect 76665 765 76699 799
rect 78965 765 78999 799
rect 75561 629 75595 663
rect 75837 629 75871 663
rect 75929 629 75963 663
rect 73905 357 73939 391
rect 74365 357 74399 391
rect 76573 357 76607 391
rect 72525 153 72559 187
rect 72617 153 72651 187
rect 73445 221 73479 255
rect 73537 221 73571 255
rect 73721 221 73755 255
rect 76481 153 76515 187
rect 76573 153 76607 187
rect 76665 357 76699 391
rect 14473 17 14507 51
rect 83105 1309 83139 1343
rect 83197 1309 83231 1343
rect 83381 1309 83415 1343
rect 83565 1309 83599 1343
rect 82829 1173 82863 1207
rect 83013 1173 83047 1207
rect 82737 1105 82771 1139
rect 83289 1105 83323 1139
rect 82829 969 82863 1003
rect 82921 901 82955 935
rect 83013 765 83047 799
rect 83105 901 83139 935
rect 83473 969 83507 1003
rect 83565 969 83599 1003
rect 83381 833 83415 867
rect 82277 629 82311 663
rect 82737 629 82771 663
rect 83381 153 83415 187
rect 84117 1377 84151 1411
rect 84117 833 84151 867
rect 84209 1377 84243 1411
rect 85957 1377 85991 1411
rect 86049 1377 86083 1411
rect 84853 1173 84887 1207
rect 84853 833 84887 867
rect 84393 153 84427 187
rect 84577 153 84611 187
rect 85773 1173 85807 1207
rect 87429 1377 87463 1411
rect 87521 1513 87555 1547
rect 87521 1377 87555 1411
rect 87061 1309 87095 1343
rect 87613 1309 87647 1343
rect 87705 1445 87739 1479
rect 85865 833 85899 867
rect 86417 833 86451 867
rect 92765 1445 92799 1479
rect 91845 1377 91879 1411
rect 92581 1377 92615 1411
rect 93041 1377 93075 1411
rect 92397 1309 92431 1343
rect 93133 1309 93167 1343
rect 87889 1173 87923 1207
rect 87797 833 87831 867
rect 89637 357 89671 391
rect 87797 153 87831 187
rect 91661 1173 91695 1207
rect 91753 1173 91787 1207
rect 91845 1241 91879 1275
rect 92121 1173 92155 1207
rect 92305 1105 92339 1139
rect 92673 1105 92707 1139
rect 91845 1037 91879 1071
rect 91937 1037 91971 1071
rect 92581 765 92615 799
rect 92949 765 92983 799
rect 91569 697 91603 731
rect 91661 697 91695 731
rect 92121 629 92155 663
rect 92489 629 92523 663
rect 106013 1785 106047 1819
rect 106105 1785 106139 1819
rect 93317 1173 93351 1207
rect 101413 1513 101447 1547
rect 101505 1445 101539 1479
rect 101597 1445 101631 1479
rect 102425 1513 102459 1547
rect 102333 1445 102367 1479
rect 102057 1377 102091 1411
rect 93225 1105 93259 1139
rect 101873 1309 101907 1343
rect 102241 1309 102275 1343
rect 103437 1513 103471 1547
rect 93133 765 93167 799
rect 100401 1241 100435 1275
rect 100677 1241 100711 1275
rect 100769 1241 100803 1275
rect 102057 1241 102091 1275
rect 102425 1241 102459 1275
rect 97365 901 97399 935
rect 93409 833 93443 867
rect 93961 833 93995 867
rect 96353 833 96387 867
rect 96445 833 96479 867
rect 96997 833 97031 867
rect 93409 561 93443 595
rect 94145 561 94179 595
rect 97365 697 97399 731
rect 93225 493 93259 527
rect 94329 493 94363 527
rect 97365 493 97399 527
rect 97457 697 97491 731
rect 92673 357 92707 391
rect 92857 357 92891 391
rect 94329 357 94363 391
rect 95709 425 95743 459
rect 96721 425 96755 459
rect 95801 357 95835 391
rect 97181 425 97215 459
rect 100861 1037 100895 1071
rect 100953 1037 100987 1071
rect 102701 1241 102735 1275
rect 103253 1241 103287 1275
rect 100585 765 100619 799
rect 100861 765 100895 799
rect 101045 901 101079 935
rect 101321 901 101355 935
rect 101873 901 101907 935
rect 102885 901 102919 935
rect 101137 833 101171 867
rect 101229 833 101263 867
rect 102241 765 102275 799
rect 98193 561 98227 595
rect 98285 561 98319 595
rect 91477 153 91511 187
rect 91569 153 91603 187
rect 92121 85 92155 119
rect 92489 85 92523 119
rect 100125 697 100159 731
rect 100493 697 100527 731
rect 100677 697 100711 731
rect 102333 697 102367 731
rect 100309 493 100343 527
rect 100677 493 100711 527
rect 102333 561 102367 595
rect 102425 561 102459 595
rect 103529 1105 103563 1139
rect 103805 1513 103839 1547
rect 104357 1513 104391 1547
rect 104541 1513 104575 1547
rect 104541 1173 104575 1207
rect 105921 1377 105955 1411
rect 106013 1377 106047 1411
rect 106289 1173 106323 1207
rect 103713 1105 103747 1139
rect 104081 1105 104115 1139
rect 104909 1105 104943 1139
rect 105921 1105 105955 1139
rect 103529 833 103563 867
rect 106841 1785 106875 1819
rect 107025 1717 107059 1751
rect 106841 1445 106875 1479
rect 109969 1377 110003 1411
rect 106381 833 106415 867
rect 106565 833 106599 867
rect 107301 833 107335 867
rect 109325 833 109359 867
rect 111625 1717 111659 1751
rect 109049 765 109083 799
rect 102609 697 102643 731
rect 110705 1445 110739 1479
rect 103161 561 103195 595
rect 107025 289 107059 323
rect 106841 221 106875 255
rect 110797 1445 110831 1479
rect 110797 833 110831 867
rect 110889 833 110923 867
rect 110889 561 110923 595
rect 111073 1445 111107 1479
rect 111257 1581 111291 1615
rect 111165 1377 111199 1411
rect 111441 1581 111475 1615
rect 111257 1241 111291 1275
rect 111349 1377 111383 1411
rect 111073 765 111107 799
rect 111165 765 111199 799
rect 111809 1581 111843 1615
rect 112361 1581 112395 1615
rect 111533 1377 111567 1411
rect 111809 1241 111843 1275
rect 111993 1173 112027 1207
rect 112085 1173 112119 1207
rect 111809 1037 111843 1071
rect 112085 1037 112119 1071
rect 111809 833 111843 867
rect 112545 833 112579 867
rect 115121 1581 115155 1615
rect 114845 1445 114879 1479
rect 114937 1445 114971 1479
rect 114937 1241 114971 1275
rect 115029 1241 115063 1275
rect 114753 833 114787 867
rect 114845 833 114879 867
rect 115305 1377 115339 1411
rect 115857 1105 115891 1139
rect 116133 1785 116167 1819
rect 116225 1785 116259 1819
rect 121561 1717 121595 1751
rect 116225 1377 116259 1411
rect 116317 1377 116351 1411
rect 121377 1649 121411 1683
rect 116501 1581 116535 1615
rect 116593 1581 116627 1615
rect 116593 1173 116627 1207
rect 116685 1241 116719 1275
rect 116869 1173 116903 1207
rect 116409 1037 116443 1071
rect 116501 1037 116535 1071
rect 111717 765 111751 799
rect 111993 765 112027 799
rect 112913 765 112947 799
rect 116133 969 116167 1003
rect 116685 901 116719 935
rect 120457 1377 120491 1411
rect 119261 1173 119295 1207
rect 119445 1173 119479 1207
rect 119537 1173 119571 1207
rect 120917 1377 120951 1411
rect 121009 1241 121043 1275
rect 121101 1241 121135 1275
rect 117053 901 117087 935
rect 120181 969 120215 1003
rect 110981 561 111015 595
rect 111717 629 111751 663
rect 112177 629 112211 663
rect 111441 561 111475 595
rect 112453 561 112487 595
rect 111993 493 112027 527
rect 112177 493 112211 527
rect 111809 425 111843 459
rect 112269 425 112303 459
rect 111993 289 112027 323
rect 112269 221 112303 255
rect 111809 153 111843 187
rect 111901 153 111935 187
rect 112361 153 112395 187
rect 120733 765 120767 799
rect 121285 1037 121319 1071
rect 122113 1445 122147 1479
rect 121929 1377 121963 1411
rect 122297 1377 122331 1411
rect 122113 1241 122147 1275
rect 122665 1445 122699 1479
rect 124689 1649 124723 1683
rect 121377 969 121411 1003
rect 121469 969 121503 1003
rect 121837 969 121871 1003
rect 121929 969 121963 1003
rect 121377 833 121411 867
rect 121285 765 121319 799
rect 121469 765 121503 799
rect 121469 629 121503 663
rect 121561 629 121595 663
rect 123033 1037 123067 1071
rect 122389 969 122423 1003
rect 124045 969 124079 1003
rect 124321 969 124355 1003
rect 122665 901 122699 935
rect 122113 629 122147 663
rect 125333 1581 125367 1615
rect 125609 1785 125643 1819
rect 125609 1649 125643 1683
rect 125701 1785 125735 1819
rect 125701 1581 125735 1615
rect 125425 1241 125459 1275
rect 125517 1445 125551 1479
rect 125517 1241 125551 1275
rect 125609 1445 125643 1479
rect 125885 1445 125919 1479
rect 125977 1581 126011 1615
rect 126069 1581 126103 1615
rect 127357 1581 127391 1615
rect 127449 1581 127483 1615
rect 128093 1717 128127 1751
rect 128461 1785 128495 1819
rect 130485 1785 130519 1819
rect 134257 1785 134291 1819
rect 134349 1785 134383 1819
rect 134625 1785 134659 1819
rect 128277 1717 128311 1751
rect 128093 1581 128127 1615
rect 128185 1581 128219 1615
rect 128093 1445 128127 1479
rect 128369 1445 128403 1479
rect 128645 1649 128679 1683
rect 129565 1717 129599 1751
rect 130301 1717 130335 1751
rect 134441 1717 134475 1751
rect 140513 1717 140547 1751
rect 129381 1649 129415 1683
rect 134625 1649 134659 1683
rect 128645 1445 128679 1479
rect 128737 1445 128771 1479
rect 129289 1445 129323 1479
rect 129749 1445 129783 1479
rect 131773 1377 131807 1411
rect 132601 1377 132635 1411
rect 126069 1241 126103 1275
rect 128185 1309 128219 1343
rect 128737 1309 128771 1343
rect 128921 1309 128955 1343
rect 128001 1241 128035 1275
rect 128093 1241 128127 1275
rect 128829 1241 128863 1275
rect 129197 1241 129231 1275
rect 129381 1241 129415 1275
rect 131957 1309 131991 1343
rect 132785 1377 132819 1411
rect 134165 1445 134199 1479
rect 134441 1377 134475 1411
rect 141617 1717 141651 1751
rect 141709 1717 141743 1751
rect 135085 1649 135119 1683
rect 137293 1649 137327 1683
rect 138489 1649 138523 1683
rect 138581 1649 138615 1683
rect 140329 1649 140363 1683
rect 140881 1649 140915 1683
rect 136557 1581 136591 1615
rect 137017 1581 137051 1615
rect 141065 1581 141099 1615
rect 134717 1377 134751 1411
rect 136649 1513 136683 1547
rect 136833 1513 136867 1547
rect 135913 1377 135947 1411
rect 138673 1377 138707 1411
rect 134441 1241 134475 1275
rect 134717 1241 134751 1275
rect 135361 1241 135395 1275
rect 134901 1105 134935 1139
rect 125517 969 125551 1003
rect 128921 969 128955 1003
rect 131773 969 131807 1003
rect 129105 901 129139 935
rect 129289 901 129323 935
rect 124505 629 124539 663
rect 124689 629 124723 663
rect 129565 901 129599 935
rect 134625 901 134659 935
rect 134809 901 134843 935
rect 135269 901 135303 935
rect 135361 901 135395 935
rect 135545 1241 135579 1275
rect 140881 1241 140915 1275
rect 139317 1173 139351 1207
rect 139409 1173 139443 1207
rect 139593 1173 139627 1207
rect 140697 1105 140731 1139
rect 136097 901 136131 935
rect 136189 901 136223 935
rect 140053 1037 140087 1071
rect 140605 1037 140639 1071
rect 140697 969 140731 1003
rect 140881 969 140915 1003
rect 140421 901 140455 935
rect 140513 901 140547 935
rect 141157 901 141191 935
rect 141249 1377 141283 1411
rect 142445 1513 142479 1547
rect 142997 1513 143031 1547
rect 144101 1513 144135 1547
rect 144377 1513 144411 1547
rect 143089 1377 143123 1411
rect 143641 1377 143675 1411
rect 142905 1241 142939 1275
rect 142261 1105 142295 1139
rect 144009 1445 144043 1479
rect 144285 1445 144319 1479
rect 144837 1717 144871 1751
rect 144837 1581 144871 1615
rect 145113 1513 145147 1547
rect 145205 1513 145239 1547
rect 145021 1445 145055 1479
rect 146861 1785 146895 1819
rect 147137 1785 147171 1819
rect 147229 1785 147263 1819
rect 147873 1785 147907 1819
rect 147965 1785 147999 1819
rect 148057 1785 148091 1819
rect 148425 1717 148459 1751
rect 148517 1785 148551 1819
rect 149069 1785 149103 1819
rect 149161 1785 149195 1819
rect 148977 1717 149011 1751
rect 150081 1717 150115 1751
rect 148885 1581 148919 1615
rect 149069 1581 149103 1615
rect 149161 1581 149195 1615
rect 149529 1581 149563 1615
rect 145573 1445 145607 1479
rect 145665 1445 145699 1479
rect 144101 1377 144135 1411
rect 147413 1445 147447 1479
rect 147781 1377 147815 1411
rect 149345 1445 149379 1479
rect 149529 1445 149563 1479
rect 149621 1581 149655 1615
rect 148793 1377 148827 1411
rect 150265 1785 150299 1819
rect 150357 1785 150391 1819
rect 150449 1717 150483 1751
rect 150449 1581 150483 1615
rect 150449 1445 150483 1479
rect 150541 1445 150575 1479
rect 149529 1173 149563 1207
rect 149897 1173 149931 1207
rect 145573 969 145607 1003
rect 142353 901 142387 935
rect 143181 901 143215 935
rect 143273 901 143307 935
rect 145757 901 145791 935
rect 147413 1037 147447 1071
rect 147781 1037 147815 1071
rect 147965 1105 147999 1139
rect 149713 1105 149747 1139
rect 150081 1105 150115 1139
rect 148149 1037 148183 1071
rect 148977 1037 149011 1071
rect 149345 1037 149379 1071
rect 149437 1037 149471 1071
rect 146309 901 146343 935
rect 147321 901 147355 935
rect 147413 901 147447 935
rect 149437 901 149471 935
rect 150081 901 150115 935
rect 150173 901 150207 935
rect 150449 1241 150483 1275
rect 151277 1717 151311 1751
rect 151369 1717 151403 1751
rect 151461 1785 151495 1819
rect 151093 1241 151127 1275
rect 151185 1581 151219 1615
rect 151645 1785 151679 1819
rect 152013 1717 152047 1751
rect 152105 1717 152139 1751
rect 152289 1785 152323 1819
rect 151461 1513 151495 1547
rect 151553 1581 151587 1615
rect 151277 1241 151311 1275
rect 151369 1377 151403 1411
rect 151461 1377 151495 1411
rect 151461 1105 151495 1139
rect 151553 1105 151587 1139
rect 151645 1581 151679 1615
rect 152289 1581 152323 1615
rect 152381 1785 152415 1819
rect 151921 1513 151955 1547
rect 153301 1785 153335 1819
rect 153393 1785 153427 1819
rect 154221 1785 154255 1819
rect 152105 1513 152139 1547
rect 152657 1581 152691 1615
rect 152749 1581 152783 1615
rect 154497 1785 154531 1819
rect 156153 1785 156187 1819
rect 152657 1445 152691 1479
rect 153209 1513 153243 1547
rect 153301 1513 153335 1547
rect 153577 1581 153611 1615
rect 153761 1513 153795 1547
rect 151737 1241 151771 1275
rect 152565 1241 152599 1275
rect 152749 1377 152783 1411
rect 152749 1241 152783 1275
rect 152841 1377 152875 1411
rect 152013 969 152047 1003
rect 152289 969 152323 1003
rect 152841 1105 152875 1139
rect 152473 901 152507 935
rect 153025 1241 153059 1275
rect 152013 765 152047 799
rect 149713 629 149747 663
rect 135361 425 135395 459
rect 144837 425 144871 459
rect 149897 561 149931 595
rect 150081 629 150115 663
rect 152289 697 152323 731
rect 150265 629 150299 663
rect 150449 561 150483 595
rect 151369 561 151403 595
rect 151461 561 151495 595
rect 153301 1241 153335 1275
rect 153577 1241 153611 1275
rect 154589 1241 154623 1275
rect 155049 1241 155083 1275
rect 153393 1105 153427 1139
rect 153761 1105 153795 1139
rect 154037 1105 154071 1139
rect 154129 1105 154163 1139
rect 153301 833 153335 867
rect 153209 765 153243 799
rect 153393 765 153427 799
rect 153853 765 153887 799
rect 153945 765 153979 799
rect 154313 1105 154347 1139
rect 154313 765 154347 799
rect 154405 765 154439 799
rect 154681 697 154715 731
rect 153393 629 153427 663
rect 154497 629 154531 663
rect 154589 629 154623 663
rect 153301 357 153335 391
rect 153853 357 153887 391
rect 151277 221 151311 255
rect 151829 221 151863 255
rect 154589 357 154623 391
rect 155233 901 155267 935
rect 156521 1785 156555 1819
rect 156337 1717 156371 1751
rect 156337 1513 156371 1547
rect 156521 1513 156555 1547
rect 157257 1785 157291 1819
rect 157441 1717 157475 1751
rect 157809 1717 157843 1751
rect 156981 1581 157015 1615
rect 156889 1513 156923 1547
rect 157165 1513 157199 1547
rect 156521 1377 156555 1411
rect 156521 1241 156555 1275
rect 156613 1377 156647 1411
rect 156613 697 156647 731
rect 157165 901 157199 935
rect 156889 765 156923 799
rect 156797 697 156831 731
rect 157165 697 157199 731
rect 156705 629 156739 663
rect 157441 1581 157475 1615
rect 157625 1581 157659 1615
rect 158729 1581 158763 1615
rect 157349 1513 157383 1547
rect 157349 1241 157383 1275
rect 157901 1513 157935 1547
rect 158269 1241 158303 1275
rect 158729 1241 158763 1275
rect 159005 1649 159039 1683
rect 159005 1513 159039 1547
rect 159281 1581 159315 1615
rect 159189 1513 159223 1547
rect 157441 1105 157475 1139
rect 157441 833 157475 867
rect 158269 1105 158303 1139
rect 157809 765 157843 799
rect 157993 765 158027 799
rect 157625 629 157659 663
rect 159005 1241 159039 1275
rect 158361 901 158395 935
rect 159005 629 159039 663
rect 159557 1241 159591 1275
rect 160385 1649 160419 1683
rect 160477 1649 160511 1683
rect 161029 1649 161063 1683
rect 160845 1581 160879 1615
rect 161121 1581 161155 1615
rect 160385 1513 160419 1547
rect 159649 901 159683 935
rect 159281 629 159315 663
rect 156521 493 156555 527
rect 156981 493 157015 527
rect 157165 357 157199 391
rect 159741 629 159775 663
rect 160845 901 160879 935
rect 161213 901 161247 935
rect 161673 1717 161707 1751
rect 161489 1241 161523 1275
rect 161765 1241 161799 1275
rect 169677 1717 169711 1751
rect 169217 1649 169251 1683
rect 161949 1377 161983 1411
rect 164065 1445 164099 1479
rect 164157 1445 164191 1479
rect 162133 1377 162167 1411
rect 162961 1377 162995 1411
rect 164525 1445 164559 1479
rect 164617 1445 164651 1479
rect 164801 1377 164835 1411
rect 164893 1377 164927 1411
rect 160569 765 160603 799
rect 159925 697 159959 731
rect 160017 697 160051 731
rect 160661 697 160695 731
rect 161029 833 161063 867
rect 161305 833 161339 867
rect 162409 1241 162443 1275
rect 162409 901 162443 935
rect 162501 901 162535 935
rect 161121 765 161155 799
rect 161213 765 161247 799
rect 161029 629 161063 663
rect 162685 901 162719 935
rect 162225 629 162259 663
rect 162317 629 162351 663
rect 163605 1241 163639 1275
rect 170045 1785 170079 1819
rect 170229 1717 170263 1751
rect 175565 1785 175599 1819
rect 174185 1717 174219 1751
rect 175381 1717 175415 1751
rect 175749 1717 175783 1751
rect 169309 1445 169343 1479
rect 166733 1377 166767 1411
rect 169493 1377 169527 1411
rect 167009 1105 167043 1139
rect 163053 901 163087 935
rect 163145 901 163179 935
rect 164341 901 164375 935
rect 164525 833 164559 867
rect 165905 833 165939 867
rect 163053 765 163087 799
rect 166089 765 166123 799
rect 163053 629 163087 663
rect 166089 629 166123 663
rect 166273 629 166307 663
rect 167101 629 167135 663
rect 167193 629 167227 663
rect 170045 1241 170079 1275
rect 168941 1105 168975 1139
rect 169585 1105 169619 1139
rect 169677 1105 169711 1139
rect 169125 697 169159 731
rect 168941 629 168975 663
rect 171609 1445 171643 1479
rect 175749 1513 175783 1547
rect 175841 1513 175875 1547
rect 177773 1717 177807 1751
rect 173449 1445 173483 1479
rect 173541 1445 173575 1479
rect 173725 1445 173759 1479
rect 176577 1513 176611 1547
rect 175749 1309 175783 1343
rect 175933 1309 175967 1343
rect 176485 1377 176519 1411
rect 176577 1377 176611 1411
rect 176853 1377 176887 1411
rect 175841 1241 175875 1275
rect 177589 1377 177623 1411
rect 176945 1241 176979 1275
rect 177681 1241 177715 1275
rect 177865 1581 177899 1615
rect 177957 1581 177991 1615
rect 178877 1717 178911 1751
rect 178601 1649 178635 1683
rect 178785 1581 178819 1615
rect 178969 1581 179003 1615
rect 178049 1445 178083 1479
rect 177957 1377 177991 1411
rect 178969 1445 179003 1479
rect 178693 1377 178727 1411
rect 177865 1241 177899 1275
rect 169953 697 169987 731
rect 170045 697 170079 731
rect 176577 697 176611 731
rect 170229 629 170263 663
rect 170321 629 170355 663
rect 176209 629 176243 663
rect 177313 697 177347 731
rect 177037 629 177071 663
rect 177405 629 177439 663
rect 177589 629 177623 663
rect 268393 3077 268427 3111
rect 179245 1649 179279 1683
rect 179705 1717 179739 1751
rect 179153 1445 179187 1479
rect 179337 1037 179371 1071
rect 179613 1037 179647 1071
rect 179245 969 179279 1003
rect 179429 969 179463 1003
rect 179337 901 179371 935
rect 179521 901 179555 935
rect 180441 1717 180475 1751
rect 180533 1717 180567 1751
rect 179889 1513 179923 1547
rect 180441 1445 180475 1479
rect 179889 1377 179923 1411
rect 180073 1377 180107 1411
rect 180073 1173 180107 1207
rect 180165 1173 180199 1207
rect 180533 1173 180567 1207
rect 183569 1785 183603 1819
rect 184029 1581 184063 1615
rect 184121 1513 184155 1547
rect 189457 1513 189491 1547
rect 189549 1513 189583 1547
rect 180625 1173 180659 1207
rect 180717 1445 180751 1479
rect 180809 1445 180843 1479
rect 182557 1445 182591 1479
rect 180073 833 180107 867
rect 178049 629 178083 663
rect 175657 561 175691 595
rect 175933 561 175967 595
rect 176393 561 176427 595
rect 175841 493 175875 527
rect 176209 493 176243 527
rect 176485 493 176519 527
rect 175933 357 175967 391
rect 176301 357 176335 391
rect 176393 357 176427 391
rect 180257 833 180291 867
rect 183845 1173 183879 1207
rect 189733 1241 189767 1275
rect 189825 1377 189859 1411
rect 190009 1377 190043 1411
rect 190285 1717 190319 1751
rect 191205 1717 191239 1751
rect 191297 1717 191331 1751
rect 190837 1581 190871 1615
rect 190377 1445 190411 1479
rect 190653 1445 190687 1479
rect 191113 1445 191147 1479
rect 190469 1377 190503 1411
rect 190561 1377 190595 1411
rect 190653 1309 190687 1343
rect 190745 1241 190779 1275
rect 191021 1309 191055 1343
rect 191113 1309 191147 1343
rect 191021 1173 191055 1207
rect 191389 1445 191423 1479
rect 191389 1309 191423 1343
rect 191297 1241 191331 1275
rect 183661 765 183695 799
rect 183937 697 183971 731
rect 183477 629 183511 663
rect 183753 629 183787 663
rect 183845 561 183879 595
rect 183661 493 183695 527
rect 183477 425 183511 459
rect 183569 357 183603 391
rect 183661 357 183695 391
rect 190193 765 190227 799
rect 190285 765 190319 799
rect 191665 1717 191699 1751
rect 196633 1649 196667 1683
rect 196909 1717 196943 1751
rect 196817 1649 196851 1683
rect 197001 1649 197035 1683
rect 197185 1717 197219 1751
rect 191573 1445 191607 1479
rect 191665 1445 191699 1479
rect 191941 1445 191975 1479
rect 196633 1445 196667 1479
rect 195345 1309 195379 1343
rect 196633 1309 196667 1343
rect 197369 1717 197403 1751
rect 220277 1785 220311 1819
rect 220737 1785 220771 1819
rect 197921 1513 197955 1547
rect 196909 1445 196943 1479
rect 198749 1513 198783 1547
rect 199209 1513 199243 1547
rect 196817 1309 196851 1343
rect 197185 1309 197219 1343
rect 198565 1309 198599 1343
rect 197001 629 197035 663
rect 197093 629 197127 663
rect 193413 425 193447 459
rect 183753 289 183787 323
rect 183845 289 183879 323
rect 183569 221 183603 255
rect 184213 221 184247 255
rect 193321 357 193355 391
rect 183753 153 183787 187
rect 184305 153 184339 187
rect 198473 425 198507 459
rect 199025 629 199059 663
rect 199117 1309 199151 1343
rect 199209 1309 199243 1343
rect 200405 1309 200439 1343
rect 214113 1581 214147 1615
rect 214389 1581 214423 1615
rect 200865 1445 200899 1479
rect 202889 1513 202923 1547
rect 211077 1513 211111 1547
rect 211169 1513 211203 1547
rect 211445 1445 211479 1479
rect 202889 1309 202923 1343
rect 211261 1309 211295 1343
rect 214205 1309 214239 1343
rect 214297 1309 214331 1343
rect 208041 765 208075 799
rect 199117 629 199151 663
rect 204269 697 204303 731
rect 204545 697 204579 731
rect 198933 425 198967 459
rect 196541 357 196575 391
rect 196909 357 196943 391
rect 198289 357 198323 391
rect 198657 357 198691 391
rect 204453 629 204487 663
rect 208133 697 208167 731
rect 208777 697 208811 731
rect 212549 629 212583 663
rect 214481 1309 214515 1343
rect 214849 1581 214883 1615
rect 214849 1309 214883 1343
rect 220369 1581 220403 1615
rect 220645 1581 220679 1615
rect 220737 1581 220771 1615
rect 220921 1581 220955 1615
rect 217793 1377 217827 1411
rect 220829 1513 220863 1547
rect 218345 1377 218379 1411
rect 220185 1445 220219 1479
rect 220369 1445 220403 1479
rect 218713 1377 218747 1411
rect 218621 1309 218655 1343
rect 231593 1785 231627 1819
rect 231685 1785 231719 1819
rect 231501 1717 231535 1751
rect 224049 1649 224083 1683
rect 224601 1649 224635 1683
rect 224693 1649 224727 1683
rect 231777 1649 231811 1683
rect 222025 1581 222059 1615
rect 222117 1581 222151 1615
rect 224417 1581 224451 1615
rect 224969 1581 225003 1615
rect 224325 1513 224359 1547
rect 224509 1377 224543 1411
rect 225061 1377 225095 1411
rect 224601 1309 224635 1343
rect 225429 1309 225463 1343
rect 228189 1309 228223 1343
rect 228281 1309 228315 1343
rect 213745 765 213779 799
rect 213929 697 213963 731
rect 214297 697 214331 731
rect 212733 629 212767 663
rect 214021 629 214055 663
rect 214941 629 214975 663
rect 217701 629 217735 663
rect 217609 493 217643 527
rect 217885 1105 217919 1139
rect 223865 1105 223899 1139
rect 218345 969 218379 1003
rect 218529 969 218563 1003
rect 218069 901 218103 935
rect 218437 901 218471 935
rect 224141 1173 224175 1207
rect 224233 1173 224267 1207
rect 224417 1241 224451 1275
rect 224969 1241 225003 1275
rect 225153 1105 225187 1139
rect 225521 1105 225555 1139
rect 225613 1105 225647 1139
rect 228281 1173 228315 1207
rect 228373 1173 228407 1207
rect 231685 1105 231719 1139
rect 231777 1105 231811 1139
rect 224969 1037 225003 1071
rect 225429 1037 225463 1071
rect 223865 765 223899 799
rect 224233 765 224267 799
rect 221473 697 221507 731
rect 232145 1785 232179 1819
rect 232145 1649 232179 1683
rect 232421 1717 232455 1751
rect 232605 1785 232639 1819
rect 232605 1581 232639 1615
rect 236745 1785 236779 1819
rect 233341 1649 233375 1683
rect 231961 1445 231995 1479
rect 233249 1445 233283 1479
rect 232237 1241 232271 1275
rect 233985 1717 234019 1751
rect 233985 1581 234019 1615
rect 239137 1717 239171 1751
rect 236561 1445 236595 1479
rect 236653 1445 236687 1479
rect 236653 1173 236687 1207
rect 236745 1173 236779 1207
rect 239045 1445 239079 1479
rect 239321 1717 239355 1751
rect 240057 1717 240091 1751
rect 241621 1717 241655 1751
rect 250085 1717 250119 1751
rect 250821 1717 250855 1751
rect 241437 1445 241471 1479
rect 249809 1445 249843 1479
rect 250821 1445 250855 1479
rect 250913 1717 250947 1751
rect 251465 1717 251499 1751
rect 251557 1717 251591 1751
rect 237941 1173 237975 1207
rect 238217 1241 238251 1275
rect 231961 765 231995 799
rect 232053 765 232087 799
rect 232881 765 232915 799
rect 233433 765 233467 799
rect 238401 765 238435 799
rect 221013 629 221047 663
rect 224141 629 224175 663
rect 224325 629 224359 663
rect 225061 697 225095 731
rect 225153 697 225187 731
rect 224417 629 224451 663
rect 231777 697 231811 731
rect 225429 629 225463 663
rect 217885 493 217919 527
rect 231593 629 231627 663
rect 238677 1241 238711 1275
rect 239137 1241 239171 1275
rect 239321 1241 239355 1275
rect 238769 1173 238803 1207
rect 239597 1241 239631 1275
rect 251465 1241 251499 1275
rect 251557 1241 251591 1275
rect 239045 1037 239079 1071
rect 239229 1037 239263 1071
rect 239321 1037 239355 1071
rect 239045 833 239079 867
rect 239413 833 239447 867
rect 252569 1717 252603 1751
rect 252661 1717 252695 1751
rect 251189 1173 251223 1207
rect 247325 1105 247359 1139
rect 247601 1105 247635 1139
rect 245485 1037 245519 1071
rect 248337 1037 248371 1071
rect 241805 969 241839 1003
rect 242081 969 242115 1003
rect 241897 901 241931 935
rect 242173 901 242207 935
rect 241713 833 241747 867
rect 242081 833 242115 867
rect 238769 765 238803 799
rect 241897 765 241931 799
rect 241529 493 241563 527
rect 252569 629 252603 663
rect 258457 1785 258491 1819
rect 258549 1785 258583 1819
rect 262045 1785 262079 1819
rect 253581 1717 253615 1751
rect 257169 1717 257203 1751
rect 258181 1717 258215 1751
rect 258365 1717 258399 1751
rect 258273 1649 258307 1683
rect 261861 1717 261895 1751
rect 262321 1717 262355 1751
rect 262505 1717 262539 1751
rect 260665 1649 260699 1683
rect 261401 1649 261435 1683
rect 262873 1649 262907 1683
rect 260297 1581 260331 1615
rect 260849 1581 260883 1615
rect 262229 1581 262263 1615
rect 262413 1581 262447 1615
rect 262781 1581 262815 1615
rect 263241 1785 263275 1819
rect 260573 1445 260607 1479
rect 258365 1377 258399 1411
rect 258457 1377 258491 1411
rect 263149 1445 263183 1479
rect 261033 1377 261067 1411
rect 260757 1173 260791 1207
rect 259377 629 259411 663
rect 261309 697 261343 731
rect 268945 1785 268979 1819
rect 268761 1717 268795 1751
rect 279985 1717 280019 1751
rect 280169 1717 280203 1751
rect 270509 1581 270543 1615
rect 280353 1581 280387 1615
rect 265081 1445 265115 1479
rect 265265 1445 265299 1479
rect 265449 1445 265483 1479
rect 268853 1445 268887 1479
rect 271429 1445 271463 1479
rect 270693 1241 270727 1275
rect 272349 1241 272383 1275
rect 274005 1445 274039 1479
rect 280629 1581 280663 1615
rect 274557 1445 274591 1479
rect 279525 1445 279559 1479
rect 273821 1241 273855 1275
rect 279985 1241 280019 1275
rect 280077 1173 280111 1207
rect 273269 697 273303 731
rect 279341 697 279375 731
rect 279801 697 279835 731
rect 267105 629 267139 663
rect 267289 629 267323 663
rect 279985 629 280019 663
rect 289737 1717 289771 1751
rect 290473 1717 290507 1751
rect 290473 1581 290507 1615
rect 293877 1717 293911 1751
rect 285873 1513 285907 1547
rect 289645 1513 289679 1547
rect 281917 1445 281951 1479
rect 285597 1445 285631 1479
rect 285689 1445 285723 1479
rect 285965 1445 285999 1479
rect 289277 1445 289311 1479
rect 289553 1445 289587 1479
rect 281549 1173 281583 1207
rect 282009 1173 282043 1207
rect 282101 1173 282135 1207
rect 285137 1377 285171 1411
rect 281457 697 281491 731
rect 281733 697 281767 731
rect 281641 629 281675 663
rect 247601 493 247635 527
rect 251649 493 251683 527
rect 259653 493 259687 527
rect 260849 493 260883 527
rect 265541 493 265575 527
rect 268853 493 268887 527
rect 270417 493 270451 527
rect 270509 493 270543 527
rect 270785 493 270819 527
rect 279801 493 279835 527
rect 199301 357 199335 391
rect 199393 425 199427 459
rect 203073 425 203107 459
rect 212457 425 212491 459
rect 241621 425 241655 459
rect 251005 425 251039 459
rect 251373 425 251407 459
rect 260665 425 260699 459
rect 260941 425 260975 459
rect 265081 425 265115 459
rect 268945 425 268979 459
rect 270325 425 270359 459
rect 270601 425 270635 459
rect 279985 425 280019 459
rect 280261 425 280295 459
rect 281641 425 281675 459
rect 199485 357 199519 391
rect 251557 357 251591 391
rect 259837 357 259871 391
rect 270509 357 270543 391
rect 280077 357 280111 391
rect 285781 1377 285815 1411
rect 287345 1377 287379 1411
rect 285505 697 285539 731
rect 285781 697 285815 731
rect 286149 833 286183 867
rect 286149 629 286183 663
rect 285505 425 285539 459
rect 285781 425 285815 459
rect 290289 1173 290323 1207
rect 290657 1173 290691 1207
rect 287437 833 287471 867
rect 289737 833 289771 867
rect 289645 629 289679 663
rect 290197 629 290231 663
rect 290657 629 290691 663
rect 291025 1581 291059 1615
rect 293785 1581 293819 1615
rect 293877 1445 293911 1479
rect 290933 1241 290967 1275
rect 291117 1241 291151 1275
rect 290841 1173 290875 1207
rect 295165 1717 295199 1751
rect 295257 1717 295291 1751
rect 296913 1649 296947 1683
rect 296729 1445 296763 1479
rect 296821 1241 296855 1275
rect 293877 833 293911 867
rect 293969 1173 294003 1207
rect 294061 1173 294095 1207
rect 295257 1173 295291 1207
rect 295349 1173 295383 1207
rect 296821 969 296855 1003
rect 295257 697 295291 731
rect 298385 1649 298419 1683
rect 298477 1649 298511 1683
rect 368397 1785 368431 1819
rect 300041 1649 300075 1683
rect 304089 1649 304123 1683
rect 298845 1581 298879 1615
rect 298477 1513 298511 1547
rect 298661 1513 298695 1547
rect 296913 629 296947 663
rect 300041 1445 300075 1479
rect 297925 1241 297959 1275
rect 298109 1173 298143 1207
rect 293969 493 294003 527
rect 296729 493 296763 527
rect 297465 493 297499 527
rect 297557 493 297591 527
rect 289921 425 289955 459
rect 289829 357 289863 391
rect 285781 289 285815 323
rect 285873 289 285907 323
rect 289185 289 289219 323
rect 297005 425 297039 459
rect 297557 357 297591 391
rect 297649 357 297683 391
rect 304181 1649 304215 1683
rect 304181 1513 304215 1547
rect 304273 1513 304307 1547
rect 309149 1445 309183 1479
rect 314669 1649 314703 1683
rect 309425 1377 309459 1411
rect 309701 1377 309735 1411
rect 309241 1241 309275 1275
rect 300777 1173 300811 1207
rect 309425 1173 309459 1207
rect 306849 969 306883 1003
rect 306849 833 306883 867
rect 337945 1717 337979 1751
rect 319821 1649 319855 1683
rect 318993 1513 319027 1547
rect 319361 1513 319395 1547
rect 319453 1513 319487 1547
rect 318441 1445 318475 1479
rect 318625 1445 318659 1479
rect 318625 1241 318659 1275
rect 314669 765 314703 799
rect 314761 765 314795 799
rect 318717 969 318751 1003
rect 317521 765 317555 799
rect 317613 901 317647 935
rect 317613 765 317647 799
rect 320189 1445 320223 1479
rect 329665 1445 329699 1479
rect 319637 1377 319671 1411
rect 319637 833 319671 867
rect 319729 1377 319763 1411
rect 319453 765 319487 799
rect 319361 629 319395 663
rect 327089 1241 327123 1275
rect 326905 1173 326939 1207
rect 327457 1241 327491 1275
rect 329757 1241 329791 1275
rect 335829 1241 335863 1275
rect 318809 493 318843 527
rect 321845 493 321879 527
rect 322949 493 322983 527
rect 323409 901 323443 935
rect 323501 901 323535 935
rect 323409 493 323443 527
rect 336013 1173 336047 1207
rect 335461 561 335495 595
rect 335737 561 335771 595
rect 328009 493 328043 527
rect 335553 493 335587 527
rect 336013 493 336047 527
rect 337577 1241 337611 1275
rect 348985 1717 349019 1751
rect 345765 1649 345799 1683
rect 338865 1241 338899 1275
rect 337945 969 337979 1003
rect 338773 969 338807 1003
rect 336105 493 336139 527
rect 337485 493 337519 527
rect 337577 493 337611 527
rect 338773 493 338807 527
rect 345397 1241 345431 1275
rect 342177 1037 342211 1071
rect 345397 1037 345431 1071
rect 345765 969 345799 1003
rect 348525 1173 348559 1207
rect 348985 1173 349019 1207
rect 349445 1717 349479 1751
rect 343189 901 343223 935
rect 348249 901 348283 935
rect 347329 561 347363 595
rect 347513 561 347547 595
rect 338865 493 338899 527
rect 309241 425 309275 459
rect 318625 425 318659 459
rect 323225 425 323259 459
rect 335737 425 335771 459
rect 337945 425 337979 459
rect 300685 357 300719 391
rect 300777 357 300811 391
rect 322949 357 322983 391
rect 323409 357 323443 391
rect 352849 1717 352883 1751
rect 349445 901 349479 935
rect 352665 1037 352699 1071
rect 348249 357 348283 391
rect 348341 493 348375 527
rect 348525 493 348559 527
rect 352665 493 352699 527
rect 358093 1649 358127 1683
rect 356437 1445 356471 1479
rect 352849 493 352883 527
rect 354137 1173 354171 1207
rect 348341 357 348375 391
rect 351929 289 351963 323
rect 355977 1173 356011 1207
rect 356161 1173 356195 1207
rect 356161 901 356195 935
rect 358093 1377 358127 1411
rect 367293 1377 367327 1411
rect 357909 1241 357943 1275
rect 367293 1241 367327 1275
rect 357081 1173 357115 1207
rect 357081 1037 357115 1071
rect 374837 1785 374871 1819
rect 367017 1173 367051 1207
rect 367109 1173 367143 1207
rect 368397 1173 368431 1207
rect 368489 1377 368523 1411
rect 357909 1037 357943 1071
rect 364165 1037 364199 1071
rect 364257 1037 364291 1071
rect 364257 901 364291 935
rect 364349 901 364383 935
rect 374653 1377 374687 1411
rect 374653 1241 374687 1275
rect 374745 1377 374779 1411
rect 374745 1173 374779 1207
rect 388453 1785 388487 1819
rect 374837 1173 374871 1207
rect 376033 1717 376067 1751
rect 372721 969 372755 1003
rect 386521 1445 386555 1479
rect 386429 1241 386463 1275
rect 376033 1037 376067 1071
rect 378425 1037 378459 1071
rect 373089 969 373123 1003
rect 368489 901 368523 935
rect 356437 765 356471 799
rect 372813 833 372847 867
rect 378425 833 378459 867
rect 391581 1785 391615 1819
rect 388453 1377 388487 1411
rect 391213 1445 391247 1479
rect 390385 1309 390419 1343
rect 390753 1309 390787 1343
rect 386521 1173 386555 1207
rect 568313 1717 568347 1751
rect 528201 1649 528235 1683
rect 412189 1581 412223 1615
rect 391581 1377 391615 1411
rect 393605 1445 393639 1479
rect 391213 1173 391247 1207
rect 390661 1105 390695 1139
rect 390845 1105 390879 1139
rect 393605 1037 393639 1071
rect 404277 1241 404311 1275
rect 386521 833 386555 867
rect 404277 833 404311 867
rect 372445 765 372479 799
rect 386337 765 386371 799
rect 356529 493 356563 527
rect 356621 493 356655 527
rect 356621 357 356655 391
rect 386429 765 386463 799
rect 395997 765 396031 799
rect 432245 1513 432279 1547
rect 500969 1513 501003 1547
rect 432245 1241 432279 1275
rect 459569 1445 459603 1479
rect 459569 1241 459603 1275
rect 473185 1445 473219 1479
rect 473185 1241 473219 1275
rect 473369 1241 473403 1275
rect 500969 1241 501003 1275
rect 509525 1513 509559 1547
rect 509525 1241 509559 1275
rect 473369 1037 473403 1071
rect 493885 1105 493919 1139
rect 521669 1105 521703 1139
rect 521761 1105 521795 1139
rect 494069 1037 494103 1071
rect 516793 1037 516827 1071
rect 516793 901 516827 935
rect 556169 1581 556203 1615
rect 555433 1445 555467 1479
rect 555433 1241 555467 1275
rect 560217 1445 560251 1479
rect 560217 1309 560251 1343
rect 556169 1241 556203 1275
rect 528201 901 528235 935
rect 538229 1105 538263 1139
rect 412189 697 412223 731
rect 425069 833 425103 867
rect 386429 493 386463 527
rect 386521 493 386555 527
rect 395997 493 396031 527
rect 430865 833 430899 867
rect 425069 493 425103 527
rect 430773 765 430807 799
rect 372629 425 372663 459
rect 356713 357 356747 391
rect 367109 357 367143 391
rect 355977 289 356011 323
rect 368581 289 368615 323
rect 372813 357 372847 391
rect 373181 357 373215 391
rect 372353 289 372387 323
rect 372537 221 372571 255
rect 372997 221 373031 255
rect 335369 153 335403 187
rect 335645 153 335679 187
rect 347513 153 347547 187
rect 347697 153 347731 187
rect 372353 153 372387 187
rect 373273 153 373307 187
rect 376769 153 376803 187
rect 376953 153 376987 187
rect 481097 833 481131 867
rect 430865 493 430899 527
rect 436109 765 436143 799
rect 183569 85 183603 119
rect 184029 85 184063 119
rect 335553 85 335587 119
rect 335737 85 335771 119
rect 347421 85 347455 119
rect 347605 85 347639 119
rect 372445 85 372479 119
rect 372721 85 372755 119
rect 430773 85 430807 119
rect 463709 765 463743 799
rect 463709 493 463743 527
rect 473185 765 473219 799
rect 473369 765 473403 799
rect 473369 629 473403 663
rect 473461 561 473495 595
rect 473553 561 473587 595
rect 473185 493 473219 527
rect 473369 493 473403 527
rect 473645 493 473679 527
rect 481097 493 481131 527
rect 508881 833 508915 867
rect 538229 833 538263 867
rect 543105 1105 543139 1139
rect 549269 1105 549303 1139
rect 549361 1105 549395 1139
rect 559481 1105 559515 1139
rect 559481 901 559515 935
rect 543105 833 543139 867
rect 508881 493 508915 527
rect 514769 765 514803 799
rect 514769 493 514803 527
rect 459569 425 459603 459
rect 459753 425 459787 459
rect 473461 425 473495 459
rect 473553 425 473587 459
rect 473369 357 473403 391
rect 473645 357 473679 391
rect 507777 357 507811 391
rect 507869 357 507903 391
rect 473461 289 473495 323
rect 473737 289 473771 323
rect 473461 153 473495 187
rect 473645 153 473679 187
rect 436109 85 436143 119
rect 335461 17 335495 51
rect 335645 17 335679 51
rect 347329 17 347363 51
rect 347697 17 347731 51
rect 568313 17 568347 51
<< metal1 >>
rect 129642 700680 129648 700732
rect 129700 700720 129706 700732
rect 170306 700720 170312 700732
rect 129700 700692 170312 700720
rect 129700 700680 129706 700692
rect 170306 700680 170312 700692
rect 170364 700680 170370 700732
rect 105446 700612 105452 700664
rect 105504 700652 105510 700664
rect 106182 700652 106188 700664
rect 105504 700624 106188 700652
rect 105504 700612 105510 700624
rect 106182 700612 106188 700624
rect 106240 700612 106246 700664
rect 110322 700612 110328 700664
rect 110380 700652 110386 700664
rect 235166 700652 235172 700664
rect 110380 700624 235172 700652
rect 110380 700612 110386 700624
rect 235166 700612 235172 700624
rect 235224 700612 235230 700664
rect 89622 700544 89628 700596
rect 89680 700584 89686 700596
rect 300118 700584 300124 700596
rect 89680 700556 300124 700584
rect 89680 700544 89686 700556
rect 300118 700544 300124 700556
rect 300176 700544 300182 700596
rect 40494 700476 40500 700528
rect 40552 700516 40558 700528
rect 41322 700516 41328 700528
rect 40552 700488 41328 700516
rect 40552 700476 40558 700488
rect 41322 700476 41328 700488
rect 41380 700476 41386 700528
rect 70302 700476 70308 700528
rect 70360 700516 70366 700528
rect 364978 700516 364984 700528
rect 70360 700488 364984 700516
rect 70360 700476 70366 700488
rect 364978 700476 364984 700488
rect 365036 700476 365042 700528
rect 50982 700408 50988 700460
rect 51040 700448 51046 700460
rect 429838 700448 429844 700460
rect 51040 700420 429844 700448
rect 51040 700408 51046 700420
rect 429838 700408 429844 700420
rect 429896 700408 429902 700460
rect 31662 700340 31668 700392
rect 31720 700380 31726 700392
rect 494790 700380 494796 700392
rect 31720 700352 494796 700380
rect 31720 700340 31726 700352
rect 494790 700340 494796 700352
rect 494848 700340 494854 700392
rect 10962 700272 10968 700324
rect 11020 700312 11026 700324
rect 559650 700312 559656 700324
rect 11020 700284 559656 700312
rect 11020 700272 11026 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 30374 684428 30380 684480
rect 30432 684468 30438 684480
rect 31662 684468 31668 684480
rect 30432 684440 31668 684468
rect 30432 684428 30438 684440
rect 31662 684428 31668 684440
rect 31720 684428 31726 684480
rect 50062 684428 50068 684480
rect 50120 684468 50126 684480
rect 50982 684468 50988 684480
rect 50120 684440 50988 684468
rect 50120 684428 50126 684440
rect 50982 684428 50988 684440
rect 51040 684428 51046 684480
rect 128630 684428 128636 684480
rect 128688 684468 128694 684480
rect 129642 684468 129648 684480
rect 128688 684440 129648 684468
rect 128688 684428 128694 684440
rect 129642 684428 129648 684440
rect 129700 684428 129706 684480
rect 109034 684020 109040 684072
rect 109092 684060 109098 684072
rect 110322 684060 110328 684072
rect 109092 684032 110328 684060
rect 109092 684020 109098 684032
rect 110322 684020 110328 684032
rect 110380 684020 110386 684072
rect 106182 683816 106188 683868
rect 106240 683856 106246 683868
rect 148318 683856 148324 683868
rect 106240 683828 148324 683856
rect 106240 683816 106246 683828
rect 148318 683816 148324 683828
rect 148376 683816 148382 683868
rect 41322 683748 41328 683800
rect 41380 683788 41386 683800
rect 168006 683788 168012 683800
rect 41380 683760 168012 683788
rect 41380 683748 41386 683760
rect 168006 683748 168012 683760
rect 168064 683748 168070 683800
rect 285950 683204 285956 683256
rect 286008 683244 286014 683256
rect 295242 683244 295248 683256
rect 286008 683216 295248 683244
rect 286008 683204 286014 683216
rect 295242 683204 295248 683216
rect 295300 683204 295306 683256
rect 364518 683204 364524 683256
rect 364576 683244 364582 683256
rect 375374 683244 375380 683256
rect 364576 683216 375380 683244
rect 364576 683204 364582 683216
rect 375374 683204 375380 683216
rect 375432 683204 375438 683256
rect 384206 683204 384212 683256
rect 384264 683244 384270 683256
rect 391198 683244 391204 683256
rect 384264 683216 391204 683244
rect 384264 683204 384270 683216
rect 391198 683204 391204 683216
rect 391256 683204 391262 683256
rect 403894 683204 403900 683256
rect 403952 683244 403958 683256
rect 408402 683244 408408 683256
rect 403952 683216 408408 683244
rect 403952 683204 403958 683216
rect 408402 683204 408408 683216
rect 408460 683204 408466 683256
rect 462866 683204 462872 683256
rect 462924 683244 462930 683256
rect 471974 683244 471980 683256
rect 462924 683216 471980 683244
rect 462924 683204 462930 683216
rect 471974 683204 471980 683216
rect 472032 683204 472038 683256
rect 482462 683204 482468 683256
rect 482520 683244 482526 683256
rect 494054 683244 494060 683256
rect 482520 683216 494060 683244
rect 482520 683204 482526 683216
rect 494054 683204 494060 683216
rect 494112 683204 494118 683256
rect 187602 683136 187608 683188
rect 187660 683176 187666 683188
rect 569862 683176 569868 683188
rect 187660 683148 569868 683176
rect 187660 683136 187666 683148
rect 569862 683136 569868 683148
rect 569920 683136 569926 683188
rect 305914 680960 305920 681012
rect 305972 681000 305978 681012
rect 327626 681000 327632 681012
rect 305972 680972 327632 681000
rect 305972 680960 305978 680972
rect 327626 680960 327632 680972
rect 327684 680960 327690 681012
rect 379422 680552 379428 680604
rect 379480 680592 379486 680604
rect 381630 680592 381636 680604
rect 379480 680564 381636 680592
rect 379480 680552 379486 680564
rect 381630 680552 381636 680564
rect 381688 680552 381694 680604
rect 557442 680552 557448 680604
rect 557500 680592 557506 680604
rect 563238 680592 563244 680604
rect 557500 680564 563244 680592
rect 557500 680552 557506 680564
rect 563238 680552 563244 680564
rect 563296 680552 563302 680604
rect 408328 680428 408540 680456
rect 216585 680391 216643 680397
rect 216585 680357 216597 680391
rect 216631 680388 216643 680391
rect 226702 680388 226708 680400
rect 216631 680360 226708 680388
rect 216631 680357 216643 680360
rect 216585 680351 216643 680357
rect 226702 680348 226708 680360
rect 226760 680348 226766 680400
rect 231949 680391 232007 680397
rect 231949 680357 231961 680391
rect 231995 680388 232007 680391
rect 246206 680388 246212 680400
rect 231995 680360 246212 680388
rect 231995 680357 232007 680360
rect 231949 680351 232007 680357
rect 246206 680348 246212 680360
rect 246264 680348 246270 680400
rect 265894 680388 265900 680400
rect 253952 680360 265900 680388
rect 207014 680320 207020 680332
rect 206975 680292 207020 680320
rect 207014 680280 207020 680292
rect 207072 680280 207078 680332
rect 1946 679804 1952 679856
rect 2004 679844 2010 679856
rect 11701 679847 11759 679853
rect 11701 679844 11713 679847
rect 2004 679816 11713 679844
rect 2004 679804 2010 679816
rect 11701 679813 11713 679816
rect 11747 679813 11759 679847
rect 11701 679807 11759 679813
rect 16577 679847 16635 679853
rect 16577 679813 16589 679847
rect 16623 679844 16635 679847
rect 31021 679847 31079 679853
rect 31021 679844 31033 679847
rect 16623 679816 31033 679844
rect 16623 679813 16635 679816
rect 16577 679807 16635 679813
rect 31021 679813 31033 679816
rect 31067 679813 31079 679847
rect 31021 679807 31079 679813
rect 35897 679847 35955 679853
rect 35897 679813 35909 679847
rect 35943 679844 35955 679847
rect 50341 679847 50399 679853
rect 50341 679844 50353 679847
rect 35943 679816 50353 679844
rect 35943 679813 35955 679816
rect 35897 679807 35955 679813
rect 50341 679813 50353 679816
rect 50387 679813 50399 679847
rect 50341 679807 50399 679813
rect 55217 679847 55275 679853
rect 55217 679813 55229 679847
rect 55263 679844 55275 679847
rect 69661 679847 69719 679853
rect 69661 679844 69673 679847
rect 55263 679816 69673 679844
rect 55263 679813 55275 679816
rect 55217 679807 55275 679813
rect 69661 679813 69673 679816
rect 69707 679813 69719 679847
rect 69661 679807 69719 679813
rect 74537 679847 74595 679853
rect 74537 679813 74549 679847
rect 74583 679844 74595 679847
rect 88981 679847 89039 679853
rect 88981 679844 88993 679847
rect 74583 679816 88993 679844
rect 74583 679813 74595 679816
rect 74537 679807 74595 679813
rect 88981 679813 88993 679816
rect 89027 679813 89039 679847
rect 88981 679807 89039 679813
rect 93857 679847 93915 679853
rect 93857 679813 93869 679847
rect 93903 679844 93915 679847
rect 108301 679847 108359 679853
rect 108301 679844 108313 679847
rect 93903 679816 108313 679844
rect 93903 679813 93915 679816
rect 93857 679807 93915 679813
rect 108301 679813 108313 679816
rect 108347 679813 108359 679847
rect 108301 679807 108359 679813
rect 113177 679847 113235 679853
rect 113177 679813 113189 679847
rect 113223 679844 113235 679847
rect 127621 679847 127679 679853
rect 127621 679844 127633 679847
rect 113223 679816 127633 679844
rect 113223 679813 113235 679816
rect 113177 679807 113235 679813
rect 127621 679813 127633 679816
rect 127667 679813 127679 679847
rect 127621 679807 127679 679813
rect 132497 679847 132555 679853
rect 132497 679813 132509 679847
rect 132543 679844 132555 679847
rect 146941 679847 146999 679853
rect 146941 679844 146953 679847
rect 132543 679816 146953 679844
rect 132543 679813 132555 679816
rect 132497 679807 132555 679813
rect 146941 679813 146953 679816
rect 146987 679813 146999 679847
rect 146941 679807 146999 679813
rect 151817 679847 151875 679853
rect 151817 679813 151829 679847
rect 151863 679844 151875 679847
rect 166261 679847 166319 679853
rect 166261 679844 166273 679847
rect 151863 679816 166273 679844
rect 151863 679813 151875 679816
rect 151817 679807 151875 679813
rect 166261 679813 166273 679816
rect 166307 679813 166319 679847
rect 166261 679807 166319 679813
rect 171137 679847 171195 679853
rect 171137 679813 171149 679847
rect 171183 679844 171195 679847
rect 185581 679847 185639 679853
rect 185581 679844 185593 679847
rect 171183 679816 185593 679844
rect 171183 679813 171195 679816
rect 171137 679807 171195 679813
rect 185581 679813 185593 679816
rect 185627 679813 185639 679847
rect 185581 679807 185639 679813
rect 190457 679847 190515 679853
rect 190457 679813 190469 679847
rect 190503 679844 190515 679847
rect 204901 679847 204959 679853
rect 204901 679844 204913 679847
rect 190503 679816 204913 679844
rect 190503 679813 190515 679816
rect 190457 679807 190515 679813
rect 204901 679813 204913 679816
rect 204947 679813 204959 679847
rect 204901 679807 204959 679813
rect 209777 679847 209835 679853
rect 209777 679813 209789 679847
rect 209823 679844 209835 679847
rect 222013 679847 222071 679853
rect 222013 679844 222025 679847
rect 209823 679816 222025 679844
rect 209823 679813 209835 679816
rect 209777 679807 209835 679813
rect 222013 679813 222025 679816
rect 222059 679813 222071 679847
rect 222013 679807 222071 679813
rect 3418 679736 3424 679788
rect 3476 679776 3482 679788
rect 216585 679779 216643 679785
rect 216585 679776 216597 679779
rect 3476 679748 216597 679776
rect 3476 679736 3482 679748
rect 216585 679745 216597 679748
rect 216631 679745 216643 679779
rect 216585 679739 216643 679745
rect 222105 679779 222163 679785
rect 222105 679745 222117 679779
rect 222151 679745 222163 679779
rect 222105 679739 222163 679745
rect 231765 679779 231823 679785
rect 231765 679745 231777 679779
rect 231811 679776 231823 679779
rect 231949 679779 232007 679785
rect 231949 679776 231961 679779
rect 231811 679748 231961 679776
rect 231811 679745 231823 679748
rect 231765 679739 231823 679745
rect 231949 679745 231961 679748
rect 231995 679745 232007 679779
rect 231949 679739 232007 679745
rect 11701 679711 11759 679717
rect 11701 679677 11713 679711
rect 11747 679708 11759 679711
rect 16577 679711 16635 679717
rect 16577 679708 16589 679711
rect 11747 679680 16589 679708
rect 11747 679677 11759 679680
rect 11701 679671 11759 679677
rect 16577 679677 16589 679680
rect 16623 679677 16635 679711
rect 16577 679671 16635 679677
rect 31021 679711 31079 679717
rect 31021 679677 31033 679711
rect 31067 679708 31079 679711
rect 35897 679711 35955 679717
rect 35897 679708 35909 679711
rect 31067 679680 35909 679708
rect 31067 679677 31079 679680
rect 31021 679671 31079 679677
rect 35897 679677 35909 679680
rect 35943 679677 35955 679711
rect 35897 679671 35955 679677
rect 50341 679711 50399 679717
rect 50341 679677 50353 679711
rect 50387 679708 50399 679711
rect 55217 679711 55275 679717
rect 55217 679708 55229 679711
rect 50387 679680 55229 679708
rect 50387 679677 50399 679680
rect 50341 679671 50399 679677
rect 55217 679677 55229 679680
rect 55263 679677 55275 679711
rect 55217 679671 55275 679677
rect 69661 679711 69719 679717
rect 69661 679677 69673 679711
rect 69707 679708 69719 679711
rect 74537 679711 74595 679717
rect 74537 679708 74549 679711
rect 69707 679680 74549 679708
rect 69707 679677 69719 679680
rect 69661 679671 69719 679677
rect 74537 679677 74549 679680
rect 74583 679677 74595 679711
rect 74537 679671 74595 679677
rect 88981 679711 89039 679717
rect 88981 679677 88993 679711
rect 89027 679708 89039 679711
rect 93857 679711 93915 679717
rect 93857 679708 93869 679711
rect 89027 679680 93869 679708
rect 89027 679677 89039 679680
rect 88981 679671 89039 679677
rect 93857 679677 93869 679680
rect 93903 679677 93915 679711
rect 93857 679671 93915 679677
rect 108301 679711 108359 679717
rect 108301 679677 108313 679711
rect 108347 679708 108359 679711
rect 113177 679711 113235 679717
rect 113177 679708 113189 679711
rect 108347 679680 113189 679708
rect 108347 679677 108359 679680
rect 108301 679671 108359 679677
rect 113177 679677 113189 679680
rect 113223 679677 113235 679711
rect 113177 679671 113235 679677
rect 127621 679711 127679 679717
rect 127621 679677 127633 679711
rect 127667 679708 127679 679711
rect 132497 679711 132555 679717
rect 132497 679708 132509 679711
rect 127667 679680 132509 679708
rect 127667 679677 127679 679680
rect 127621 679671 127679 679677
rect 132497 679677 132509 679680
rect 132543 679677 132555 679711
rect 132497 679671 132555 679677
rect 146941 679711 146999 679717
rect 146941 679677 146953 679711
rect 146987 679708 146999 679711
rect 151817 679711 151875 679717
rect 151817 679708 151829 679711
rect 146987 679680 151829 679708
rect 146987 679677 146999 679680
rect 146941 679671 146999 679677
rect 151817 679677 151829 679680
rect 151863 679677 151875 679711
rect 151817 679671 151875 679677
rect 166261 679711 166319 679717
rect 166261 679677 166273 679711
rect 166307 679708 166319 679711
rect 171137 679711 171195 679717
rect 171137 679708 171149 679711
rect 166307 679680 171149 679708
rect 166307 679677 166319 679680
rect 166261 679671 166319 679677
rect 171137 679677 171149 679680
rect 171183 679677 171195 679711
rect 171137 679671 171195 679677
rect 185581 679711 185639 679717
rect 185581 679677 185593 679711
rect 185627 679708 185639 679711
rect 190457 679711 190515 679717
rect 190457 679708 190469 679711
rect 185627 679680 190469 679708
rect 185627 679677 185639 679680
rect 185581 679671 185639 679677
rect 190457 679677 190469 679680
rect 190503 679677 190515 679711
rect 190457 679671 190515 679677
rect 204901 679711 204959 679717
rect 204901 679677 204913 679711
rect 204947 679708 204959 679711
rect 209777 679711 209835 679717
rect 209777 679708 209789 679711
rect 204947 679680 209789 679708
rect 204947 679677 204959 679680
rect 204901 679671 204959 679677
rect 209777 679677 209789 679680
rect 209823 679677 209835 679711
rect 222120 679708 222148 679739
rect 222197 679711 222255 679717
rect 222197 679708 222209 679711
rect 222120 679680 222209 679708
rect 209777 679671 209835 679677
rect 222197 679677 222209 679680
rect 222243 679677 222255 679711
rect 222197 679671 222255 679677
rect 2498 679600 2504 679652
rect 2556 679640 2562 679652
rect 253952 679640 253980 680360
rect 265894 680348 265900 680360
rect 265952 680348 265958 680400
rect 380066 680388 380072 680400
rect 380027 680360 380072 680388
rect 380066 680348 380072 680360
rect 380124 680348 380130 680400
rect 391198 680348 391204 680400
rect 391256 680388 391262 680400
rect 394513 680391 394571 680397
rect 394513 680388 394525 680391
rect 391256 680360 394525 680388
rect 391256 680348 391262 680360
rect 394513 680357 394525 680360
rect 394559 680357 394571 680391
rect 394694 680388 394700 680400
rect 394655 680360 394700 680388
rect 394513 680351 394571 680357
rect 394694 680348 394700 680360
rect 394752 680348 394758 680400
rect 403158 680388 403164 680400
rect 403119 680360 403164 680388
rect 403158 680348 403164 680360
rect 403216 680348 403222 680400
rect 295242 680280 295248 680332
rect 295300 680320 295306 680332
rect 296714 680320 296720 680332
rect 295300 680292 296720 680320
rect 295300 680280 295306 680292
rect 296714 680280 296720 680292
rect 296772 680280 296778 680332
rect 327626 680280 327632 680332
rect 327684 680280 327690 680332
rect 364794 680320 364800 680332
rect 364755 680292 364800 680320
rect 364794 680280 364800 680292
rect 364852 680280 364858 680332
rect 370222 680320 370228 680332
rect 370183 680292 370228 680320
rect 370222 680280 370228 680292
rect 370280 680280 370286 680332
rect 375374 680280 375380 680332
rect 375432 680320 375438 680332
rect 408328 680320 408356 680428
rect 375432 680292 408356 680320
rect 375432 680280 375438 680292
rect 408402 680280 408408 680332
rect 408460 680280 408466 680332
rect 408512 680320 408540 680428
rect 463786 680416 463792 680468
rect 463844 680456 463850 680468
rect 466638 680456 466644 680468
rect 463844 680428 466644 680456
rect 463844 680416 463850 680428
rect 466638 680416 466644 680428
rect 466696 680416 466702 680468
rect 557721 680459 557779 680465
rect 557721 680425 557733 680459
rect 557767 680456 557779 680459
rect 559374 680456 559380 680468
rect 557767 680428 559380 680456
rect 557767 680425 557779 680428
rect 557721 680419 557779 680425
rect 559374 680416 559380 680428
rect 559432 680416 559438 680468
rect 412726 680388 412732 680400
rect 412687 680360 412732 680388
rect 412726 680348 412732 680360
rect 412784 680348 412790 680400
rect 418614 680388 418620 680400
rect 418575 680360 418620 680388
rect 418614 680348 418620 680360
rect 418672 680348 418678 680400
rect 423582 680348 423588 680400
rect 423640 680388 423646 680400
rect 428001 680391 428059 680397
rect 428001 680388 428013 680391
rect 423640 680360 428013 680388
rect 423640 680348 423646 680360
rect 428001 680357 428013 680360
rect 428047 680357 428059 680391
rect 428182 680388 428188 680400
rect 428143 680360 428188 680388
rect 428001 680351 428059 680357
rect 428182 680348 428188 680360
rect 428240 680348 428246 680400
rect 437750 680388 437756 680400
rect 437711 680360 437756 680388
rect 437750 680348 437756 680360
rect 437808 680348 437814 680400
rect 443546 680388 443552 680400
rect 443507 680360 443552 680388
rect 443546 680348 443552 680360
rect 443604 680348 443610 680400
rect 451366 680388 451372 680400
rect 451327 680360 451372 680388
rect 451366 680348 451372 680360
rect 451424 680348 451430 680400
rect 457162 680388 457168 680400
rect 457123 680360 457168 680388
rect 457162 680348 457168 680360
rect 457220 680348 457226 680400
rect 466546 680388 466552 680400
rect 466507 680360 466552 680388
rect 466546 680348 466552 680360
rect 466604 680348 466610 680400
rect 471974 680348 471980 680400
rect 472032 680388 472038 680400
rect 474737 680391 474795 680397
rect 474737 680388 474749 680391
rect 472032 680360 474749 680388
rect 472032 680348 472038 680360
rect 474737 680357 474749 680360
rect 474783 680357 474795 680391
rect 494054 680388 494060 680400
rect 494015 680360 494060 680388
rect 474737 680351 474795 680357
rect 494054 680348 494060 680360
rect 494112 680348 494118 680400
rect 495434 680348 495440 680400
rect 495492 680388 495498 680400
rect 502242 680388 502248 680400
rect 495492 680360 495537 680388
rect 502203 680360 502248 680388
rect 495492 680348 495498 680360
rect 502242 680348 502248 680360
rect 502300 680348 502306 680400
rect 505922 680388 505928 680400
rect 505883 680360 505928 680388
rect 505922 680348 505928 680360
rect 505980 680348 505986 680400
rect 515398 680388 515404 680400
rect 515359 680360 515404 680388
rect 515398 680348 515404 680360
rect 515456 680348 515462 680400
rect 522114 680388 522120 680400
rect 522075 680360 522120 680388
rect 522114 680348 522120 680360
rect 522172 680348 522178 680400
rect 524414 680348 524420 680400
rect 524472 680388 524478 680400
rect 534350 680388 534356 680400
rect 524472 680360 524517 680388
rect 534311 680360 534356 680388
rect 524472 680348 524478 680360
rect 534350 680348 534356 680360
rect 534408 680348 534414 680400
rect 541802 680348 541808 680400
rect 541860 680388 541866 680400
rect 543737 680391 543795 680397
rect 543737 680388 543749 680391
rect 541860 680360 543749 680388
rect 541860 680348 541866 680360
rect 543737 680357 543749 680360
rect 543783 680357 543795 680391
rect 544010 680388 544016 680400
rect 543971 680360 544016 680388
rect 543737 680351 543795 680357
rect 544010 680348 544016 680360
rect 544068 680348 544074 680400
rect 480993 680323 481051 680329
rect 480993 680320 481005 680323
rect 408512 680292 481005 680320
rect 480993 680289 481005 680292
rect 481039 680289 481051 680323
rect 481174 680320 481180 680332
rect 481135 680292 481180 680320
rect 480993 680283 481051 680289
rect 481174 680280 481180 680292
rect 481232 680280 481238 680332
rect 485774 680280 485780 680332
rect 485832 680320 485838 680332
rect 489733 680323 489791 680329
rect 485832 680292 485877 680320
rect 485832 680280 485838 680292
rect 489733 680289 489745 680323
rect 489779 680320 489791 680323
rect 553489 680323 553547 680329
rect 553489 680320 553501 680323
rect 489779 680292 553501 680320
rect 489779 680289 489791 680292
rect 489733 680283 489791 680289
rect 553489 680289 553501 680292
rect 553535 680289 553547 680323
rect 553489 680283 553547 680289
rect 554774 680280 554780 680332
rect 554832 680280 554838 680332
rect 554866 680280 554872 680332
rect 554924 680320 554930 680332
rect 554924 680292 554969 680320
rect 554924 680280 554930 680292
rect 558546 680280 558552 680332
rect 558604 680280 558610 680332
rect 559190 680320 559196 680332
rect 559151 680292 559196 680320
rect 559190 680280 559196 680292
rect 559248 680280 559254 680332
rect 560754 680320 560760 680332
rect 560715 680292 560760 680320
rect 560754 680280 560760 680292
rect 560812 680280 560818 680332
rect 561582 680320 561588 680332
rect 561543 680292 561588 680320
rect 561582 680280 561588 680292
rect 561640 680280 561646 680332
rect 561766 680320 561772 680332
rect 561727 680292 561772 680320
rect 561766 680280 561772 680292
rect 561824 680280 561830 680332
rect 561858 680280 561864 680332
rect 561916 680320 561922 680332
rect 562502 680320 562508 680332
rect 561916 680292 561961 680320
rect 562463 680292 562508 680320
rect 561916 680280 561922 680292
rect 562502 680280 562508 680292
rect 562560 680280 562566 680332
rect 566366 680280 566372 680332
rect 566424 680280 566430 680332
rect 327644 680252 327672 680280
rect 394513 680255 394571 680261
rect 327644 680224 330524 680252
rect 2556 679612 253980 679640
rect 330496 679640 330524 680224
rect 394513 680221 394525 680255
rect 394559 680252 394571 680255
rect 408420 680252 408448 680280
rect 412637 680255 412695 680261
rect 394559 680224 407804 680252
rect 408420 680224 408540 680252
rect 394559 680221 394571 680224
rect 394513 680215 394571 680221
rect 407776 680048 407804 680224
rect 408512 680184 408540 680224
rect 412637 680221 412649 680255
rect 412683 680252 412695 680255
rect 451277 680255 451335 680261
rect 451277 680252 451289 680255
rect 412683 680224 451289 680252
rect 412683 680221 412695 680224
rect 412637 680215 412695 680221
rect 451277 680221 451289 680224
rect 451323 680221 451335 680255
rect 451277 680215 451335 680221
rect 461581 680255 461639 680261
rect 461581 680221 461593 680255
rect 461627 680252 461639 680255
rect 469585 680255 469643 680261
rect 469585 680252 469597 680255
rect 461627 680224 469597 680252
rect 461627 680221 461639 680224
rect 461581 680215 461639 680221
rect 469585 680221 469597 680224
rect 469631 680221 469643 680255
rect 490469 680255 490527 680261
rect 490469 680252 490481 680255
rect 469585 680215 469643 680221
rect 478064 680224 490481 680252
rect 477957 680187 478015 680193
rect 477957 680184 477969 680187
rect 408512 680156 477969 680184
rect 477957 680153 477969 680156
rect 478003 680153 478015 680187
rect 477957 680147 478015 680153
rect 444285 680119 444343 680125
rect 444285 680085 444297 680119
rect 444331 680116 444343 680119
rect 469585 680119 469643 680125
rect 444331 680088 469536 680116
rect 444331 680085 444343 680088
rect 444285 680079 444343 680085
rect 412637 680051 412695 680057
rect 412637 680048 412649 680051
rect 407776 680020 412649 680048
rect 412637 680017 412649 680020
rect 412683 680017 412695 680051
rect 412637 680011 412695 680017
rect 428001 679983 428059 679989
rect 428001 679949 428013 679983
rect 428047 679980 428059 679983
rect 434717 679983 434775 679989
rect 434717 679980 434729 679983
rect 428047 679952 434729 679980
rect 428047 679949 428059 679952
rect 428001 679943 428059 679949
rect 434717 679949 434729 679952
rect 434763 679949 434775 679983
rect 434717 679943 434775 679949
rect 451277 679983 451335 679989
rect 451277 679949 451289 679983
rect 451323 679980 451335 679983
rect 461581 679983 461639 679989
rect 461581 679980 461593 679983
rect 451323 679952 461593 679980
rect 451323 679949 451335 679952
rect 451277 679943 451335 679949
rect 461581 679949 461593 679952
rect 461627 679949 461639 679983
rect 461581 679943 461639 679949
rect 469508 679912 469536 680088
rect 469585 680085 469597 680119
rect 469631 680116 469643 680119
rect 478064 680116 478092 680224
rect 490469 680221 490481 680224
rect 490515 680221 490527 680255
rect 490469 680215 490527 680221
rect 500221 680255 500279 680261
rect 500221 680221 500233 680255
rect 500267 680252 500279 680255
rect 509789 680255 509847 680261
rect 509789 680252 509801 680255
rect 500267 680224 509801 680252
rect 500267 680221 500279 680224
rect 500221 680215 500279 680221
rect 509789 680221 509801 680224
rect 509835 680221 509847 680255
rect 509789 680215 509847 680221
rect 533985 680255 534043 680261
rect 533985 680221 533997 680255
rect 534031 680252 534043 680255
rect 538861 680255 538919 680261
rect 538861 680252 538873 680255
rect 534031 680224 538873 680252
rect 534031 680221 534043 680224
rect 533985 680215 534043 680221
rect 538861 680221 538873 680224
rect 538907 680221 538919 680255
rect 538861 680215 538919 680221
rect 546865 680255 546923 680261
rect 546865 680221 546877 680255
rect 546911 680252 546923 680255
rect 553397 680255 553455 680261
rect 553397 680252 553409 680255
rect 546911 680224 553409 680252
rect 546911 680221 546923 680224
rect 546865 680215 546923 680221
rect 553397 680221 553409 680224
rect 553443 680221 553455 680255
rect 553397 680215 553455 680221
rect 478141 680187 478199 680193
rect 478141 680153 478153 680187
rect 478187 680184 478199 680187
rect 519541 680187 519599 680193
rect 519541 680184 519553 680187
rect 478187 680156 519553 680184
rect 478187 680153 478199 680156
rect 478141 680147 478199 680153
rect 519541 680153 519553 680156
rect 519587 680153 519599 680187
rect 519541 680147 519599 680153
rect 529109 680187 529167 680193
rect 529109 680153 529121 680187
rect 529155 680184 529167 680187
rect 554792 680184 554820 680280
rect 529155 680156 554820 680184
rect 529155 680153 529167 680156
rect 529109 680147 529167 680153
rect 469631 680088 478092 680116
rect 485685 680119 485743 680125
rect 469631 680085 469643 680088
rect 469585 680079 469643 680085
rect 485685 680085 485697 680119
rect 485731 680116 485743 680119
rect 506477 680119 506535 680125
rect 506477 680116 506489 680119
rect 485731 680088 506489 680116
rect 485731 680085 485743 680088
rect 485685 680079 485743 680085
rect 506477 680085 506489 680088
rect 506523 680085 506535 680119
rect 506477 680079 506535 680085
rect 516321 680119 516379 680125
rect 516321 680085 516333 680119
rect 516367 680116 516379 680119
rect 529017 680119 529075 680125
rect 529017 680116 529029 680119
rect 516367 680088 529029 680116
rect 516367 680085 516379 680088
rect 516321 680079 516379 680085
rect 529017 680085 529029 680088
rect 529063 680085 529075 680119
rect 529017 680079 529075 680085
rect 529201 680119 529259 680125
rect 529201 680085 529213 680119
rect 529247 680116 529259 680119
rect 557721 680119 557779 680125
rect 557721 680116 557733 680119
rect 529247 680088 557733 680116
rect 529247 680085 529259 680088
rect 529201 680079 529259 680085
rect 557721 680085 557733 680088
rect 557767 680085 557779 680119
rect 557721 680079 557779 680085
rect 474737 680051 474795 680057
rect 474737 680017 474749 680051
rect 474783 680048 474795 680051
rect 558564 680048 558592 680280
rect 474783 680020 558592 680048
rect 474783 680017 474795 680020
rect 474737 680011 474795 680017
rect 481085 679983 481143 679989
rect 481085 679949 481097 679983
rect 481131 679980 481143 679983
rect 489733 679983 489791 679989
rect 489733 679980 489745 679983
rect 481131 679952 489745 679980
rect 481131 679949 481143 679952
rect 481085 679943 481143 679949
rect 489733 679949 489745 679952
rect 489779 679949 489791 679983
rect 489733 679943 489791 679949
rect 494057 679983 494115 679989
rect 494057 679949 494069 679983
rect 494103 679980 494115 679983
rect 559193 679983 559251 679989
rect 559193 679980 559205 679983
rect 494103 679952 559205 679980
rect 494103 679949 494115 679952
rect 494057 679943 494115 679949
rect 559193 679949 559205 679952
rect 559239 679949 559251 679983
rect 559193 679943 559251 679949
rect 485593 679915 485651 679921
rect 485593 679912 485605 679915
rect 469508 679884 485605 679912
rect 485593 679881 485605 679884
rect 485639 679881 485651 679915
rect 485593 679875 485651 679881
rect 506477 679915 506535 679921
rect 506477 679881 506489 679915
rect 506523 679912 506535 679915
rect 529201 679915 529259 679921
rect 529201 679912 529213 679915
rect 506523 679884 529213 679912
rect 506523 679881 506535 679884
rect 506477 679875 506535 679881
rect 529201 679881 529213 679884
rect 529247 679881 529259 679915
rect 529201 679875 529259 679881
rect 538861 679915 538919 679921
rect 538861 679881 538873 679915
rect 538907 679912 538919 679915
rect 546865 679915 546923 679921
rect 546865 679912 546877 679915
rect 538907 679884 546877 679912
rect 538907 679881 538919 679884
rect 538861 679875 538919 679881
rect 546865 679881 546877 679884
rect 546911 679881 546923 679915
rect 561585 679915 561643 679921
rect 561585 679912 561597 679915
rect 546865 679875 546923 679881
rect 546972 679884 561597 679912
rect 434717 679847 434775 679853
rect 434717 679813 434729 679847
rect 434763 679844 434775 679847
rect 444285 679847 444343 679853
rect 444285 679844 444297 679847
rect 434763 679816 444297 679844
rect 434763 679813 434775 679816
rect 434717 679807 434775 679813
rect 444285 679813 444297 679816
rect 444331 679813 444343 679847
rect 444285 679807 444343 679813
rect 490469 679847 490527 679853
rect 490469 679813 490481 679847
rect 490515 679844 490527 679847
rect 500221 679847 500279 679853
rect 500221 679844 500233 679847
rect 490515 679816 500233 679844
rect 490515 679813 490527 679816
rect 490469 679807 490527 679813
rect 500221 679813 500233 679816
rect 500267 679813 500279 679847
rect 500221 679807 500279 679813
rect 519541 679847 519599 679853
rect 519541 679813 519553 679847
rect 519587 679844 519599 679847
rect 529109 679847 529167 679853
rect 529109 679844 529121 679847
rect 519587 679816 529121 679844
rect 519587 679813 519599 679816
rect 519541 679807 519599 679813
rect 529109 679813 529121 679816
rect 529155 679813 529167 679847
rect 529109 679807 529167 679813
rect 509789 679779 509847 679785
rect 509789 679745 509801 679779
rect 509835 679776 509847 679779
rect 516321 679779 516379 679785
rect 516321 679776 516333 679779
rect 509835 679748 516333 679776
rect 509835 679745 509847 679748
rect 509789 679739 509847 679745
rect 516321 679745 516333 679748
rect 516367 679745 516379 679779
rect 516321 679739 516379 679745
rect 529017 679779 529075 679785
rect 529017 679745 529029 679779
rect 529063 679776 529075 679779
rect 533985 679779 534043 679785
rect 533985 679776 533997 679779
rect 529063 679748 533997 679776
rect 529063 679745 529075 679748
rect 529017 679739 529075 679745
rect 533985 679745 533997 679748
rect 534031 679745 534043 679779
rect 533985 679739 534043 679745
rect 543737 679779 543795 679785
rect 543737 679745 543749 679779
rect 543783 679776 543795 679779
rect 546972 679776 547000 679884
rect 561585 679881 561597 679884
rect 561631 679881 561643 679915
rect 561585 679875 561643 679881
rect 553489 679847 553547 679853
rect 553489 679813 553501 679847
rect 553535 679844 553547 679847
rect 561769 679847 561827 679853
rect 561769 679844 561781 679847
rect 553535 679816 561781 679844
rect 553535 679813 553547 679816
rect 553489 679807 553547 679813
rect 561769 679813 561781 679816
rect 561815 679813 561827 679847
rect 561769 679807 561827 679813
rect 543783 679748 547000 679776
rect 553397 679779 553455 679785
rect 543783 679745 543795 679748
rect 543737 679739 543795 679745
rect 553397 679745 553409 679779
rect 553443 679776 553455 679779
rect 566384 679776 566412 680280
rect 553443 679748 566412 679776
rect 553443 679745 553455 679748
rect 553397 679739 553455 679745
rect 568390 679640 568396 679652
rect 330496 679612 568396 679640
rect 2556 679600 2562 679612
rect 568390 679600 568396 679612
rect 568448 679600 568454 679652
rect 222197 679575 222255 679581
rect 222197 679541 222209 679575
rect 222243 679572 222255 679575
rect 231765 679575 231823 679581
rect 231765 679572 231777 679575
rect 222243 679544 231777 679572
rect 222243 679541 222255 679544
rect 222197 679535 222255 679541
rect 231765 679541 231777 679544
rect 231811 679541 231823 679575
rect 231765 679535 231823 679541
rect 364797 679575 364855 679581
rect 364797 679541 364809 679575
rect 364843 679572 364855 679575
rect 370225 679575 370283 679581
rect 370225 679572 370237 679575
rect 364843 679544 370237 679572
rect 364843 679541 364855 679544
rect 364797 679535 364855 679541
rect 370225 679541 370237 679544
rect 370271 679541 370283 679575
rect 370225 679535 370283 679541
rect 380069 679575 380127 679581
rect 380069 679541 380081 679575
rect 380115 679572 380127 679575
rect 394697 679575 394755 679581
rect 394697 679572 394709 679575
rect 380115 679544 394709 679572
rect 380115 679541 380127 679544
rect 380069 679535 380127 679541
rect 394697 679541 394709 679544
rect 394743 679541 394755 679575
rect 394697 679535 394755 679541
rect 403161 679575 403219 679581
rect 403161 679541 403173 679575
rect 403207 679572 403219 679575
rect 412729 679575 412787 679581
rect 412729 679572 412741 679575
rect 403207 679544 412741 679572
rect 403207 679541 403219 679544
rect 403161 679535 403219 679541
rect 412729 679541 412741 679544
rect 412775 679541 412787 679575
rect 412729 679535 412787 679541
rect 418617 679575 418675 679581
rect 418617 679541 418629 679575
rect 418663 679572 418675 679575
rect 428185 679575 428243 679581
rect 428185 679572 428197 679575
rect 418663 679544 428197 679572
rect 418663 679541 418675 679544
rect 418617 679535 418675 679541
rect 428185 679541 428197 679544
rect 428231 679541 428243 679575
rect 428185 679535 428243 679541
rect 437753 679575 437811 679581
rect 437753 679541 437765 679575
rect 437799 679572 437811 679575
rect 451369 679575 451427 679581
rect 451369 679572 451381 679575
rect 437799 679544 451381 679572
rect 437799 679541 437811 679544
rect 437753 679535 437811 679541
rect 451369 679541 451381 679544
rect 451415 679541 451427 679575
rect 451369 679535 451427 679541
rect 457165 679575 457223 679581
rect 457165 679541 457177 679575
rect 457211 679572 457223 679575
rect 466549 679575 466607 679581
rect 466549 679572 466561 679575
rect 457211 679544 466561 679572
rect 457211 679541 457223 679544
rect 457165 679535 457223 679541
rect 466549 679541 466561 679544
rect 466595 679541 466607 679575
rect 466549 679535 466607 679541
rect 481177 679575 481235 679581
rect 481177 679541 481189 679575
rect 481223 679572 481235 679575
rect 485777 679575 485835 679581
rect 485777 679572 485789 679575
rect 481223 679544 485789 679572
rect 481223 679541 481235 679544
rect 481177 679535 481235 679541
rect 485777 679541 485789 679544
rect 485823 679541 485835 679575
rect 485777 679535 485835 679541
rect 495437 679575 495495 679581
rect 495437 679541 495449 679575
rect 495483 679572 495495 679575
rect 505925 679575 505983 679581
rect 505925 679572 505937 679575
rect 495483 679544 505937 679572
rect 495483 679541 495495 679544
rect 495437 679535 495495 679541
rect 505925 679541 505937 679544
rect 505971 679541 505983 679575
rect 505925 679535 505983 679541
rect 515401 679575 515459 679581
rect 515401 679541 515413 679575
rect 515447 679572 515459 679575
rect 524417 679575 524475 679581
rect 524417 679572 524429 679575
rect 515447 679544 524429 679572
rect 515447 679541 515459 679544
rect 515401 679535 515459 679541
rect 524417 679541 524429 679544
rect 524463 679541 524475 679575
rect 524417 679535 524475 679541
rect 534353 679575 534411 679581
rect 534353 679541 534365 679575
rect 534399 679572 534411 679575
rect 544013 679575 544071 679581
rect 544013 679572 544025 679575
rect 534399 679544 544025 679572
rect 534399 679541 534411 679544
rect 534353 679535 534411 679541
rect 544013 679541 544025 679544
rect 544059 679541 544071 679575
rect 544013 679535 544071 679541
rect 522117 679303 522175 679309
rect 522117 679269 522129 679303
rect 522163 679300 522175 679303
rect 561861 679303 561919 679309
rect 561861 679300 561873 679303
rect 522163 679272 561873 679300
rect 522163 679269 522175 679272
rect 522117 679263 522175 679269
rect 561861 679269 561873 679272
rect 561907 679269 561919 679303
rect 561861 679263 561919 679269
rect 502245 679235 502303 679241
rect 502245 679201 502257 679235
rect 502291 679232 502303 679235
rect 562505 679235 562563 679241
rect 562505 679232 562517 679235
rect 502291 679204 562517 679232
rect 502291 679201 502303 679204
rect 502245 679195 502303 679201
rect 562505 679201 562517 679204
rect 562551 679201 562563 679235
rect 562505 679195 562563 679201
rect 3694 679124 3700 679176
rect 3752 679164 3758 679176
rect 207017 679167 207075 679173
rect 207017 679164 207029 679167
rect 3752 679136 207029 679164
rect 3752 679124 3758 679136
rect 207017 679133 207029 679136
rect 207063 679133 207075 679167
rect 207017 679127 207075 679133
rect 443549 679167 443607 679173
rect 443549 679133 443561 679167
rect 443595 679164 443607 679167
rect 554869 679167 554927 679173
rect 554869 679164 554881 679167
rect 443595 679136 554881 679164
rect 443595 679133 443607 679136
rect 443549 679127 443607 679133
rect 554869 679133 554881 679136
rect 554915 679133 554927 679167
rect 554869 679127 554927 679133
rect 560757 679167 560815 679173
rect 560757 679133 560769 679167
rect 560803 679164 560815 679167
rect 572714 679164 572720 679176
rect 560803 679136 572720 679164
rect 560803 679133 560815 679136
rect 560757 679127 560815 679133
rect 572714 679124 572720 679136
rect 572772 679124 572778 679176
rect 2222 679056 2228 679108
rect 2280 679096 2286 679108
rect 569218 679096 569224 679108
rect 2280 679068 569224 679096
rect 2280 679056 2286 679068
rect 569218 679056 569224 679068
rect 569276 679056 569282 679108
rect 1854 678988 1860 679040
rect 1912 679028 1918 679040
rect 571426 679028 571432 679040
rect 1912 679000 571432 679028
rect 1912 678988 1918 679000
rect 571426 678988 571432 679000
rect 571484 678988 571490 679040
rect 198 677492 204 677544
rect 256 677532 262 677544
rect 1394 677532 1400 677544
rect 256 677504 1400 677532
rect 256 677492 262 677504
rect 1394 677492 1400 677504
rect 1452 677492 1458 677544
rect 571426 677492 571432 677544
rect 571484 677532 571490 677544
rect 578142 677532 578148 677544
rect 571484 677504 578148 677532
rect 571484 677492 571490 677504
rect 578142 677492 578148 677504
rect 578200 677492 578206 677544
rect 1946 676132 1952 676184
rect 2004 676132 2010 676184
rect 1964 676048 1992 676132
rect 1946 675996 1952 676048
rect 2004 675996 2010 676048
rect 578142 674772 578148 674824
rect 578200 674812 578206 674824
rect 580166 674812 580172 674824
rect 578200 674784 580172 674812
rect 578200 674772 578206 674784
rect 580166 674772 580172 674784
rect 580224 674772 580230 674824
rect 569954 659240 569960 659252
rect 569915 659212 569960 659240
rect 569954 659200 569960 659212
rect 570012 659200 570018 659252
rect 569954 654168 569960 654220
rect 570012 654208 570018 654220
rect 577498 654208 577504 654220
rect 570012 654180 577504 654208
rect 570012 654168 570018 654180
rect 577498 654168 577504 654180
rect 577556 654168 577562 654220
rect 569954 654072 569960 654084
rect 569915 654044 569960 654072
rect 569954 654032 569960 654044
rect 570012 654032 570018 654084
rect 1854 648592 1860 648644
rect 1912 648632 1918 648644
rect 1946 648632 1952 648644
rect 1912 648604 1952 648632
rect 1912 648592 1918 648604
rect 1946 648592 1952 648604
rect 2004 648592 2010 648644
rect 1946 648088 1952 648100
rect 1907 648060 1952 648088
rect 1946 648048 1952 648060
rect 2004 648048 2010 648100
rect 1857 642651 1915 642657
rect 1857 642617 1869 642651
rect 1903 642648 1915 642651
rect 1946 642648 1952 642660
rect 1903 642620 1952 642648
rect 1903 642617 1915 642620
rect 1857 642611 1915 642617
rect 1946 642608 1952 642620
rect 2004 642608 2010 642660
rect 1946 641792 1952 641844
rect 2004 641792 2010 641844
rect 1964 641640 1992 641792
rect 1946 641588 1952 641640
rect 2004 641588 2010 641640
rect 1946 639316 1952 639328
rect 1907 639288 1952 639316
rect 1946 639276 1952 639288
rect 2004 639276 2010 639328
rect 1854 633468 1860 633480
rect 1815 633440 1860 633468
rect 1854 633428 1860 633440
rect 1912 633428 1918 633480
rect 569954 630164 569960 630216
rect 570012 630204 570018 630216
rect 572714 630204 572720 630216
rect 570012 630176 572720 630204
rect 570012 630164 570018 630176
rect 572714 630164 572720 630176
rect 572772 630164 572778 630216
rect 577498 627852 577504 627904
rect 577556 627892 577562 627904
rect 579706 627892 579712 627904
rect 577556 627864 579712 627892
rect 577556 627852 577562 627864
rect 579706 627852 579712 627864
rect 579764 627852 579770 627904
rect 1578 618264 1584 618316
rect 1636 618304 1642 618316
rect 1670 618304 1676 618316
rect 1636 618276 1676 618304
rect 1636 618264 1642 618276
rect 1670 618264 1676 618276
rect 1728 618264 1734 618316
rect 1854 618264 1860 618316
rect 1912 618304 1918 618316
rect 1946 618304 1952 618316
rect 1912 618276 1952 618304
rect 1912 618264 1918 618276
rect 1946 618264 1952 618276
rect 2004 618264 2010 618316
rect 569954 609628 569960 609680
rect 570012 609668 570018 609680
rect 570322 609668 570328 609680
rect 570012 609640 570328 609668
rect 570012 609628 570018 609640
rect 570322 609628 570328 609640
rect 570380 609628 570386 609680
rect 569954 609220 569960 609272
rect 570012 609260 570018 609272
rect 570046 609260 570052 609272
rect 570012 609232 570052 609260
rect 570012 609220 570018 609232
rect 570046 609220 570052 609232
rect 570104 609220 570110 609272
rect 1946 608716 1952 608728
rect 1872 608688 1952 608716
rect 1872 608592 1900 608688
rect 1946 608676 1952 608688
rect 2004 608676 2010 608728
rect 1854 608540 1860 608592
rect 1912 608540 1918 608592
rect 1857 602395 1915 602401
rect 1857 602361 1869 602395
rect 1903 602392 1915 602395
rect 1946 602392 1952 602404
rect 1903 602364 1952 602392
rect 1903 602361 1915 602364
rect 1857 602355 1915 602361
rect 1946 602352 1952 602364
rect 2004 602352 2010 602404
rect 1946 602120 1952 602132
rect 1907 602092 1952 602120
rect 1946 602080 1952 602092
rect 2004 602080 2010 602132
rect 1765 601987 1823 601993
rect 1765 601953 1777 601987
rect 1811 601984 1823 601987
rect 1946 601984 1952 601996
rect 1811 601956 1952 601984
rect 1811 601953 1823 601956
rect 1765 601947 1823 601953
rect 1946 601944 1952 601956
rect 2004 601944 2010 601996
rect 1673 601103 1731 601109
rect 1673 601069 1685 601103
rect 1719 601100 1731 601103
rect 1946 601100 1952 601112
rect 1719 601072 1952 601100
rect 1719 601069 1731 601072
rect 1673 601063 1731 601069
rect 1946 601060 1952 601072
rect 2004 601060 2010 601112
rect 1578 600924 1584 600976
rect 1636 600964 1642 600976
rect 1946 600964 1952 600976
rect 1636 600936 1952 600964
rect 1636 600924 1642 600936
rect 1946 600924 1952 600936
rect 2004 600924 2010 600976
rect 1673 600559 1731 600565
rect 1673 600525 1685 600559
rect 1719 600556 1731 600559
rect 1946 600556 1952 600568
rect 1719 600528 1952 600556
rect 1719 600525 1731 600528
rect 1673 600519 1731 600525
rect 1946 600516 1952 600528
rect 2004 600516 2010 600568
rect 1946 599876 1952 599888
rect 1907 599848 1952 599876
rect 1946 599836 1952 599848
rect 2004 599836 2010 599888
rect 1765 599743 1823 599749
rect 1765 599709 1777 599743
rect 1811 599740 1823 599743
rect 1946 599740 1952 599752
rect 1811 599712 1952 599740
rect 1811 599709 1823 599712
rect 1765 599703 1823 599709
rect 1946 599700 1952 599712
rect 2004 599700 2010 599752
rect 1857 597023 1915 597029
rect 1857 596989 1869 597023
rect 1903 597020 1915 597023
rect 1946 597020 1952 597032
rect 1903 596992 1952 597020
rect 1903 596989 1915 596992
rect 1857 596983 1915 596989
rect 1946 596980 1952 596992
rect 2004 596980 2010 597032
rect 1670 591948 1676 592000
rect 1728 591988 1734 592000
rect 1854 591988 1860 592000
rect 1728 591960 1860 591988
rect 1728 591948 1734 591960
rect 1854 591948 1860 591960
rect 1912 591948 1918 592000
rect 1857 580499 1915 580505
rect 1857 580465 1869 580499
rect 1903 580496 1915 580499
rect 1946 580496 1952 580508
rect 1903 580468 1952 580496
rect 1903 580465 1915 580468
rect 1857 580459 1915 580465
rect 1946 580456 1952 580468
rect 2004 580456 2010 580508
rect 1946 580224 1952 580236
rect 1907 580196 1952 580224
rect 1946 580184 1952 580196
rect 2004 580184 2010 580236
rect 1578 577260 1584 577312
rect 1636 577300 1642 577312
rect 1946 577300 1952 577312
rect 1636 577272 1952 577300
rect 1636 577260 1642 577272
rect 1946 577260 1952 577272
rect 2004 577260 2010 577312
rect 574738 574744 574744 574796
rect 574796 574784 574802 574796
rect 580258 574784 580264 574796
rect 574796 574756 580264 574784
rect 574796 574744 574802 574756
rect 580258 574744 580264 574756
rect 580316 574744 580322 574796
rect 569954 571344 569960 571396
rect 570012 571384 570018 571396
rect 572714 571384 572720 571396
rect 570012 571356 572720 571384
rect 570012 571344 570018 571356
rect 572714 571344 572720 571356
rect 572772 571344 572778 571396
rect 1946 569304 1952 569356
rect 2004 569304 2010 569356
rect 1762 569100 1768 569152
rect 1820 569140 1826 569152
rect 1964 569140 1992 569304
rect 1820 569112 1992 569140
rect 1820 569100 1826 569112
rect 1854 566624 1860 566636
rect 1815 566596 1860 566624
rect 1854 566584 1860 566596
rect 1912 566584 1918 566636
rect 1765 565539 1823 565545
rect 1765 565505 1777 565539
rect 1811 565536 1823 565539
rect 1946 565536 1952 565548
rect 1811 565508 1952 565536
rect 1811 565505 1823 565508
rect 1765 565499 1823 565505
rect 1946 565496 1952 565508
rect 2004 565496 2010 565548
rect 1673 564451 1731 564457
rect 1673 564417 1685 564451
rect 1719 564448 1731 564451
rect 1946 564448 1952 564460
rect 1719 564420 1952 564448
rect 1719 564417 1731 564420
rect 1673 564411 1731 564417
rect 1946 564408 1952 564420
rect 2004 564408 2010 564460
rect 1302 564068 1308 564120
rect 1360 564108 1366 564120
rect 1946 564108 1952 564120
rect 1360 564080 1952 564108
rect 1360 564068 1366 564080
rect 1946 564068 1952 564080
rect 2004 564068 2010 564120
rect 1854 563728 1860 563780
rect 1912 563768 1918 563780
rect 1949 563771 2007 563777
rect 1949 563768 1961 563771
rect 1912 563740 1961 563768
rect 1912 563728 1918 563740
rect 1949 563737 1961 563740
rect 1995 563737 2007 563771
rect 1949 563731 2007 563737
rect 1673 563431 1731 563437
rect 1673 563397 1685 563431
rect 1719 563428 1731 563431
rect 1946 563428 1952 563440
rect 1719 563400 1952 563428
rect 1719 563397 1731 563400
rect 1673 563391 1731 563397
rect 1946 563388 1952 563400
rect 2004 563388 2010 563440
rect 1765 563159 1823 563165
rect 1765 563125 1777 563159
rect 1811 563156 1823 563159
rect 1946 563156 1952 563168
rect 1811 563128 1952 563156
rect 1811 563125 1823 563128
rect 1765 563119 1823 563125
rect 1946 563116 1952 563128
rect 2004 563116 2010 563168
rect 569954 563048 569960 563100
rect 570012 563088 570018 563100
rect 574738 563088 574744 563100
rect 570012 563060 574744 563088
rect 570012 563048 570018 563060
rect 574738 563048 574744 563060
rect 574796 563048 574802 563100
rect 1857 561119 1915 561125
rect 1857 561085 1869 561119
rect 1903 561116 1915 561119
rect 1946 561116 1952 561128
rect 1903 561088 1952 561116
rect 1903 561085 1915 561088
rect 1857 561079 1915 561085
rect 1946 561076 1952 561088
rect 2004 561076 2010 561128
rect 1578 556180 1584 556232
rect 1636 556220 1642 556232
rect 1946 556220 1952 556232
rect 1636 556192 1952 556220
rect 1636 556180 1642 556192
rect 1946 556180 1952 556192
rect 2004 556180 2010 556232
rect 569954 552072 569960 552084
rect 569915 552044 569960 552072
rect 569954 552032 569960 552044
rect 570012 552032 570018 552084
rect 569954 551828 569960 551880
rect 570012 551868 570018 551880
rect 572714 551868 572720 551880
rect 570012 551840 572720 551868
rect 570012 551828 570018 551840
rect 572714 551828 572720 551840
rect 572772 551828 572778 551880
rect 569954 551052 569960 551064
rect 569915 551024 569960 551052
rect 569954 551012 569960 551024
rect 570012 551012 570018 551064
rect 1854 547680 1860 547732
rect 1912 547720 1918 547732
rect 1949 547723 2007 547729
rect 1949 547720 1961 547723
rect 1912 547692 1961 547720
rect 1912 547680 1918 547692
rect 1949 547689 1961 547692
rect 1995 547689 2007 547723
rect 1949 547683 2007 547689
rect 1854 534012 1860 534064
rect 1912 534012 1918 534064
rect 1872 533860 1900 534012
rect 1854 533808 1860 533860
rect 1912 533808 1918 533860
rect 573358 532720 573364 532772
rect 573416 532760 573422 532772
rect 580166 532760 580172 532772
rect 573416 532732 580172 532760
rect 573416 532720 573422 532732
rect 580166 532720 580172 532732
rect 580224 532720 580230 532772
rect 569954 531088 569960 531140
rect 570012 531128 570018 531140
rect 570049 531131 570107 531137
rect 570049 531128 570061 531131
rect 570012 531100 570061 531128
rect 570012 531088 570018 531100
rect 570049 531097 570061 531100
rect 570095 531097 570107 531131
rect 570049 531091 570107 531097
rect 569954 530992 569960 531004
rect 569915 530964 569960 530992
rect 569954 530952 569960 530964
rect 570012 530952 570018 531004
rect 1946 529224 1952 529236
rect 1907 529196 1952 529224
rect 1946 529184 1952 529196
rect 2004 529184 2010 529236
rect 569954 528884 569960 528896
rect 569915 528856 569960 528884
rect 569954 528844 569960 528856
rect 570012 528844 570018 528896
rect 569954 528708 569960 528760
rect 570012 528748 570018 528760
rect 570049 528751 570107 528757
rect 570049 528748 570061 528751
rect 570012 528720 570061 528748
rect 570012 528708 570018 528720
rect 570049 528717 570061 528720
rect 570095 528717 570107 528751
rect 570049 528711 570107 528717
rect 1857 527731 1915 527737
rect 1857 527697 1869 527731
rect 1903 527728 1915 527731
rect 1946 527728 1952 527740
rect 1903 527700 1952 527728
rect 1903 527697 1915 527700
rect 1857 527691 1915 527697
rect 1946 527688 1952 527700
rect 2004 527688 2010 527740
rect 1765 527187 1823 527193
rect 1765 527153 1777 527187
rect 1811 527184 1823 527187
rect 1946 527184 1952 527196
rect 1811 527156 1952 527184
rect 1811 527153 1823 527156
rect 1765 527147 1823 527153
rect 1946 527144 1952 527156
rect 2004 527144 2010 527196
rect 1670 527116 1676 527128
rect 1631 527088 1676 527116
rect 1670 527076 1676 527088
rect 1728 527076 1734 527128
rect 1673 526983 1731 526989
rect 1673 526949 1685 526983
rect 1719 526980 1731 526983
rect 1762 526980 1768 526992
rect 1719 526952 1768 526980
rect 1719 526949 1731 526952
rect 1673 526943 1731 526949
rect 1762 526940 1768 526952
rect 1820 526940 1826 526992
rect 1673 526507 1731 526513
rect 1673 526473 1685 526507
rect 1719 526504 1731 526507
rect 1946 526504 1952 526516
rect 1719 526476 1952 526504
rect 1719 526473 1731 526476
rect 1673 526467 1731 526473
rect 1946 526464 1952 526476
rect 2004 526464 2010 526516
rect 1578 526328 1584 526380
rect 1636 526368 1642 526380
rect 1946 526368 1952 526380
rect 1636 526340 1952 526368
rect 1636 526328 1642 526340
rect 1946 526328 1952 526340
rect 2004 526328 2010 526380
rect 1673 526167 1731 526173
rect 1673 526133 1685 526167
rect 1719 526164 1731 526167
rect 1946 526164 1952 526176
rect 1719 526136 1952 526164
rect 1719 526133 1731 526136
rect 1673 526127 1731 526133
rect 1946 526124 1952 526136
rect 2004 526124 2010 526176
rect 569954 522628 569960 522640
rect 569915 522600 569960 522628
rect 569954 522588 569960 522600
rect 570012 522588 570018 522640
rect 1765 522495 1823 522501
rect 1765 522461 1777 522495
rect 1811 522492 1823 522495
rect 1946 522492 1952 522504
rect 1811 522464 1952 522492
rect 1811 522461 1823 522464
rect 1765 522455 1823 522461
rect 1946 522452 1952 522464
rect 2004 522452 2010 522504
rect 569954 522452 569960 522504
rect 570012 522492 570018 522504
rect 570049 522495 570107 522501
rect 570049 522492 570061 522495
rect 570012 522464 570061 522492
rect 570012 522452 570018 522464
rect 570049 522461 570061 522464
rect 570095 522461 570107 522495
rect 570049 522455 570107 522461
rect 1857 522359 1915 522365
rect 1857 522325 1869 522359
rect 1903 522356 1915 522359
rect 1946 522356 1952 522368
rect 1903 522328 1952 522356
rect 1903 522325 1915 522328
rect 1857 522319 1915 522325
rect 1946 522316 1952 522328
rect 2004 522316 2010 522368
rect 569954 522316 569960 522368
rect 570012 522356 570018 522368
rect 573358 522356 573364 522368
rect 570012 522328 573364 522356
rect 570012 522316 570018 522328
rect 573358 522316 573364 522328
rect 573416 522316 573422 522368
rect 569954 521024 569960 521076
rect 570012 521064 570018 521076
rect 570049 521067 570107 521073
rect 570049 521064 570061 521067
rect 570012 521036 570061 521064
rect 570012 521024 570018 521036
rect 570049 521033 570061 521036
rect 570095 521033 570107 521067
rect 570049 521027 570107 521033
rect 569954 518480 569960 518492
rect 569915 518452 569960 518480
rect 569954 518440 569960 518452
rect 570012 518440 570018 518492
rect 1946 510660 1952 510672
rect 1907 510632 1952 510660
rect 1946 510620 1952 510632
rect 2004 510620 2010 510672
rect 1946 510048 1952 510060
rect 1907 510020 1952 510048
rect 1946 510008 1952 510020
rect 2004 510008 2010 510060
rect 1762 509912 1768 509924
rect 1688 509884 1768 509912
rect 1688 509584 1716 509884
rect 1762 509872 1768 509884
rect 1820 509872 1826 509924
rect 1857 509915 1915 509921
rect 1857 509881 1869 509915
rect 1903 509912 1915 509915
rect 1946 509912 1952 509924
rect 1903 509884 1952 509912
rect 1903 509881 1915 509884
rect 1857 509875 1915 509881
rect 1946 509872 1952 509884
rect 2004 509872 2010 509924
rect 1670 509532 1676 509584
rect 1728 509532 1734 509584
rect 1581 507331 1639 507337
rect 1581 507297 1593 507331
rect 1627 507328 1639 507331
rect 1946 507328 1952 507340
rect 1627 507300 1952 507328
rect 1627 507297 1639 507300
rect 1581 507291 1639 507297
rect 1946 507288 1952 507300
rect 2004 507288 2010 507340
rect 1489 507195 1547 507201
rect 1489 507161 1501 507195
rect 1535 507192 1547 507195
rect 1946 507192 1952 507204
rect 1535 507164 1952 507192
rect 1535 507161 1547 507164
rect 1489 507155 1547 507161
rect 1946 507152 1952 507164
rect 2004 507152 2010 507204
rect 1765 506107 1823 506113
rect 1765 506073 1777 506107
rect 1811 506104 1823 506107
rect 1946 506104 1952 506116
rect 1811 506076 1952 506104
rect 1811 506073 1823 506076
rect 1765 506067 1823 506073
rect 1946 506064 1952 506076
rect 2004 506064 2010 506116
rect 1578 505180 1584 505232
rect 1636 505220 1642 505232
rect 1946 505220 1952 505232
rect 1636 505192 1952 505220
rect 1636 505180 1642 505192
rect 1946 505180 1952 505192
rect 2004 505180 2010 505232
rect 569954 505152 569960 505164
rect 569915 505124 569960 505152
rect 569954 505112 569960 505124
rect 570012 505112 570018 505164
rect 1765 504883 1823 504889
rect 1765 504849 1777 504883
rect 1811 504880 1823 504883
rect 1811 504852 1992 504880
rect 1811 504849 1823 504852
rect 1765 504843 1823 504849
rect 1964 504824 1992 504852
rect 1946 504772 1952 504824
rect 2004 504772 2010 504824
rect 1854 504472 1860 504484
rect 1815 504444 1860 504472
rect 1854 504432 1860 504444
rect 1912 504432 1918 504484
rect 569954 504160 569960 504212
rect 570012 504200 570018 504212
rect 570049 504203 570107 504209
rect 570049 504200 570061 504203
rect 570012 504172 570061 504200
rect 570012 504160 570018 504172
rect 570049 504169 570061 504172
rect 570095 504169 570107 504203
rect 570049 504163 570107 504169
rect 1762 504132 1768 504144
rect 1723 504104 1768 504132
rect 1762 504092 1768 504104
rect 1820 504092 1826 504144
rect 569954 503140 569960 503192
rect 570012 503180 570018 503192
rect 570049 503183 570107 503189
rect 570049 503180 570061 503183
rect 570012 503152 570061 503180
rect 570012 503140 570018 503152
rect 570049 503149 570061 503152
rect 570095 503149 570107 503183
rect 570049 503143 570107 503149
rect 569954 503044 569960 503056
rect 569915 503016 569960 503044
rect 569954 503004 569960 503016
rect 570012 503004 570018 503056
rect 1670 502296 1676 502308
rect 1631 502268 1676 502296
rect 1670 502256 1676 502268
rect 1728 502256 1734 502308
rect 1489 502231 1547 502237
rect 1489 502197 1501 502231
rect 1535 502228 1547 502231
rect 1946 502228 1952 502240
rect 1535 502200 1952 502228
rect 1535 502197 1547 502200
rect 1489 502191 1547 502197
rect 1946 502188 1952 502200
rect 2004 502188 2010 502240
rect 1581 501823 1639 501829
rect 1581 501789 1593 501823
rect 1627 501820 1639 501823
rect 1946 501820 1952 501832
rect 1627 501792 1952 501820
rect 1627 501789 1639 501792
rect 1581 501783 1639 501789
rect 1946 501780 1952 501792
rect 2004 501780 2010 501832
rect 1762 497536 1768 497548
rect 1723 497508 1768 497536
rect 1762 497496 1768 497508
rect 1820 497496 1826 497548
rect 1946 497536 1952 497548
rect 1907 497508 1952 497536
rect 1946 497496 1952 497508
rect 2004 497496 2010 497548
rect 1673 493391 1731 493397
rect 1673 493357 1685 493391
rect 1719 493388 1731 493391
rect 1854 493388 1860 493400
rect 1719 493360 1860 493388
rect 1719 493357 1731 493360
rect 1673 493351 1731 493357
rect 1854 493348 1860 493360
rect 1912 493348 1918 493400
rect 569954 487092 569960 487144
rect 570012 487132 570018 487144
rect 579798 487132 579804 487144
rect 570012 487104 579804 487132
rect 570012 487092 570018 487104
rect 579798 487092 579804 487104
rect 579856 487092 579862 487144
rect 569954 486956 569960 487008
rect 570012 486996 570018 487008
rect 570138 486996 570144 487008
rect 570012 486968 570144 486996
rect 570012 486956 570018 486968
rect 570138 486956 570144 486968
rect 570196 486956 570202 487008
rect 1673 483735 1731 483741
rect 1673 483701 1685 483735
rect 1719 483732 1731 483735
rect 1762 483732 1768 483744
rect 1719 483704 1768 483732
rect 1719 483701 1731 483704
rect 1673 483695 1731 483701
rect 1762 483692 1768 483704
rect 1820 483692 1826 483744
rect 1946 479544 1952 479596
rect 2004 479544 2010 479596
rect 1964 479392 1992 479544
rect 1946 479340 1952 479392
rect 2004 479340 2010 479392
rect 1946 474688 1952 474700
rect 1907 474660 1952 474688
rect 1946 474648 1952 474660
rect 2004 474648 2010 474700
rect 1854 474076 1860 474088
rect 1815 474048 1860 474076
rect 1854 474036 1860 474048
rect 1912 474036 1918 474088
rect 1670 472744 1676 472796
rect 1728 472784 1734 472796
rect 1946 472784 1952 472796
rect 1728 472756 1952 472784
rect 1728 472744 1734 472756
rect 1946 472744 1952 472756
rect 2004 472744 2010 472796
rect 1762 472104 1768 472116
rect 1723 472076 1768 472104
rect 1762 472064 1768 472076
rect 1820 472064 1826 472116
rect 1026 469752 1032 469804
rect 1084 469792 1090 469804
rect 1946 469792 1952 469804
rect 1084 469764 1952 469792
rect 1084 469752 1090 469764
rect 1946 469752 1952 469764
rect 2004 469752 2010 469804
rect 569954 468568 569960 468580
rect 569915 468540 569960 468568
rect 569954 468528 569960 468540
rect 570012 468528 570018 468580
rect 1946 468256 1952 468308
rect 2004 468256 2010 468308
rect 569954 468256 569960 468308
rect 570012 468296 570018 468308
rect 570141 468299 570199 468305
rect 570141 468296 570153 468299
rect 570012 468268 570153 468296
rect 570012 468256 570018 468268
rect 570141 468265 570153 468268
rect 570187 468265 570199 468299
rect 570141 468259 570199 468265
rect 1964 468104 1992 468256
rect 1946 468052 1952 468104
rect 2004 468052 2010 468104
rect 1857 467619 1915 467625
rect 1857 467585 1869 467619
rect 1903 467616 1915 467619
rect 1946 467616 1952 467628
rect 1903 467588 1952 467616
rect 1903 467585 1915 467588
rect 1857 467579 1915 467585
rect 1946 467576 1952 467588
rect 2004 467576 2010 467628
rect 569954 467576 569960 467628
rect 570012 467616 570018 467628
rect 570233 467619 570291 467625
rect 570233 467616 570245 467619
rect 570012 467588 570245 467616
rect 570012 467576 570018 467588
rect 570233 467585 570245 467588
rect 570279 467585 570291 467619
rect 570233 467579 570291 467585
rect 570046 467072 570052 467084
rect 570007 467044 570052 467072
rect 570046 467032 570052 467044
rect 570104 467032 570110 467084
rect 570046 466828 570052 466880
rect 570104 466868 570110 466880
rect 570141 466871 570199 466877
rect 570141 466868 570153 466871
rect 570104 466840 570153 466868
rect 570104 466828 570110 466840
rect 570141 466837 570153 466840
rect 570187 466837 570199 466871
rect 570141 466831 570199 466837
rect 569957 466599 570015 466605
rect 569957 466565 569969 466599
rect 570003 466596 570015 466599
rect 570233 466599 570291 466605
rect 570233 466596 570245 466599
rect 570003 466568 570245 466596
rect 570003 466565 570015 466568
rect 569957 466559 570015 466565
rect 570233 466565 570245 466568
rect 570279 466565 570291 466599
rect 570233 466559 570291 466565
rect 570049 465511 570107 465517
rect 570049 465477 570061 465511
rect 570095 465508 570107 465511
rect 570325 465511 570383 465517
rect 570325 465508 570337 465511
rect 570095 465480 570337 465508
rect 570095 465477 570107 465480
rect 570049 465471 570107 465477
rect 570325 465477 570337 465480
rect 570371 465477 570383 465511
rect 570325 465471 570383 465477
rect 570046 465332 570052 465384
rect 570104 465372 570110 465384
rect 570141 465375 570199 465381
rect 570141 465372 570153 465375
rect 570104 465344 570153 465372
rect 570104 465332 570110 465344
rect 570141 465341 570153 465344
rect 570187 465341 570199 465375
rect 570141 465335 570199 465341
rect 569954 465196 569960 465248
rect 570012 465236 570018 465248
rect 570049 465239 570107 465245
rect 570049 465236 570061 465239
rect 570012 465208 570061 465236
rect 570012 465196 570018 465208
rect 570049 465205 570061 465208
rect 570095 465205 570107 465239
rect 570049 465199 570107 465205
rect 570138 465196 570144 465248
rect 570196 465196 570202 465248
rect 570156 465112 570184 465196
rect 570138 465060 570144 465112
rect 570196 465060 570202 465112
rect 1673 464967 1731 464973
rect 1673 464933 1685 464967
rect 1719 464964 1731 464967
rect 1946 464964 1952 464976
rect 1719 464936 1952 464964
rect 1719 464933 1731 464936
rect 1673 464927 1731 464933
rect 1946 464924 1952 464936
rect 2004 464924 2010 464976
rect 569862 464244 569868 464296
rect 569920 464244 569926 464296
rect 569880 464148 569908 464244
rect 570046 464148 570052 464160
rect 569880 464120 570052 464148
rect 570046 464108 570052 464120
rect 570104 464108 570110 464160
rect 569954 464012 569960 464024
rect 569880 463984 569960 464012
rect 569880 463740 569908 463984
rect 569954 463972 569960 463984
rect 570012 463972 570018 464024
rect 569954 463836 569960 463888
rect 570012 463876 570018 463888
rect 570325 463879 570383 463885
rect 570325 463876 570337 463879
rect 570012 463848 570337 463876
rect 570012 463836 570018 463848
rect 570325 463845 570337 463848
rect 570371 463845 570383 463879
rect 570325 463839 570383 463845
rect 569954 463740 569960 463752
rect 569880 463712 569960 463740
rect 569954 463700 569960 463712
rect 570012 463700 570018 463752
rect 569954 463564 569960 463616
rect 570012 463604 570018 463616
rect 570049 463607 570107 463613
rect 570049 463604 570061 463607
rect 570012 463576 570061 463604
rect 570012 463564 570018 463576
rect 570049 463573 570061 463576
rect 570095 463573 570107 463607
rect 570049 463567 570107 463573
rect 570046 462748 570052 462800
rect 570104 462788 570110 462800
rect 570141 462791 570199 462797
rect 570141 462788 570153 462791
rect 570104 462760 570153 462788
rect 570104 462748 570110 462760
rect 570141 462757 570153 462760
rect 570187 462757 570199 462791
rect 570141 462751 570199 462757
rect 1946 462380 1952 462392
rect 1907 462352 1952 462380
rect 1946 462340 1952 462352
rect 2004 462340 2010 462392
rect 569954 461700 569960 461712
rect 569915 461672 569960 461700
rect 569954 461660 569960 461672
rect 570012 461660 570018 461712
rect 569954 461428 569960 461440
rect 569915 461400 569960 461428
rect 569954 461388 569960 461400
rect 570012 461388 570018 461440
rect 1394 459824 1400 459876
rect 1452 459864 1458 459876
rect 1854 459864 1860 459876
rect 1452 459836 1860 459864
rect 1452 459824 1458 459836
rect 1854 459824 1860 459836
rect 1912 459824 1918 459876
rect 1946 454628 1952 454640
rect 1907 454600 1952 454628
rect 1946 454588 1952 454600
rect 2004 454588 2010 454640
rect 1762 450848 1768 450900
rect 1820 450888 1826 450900
rect 1946 450888 1952 450900
rect 1820 450860 1952 450888
rect 1820 450848 1826 450860
rect 1946 450848 1952 450860
rect 2004 450848 2010 450900
rect 1581 450755 1639 450761
rect 1581 450721 1593 450755
rect 1627 450752 1639 450755
rect 1946 450752 1952 450764
rect 1627 450724 1952 450752
rect 1627 450721 1639 450724
rect 1581 450715 1639 450721
rect 1946 450712 1952 450724
rect 2004 450712 2010 450764
rect 1765 450075 1823 450081
rect 1765 450041 1777 450075
rect 1811 450072 1823 450075
rect 1946 450072 1952 450084
rect 1811 450044 1952 450072
rect 1811 450041 1823 450044
rect 1765 450035 1823 450041
rect 1946 450032 1952 450044
rect 2004 450032 2010 450084
rect 1397 449939 1455 449945
rect 1397 449905 1409 449939
rect 1443 449936 1455 449939
rect 1946 449936 1952 449948
rect 1443 449908 1952 449936
rect 1443 449905 1455 449908
rect 1397 449899 1455 449905
rect 1946 449896 1952 449908
rect 2004 449896 2010 449948
rect 569954 449352 569960 449404
rect 570012 449352 570018 449404
rect 569972 449200 570000 449352
rect 1854 449188 1860 449200
rect 1815 449160 1860 449188
rect 1854 449148 1860 449160
rect 1912 449148 1918 449200
rect 569954 449148 569960 449200
rect 570012 449148 570018 449200
rect 1581 449055 1639 449061
rect 1581 449021 1593 449055
rect 1627 449052 1639 449055
rect 1854 449052 1860 449064
rect 1627 449024 1860 449052
rect 1627 449021 1639 449024
rect 1581 449015 1639 449021
rect 1854 449012 1860 449024
rect 1912 449012 1918 449064
rect 1581 448783 1639 448789
rect 1581 448749 1593 448783
rect 1627 448780 1639 448783
rect 1946 448780 1952 448792
rect 1627 448752 1952 448780
rect 1627 448749 1639 448752
rect 1581 448743 1639 448749
rect 1946 448740 1952 448752
rect 2004 448740 2010 448792
rect 1670 448712 1676 448724
rect 1631 448684 1676 448712
rect 1670 448672 1676 448684
rect 1728 448672 1734 448724
rect 1394 448604 1400 448656
rect 1452 448644 1458 448656
rect 1946 448644 1952 448656
rect 1452 448616 1952 448644
rect 1452 448604 1458 448616
rect 1946 448604 1952 448616
rect 2004 448604 2010 448656
rect 1581 448511 1639 448517
rect 1581 448477 1593 448511
rect 1627 448508 1639 448511
rect 1946 448508 1952 448520
rect 1627 448480 1952 448508
rect 1627 448477 1639 448480
rect 1581 448471 1639 448477
rect 1946 448468 1952 448480
rect 2004 448468 2010 448520
rect 1397 447967 1455 447973
rect 1397 447933 1409 447967
rect 1443 447964 1455 447967
rect 1946 447964 1952 447976
rect 1443 447936 1952 447964
rect 1443 447933 1455 447936
rect 1397 447927 1455 447933
rect 1946 447924 1952 447936
rect 2004 447924 2010 447976
rect 1765 447831 1823 447837
rect 1765 447797 1777 447831
rect 1811 447828 1823 447831
rect 1946 447828 1952 447840
rect 1811 447800 1952 447828
rect 1811 447797 1823 447800
rect 1765 447791 1823 447797
rect 1946 447788 1952 447800
rect 2004 447788 2010 447840
rect 1765 442323 1823 442329
rect 1765 442289 1777 442323
rect 1811 442320 1823 442323
rect 1854 442320 1860 442332
rect 1811 442292 1860 442320
rect 1811 442289 1823 442292
rect 1765 442283 1823 442289
rect 1854 442280 1860 442292
rect 1912 442280 1918 442332
rect 569954 441600 569960 441652
rect 570012 441640 570018 441652
rect 570049 441643 570107 441649
rect 570049 441640 570061 441643
rect 570012 441612 570061 441640
rect 570012 441600 570018 441612
rect 570049 441609 570061 441612
rect 570095 441609 570107 441643
rect 570049 441603 570107 441609
rect 1765 441439 1823 441445
rect 1765 441405 1777 441439
rect 1811 441436 1823 441439
rect 1946 441436 1952 441448
rect 1811 441408 1952 441436
rect 1811 441405 1823 441408
rect 1765 441399 1823 441405
rect 1946 441396 1952 441408
rect 2004 441396 2010 441448
rect 1854 440960 1860 440972
rect 1815 440932 1860 440960
rect 1854 440920 1860 440932
rect 1912 440920 1918 440972
rect 1946 439192 1952 439204
rect 1907 439164 1952 439192
rect 1946 439152 1952 439164
rect 2004 439152 2010 439204
rect 574738 438880 574744 438932
rect 574796 438920 574802 438932
rect 580166 438920 580172 438932
rect 574796 438892 580172 438920
rect 574796 438880 574802 438892
rect 580166 438880 580172 438892
rect 580224 438880 580230 438932
rect 570046 436812 570052 436824
rect 570007 436784 570052 436812
rect 570046 436772 570052 436784
rect 570104 436772 570110 436824
rect 1946 434228 1952 434240
rect 1907 434200 1952 434228
rect 1946 434188 1952 434200
rect 2004 434188 2010 434240
rect 569954 432528 569960 432540
rect 569915 432500 569960 432528
rect 569954 432488 569960 432500
rect 570012 432488 570018 432540
rect 1670 432216 1676 432268
rect 1728 432256 1734 432268
rect 1946 432256 1952 432268
rect 1728 432228 1952 432256
rect 1728 432216 1734 432228
rect 1946 432216 1952 432228
rect 2004 432216 2010 432268
rect 1946 425728 1952 425740
rect 1907 425700 1952 425728
rect 1946 425688 1952 425700
rect 2004 425688 2010 425740
rect 1394 425552 1400 425604
rect 1452 425592 1458 425604
rect 1762 425592 1768 425604
rect 1452 425564 1768 425592
rect 1452 425552 1458 425564
rect 1762 425552 1768 425564
rect 1820 425552 1826 425604
rect 1394 419840 1400 419892
rect 1452 419880 1458 419892
rect 1670 419880 1676 419892
rect 1452 419852 1676 419880
rect 1452 419840 1458 419852
rect 1670 419840 1676 419852
rect 1728 419840 1734 419892
rect 569954 418276 569960 418328
rect 570012 418316 570018 418328
rect 570012 418288 570092 418316
rect 570012 418276 570018 418288
rect 569954 418180 569960 418192
rect 569915 418152 569960 418180
rect 569954 418140 569960 418152
rect 570012 418140 570018 418192
rect 569957 418047 570015 418053
rect 569957 418013 569969 418047
rect 570003 418044 570015 418047
rect 570064 418044 570092 418288
rect 570003 418016 570092 418044
rect 570003 418013 570015 418016
rect 569957 418007 570015 418013
rect 1854 414944 1860 414996
rect 1912 414944 1918 414996
rect 1946 414944 1952 414996
rect 2004 414984 2010 414996
rect 2004 414956 2049 414984
rect 2004 414944 2010 414956
rect 1872 414792 1900 414944
rect 1854 414740 1860 414792
rect 1912 414740 1918 414792
rect 1394 414604 1400 414656
rect 1452 414644 1458 414656
rect 1670 414644 1676 414656
rect 1452 414616 1676 414644
rect 1452 414604 1458 414616
rect 1670 414604 1676 414616
rect 1728 414604 1734 414656
rect 570598 411952 570604 412004
rect 570656 411992 570662 412004
rect 572714 411992 572720 412004
rect 570656 411964 572720 411992
rect 570656 411952 570662 411964
rect 572714 411952 572720 411964
rect 572772 411952 572778 412004
rect 1946 407300 1952 407312
rect 1907 407272 1952 407300
rect 1946 407260 1952 407272
rect 2004 407260 2010 407312
rect 569954 407056 569960 407108
rect 570012 407096 570018 407108
rect 570046 407096 570052 407108
rect 570012 407068 570052 407096
rect 570012 407056 570018 407068
rect 570046 407056 570052 407068
rect 570104 407056 570110 407108
rect 1946 405668 1952 405680
rect 1907 405640 1952 405668
rect 1946 405628 1952 405640
rect 2004 405628 2010 405680
rect 1854 405600 1860 405612
rect 1815 405572 1860 405600
rect 1854 405560 1860 405572
rect 1912 405560 1918 405612
rect 1394 405424 1400 405476
rect 1452 405464 1458 405476
rect 1762 405464 1768 405476
rect 1452 405436 1768 405464
rect 1452 405424 1458 405436
rect 1762 405424 1768 405436
rect 1820 405424 1826 405476
rect 569954 402268 569960 402280
rect 569915 402240 569960 402268
rect 569954 402228 569960 402240
rect 570012 402228 570018 402280
rect 569954 401616 569960 401668
rect 570012 401656 570018 401668
rect 570598 401656 570604 401668
rect 570012 401628 570604 401656
rect 570012 401616 570018 401628
rect 570598 401616 570604 401628
rect 570656 401616 570662 401668
rect 569957 399551 570015 399557
rect 569957 399517 569969 399551
rect 570003 399548 570015 399551
rect 570046 399548 570052 399560
rect 570003 399520 570052 399548
rect 570003 399517 570015 399520
rect 569957 399511 570015 399517
rect 570046 399508 570052 399520
rect 570104 399508 570110 399560
rect 1394 398420 1400 398472
rect 1452 398460 1458 398472
rect 1762 398460 1768 398472
rect 1452 398432 1768 398460
rect 1452 398420 1458 398432
rect 1762 398420 1768 398432
rect 1820 398420 1826 398472
rect 569954 396788 569960 396840
rect 570012 396828 570018 396840
rect 570049 396831 570107 396837
rect 570049 396828 570061 396831
rect 570012 396800 570061 396828
rect 570012 396788 570018 396800
rect 570049 396797 570061 396800
rect 570095 396797 570107 396831
rect 570049 396791 570107 396797
rect 569954 394952 569960 395004
rect 570012 394992 570018 395004
rect 570233 394995 570291 395001
rect 570233 394992 570245 394995
rect 570012 394964 570245 394992
rect 570012 394952 570018 394964
rect 570233 394961 570245 394964
rect 570279 394961 570291 394995
rect 570233 394955 570291 394961
rect 570046 394612 570052 394664
rect 570104 394652 570110 394664
rect 570230 394652 570236 394664
rect 570104 394624 570236 394652
rect 570104 394612 570110 394624
rect 570230 394612 570236 394624
rect 570288 394612 570294 394664
rect 1854 393972 1860 393984
rect 1815 393944 1860 393972
rect 1854 393932 1860 393944
rect 1912 393932 1918 393984
rect 569954 393796 569960 393848
rect 570012 393836 570018 393848
rect 570141 393839 570199 393845
rect 570141 393836 570153 393839
rect 570012 393808 570153 393836
rect 570012 393796 570018 393808
rect 570141 393805 570153 393808
rect 570187 393805 570199 393839
rect 570141 393799 570199 393805
rect 569954 393700 569960 393712
rect 569915 393672 569960 393700
rect 569954 393660 569960 393672
rect 570012 393660 570018 393712
rect 1946 393496 1952 393508
rect 1907 393468 1952 393496
rect 1946 393456 1952 393468
rect 2004 393456 2010 393508
rect 569954 393116 569960 393168
rect 570012 393156 570018 393168
rect 570325 393159 570383 393165
rect 570325 393156 570337 393159
rect 570012 393128 570337 393156
rect 570012 393116 570018 393128
rect 570325 393125 570337 393128
rect 570371 393125 570383 393159
rect 570325 393119 570383 393125
rect 569954 392912 569960 392964
rect 570012 392912 570018 392964
rect 569972 392760 570000 392912
rect 569954 392708 569960 392760
rect 570012 392708 570018 392760
rect 569954 392572 569960 392624
rect 570012 392612 570018 392624
rect 570322 392612 570328 392624
rect 570012 392584 570328 392612
rect 570012 392572 570018 392584
rect 570322 392572 570328 392584
rect 570380 392572 570386 392624
rect 569954 392300 569960 392352
rect 570012 392340 570018 392352
rect 570049 392343 570107 392349
rect 570049 392340 570061 392343
rect 570012 392312 570061 392340
rect 570012 392300 570018 392312
rect 570049 392309 570061 392312
rect 570095 392309 570107 392343
rect 570049 392303 570107 392309
rect 574830 391960 574836 392012
rect 574888 392000 574894 392012
rect 580166 392000 580172 392012
rect 574888 391972 580172 392000
rect 574888 391960 574894 391972
rect 580166 391960 580172 391972
rect 580224 391960 580230 392012
rect 569954 389988 569960 390040
rect 570012 390028 570018 390040
rect 570325 390031 570383 390037
rect 570325 390028 570337 390031
rect 570012 390000 570337 390028
rect 570012 389988 570018 390000
rect 570325 389997 570337 390000
rect 570371 389997 570383 390031
rect 570325 389991 570383 389997
rect 569954 389892 569960 389904
rect 569915 389864 569960 389892
rect 569954 389852 569960 389864
rect 570012 389852 570018 389904
rect 569954 389036 569960 389088
rect 570012 389076 570018 389088
rect 570141 389079 570199 389085
rect 570141 389076 570153 389079
rect 570012 389048 570153 389076
rect 570012 389036 570018 389048
rect 570141 389045 570153 389048
rect 570187 389045 570199 389079
rect 570141 389039 570199 389045
rect 569954 388492 569960 388544
rect 570012 388532 570018 388544
rect 570233 388535 570291 388541
rect 570233 388532 570245 388535
rect 570012 388504 570245 388532
rect 570012 388492 570018 388504
rect 570233 388501 570245 388504
rect 570279 388501 570291 388535
rect 570233 388495 570291 388501
rect 569954 388356 569960 388408
rect 570012 388396 570018 388408
rect 570230 388396 570236 388408
rect 570012 388368 570236 388396
rect 570012 388356 570018 388368
rect 570230 388356 570236 388368
rect 570288 388356 570294 388408
rect 1765 387379 1823 387385
rect 1765 387345 1777 387379
rect 1811 387376 1823 387379
rect 1946 387376 1952 387388
rect 1811 387348 1952 387376
rect 1811 387345 1823 387348
rect 1765 387339 1823 387345
rect 1946 387336 1952 387348
rect 2004 387336 2010 387388
rect 1857 387243 1915 387249
rect 1857 387209 1869 387243
rect 1903 387240 1915 387243
rect 1946 387240 1952 387252
rect 1903 387212 1952 387240
rect 1903 387209 1915 387212
rect 1857 387203 1915 387209
rect 1946 387200 1952 387212
rect 2004 387200 2010 387252
rect 1394 387104 1400 387116
rect 1355 387076 1400 387104
rect 1394 387064 1400 387076
rect 1452 387064 1458 387116
rect 1762 387064 1768 387116
rect 1820 387064 1826 387116
rect 1946 387104 1952 387116
rect 1907 387076 1952 387104
rect 1946 387064 1952 387076
rect 2004 387064 2010 387116
rect 1780 387036 1808 387064
rect 1412 387008 1808 387036
rect 1412 386980 1440 387008
rect 1394 386928 1400 386980
rect 1452 386928 1458 386980
rect 1762 386928 1768 386980
rect 1820 386968 1826 386980
rect 1946 386968 1952 386980
rect 1820 386940 1952 386968
rect 1820 386928 1826 386940
rect 1946 386928 1952 386940
rect 2004 386928 2010 386980
rect 569954 382820 569960 382832
rect 569915 382792 569960 382820
rect 569954 382780 569960 382792
rect 570012 382780 570018 382832
rect 569865 382687 569923 382693
rect 569865 382653 569877 382687
rect 569911 382684 569923 382687
rect 569954 382684 569960 382696
rect 569911 382656 569960 382684
rect 569911 382653 569923 382656
rect 569865 382647 569923 382653
rect 569954 382644 569960 382656
rect 570012 382644 570018 382696
rect 569954 381828 569960 381880
rect 570012 381868 570018 381880
rect 570049 381871 570107 381877
rect 570049 381868 570061 381871
rect 570012 381840 570061 381868
rect 570012 381828 570018 381840
rect 570049 381837 570061 381840
rect 570095 381837 570107 381871
rect 570049 381831 570107 381837
rect 1581 381463 1639 381469
rect 1581 381429 1593 381463
rect 1627 381460 1639 381463
rect 1949 381463 2007 381469
rect 1949 381460 1961 381463
rect 1627 381432 1961 381460
rect 1627 381429 1639 381432
rect 1581 381423 1639 381429
rect 1949 381429 1961 381432
rect 1995 381429 2007 381463
rect 1949 381423 2007 381429
rect 1397 381191 1455 381197
rect 1397 381157 1409 381191
rect 1443 381188 1455 381191
rect 1946 381188 1952 381200
rect 1443 381160 1952 381188
rect 1443 381157 1455 381160
rect 1397 381151 1455 381157
rect 1946 381148 1952 381160
rect 2004 381148 2010 381200
rect 1673 380715 1731 380721
rect 1673 380681 1685 380715
rect 1719 380712 1731 380715
rect 1762 380712 1768 380724
rect 1719 380684 1768 380712
rect 1719 380681 1731 380684
rect 1673 380675 1731 380681
rect 1762 380672 1768 380684
rect 1820 380672 1826 380724
rect 1857 380715 1915 380721
rect 1857 380681 1869 380715
rect 1903 380712 1915 380715
rect 1946 380712 1952 380724
rect 1903 380684 1952 380712
rect 1903 380681 1915 380684
rect 1857 380675 1915 380681
rect 1946 380672 1952 380684
rect 2004 380672 2010 380724
rect 1394 380536 1400 380588
rect 1452 380576 1458 380588
rect 1762 380576 1768 380588
rect 1452 380548 1768 380576
rect 1452 380536 1458 380548
rect 1762 380536 1768 380548
rect 1820 380536 1826 380588
rect 1581 379151 1639 379157
rect 1581 379117 1593 379151
rect 1627 379148 1639 379151
rect 1946 379148 1952 379160
rect 1627 379120 1952 379148
rect 1627 379117 1639 379120
rect 1581 379111 1639 379117
rect 1946 379108 1952 379120
rect 2004 379108 2010 379160
rect 1673 379015 1731 379021
rect 1673 378981 1685 379015
rect 1719 379012 1731 379015
rect 1946 379012 1952 379024
rect 1719 378984 1952 379012
rect 1719 378981 1731 378984
rect 1673 378975 1731 378981
rect 1946 378972 1952 378984
rect 2004 378972 2010 379024
rect 1765 376771 1823 376777
rect 1765 376737 1777 376771
rect 1811 376768 1823 376771
rect 1946 376768 1952 376780
rect 1811 376740 1952 376768
rect 1811 376737 1823 376740
rect 1765 376731 1823 376737
rect 1946 376728 1952 376740
rect 2004 376728 2010 376780
rect 569954 376700 569960 376712
rect 569915 376672 569960 376700
rect 569954 376660 569960 376672
rect 570012 376660 570018 376712
rect 570138 376660 570144 376712
rect 570196 376700 570202 376712
rect 570233 376703 570291 376709
rect 570233 376700 570245 376703
rect 570196 376672 570245 376700
rect 570196 376660 570202 376672
rect 570233 376669 570245 376672
rect 570279 376669 570291 376703
rect 570233 376663 570291 376669
rect 569954 376524 569960 376576
rect 570012 376564 570018 376576
rect 570049 376567 570107 376573
rect 570049 376564 570061 376567
rect 570012 376536 570061 376564
rect 570012 376524 570018 376536
rect 570049 376533 570061 376536
rect 570095 376533 570107 376567
rect 570049 376527 570107 376533
rect 1946 370648 1952 370660
rect 1907 370620 1952 370648
rect 1946 370608 1952 370620
rect 2004 370608 2010 370660
rect 1670 370512 1676 370524
rect 1631 370484 1676 370512
rect 1670 370472 1676 370484
rect 1728 370472 1734 370524
rect 1857 370379 1915 370385
rect 1857 370345 1869 370379
rect 1903 370376 1915 370379
rect 1946 370376 1952 370388
rect 1903 370348 1952 370376
rect 1903 370345 1915 370348
rect 1857 370339 1915 370345
rect 1946 370336 1952 370348
rect 2004 370336 2010 370388
rect 1765 370243 1823 370249
rect 1765 370209 1777 370243
rect 1811 370240 1823 370243
rect 1946 370240 1952 370252
rect 1811 370212 1952 370240
rect 1811 370209 1823 370212
rect 1765 370203 1823 370209
rect 1946 370200 1952 370212
rect 2004 370200 2010 370252
rect 569954 369724 569960 369776
rect 570012 369764 570018 369776
rect 570141 369767 570199 369773
rect 570141 369764 570153 369767
rect 570012 369736 570153 369764
rect 570012 369724 570018 369736
rect 570141 369733 570153 369736
rect 570187 369733 570199 369767
rect 570141 369727 570199 369733
rect 569954 369424 569960 369436
rect 569915 369396 569960 369424
rect 569954 369384 569960 369396
rect 570012 369384 570018 369436
rect 1397 369291 1455 369297
rect 1397 369257 1409 369291
rect 1443 369288 1455 369291
rect 1946 369288 1952 369300
rect 1443 369260 1952 369288
rect 1443 369257 1455 369260
rect 1397 369251 1455 369257
rect 1946 369248 1952 369260
rect 2004 369248 2010 369300
rect 569954 368336 569960 368348
rect 569915 368308 569960 368336
rect 569954 368296 569960 368308
rect 570012 368296 570018 368348
rect 569954 368024 569960 368076
rect 570012 368064 570018 368076
rect 570138 368064 570144 368076
rect 570012 368036 570144 368064
rect 570012 368024 570018 368036
rect 570138 368024 570144 368036
rect 570196 368024 570202 368076
rect 1670 367792 1676 367804
rect 1631 367764 1676 367792
rect 1670 367752 1676 367764
rect 1728 367752 1734 367804
rect 569954 367752 569960 367804
rect 570012 367792 570018 367804
rect 570417 367795 570475 367801
rect 570417 367792 570429 367795
rect 570012 367764 570429 367792
rect 570012 367752 570018 367764
rect 570417 367761 570429 367764
rect 570463 367761 570475 367795
rect 570417 367755 570475 367761
rect 570046 362312 570052 362364
rect 570104 362352 570110 362364
rect 570230 362352 570236 362364
rect 570104 362324 570236 362352
rect 570104 362312 570110 362324
rect 570230 362312 570236 362324
rect 570288 362312 570294 362364
rect 569954 360000 569960 360052
rect 570012 360040 570018 360052
rect 570322 360040 570328 360052
rect 570012 360012 570328 360040
rect 570012 360000 570018 360012
rect 570322 360000 570328 360012
rect 570380 360000 570386 360052
rect 569954 359864 569960 359916
rect 570012 359904 570018 359916
rect 570325 359907 570383 359913
rect 570325 359904 570337 359907
rect 570012 359876 570337 359904
rect 570012 359864 570018 359876
rect 570325 359873 570337 359876
rect 570371 359873 570383 359907
rect 570325 359867 570383 359873
rect 569954 359524 569960 359576
rect 570012 359564 570018 359576
rect 570049 359567 570107 359573
rect 570049 359564 570061 359567
rect 570012 359536 570061 359564
rect 570012 359524 570018 359536
rect 570049 359533 570061 359536
rect 570095 359533 570107 359567
rect 570049 359527 570107 359533
rect 569954 359116 569960 359168
rect 570012 359156 570018 359168
rect 570509 359159 570567 359165
rect 570509 359156 570521 359159
rect 570012 359128 570521 359156
rect 570012 359116 570018 359128
rect 570509 359125 570521 359128
rect 570555 359125 570567 359159
rect 570509 359119 570567 359125
rect 569954 358884 569960 358896
rect 569880 358856 569960 358884
rect 569880 358612 569908 358856
rect 569954 358844 569960 358856
rect 570012 358844 570018 358896
rect 569954 358708 569960 358760
rect 570012 358748 570018 358760
rect 570230 358748 570236 358760
rect 570012 358720 570236 358748
rect 570012 358708 570018 358720
rect 570230 358708 570236 358720
rect 570288 358708 570294 358760
rect 569954 358612 569960 358624
rect 569880 358584 569960 358612
rect 569954 358572 569960 358584
rect 570012 358572 570018 358624
rect 1394 358368 1400 358420
rect 1452 358408 1458 358420
rect 1762 358408 1768 358420
rect 1452 358380 1768 358408
rect 1452 358368 1458 358380
rect 1762 358368 1768 358380
rect 1820 358368 1826 358420
rect 1765 358275 1823 358281
rect 1765 358241 1777 358275
rect 1811 358272 1823 358275
rect 1854 358272 1860 358284
rect 1811 358244 1860 358272
rect 1811 358241 1823 358244
rect 1765 358235 1823 358241
rect 1854 358232 1860 358244
rect 1912 358232 1918 358284
rect 569954 358232 569960 358284
rect 570012 358272 570018 358284
rect 570049 358275 570107 358281
rect 570049 358272 570061 358275
rect 570012 358244 570061 358272
rect 570012 358232 570018 358244
rect 570049 358241 570061 358244
rect 570095 358241 570107 358275
rect 570049 358235 570107 358241
rect 1854 358136 1860 358148
rect 1815 358108 1860 358136
rect 1854 358096 1860 358108
rect 1912 358096 1918 358148
rect 569957 358139 570015 358145
rect 569957 358136 569969 358139
rect 569880 358108 569969 358136
rect 1397 358071 1455 358077
rect 1397 358037 1409 358071
rect 1443 358068 1455 358071
rect 1762 358068 1768 358080
rect 1443 358040 1768 358068
rect 1443 358037 1455 358040
rect 1397 358031 1455 358037
rect 1762 358028 1768 358040
rect 1820 358028 1826 358080
rect 569880 357864 569908 358108
rect 569957 358105 569969 358108
rect 570003 358105 570015 358139
rect 569957 358099 570015 358105
rect 570046 358096 570052 358148
rect 570104 358096 570110 358148
rect 570138 358096 570144 358148
rect 570196 358096 570202 358148
rect 570064 357944 570092 358096
rect 570156 357944 570184 358096
rect 570230 358028 570236 358080
rect 570288 358068 570294 358080
rect 570325 358071 570383 358077
rect 570325 358068 570337 358071
rect 570288 358040 570337 358068
rect 570288 358028 570294 358040
rect 570325 358037 570337 358040
rect 570371 358037 570383 358071
rect 570325 358031 570383 358037
rect 570046 357892 570052 357944
rect 570104 357892 570110 357944
rect 570138 357892 570144 357944
rect 570196 357892 570202 357944
rect 569954 357864 569960 357876
rect 569880 357836 569960 357864
rect 569954 357824 569960 357836
rect 570012 357824 570018 357876
rect 569957 357663 570015 357669
rect 569957 357629 569969 357663
rect 570003 357660 570015 357663
rect 570233 357663 570291 357669
rect 570233 357660 570245 357663
rect 570003 357632 570245 357660
rect 570003 357629 570015 357632
rect 569957 357623 570015 357629
rect 570233 357629 570245 357632
rect 570279 357629 570291 357663
rect 570233 357623 570291 357629
rect 569954 353948 569960 354000
rect 570012 353988 570018 354000
rect 570012 353960 570057 353988
rect 570012 353948 570018 353960
rect 569954 353744 569960 353796
rect 570012 353744 570018 353796
rect 569972 353716 570000 353744
rect 570509 353719 570567 353725
rect 570509 353716 570521 353719
rect 569972 353688 570521 353716
rect 570509 353685 570521 353688
rect 570555 353685 570567 353719
rect 570509 353679 570567 353685
rect 569954 353608 569960 353660
rect 570012 353648 570018 353660
rect 570012 353620 570057 353648
rect 570012 353608 570018 353620
rect 570322 353308 570328 353320
rect 569880 353280 570328 353308
rect 569880 353252 569908 353280
rect 570322 353268 570328 353280
rect 570380 353268 570386 353320
rect 1857 353243 1915 353249
rect 1857 353209 1869 353243
rect 1903 353240 1915 353243
rect 1946 353240 1952 353252
rect 1903 353212 1952 353240
rect 1903 353209 1915 353212
rect 1857 353203 1915 353209
rect 1946 353200 1952 353212
rect 2004 353200 2010 353252
rect 569862 353200 569868 353252
rect 569920 353200 569926 353252
rect 1762 353064 1768 353116
rect 1820 353104 1826 353116
rect 1946 353104 1952 353116
rect 1820 353076 1952 353104
rect 1820 353064 1826 353076
rect 1946 353064 1952 353076
rect 2004 353064 2010 353116
rect 1394 352928 1400 352980
rect 1452 352968 1458 352980
rect 1762 352968 1768 352980
rect 1452 352940 1768 352968
rect 1452 352928 1458 352940
rect 1762 352928 1768 352940
rect 1820 352928 1826 352980
rect 1857 352971 1915 352977
rect 1857 352937 1869 352971
rect 1903 352968 1915 352971
rect 1946 352968 1952 352980
rect 1903 352940 1952 352968
rect 1903 352937 1915 352940
rect 1857 352931 1915 352937
rect 1946 352928 1952 352940
rect 2004 352928 2010 352980
rect 569957 352631 570015 352637
rect 569957 352597 569969 352631
rect 570003 352628 570015 352631
rect 570046 352628 570052 352640
rect 570003 352600 570052 352628
rect 570003 352597 570015 352600
rect 569957 352591 570015 352597
rect 570046 352588 570052 352600
rect 570104 352588 570110 352640
rect 570049 352495 570107 352501
rect 570049 352461 570061 352495
rect 570095 352492 570107 352495
rect 570233 352495 570291 352501
rect 570233 352492 570245 352495
rect 570095 352464 570245 352492
rect 570095 352461 570107 352464
rect 570049 352455 570107 352461
rect 570233 352461 570245 352464
rect 570279 352461 570291 352495
rect 570233 352455 570291 352461
rect 569954 352316 569960 352368
rect 570012 352356 570018 352368
rect 570417 352359 570475 352365
rect 570417 352356 570429 352359
rect 570012 352328 570429 352356
rect 570012 352316 570018 352328
rect 570417 352325 570429 352328
rect 570463 352325 570475 352359
rect 570417 352319 570475 352325
rect 569954 348956 569960 348968
rect 569915 348928 569960 348956
rect 569954 348916 569960 348928
rect 570012 348916 570018 348968
rect 569954 347964 569960 348016
rect 570012 348004 570018 348016
rect 570233 348007 570291 348013
rect 570233 348004 570245 348007
rect 570012 347976 570245 348004
rect 570012 347964 570018 347976
rect 570233 347973 570245 347976
rect 570279 347973 570291 348007
rect 570233 347967 570291 347973
rect 569954 347692 569960 347744
rect 570012 347732 570018 347744
rect 570141 347735 570199 347741
rect 570141 347732 570153 347735
rect 570012 347704 570153 347732
rect 570012 347692 570018 347704
rect 570141 347701 570153 347704
rect 570187 347701 570199 347735
rect 570141 347695 570199 347701
rect 1673 345763 1731 345769
rect 1673 345729 1685 345763
rect 1719 345760 1731 345763
rect 1946 345760 1952 345772
rect 1719 345732 1952 345760
rect 1719 345729 1731 345732
rect 1673 345723 1731 345729
rect 1946 345720 1952 345732
rect 2004 345720 2010 345772
rect 1765 345695 1823 345701
rect 1765 345661 1777 345695
rect 1811 345692 1823 345695
rect 1854 345692 1860 345704
rect 1811 345664 1860 345692
rect 1811 345661 1823 345664
rect 1765 345655 1823 345661
rect 1854 345652 1860 345664
rect 1912 345652 1918 345704
rect 574922 345040 574928 345092
rect 574980 345080 574986 345092
rect 580166 345080 580172 345092
rect 574980 345052 580172 345080
rect 574980 345040 574986 345052
rect 580166 345040 580172 345052
rect 580224 345040 580230 345092
rect 569954 344876 569960 344888
rect 569915 344848 569960 344876
rect 569954 344836 569960 344848
rect 570012 344836 570018 344888
rect 569954 342184 569960 342236
rect 570012 342224 570018 342236
rect 570012 342196 570057 342224
rect 570012 342184 570018 342196
rect 1857 340867 1915 340873
rect 1857 340833 1869 340867
rect 1903 340864 1915 340867
rect 1946 340864 1952 340876
rect 1903 340836 1952 340864
rect 1903 340833 1915 340836
rect 1857 340827 1915 340833
rect 1946 340824 1952 340836
rect 2004 340824 2010 340876
rect 1765 340731 1823 340737
rect 1765 340697 1777 340731
rect 1811 340728 1823 340731
rect 1946 340728 1952 340740
rect 1811 340700 1952 340728
rect 1811 340697 1823 340700
rect 1765 340691 1823 340697
rect 1946 340688 1952 340700
rect 2004 340688 2010 340740
rect 1946 340252 1952 340264
rect 1907 340224 1952 340252
rect 1946 340212 1952 340224
rect 2004 340212 2010 340264
rect 1394 340144 1400 340196
rect 1452 340184 1458 340196
rect 1762 340184 1768 340196
rect 1452 340156 1768 340184
rect 1452 340144 1458 340156
rect 1762 340144 1768 340156
rect 1820 340144 1826 340196
rect 1946 338076 1952 338088
rect 1907 338048 1952 338076
rect 1946 338036 1952 338048
rect 2004 338036 2010 338088
rect 1489 336039 1547 336045
rect 1489 336005 1501 336039
rect 1535 336036 1547 336039
rect 1857 336039 1915 336045
rect 1857 336036 1869 336039
rect 1535 336008 1869 336036
rect 1535 336005 1547 336008
rect 1489 335999 1547 336005
rect 1857 336005 1869 336008
rect 1903 336005 1915 336039
rect 1857 335999 1915 336005
rect 1397 334203 1455 334209
rect 1397 334169 1409 334203
rect 1443 334200 1455 334203
rect 1946 334200 1952 334212
rect 1443 334172 1952 334200
rect 1443 334169 1455 334172
rect 1397 334163 1455 334169
rect 1946 334160 1952 334172
rect 2004 334160 2010 334212
rect 1765 334067 1823 334073
rect 1765 334033 1777 334067
rect 1811 334064 1823 334067
rect 1946 334064 1952 334076
rect 1811 334036 1952 334064
rect 1811 334033 1823 334036
rect 1765 334027 1823 334033
rect 1946 334024 1952 334036
rect 2004 334024 2010 334076
rect 1302 333684 1308 333736
rect 1360 333724 1366 333736
rect 1946 333724 1952 333736
rect 1360 333696 1952 333724
rect 1360 333684 1366 333696
rect 1946 333684 1952 333696
rect 2004 333684 2010 333736
rect 1397 333455 1455 333461
rect 1397 333421 1409 333455
rect 1443 333452 1455 333455
rect 1946 333452 1952 333464
rect 1443 333424 1952 333452
rect 1443 333421 1455 333424
rect 1397 333415 1455 333421
rect 1946 333412 1952 333424
rect 2004 333412 2010 333464
rect 1765 332027 1823 332033
rect 1765 331993 1777 332027
rect 1811 332024 1823 332027
rect 1811 331996 1992 332024
rect 1811 331993 1823 331996
rect 1765 331987 1823 331993
rect 1489 331891 1547 331897
rect 1489 331857 1501 331891
rect 1535 331888 1547 331891
rect 1765 331891 1823 331897
rect 1765 331888 1777 331891
rect 1535 331860 1777 331888
rect 1535 331857 1547 331860
rect 1489 331851 1547 331857
rect 1765 331857 1777 331860
rect 1811 331857 1823 331891
rect 1765 331851 1823 331857
rect 1964 331832 1992 331996
rect 1946 331780 1952 331832
rect 2004 331780 2010 331832
rect 1394 331508 1400 331560
rect 1452 331548 1458 331560
rect 1762 331548 1768 331560
rect 1452 331520 1768 331548
rect 1452 331508 1458 331520
rect 1762 331508 1768 331520
rect 1820 331508 1826 331560
rect 569954 331276 569960 331288
rect 569915 331248 569960 331276
rect 569954 331236 569960 331248
rect 570012 331236 570018 331288
rect 569954 331072 569960 331084
rect 569915 331044 569960 331072
rect 569954 331032 569960 331044
rect 570012 331032 570018 331084
rect 569954 330488 569960 330540
rect 570012 330528 570018 330540
rect 570141 330531 570199 330537
rect 570141 330528 570153 330531
rect 570012 330500 570153 330528
rect 570012 330488 570018 330500
rect 570141 330497 570153 330500
rect 570187 330497 570199 330531
rect 570141 330491 570199 330497
rect 1673 329783 1731 329789
rect 1673 329749 1685 329783
rect 1719 329780 1731 329783
rect 1946 329780 1952 329792
rect 1719 329752 1952 329780
rect 1719 329749 1731 329752
rect 1673 329743 1731 329749
rect 1946 329740 1952 329752
rect 2004 329740 2010 329792
rect 569954 329672 569960 329724
rect 570012 329712 570018 329724
rect 570049 329715 570107 329721
rect 570049 329712 570061 329715
rect 570012 329684 570061 329712
rect 570012 329672 570018 329684
rect 570049 329681 570061 329684
rect 570095 329681 570107 329715
rect 570049 329675 570107 329681
rect 569865 329579 569923 329585
rect 569865 329545 569877 329579
rect 569911 329576 569923 329579
rect 569954 329576 569960 329588
rect 569911 329548 569960 329576
rect 569911 329545 569923 329548
rect 569865 329539 569923 329545
rect 569954 329536 569960 329548
rect 570012 329536 570018 329588
rect 569954 329400 569960 329452
rect 570012 329440 570018 329452
rect 570233 329443 570291 329449
rect 570233 329440 570245 329443
rect 570012 329412 570245 329440
rect 570012 329400 570018 329412
rect 570233 329409 570245 329412
rect 570279 329409 570291 329443
rect 570233 329403 570291 329409
rect 569954 329264 569960 329316
rect 570012 329304 570018 329316
rect 570325 329307 570383 329313
rect 570325 329304 570337 329307
rect 570012 329276 570337 329304
rect 570012 329264 570018 329276
rect 570325 329273 570337 329276
rect 570371 329273 570383 329307
rect 570325 329267 570383 329273
rect 1946 329168 1952 329180
rect 1907 329140 1952 329168
rect 1946 329128 1952 329140
rect 2004 329128 2010 329180
rect 569954 327808 569960 327820
rect 569880 327780 569960 327808
rect 569880 327196 569908 327780
rect 569954 327768 569960 327780
rect 570012 327768 570018 327820
rect 569954 327632 569960 327684
rect 570012 327672 570018 327684
rect 572714 327672 572720 327684
rect 570012 327644 572720 327672
rect 570012 327632 570018 327644
rect 572714 327632 572720 327644
rect 572772 327632 572778 327684
rect 569954 327196 569960 327208
rect 569880 327168 569960 327196
rect 569954 327156 569960 327168
rect 570012 327156 570018 327208
rect 569954 327020 569960 327072
rect 570012 327060 570018 327072
rect 570325 327063 570383 327069
rect 570325 327060 570337 327063
rect 570012 327032 570337 327060
rect 570012 327020 570018 327032
rect 570325 327029 570337 327032
rect 570371 327029 570383 327063
rect 570325 327023 570383 327029
rect 1489 326519 1547 326525
rect 1489 326485 1501 326519
rect 1535 326516 1547 326519
rect 1857 326519 1915 326525
rect 1857 326516 1869 326519
rect 1535 326488 1869 326516
rect 1535 326485 1547 326488
rect 1489 326479 1547 326485
rect 1857 326485 1869 326488
rect 1903 326485 1915 326519
rect 1857 326479 1915 326485
rect 1581 326383 1639 326389
rect 1581 326349 1593 326383
rect 1627 326380 1639 326383
rect 1857 326383 1915 326389
rect 1857 326380 1869 326383
rect 1627 326352 1869 326380
rect 1627 326349 1639 326352
rect 1581 326343 1639 326349
rect 1857 326349 1869 326352
rect 1903 326349 1915 326383
rect 1857 326343 1915 326349
rect 569954 325660 569960 325712
rect 570012 325700 570018 325712
rect 570233 325703 570291 325709
rect 570233 325700 570245 325703
rect 570012 325672 570245 325700
rect 570012 325660 570018 325672
rect 570233 325669 570245 325672
rect 570279 325669 570291 325703
rect 570233 325663 570291 325669
rect 570138 325524 570144 325576
rect 570196 325564 570202 325576
rect 570233 325567 570291 325573
rect 570233 325564 570245 325567
rect 570196 325536 570245 325564
rect 570196 325524 570202 325536
rect 570233 325533 570245 325536
rect 570279 325533 570291 325567
rect 570233 325527 570291 325533
rect 570046 325020 570052 325032
rect 570007 324992 570052 325020
rect 570046 324980 570052 324992
rect 570104 324980 570110 325032
rect 569957 321147 570015 321153
rect 569957 321144 569969 321147
rect 569880 321116 569969 321144
rect 569880 320736 569908 321116
rect 569957 321113 569969 321116
rect 570003 321113 570015 321147
rect 569957 321107 570015 321113
rect 570141 321147 570199 321153
rect 570141 321113 570153 321147
rect 570187 321144 570199 321147
rect 570325 321147 570383 321153
rect 570325 321144 570337 321147
rect 570187 321116 570337 321144
rect 570187 321113 570199 321116
rect 570141 321107 570199 321113
rect 570325 321113 570337 321116
rect 570371 321113 570383 321147
rect 570325 321107 570383 321113
rect 569954 320968 569960 321020
rect 570012 320968 570018 321020
rect 570049 321011 570107 321017
rect 570049 320977 570061 321011
rect 570095 321008 570107 321011
rect 570138 321008 570144 321020
rect 570095 320980 570144 321008
rect 570095 320977 570107 320980
rect 570049 320971 570107 320977
rect 570138 320968 570144 320980
rect 570196 320968 570202 321020
rect 569972 320940 570000 320968
rect 569972 320912 570276 320940
rect 569954 320832 569960 320884
rect 570012 320872 570018 320884
rect 570012 320844 570057 320872
rect 570012 320832 570018 320844
rect 569957 320739 570015 320745
rect 569957 320736 569969 320739
rect 569880 320708 569969 320736
rect 569957 320705 569969 320708
rect 570003 320705 570015 320739
rect 569957 320699 570015 320705
rect 570046 320696 570052 320748
rect 570104 320736 570110 320748
rect 570248 320745 570276 320912
rect 570141 320739 570199 320745
rect 570141 320736 570153 320739
rect 570104 320708 570153 320736
rect 570104 320696 570110 320708
rect 570141 320705 570153 320708
rect 570187 320705 570199 320739
rect 570141 320699 570199 320705
rect 570233 320739 570291 320745
rect 570233 320705 570245 320739
rect 570279 320705 570291 320739
rect 570233 320699 570291 320705
rect 1946 319172 1952 319184
rect 1907 319144 1952 319172
rect 1946 319132 1952 319144
rect 2004 319132 2010 319184
rect 1581 318971 1639 318977
rect 1581 318937 1593 318971
rect 1627 318968 1639 318971
rect 1946 318968 1952 318980
rect 1627 318940 1952 318968
rect 1627 318937 1639 318940
rect 1581 318931 1639 318937
rect 1946 318928 1952 318940
rect 2004 318928 2010 318980
rect 569954 317948 569960 317960
rect 569915 317920 569960 317948
rect 569954 317908 569960 317920
rect 570012 317908 570018 317960
rect 569957 315979 570015 315985
rect 569957 315945 569969 315979
rect 570003 315945 570015 315979
rect 569957 315939 570015 315945
rect 569972 315849 570000 315939
rect 569957 315843 570015 315849
rect 569957 315809 569969 315843
rect 570003 315809 570015 315843
rect 569957 315803 570015 315809
rect 570046 315800 570052 315852
rect 570104 315840 570110 315852
rect 570322 315840 570328 315852
rect 570104 315812 570328 315840
rect 570104 315800 570110 315812
rect 570322 315800 570328 315812
rect 570380 315800 570386 315852
rect 569954 315596 569960 315648
rect 570012 315636 570018 315648
rect 570012 315608 570057 315636
rect 570012 315596 570018 315608
rect 570230 315596 570236 315648
rect 570288 315596 570294 315648
rect 570046 315528 570052 315580
rect 570104 315568 570110 315580
rect 570248 315568 570276 315596
rect 570104 315540 570276 315568
rect 570104 315528 570110 315540
rect 570230 315500 570236 315512
rect 570191 315472 570236 315500
rect 570230 315460 570236 315472
rect 570288 315460 570294 315512
rect 1305 315163 1363 315169
rect 1305 315129 1317 315163
rect 1351 315160 1363 315163
rect 1946 315160 1952 315172
rect 1351 315132 1952 315160
rect 1351 315129 1363 315132
rect 1305 315123 1363 315129
rect 1946 315120 1952 315132
rect 2004 315120 2010 315172
rect 1946 315024 1952 315036
rect 1907 314996 1952 315024
rect 1946 314984 1952 314996
rect 2004 314984 2010 315036
rect 570325 314755 570383 314761
rect 570325 314721 570337 314755
rect 570371 314752 570383 314755
rect 570509 314755 570567 314761
rect 570509 314752 570521 314755
rect 570371 314724 570521 314752
rect 570371 314721 570383 314724
rect 570325 314715 570383 314721
rect 570509 314721 570521 314724
rect 570555 314721 570567 314755
rect 570509 314715 570567 314721
rect 1673 313939 1731 313945
rect 1673 313905 1685 313939
rect 1719 313936 1731 313939
rect 1857 313939 1915 313945
rect 1857 313936 1869 313939
rect 1719 313908 1869 313936
rect 1719 313905 1731 313908
rect 1673 313899 1731 313905
rect 1857 313905 1869 313908
rect 1903 313905 1915 313939
rect 1857 313899 1915 313905
rect 1489 312715 1547 312721
rect 1489 312681 1501 312715
rect 1535 312712 1547 312715
rect 1949 312715 2007 312721
rect 1949 312712 1961 312715
rect 1535 312684 1961 312712
rect 1535 312681 1547 312684
rect 1489 312675 1547 312681
rect 1949 312681 1961 312684
rect 1995 312681 2007 312715
rect 1949 312675 2007 312681
rect 1857 312579 1915 312585
rect 1857 312545 1869 312579
rect 1903 312576 1915 312579
rect 1946 312576 1952 312588
rect 1903 312548 1952 312576
rect 1903 312545 1915 312548
rect 1857 312539 1915 312545
rect 1946 312536 1952 312548
rect 2004 312536 2010 312588
rect 1489 312443 1547 312449
rect 1489 312409 1501 312443
rect 1535 312440 1547 312443
rect 1946 312440 1952 312452
rect 1535 312412 1952 312440
rect 1535 312409 1547 312412
rect 1489 312403 1547 312409
rect 1946 312400 1952 312412
rect 2004 312400 2010 312452
rect 1397 312307 1455 312313
rect 1397 312273 1409 312307
rect 1443 312304 1455 312307
rect 1946 312304 1952 312316
rect 1443 312276 1952 312304
rect 1443 312273 1455 312276
rect 1397 312267 1455 312273
rect 1946 312264 1952 312276
rect 2004 312264 2010 312316
rect 1213 312171 1271 312177
rect 1213 312137 1225 312171
rect 1259 312168 1271 312171
rect 1397 312171 1455 312177
rect 1397 312168 1409 312171
rect 1259 312140 1409 312168
rect 1259 312137 1271 312140
rect 1213 312131 1271 312137
rect 1397 312137 1409 312140
rect 1443 312137 1455 312171
rect 1397 312131 1455 312137
rect 1946 312128 1952 312180
rect 2004 312128 2010 312180
rect 1964 312100 1992 312128
rect 1412 312072 1992 312100
rect 1412 312041 1440 312072
rect 1397 312035 1455 312041
rect 1397 312001 1409 312035
rect 1443 312001 1455 312035
rect 1397 311995 1455 312001
rect 1765 312035 1823 312041
rect 1765 312001 1777 312035
rect 1811 312032 1823 312035
rect 1946 312032 1952 312044
rect 1811 312004 1952 312032
rect 1811 312001 1823 312004
rect 1765 311995 1823 312001
rect 1946 311992 1952 312004
rect 2004 311992 2010 312044
rect 1305 311831 1363 311837
rect 1305 311797 1317 311831
rect 1351 311828 1363 311831
rect 1946 311828 1952 311840
rect 1351 311800 1952 311828
rect 1351 311797 1363 311800
rect 1305 311791 1363 311797
rect 1946 311788 1952 311800
rect 2004 311788 2010 311840
rect 1581 311695 1639 311701
rect 1581 311661 1593 311695
rect 1627 311692 1639 311695
rect 1946 311692 1952 311704
rect 1627 311664 1952 311692
rect 1627 311661 1639 311664
rect 1581 311655 1639 311661
rect 1946 311652 1952 311664
rect 2004 311652 2010 311704
rect 1673 311559 1731 311565
rect 1673 311525 1685 311559
rect 1719 311556 1731 311559
rect 1946 311556 1952 311568
rect 1719 311528 1952 311556
rect 1719 311525 1731 311528
rect 1673 311519 1731 311525
rect 1946 311516 1952 311528
rect 2004 311516 2010 311568
rect 1946 309856 1952 309868
rect 1907 309828 1952 309856
rect 1946 309816 1952 309828
rect 2004 309816 2010 309868
rect 1857 309655 1915 309661
rect 1857 309621 1869 309655
rect 1903 309652 1915 309655
rect 1946 309652 1952 309664
rect 1903 309624 1952 309652
rect 1903 309621 1915 309624
rect 1857 309615 1915 309621
rect 1946 309612 1952 309624
rect 2004 309612 2010 309664
rect 570509 309247 570567 309253
rect 570509 309244 570521 309247
rect 570248 309216 570521 309244
rect 570248 309185 570276 309216
rect 570509 309213 570521 309216
rect 570555 309213 570567 309247
rect 570509 309207 570567 309213
rect 570233 309179 570291 309185
rect 570233 309145 570245 309179
rect 570279 309145 570291 309179
rect 570233 309139 570291 309145
rect 569954 309068 569960 309120
rect 570012 309108 570018 309120
rect 570049 309111 570107 309117
rect 570049 309108 570061 309111
rect 570012 309080 570061 309108
rect 570012 309068 570018 309080
rect 570049 309077 570061 309080
rect 570095 309077 570107 309111
rect 570049 309071 570107 309077
rect 569954 306960 569960 307012
rect 570012 307000 570018 307012
rect 570417 307003 570475 307009
rect 570417 307000 570429 307003
rect 570012 306972 570429 307000
rect 570012 306960 570018 306972
rect 570417 306969 570429 306972
rect 570463 306969 570475 307003
rect 570417 306963 570475 306969
rect 1946 306660 1952 306672
rect 1907 306632 1952 306660
rect 1946 306620 1952 306632
rect 2004 306620 2010 306672
rect 569954 306184 569960 306196
rect 569915 306156 569960 306184
rect 569954 306144 569960 306156
rect 570012 306144 570018 306196
rect 1673 305643 1731 305649
rect 1673 305609 1685 305643
rect 1719 305640 1731 305643
rect 1946 305640 1952 305652
rect 1719 305612 1952 305640
rect 1719 305609 1731 305612
rect 1673 305603 1731 305609
rect 1946 305600 1952 305612
rect 2004 305600 2010 305652
rect 1765 305507 1823 305513
rect 1765 305473 1777 305507
rect 1811 305504 1823 305507
rect 1946 305504 1952 305516
rect 1811 305476 1952 305504
rect 1811 305473 1823 305476
rect 1765 305467 1823 305473
rect 1946 305464 1952 305476
rect 2004 305464 2010 305516
rect 1857 305371 1915 305377
rect 1857 305337 1869 305371
rect 1903 305368 1915 305371
rect 1946 305368 1952 305380
rect 1903 305340 1952 305368
rect 1903 305337 1915 305340
rect 1857 305331 1915 305337
rect 1946 305328 1952 305340
rect 2004 305328 2010 305380
rect 570141 305031 570199 305037
rect 570141 305028 570153 305031
rect 569880 305000 570153 305028
rect 569880 304960 569908 305000
rect 570141 304997 570153 305000
rect 570187 304997 570199 305031
rect 570141 304991 570199 304997
rect 570509 304963 570567 304969
rect 570509 304960 570521 304963
rect 569880 304932 570521 304960
rect 570509 304929 570521 304932
rect 570555 304929 570567 304963
rect 570509 304923 570567 304929
rect 1305 304555 1363 304561
rect 1305 304521 1317 304555
rect 1351 304552 1363 304555
rect 1946 304552 1952 304564
rect 1351 304524 1952 304552
rect 1351 304521 1363 304524
rect 1305 304515 1363 304521
rect 1946 304512 1952 304524
rect 2004 304512 2010 304564
rect 1489 304419 1547 304425
rect 1489 304385 1501 304419
rect 1535 304416 1547 304419
rect 1946 304416 1952 304428
rect 1535 304388 1952 304416
rect 1535 304385 1547 304388
rect 1489 304379 1547 304385
rect 1946 304376 1952 304388
rect 2004 304376 2010 304428
rect 569957 304283 570015 304289
rect 569957 304249 569969 304283
rect 570003 304280 570015 304283
rect 570046 304280 570052 304292
rect 570003 304252 570052 304280
rect 570003 304249 570015 304252
rect 569957 304243 570015 304249
rect 570046 304240 570052 304252
rect 570104 304240 570110 304292
rect 1213 304147 1271 304153
rect 1213 304113 1225 304147
rect 1259 304144 1271 304147
rect 1946 304144 1952 304156
rect 1259 304116 1952 304144
rect 1259 304113 1271 304116
rect 1213 304107 1271 304113
rect 1946 304104 1952 304116
rect 2004 304104 2010 304156
rect 1397 304011 1455 304017
rect 1397 303977 1409 304011
rect 1443 304008 1455 304011
rect 1946 304008 1952 304020
rect 1443 303980 1952 304008
rect 1443 303977 1455 303980
rect 1397 303971 1455 303977
rect 1946 303968 1952 303980
rect 2004 303968 2010 304020
rect 570230 303832 570236 303884
rect 570288 303872 570294 303884
rect 570325 303875 570383 303881
rect 570325 303872 570337 303875
rect 570288 303844 570337 303872
rect 570288 303832 570294 303844
rect 570325 303841 570337 303844
rect 570371 303841 570383 303875
rect 570325 303835 570383 303841
rect 1213 303399 1271 303405
rect 1213 303365 1225 303399
rect 1259 303396 1271 303399
rect 1946 303396 1952 303408
rect 1259 303368 1952 303396
rect 1259 303365 1271 303368
rect 1213 303359 1271 303365
rect 1946 303356 1952 303368
rect 2004 303356 2010 303408
rect 1765 303263 1823 303269
rect 1765 303229 1777 303263
rect 1811 303260 1823 303263
rect 1946 303260 1952 303272
rect 1811 303232 1952 303260
rect 1811 303229 1823 303232
rect 1765 303223 1823 303229
rect 1946 303220 1952 303232
rect 2004 303220 2010 303272
rect 570049 302923 570107 302929
rect 570049 302889 570061 302923
rect 570095 302920 570107 302923
rect 570233 302923 570291 302929
rect 570233 302920 570245 302923
rect 570095 302892 570245 302920
rect 570095 302889 570107 302892
rect 570049 302883 570107 302889
rect 570233 302889 570245 302892
rect 570279 302889 570291 302923
rect 570233 302883 570291 302889
rect 569954 302744 569960 302796
rect 570012 302784 570018 302796
rect 570233 302787 570291 302793
rect 570233 302784 570245 302787
rect 570012 302756 570245 302784
rect 570012 302744 570018 302756
rect 570233 302753 570245 302756
rect 570279 302753 570291 302787
rect 570233 302747 570291 302753
rect 569957 301903 570015 301909
rect 569957 301869 569969 301903
rect 570003 301900 570015 301903
rect 570417 301903 570475 301909
rect 570417 301900 570429 301903
rect 570003 301872 570429 301900
rect 570003 301869 570015 301872
rect 569957 301863 570015 301869
rect 570417 301869 570429 301872
rect 570463 301869 570475 301903
rect 570417 301863 570475 301869
rect 3326 301792 3332 301844
rect 3384 301832 3390 301844
rect 3694 301832 3700 301844
rect 3384 301804 3700 301832
rect 3384 301792 3390 301804
rect 3694 301792 3700 301804
rect 3752 301792 3758 301844
rect 1673 301495 1731 301501
rect 1673 301461 1685 301495
rect 1719 301492 1731 301495
rect 1946 301492 1952 301504
rect 1719 301464 1952 301492
rect 1719 301461 1731 301464
rect 1673 301455 1731 301461
rect 1946 301452 1952 301464
rect 2004 301452 2010 301504
rect 569954 301112 569960 301164
rect 570012 301152 570018 301164
rect 570417 301155 570475 301161
rect 570417 301152 570429 301155
rect 570012 301124 570429 301152
rect 570012 301112 570018 301124
rect 570417 301121 570429 301124
rect 570463 301121 570475 301155
rect 570417 301115 570475 301121
rect 569954 300840 569960 300892
rect 570012 300880 570018 300892
rect 570012 300852 570057 300880
rect 570012 300840 570018 300852
rect 570325 300407 570383 300413
rect 570325 300373 570337 300407
rect 570371 300404 570383 300407
rect 570414 300404 570420 300416
rect 570371 300376 570420 300404
rect 570371 300373 570383 300376
rect 570325 300367 570383 300373
rect 570414 300364 570420 300376
rect 570472 300364 570478 300416
rect 570049 300271 570107 300277
rect 570049 300237 570061 300271
rect 570095 300268 570107 300271
rect 570322 300268 570328 300280
rect 570095 300240 570328 300268
rect 570095 300237 570107 300240
rect 570049 300231 570107 300237
rect 570322 300228 570328 300240
rect 570380 300228 570386 300280
rect 570049 300135 570107 300141
rect 570049 300101 570061 300135
rect 570095 300132 570107 300135
rect 570138 300132 570144 300144
rect 570095 300104 570144 300132
rect 570095 300101 570107 300104
rect 570049 300095 570107 300101
rect 570138 300092 570144 300104
rect 570196 300092 570202 300144
rect 569954 300064 569960 300076
rect 569915 300036 569960 300064
rect 569954 300024 569960 300036
rect 570012 300024 570018 300076
rect 569954 298568 569960 298580
rect 569915 298540 569960 298568
rect 569954 298528 569960 298540
rect 570012 298528 570018 298580
rect 569954 298392 569960 298444
rect 570012 298432 570018 298444
rect 570233 298435 570291 298441
rect 570233 298432 570245 298435
rect 570012 298404 570245 298432
rect 570012 298392 570018 298404
rect 570233 298401 570245 298404
rect 570279 298401 570291 298435
rect 570233 298395 570291 298401
rect 575014 298120 575020 298172
rect 575072 298160 575078 298172
rect 580166 298160 580172 298172
rect 575072 298132 580172 298160
rect 575072 298120 575078 298132
rect 580166 298120 580172 298132
rect 580224 298120 580230 298172
rect 1121 298095 1179 298101
rect 1121 298061 1133 298095
rect 1167 298092 1179 298095
rect 1305 298095 1363 298101
rect 1305 298092 1317 298095
rect 1167 298064 1317 298092
rect 1167 298061 1179 298064
rect 1121 298055 1179 298061
rect 1305 298061 1317 298064
rect 1351 298061 1363 298095
rect 1305 298055 1363 298061
rect 570049 296599 570107 296605
rect 570049 296565 570061 296599
rect 570095 296596 570107 296599
rect 570325 296599 570383 296605
rect 570325 296596 570337 296599
rect 570095 296568 570337 296596
rect 570095 296565 570107 296568
rect 570049 296559 570107 296565
rect 570325 296565 570337 296568
rect 570371 296565 570383 296599
rect 570325 296559 570383 296565
rect 1302 296216 1308 296268
rect 1360 296256 1366 296268
rect 1857 296259 1915 296265
rect 1857 296256 1869 296259
rect 1360 296228 1869 296256
rect 1360 296216 1366 296228
rect 1857 296225 1869 296228
rect 1903 296225 1915 296259
rect 1857 296219 1915 296225
rect 570046 296148 570052 296200
rect 570104 296188 570110 296200
rect 570141 296191 570199 296197
rect 570141 296188 570153 296191
rect 570104 296160 570153 296188
rect 570104 296148 570110 296160
rect 570141 296157 570153 296160
rect 570187 296157 570199 296191
rect 570141 296151 570199 296157
rect 1765 296123 1823 296129
rect 1765 296089 1777 296123
rect 1811 296120 1823 296123
rect 1946 296120 1952 296132
rect 1811 296092 1952 296120
rect 1811 296089 1823 296092
rect 1765 296083 1823 296089
rect 1946 296080 1952 296092
rect 2004 296080 2010 296132
rect 569954 296080 569960 296132
rect 570012 296120 570018 296132
rect 570509 296123 570567 296129
rect 570509 296120 570521 296123
rect 570012 296092 570521 296120
rect 570012 296080 570018 296092
rect 570509 296089 570521 296092
rect 570555 296089 570567 296123
rect 570509 296083 570567 296089
rect 1305 296055 1363 296061
rect 1305 296021 1317 296055
rect 1351 296052 1363 296055
rect 1581 296055 1639 296061
rect 1581 296052 1593 296055
rect 1351 296024 1593 296052
rect 1351 296021 1363 296024
rect 1305 296015 1363 296021
rect 1581 296021 1593 296024
rect 1627 296021 1639 296055
rect 1581 296015 1639 296021
rect 570141 296055 570199 296061
rect 570141 296021 570153 296055
rect 570187 296052 570199 296055
rect 570230 296052 570236 296064
rect 570187 296024 570236 296052
rect 570187 296021 570199 296024
rect 570141 296015 570199 296021
rect 570230 296012 570236 296024
rect 570288 296012 570294 296064
rect 1394 295944 1400 295996
rect 1452 295984 1458 295996
rect 1857 295987 1915 295993
rect 1857 295984 1869 295987
rect 1452 295956 1869 295984
rect 1452 295944 1458 295956
rect 1857 295953 1869 295956
rect 1903 295953 1915 295987
rect 1857 295947 1915 295953
rect 1673 295851 1731 295857
rect 1673 295817 1685 295851
rect 1719 295848 1731 295851
rect 1946 295848 1952 295860
rect 1719 295820 1952 295848
rect 1719 295817 1731 295820
rect 1673 295811 1731 295817
rect 1946 295808 1952 295820
rect 2004 295808 2010 295860
rect 570233 295171 570291 295177
rect 570233 295137 570245 295171
rect 570279 295168 570291 295171
rect 570322 295168 570328 295180
rect 570279 295140 570328 295168
rect 570279 295137 570291 295140
rect 570233 295131 570291 295137
rect 570322 295128 570328 295140
rect 570380 295128 570386 295180
rect 474 294584 480 294636
rect 532 294624 538 294636
rect 1489 294627 1547 294633
rect 1489 294624 1501 294627
rect 532 294596 1501 294624
rect 532 294584 538 294596
rect 1489 294593 1501 294596
rect 1535 294593 1547 294627
rect 1489 294587 1547 294593
rect 1121 294491 1179 294497
rect 1121 294457 1133 294491
rect 1167 294488 1179 294491
rect 1489 294491 1547 294497
rect 1489 294488 1501 294491
rect 1167 294460 1501 294488
rect 1167 294457 1179 294460
rect 1121 294451 1179 294457
rect 1489 294457 1501 294460
rect 1535 294457 1547 294491
rect 1489 294451 1547 294457
rect 1397 293403 1455 293409
rect 1397 293369 1409 293403
rect 1443 293400 1455 293403
rect 1946 293400 1952 293412
rect 1443 293372 1952 293400
rect 1443 293369 1455 293372
rect 1397 293363 1455 293369
rect 1946 293360 1952 293372
rect 2004 293360 2010 293412
rect 1213 293131 1271 293137
rect 1213 293097 1225 293131
rect 1259 293128 1271 293131
rect 1946 293128 1952 293140
rect 1259 293100 1952 293128
rect 1259 293097 1271 293100
rect 1213 293091 1271 293097
rect 1946 293088 1952 293100
rect 2004 293088 2010 293140
rect 569957 292791 570015 292797
rect 569957 292757 569969 292791
rect 570003 292788 570015 292791
rect 570230 292788 570236 292800
rect 570003 292760 570236 292788
rect 570003 292757 570015 292760
rect 569957 292751 570015 292757
rect 570230 292748 570236 292760
rect 570288 292748 570294 292800
rect 569957 292587 570015 292593
rect 569957 292553 569969 292587
rect 570003 292584 570015 292587
rect 570414 292584 570420 292596
rect 570003 292556 570420 292584
rect 570003 292553 570015 292556
rect 569957 292547 570015 292553
rect 570414 292544 570420 292556
rect 570472 292544 570478 292596
rect 569954 292408 569960 292460
rect 570012 292448 570018 292460
rect 570417 292451 570475 292457
rect 570417 292448 570429 292451
rect 570012 292420 570429 292448
rect 570012 292408 570018 292420
rect 570417 292417 570429 292420
rect 570463 292417 570475 292451
rect 570417 292411 570475 292417
rect 1305 292179 1363 292185
rect 1305 292145 1317 292179
rect 1351 292176 1363 292179
rect 1581 292179 1639 292185
rect 1581 292176 1593 292179
rect 1351 292148 1593 292176
rect 1351 292145 1363 292148
rect 1305 292139 1363 292145
rect 1581 292145 1593 292148
rect 1627 292145 1639 292179
rect 1581 292139 1639 292145
rect 570141 291975 570199 291981
rect 570141 291941 570153 291975
rect 570187 291972 570199 291975
rect 570325 291975 570383 291981
rect 570325 291972 570337 291975
rect 570187 291944 570337 291972
rect 570187 291941 570199 291944
rect 570141 291935 570199 291941
rect 570325 291941 570337 291944
rect 570371 291941 570383 291975
rect 570325 291935 570383 291941
rect 570049 289799 570107 289805
rect 570049 289765 570061 289799
rect 570095 289796 570107 289799
rect 570141 289799 570199 289805
rect 570141 289796 570153 289799
rect 570095 289768 570153 289796
rect 570095 289765 570107 289768
rect 570049 289759 570107 289765
rect 570141 289765 570153 289768
rect 570187 289765 570199 289799
rect 570141 289759 570199 289765
rect 569954 289620 569960 289672
rect 570012 289660 570018 289672
rect 570509 289663 570567 289669
rect 570509 289660 570521 289663
rect 570012 289632 570521 289660
rect 570012 289620 570018 289632
rect 570509 289629 570521 289632
rect 570555 289629 570567 289663
rect 570509 289623 570567 289629
rect 569957 288303 570015 288309
rect 569957 288269 569969 288303
rect 570003 288300 570015 288303
rect 570322 288300 570328 288312
rect 570003 288272 570328 288300
rect 570003 288269 570015 288272
rect 569957 288263 570015 288269
rect 570322 288260 570328 288272
rect 570380 288260 570386 288312
rect 570233 288167 570291 288173
rect 570233 288133 570245 288167
rect 570279 288164 570291 288167
rect 570417 288167 570475 288173
rect 570417 288164 570429 288167
rect 570279 288136 570429 288164
rect 570279 288133 570291 288136
rect 570233 288127 570291 288133
rect 570417 288133 570429 288136
rect 570463 288133 570475 288167
rect 570417 288127 570475 288133
rect 1305 287147 1363 287153
rect 1305 287113 1317 287147
rect 1351 287144 1363 287147
rect 1489 287147 1547 287153
rect 1489 287144 1501 287147
rect 1351 287116 1501 287144
rect 1351 287113 1363 287116
rect 1305 287107 1363 287113
rect 1489 287113 1501 287116
rect 1535 287113 1547 287147
rect 1489 287107 1547 287113
rect 14 286968 20 287020
rect 72 287008 78 287020
rect 1581 287011 1639 287017
rect 1581 287008 1593 287011
rect 72 286980 1593 287008
rect 72 286968 78 286980
rect 1581 286977 1593 286980
rect 1627 286977 1639 287011
rect 1581 286971 1639 286977
rect 569957 285651 570015 285657
rect 569957 285617 569969 285651
rect 570003 285648 570015 285651
rect 570233 285651 570291 285657
rect 570233 285648 570245 285651
rect 570003 285620 570245 285648
rect 570003 285617 570015 285620
rect 569957 285611 570015 285617
rect 570233 285617 570245 285620
rect 570279 285617 570291 285651
rect 570233 285611 570291 285617
rect 569957 285515 570015 285521
rect 569957 285481 569969 285515
rect 570003 285512 570015 285515
rect 570230 285512 570236 285524
rect 570003 285484 570236 285512
rect 570003 285481 570015 285484
rect 569957 285475 570015 285481
rect 570230 285472 570236 285484
rect 570288 285472 570294 285524
rect 569954 285336 569960 285388
rect 570012 285376 570018 285388
rect 570141 285379 570199 285385
rect 570141 285376 570153 285379
rect 570012 285348 570153 285376
rect 570012 285336 570018 285348
rect 570141 285345 570153 285348
rect 570187 285345 570199 285379
rect 570141 285339 570199 285345
rect 569954 285172 569960 285184
rect 569915 285144 569960 285172
rect 569954 285132 569960 285144
rect 570012 285132 570018 285184
rect 569954 284928 569960 284980
rect 570012 284968 570018 284980
rect 570325 284971 570383 284977
rect 570325 284968 570337 284971
rect 570012 284940 570337 284968
rect 570012 284928 570018 284940
rect 570325 284937 570337 284940
rect 570371 284937 570383 284971
rect 570325 284931 570383 284937
rect 569954 284792 569960 284844
rect 570012 284832 570018 284844
rect 570601 284835 570659 284841
rect 570601 284832 570613 284835
rect 570012 284804 570613 284832
rect 570012 284792 570018 284804
rect 570601 284801 570613 284804
rect 570647 284801 570659 284835
rect 570601 284795 570659 284801
rect 1397 284767 1455 284773
rect 1397 284733 1409 284767
rect 1443 284764 1455 284767
rect 1946 284764 1952 284776
rect 1443 284736 1952 284764
rect 1443 284733 1455 284736
rect 1397 284727 1455 284733
rect 1946 284724 1952 284736
rect 2004 284724 2010 284776
rect 1305 284631 1363 284637
rect 1305 284597 1317 284631
rect 1351 284628 1363 284631
rect 1946 284628 1952 284640
rect 1351 284600 1952 284628
rect 1351 284597 1363 284600
rect 1305 284591 1363 284597
rect 1946 284588 1952 284600
rect 2004 284588 2010 284640
rect 569954 284588 569960 284640
rect 570012 284628 570018 284640
rect 570506 284628 570512 284640
rect 570012 284600 570512 284628
rect 570012 284588 570018 284600
rect 570506 284588 570512 284600
rect 570564 284588 570570 284640
rect 1489 284359 1547 284365
rect 1489 284325 1501 284359
rect 1535 284356 1547 284359
rect 1946 284356 1952 284368
rect 1535 284328 1952 284356
rect 1535 284325 1547 284328
rect 1489 284319 1547 284325
rect 1946 284316 1952 284328
rect 2004 284316 2010 284368
rect 1394 283948 1400 283960
rect 1355 283920 1400 283948
rect 1394 283908 1400 283920
rect 1452 283908 1458 283960
rect 1857 283951 1915 283957
rect 1857 283917 1869 283951
rect 1903 283948 1915 283951
rect 1946 283948 1952 283960
rect 1903 283920 1952 283948
rect 1903 283917 1915 283920
rect 1857 283911 1915 283917
rect 1946 283908 1952 283920
rect 2004 283908 2010 283960
rect 569954 283840 569960 283892
rect 570012 283880 570018 283892
rect 570012 283852 570092 283880
rect 570012 283840 570018 283852
rect 569954 283744 569960 283756
rect 569915 283716 569960 283744
rect 569954 283704 569960 283716
rect 570012 283704 570018 283756
rect 570064 283676 570092 283852
rect 569880 283648 570092 283676
rect 1397 283475 1455 283481
rect 1397 283441 1409 283475
rect 1443 283472 1455 283475
rect 1857 283475 1915 283481
rect 1857 283472 1869 283475
rect 1443 283444 1869 283472
rect 1443 283441 1455 283444
rect 1397 283435 1455 283441
rect 1857 283441 1869 283444
rect 1903 283441 1915 283475
rect 1857 283435 1915 283441
rect 1765 283407 1823 283413
rect 1765 283373 1777 283407
rect 1811 283404 1823 283407
rect 1946 283404 1952 283416
rect 1811 283376 1952 283404
rect 1811 283373 1823 283376
rect 1765 283367 1823 283373
rect 1946 283364 1952 283376
rect 2004 283364 2010 283416
rect 569880 283336 569908 283648
rect 570049 283611 570107 283617
rect 570049 283577 570061 283611
rect 570095 283608 570107 283611
rect 570233 283611 570291 283617
rect 570233 283608 570245 283611
rect 570095 283580 570245 283608
rect 570095 283577 570107 283580
rect 570049 283571 570107 283577
rect 570233 283577 570245 283580
rect 570279 283577 570291 283611
rect 570233 283571 570291 283577
rect 569954 283500 569960 283552
rect 570012 283540 570018 283552
rect 570509 283543 570567 283549
rect 570509 283540 570521 283543
rect 570012 283512 570521 283540
rect 570012 283500 570018 283512
rect 570509 283509 570521 283512
rect 570555 283509 570567 283543
rect 570509 283503 570567 283509
rect 570046 283432 570052 283484
rect 570104 283472 570110 283484
rect 570233 283475 570291 283481
rect 570233 283472 570245 283475
rect 570104 283444 570245 283472
rect 570104 283432 570110 283444
rect 570233 283441 570245 283444
rect 570279 283441 570291 283475
rect 570233 283435 570291 283441
rect 569954 283364 569960 283416
rect 570012 283404 570018 283416
rect 570325 283407 570383 283413
rect 570325 283404 570337 283407
rect 570012 283376 570337 283404
rect 570012 283364 570018 283376
rect 570325 283373 570337 283376
rect 570371 283373 570383 283407
rect 570325 283367 570383 283373
rect 570046 283336 570052 283348
rect 569880 283308 570052 283336
rect 570046 283296 570052 283308
rect 570104 283296 570110 283348
rect 1581 283271 1639 283277
rect 1581 283237 1593 283271
rect 1627 283268 1639 283271
rect 1946 283268 1952 283280
rect 1627 283240 1952 283268
rect 1627 283237 1639 283240
rect 1581 283231 1639 283237
rect 1946 283228 1952 283240
rect 2004 283228 2010 283280
rect 569954 277924 569960 277976
rect 570012 277964 570018 277976
rect 570322 277964 570328 277976
rect 570012 277936 570328 277964
rect 570012 277924 570018 277936
rect 570322 277924 570328 277936
rect 570380 277924 570386 277976
rect 569954 277516 569960 277568
rect 570012 277556 570018 277568
rect 570138 277556 570144 277568
rect 570012 277528 570144 277556
rect 570012 277516 570018 277528
rect 570138 277516 570144 277528
rect 570196 277516 570202 277568
rect 569954 277244 569960 277296
rect 570012 277284 570018 277296
rect 570509 277287 570567 277293
rect 570509 277284 570521 277287
rect 570012 277256 570521 277284
rect 570012 277244 570018 277256
rect 570509 277253 570521 277256
rect 570555 277253 570567 277287
rect 570509 277247 570567 277253
rect 569954 274456 569960 274508
rect 570012 274496 570018 274508
rect 570693 274499 570751 274505
rect 570693 274496 570705 274499
rect 570012 274468 570705 274496
rect 570012 274456 570018 274468
rect 570693 274465 570705 274468
rect 570739 274465 570751 274499
rect 570693 274459 570751 274465
rect 570141 274363 570199 274369
rect 570141 274329 570153 274363
rect 570187 274360 570199 274363
rect 570325 274363 570383 274369
rect 570325 274360 570337 274363
rect 570187 274332 570337 274360
rect 570187 274329 570199 274332
rect 570141 274323 570199 274329
rect 570325 274329 570337 274332
rect 570371 274329 570383 274363
rect 570325 274323 570383 274329
rect 569954 274224 569960 274236
rect 569880 274196 569960 274224
rect 1673 273955 1731 273961
rect 1673 273921 1685 273955
rect 1719 273952 1731 273955
rect 1946 273952 1952 273964
rect 1719 273924 1952 273952
rect 1719 273921 1731 273924
rect 1673 273915 1731 273921
rect 1946 273912 1952 273924
rect 2004 273912 2010 273964
rect 569880 273748 569908 274196
rect 569954 274184 569960 274196
rect 570012 274184 570018 274236
rect 569957 274023 570015 274029
rect 569957 273989 569969 274023
rect 570003 274020 570015 274023
rect 570003 273992 570092 274020
rect 570003 273989 570015 273992
rect 569957 273983 570015 273989
rect 570064 273893 570092 273992
rect 570049 273887 570107 273893
rect 570049 273853 570061 273887
rect 570095 273853 570107 273887
rect 570049 273847 570107 273853
rect 570046 273748 570052 273760
rect 569880 273720 570052 273748
rect 570046 273708 570052 273720
rect 570104 273708 570110 273760
rect 569954 273068 569960 273080
rect 569915 273040 569960 273068
rect 569954 273028 569960 273040
rect 570012 273028 570018 273080
rect 569954 272892 569960 272944
rect 570012 272932 570018 272944
rect 570693 272935 570751 272941
rect 570693 272932 570705 272935
rect 570012 272904 570705 272932
rect 570012 272892 570018 272904
rect 570693 272901 570705 272904
rect 570739 272901 570751 272935
rect 570693 272895 570751 272901
rect 569954 272756 569960 272808
rect 570012 272796 570018 272808
rect 572714 272796 572720 272808
rect 570012 272768 572720 272796
rect 570012 272756 570018 272768
rect 572714 272756 572720 272768
rect 572772 272756 572778 272808
rect 569954 272552 569960 272604
rect 570012 272592 570018 272604
rect 570414 272592 570420 272604
rect 570012 272564 570420 272592
rect 570012 272552 570018 272564
rect 570414 272552 570420 272564
rect 570472 272552 570478 272604
rect 570601 272527 570659 272533
rect 570601 272524 570613 272527
rect 569880 272496 570613 272524
rect 569880 272400 569908 272496
rect 570601 272493 570613 272496
rect 570647 272493 570659 272527
rect 570601 272487 570659 272493
rect 569862 272348 569868 272400
rect 569920 272348 569926 272400
rect 569954 271572 569960 271584
rect 569915 271544 569960 271572
rect 569954 271532 569960 271544
rect 570012 271532 570018 271584
rect 569954 270988 569960 271040
rect 570012 271028 570018 271040
rect 570509 271031 570567 271037
rect 570509 271028 570521 271031
rect 570012 271000 570521 271028
rect 570012 270988 570018 271000
rect 570509 270997 570521 271000
rect 570555 270997 570567 271031
rect 570509 270991 570567 270997
rect 569954 270852 569960 270904
rect 570012 270892 570018 270904
rect 570138 270892 570144 270904
rect 570012 270864 570144 270892
rect 570012 270852 570018 270864
rect 570138 270852 570144 270864
rect 570196 270852 570202 270904
rect 569954 270580 569960 270632
rect 570012 270620 570018 270632
rect 570322 270620 570328 270632
rect 570012 270592 570328 270620
rect 570012 270580 570018 270592
rect 570322 270580 570328 270592
rect 570380 270580 570386 270632
rect 569954 270444 569960 270496
rect 570012 270484 570018 270496
rect 570141 270487 570199 270493
rect 570141 270484 570153 270487
rect 570012 270456 570153 270484
rect 570012 270444 570018 270456
rect 570141 270453 570153 270456
rect 570187 270453 570199 270487
rect 570141 270447 570199 270453
rect 569954 270308 569960 270360
rect 570012 270348 570018 270360
rect 570233 270351 570291 270357
rect 570233 270348 570245 270351
rect 570012 270320 570245 270348
rect 570012 270308 570018 270320
rect 570233 270317 570245 270320
rect 570279 270317 570291 270351
rect 570233 270311 570291 270317
rect 1673 270215 1731 270221
rect 1673 270181 1685 270215
rect 1719 270212 1731 270215
rect 1946 270212 1952 270224
rect 1719 270184 1952 270212
rect 1719 270181 1731 270184
rect 1673 270175 1731 270181
rect 1946 270172 1952 270184
rect 2004 270172 2010 270224
rect 569954 270172 569960 270224
rect 570012 270212 570018 270224
rect 570230 270212 570236 270224
rect 570012 270184 570236 270212
rect 570012 270172 570018 270184
rect 570230 270172 570236 270184
rect 570288 270172 570294 270224
rect 569954 270036 569960 270088
rect 570012 270076 570018 270088
rect 570325 270079 570383 270085
rect 570325 270076 570337 270079
rect 570012 270048 570337 270076
rect 570012 270036 570018 270048
rect 570325 270045 570337 270048
rect 570371 270045 570383 270079
rect 570325 270039 570383 270045
rect 569954 269900 569960 269952
rect 570012 269940 570018 269952
rect 570417 269943 570475 269949
rect 570417 269940 570429 269943
rect 570012 269912 570429 269940
rect 570012 269900 570018 269912
rect 570417 269909 570429 269912
rect 570463 269909 570475 269943
rect 570417 269903 570475 269909
rect 1765 269807 1823 269813
rect 1765 269773 1777 269807
rect 1811 269804 1823 269807
rect 1946 269804 1952 269816
rect 1811 269776 1952 269804
rect 1811 269773 1823 269776
rect 1765 269767 1823 269773
rect 1946 269764 1952 269776
rect 2004 269764 2010 269816
rect 569954 269764 569960 269816
rect 570012 269804 570018 269816
rect 570049 269807 570107 269813
rect 570049 269804 570061 269807
rect 570012 269776 570061 269804
rect 570012 269764 570018 269776
rect 570049 269773 570061 269776
rect 570095 269773 570107 269807
rect 570049 269767 570107 269773
rect 1946 269396 1952 269408
rect 1907 269368 1952 269396
rect 1946 269356 1952 269368
rect 2004 269356 2010 269408
rect 569954 267288 569960 267300
rect 569915 267260 569960 267288
rect 569954 267248 569960 267260
rect 570012 267248 570018 267300
rect 569 266611 627 266617
rect 569 266577 581 266611
rect 615 266608 627 266611
rect 1946 266608 1952 266620
rect 615 266580 1952 266608
rect 615 266577 627 266580
rect 569 266571 627 266577
rect 1946 266568 1952 266580
rect 2004 266568 2010 266620
rect 1857 266475 1915 266481
rect 1857 266441 1869 266475
rect 1903 266472 1915 266475
rect 1946 266472 1952 266484
rect 1903 266444 1952 266472
rect 1903 266441 1915 266444
rect 1857 266435 1915 266441
rect 1946 266432 1952 266444
rect 2004 266432 2010 266484
rect 569954 266364 569960 266416
rect 570012 266404 570018 266416
rect 570049 266407 570107 266413
rect 570049 266404 570061 266407
rect 570012 266376 570061 266404
rect 570012 266364 570018 266376
rect 570049 266373 570061 266376
rect 570095 266373 570107 266407
rect 570049 266367 570107 266373
rect 290 266296 296 266348
rect 348 266336 354 266348
rect 1946 266336 1952 266348
rect 348 266308 1952 266336
rect 348 266296 354 266308
rect 1946 266296 1952 266308
rect 2004 266296 2010 266348
rect 569954 265888 569960 265940
rect 570012 265928 570018 265940
rect 570141 265931 570199 265937
rect 570141 265928 570153 265931
rect 570012 265900 570153 265928
rect 570012 265888 570018 265900
rect 570141 265897 570153 265900
rect 570187 265897 570199 265931
rect 570141 265891 570199 265897
rect 1946 264704 1952 264716
rect 1907 264676 1952 264704
rect 1946 264664 1952 264676
rect 2004 264664 2010 264716
rect 382 264256 388 264308
rect 440 264296 446 264308
rect 1946 264296 1952 264308
rect 440 264268 1952 264296
rect 440 264256 446 264268
rect 1946 264256 1952 264268
rect 2004 264256 2010 264308
rect 1765 264163 1823 264169
rect 1765 264129 1777 264163
rect 1811 264160 1823 264163
rect 1946 264160 1952 264172
rect 1811 264132 1952 264160
rect 1811 264129 1823 264132
rect 1765 264123 1823 264129
rect 1946 264120 1952 264132
rect 2004 264120 2010 264172
rect 1302 263984 1308 264036
rect 1360 264024 1366 264036
rect 1946 264024 1952 264036
rect 1360 263996 1952 264024
rect 1360 263984 1366 263996
rect 1946 263984 1952 263996
rect 2004 263984 2010 264036
rect 569954 263984 569960 264036
rect 570012 264024 570018 264036
rect 570233 264027 570291 264033
rect 570233 264024 570245 264027
rect 570012 263996 570245 264024
rect 570012 263984 570018 263996
rect 570233 263993 570245 263996
rect 570279 263993 570291 264027
rect 570233 263987 570291 263993
rect 845 261579 903 261585
rect 845 261545 857 261579
rect 891 261576 903 261579
rect 1394 261576 1400 261588
rect 891 261548 1400 261576
rect 891 261545 903 261548
rect 845 261539 903 261545
rect 1394 261536 1400 261548
rect 1452 261536 1458 261588
rect 1118 261508 1124 261520
rect 1079 261480 1124 261508
rect 1118 261468 1124 261480
rect 1176 261468 1182 261520
rect 1765 261511 1823 261517
rect 1765 261477 1777 261511
rect 1811 261508 1823 261511
rect 1854 261508 1860 261520
rect 1811 261480 1860 261508
rect 1811 261477 1823 261480
rect 1765 261471 1823 261477
rect 1854 261468 1860 261480
rect 1912 261468 1918 261520
rect 1118 260720 1124 260772
rect 1176 260760 1182 260772
rect 1762 260760 1768 260772
rect 1176 260732 1768 260760
rect 1176 260720 1182 260732
rect 1762 260720 1768 260732
rect 1820 260720 1826 260772
rect 569954 259876 569960 259888
rect 569915 259848 569960 259876
rect 569954 259836 569960 259848
rect 570012 259836 570018 259888
rect 569954 259564 569960 259616
rect 570012 259604 570018 259616
rect 570233 259607 570291 259613
rect 570233 259604 570245 259607
rect 570012 259576 570245 259604
rect 570012 259564 570018 259576
rect 570233 259573 570245 259576
rect 570279 259573 570291 259607
rect 570233 259567 570291 259573
rect 1394 258204 1400 258256
rect 1452 258244 1458 258256
rect 1762 258244 1768 258256
rect 1452 258216 1768 258244
rect 1452 258204 1458 258216
rect 1762 258204 1768 258216
rect 1820 258204 1826 258256
rect 750 257388 756 257440
rect 808 257428 814 257440
rect 1394 257428 1400 257440
rect 808 257400 1400 257428
rect 808 257388 814 257400
rect 1394 257388 1400 257400
rect 1452 257388 1458 257440
rect 566 257252 572 257304
rect 624 257292 630 257304
rect 1946 257292 1952 257304
rect 624 257264 1952 257292
rect 624 257252 630 257264
rect 1946 257252 1952 257264
rect 2004 257252 2010 257304
rect 569954 256504 569960 256556
rect 570012 256544 570018 256556
rect 570230 256544 570236 256556
rect 570012 256516 570236 256544
rect 570012 256504 570018 256516
rect 570230 256504 570236 256516
rect 570288 256504 570294 256556
rect 569957 254779 570015 254785
rect 569957 254745 569969 254779
rect 570003 254776 570015 254779
rect 570046 254776 570052 254788
rect 570003 254748 570052 254776
rect 570003 254745 570015 254748
rect 569957 254739 570015 254745
rect 570046 254736 570052 254748
rect 570104 254736 570110 254788
rect 566 251852 572 251864
rect 527 251824 572 251852
rect 566 251812 572 251824
rect 624 251812 630 251864
rect 842 251852 848 251864
rect 803 251824 848 251852
rect 842 251812 848 251824
rect 900 251812 906 251864
rect 1765 251855 1823 251861
rect 1765 251821 1777 251855
rect 1811 251852 1823 251855
rect 1854 251852 1860 251864
rect 1811 251824 1860 251852
rect 1811 251821 1823 251824
rect 1765 251815 1823 251821
rect 1854 251812 1860 251824
rect 1912 251812 1918 251864
rect 569954 251744 569960 251796
rect 570012 251784 570018 251796
rect 570138 251784 570144 251796
rect 570012 251756 570144 251784
rect 570012 251744 570018 251756
rect 570138 251744 570144 251756
rect 570196 251744 570202 251796
rect 574738 251200 574744 251252
rect 574796 251240 574802 251252
rect 580166 251240 580172 251252
rect 574796 251212 580172 251240
rect 574796 251200 574802 251212
rect 580166 251200 580172 251212
rect 580224 251200 580230 251252
rect 569954 250928 569960 250980
rect 570012 250968 570018 250980
rect 570233 250971 570291 250977
rect 570233 250968 570245 250971
rect 570012 250940 570245 250968
rect 570012 250928 570018 250940
rect 570233 250937 570245 250940
rect 570279 250937 570291 250971
rect 570233 250931 570291 250937
rect 569954 250792 569960 250844
rect 570012 250832 570018 250844
rect 570322 250832 570328 250844
rect 570012 250804 570328 250832
rect 570012 250792 570018 250804
rect 570322 250792 570328 250804
rect 570380 250792 570386 250844
rect 569954 250588 569960 250640
rect 570012 250628 570018 250640
rect 570509 250631 570567 250637
rect 570509 250628 570521 250631
rect 570012 250600 570521 250628
rect 570012 250588 570018 250600
rect 570509 250597 570521 250600
rect 570555 250597 570567 250631
rect 570509 250591 570567 250597
rect 569954 250452 569960 250504
rect 570012 250492 570018 250504
rect 570049 250495 570107 250501
rect 570049 250492 570061 250495
rect 570012 250464 570061 250492
rect 570012 250452 570018 250464
rect 570049 250461 570061 250464
rect 570095 250461 570107 250495
rect 570049 250455 570107 250461
rect 1489 250291 1547 250297
rect 1489 250257 1501 250291
rect 1535 250288 1547 250291
rect 1946 250288 1952 250300
rect 1535 250260 1952 250288
rect 1535 250257 1547 250260
rect 1489 250251 1547 250257
rect 1946 250248 1952 250260
rect 2004 250248 2010 250300
rect 1946 250152 1952 250164
rect 1907 250124 1952 250152
rect 1946 250112 1952 250124
rect 2004 250112 2010 250164
rect 1302 248956 1308 249008
rect 1360 248996 1366 249008
rect 1946 248996 1952 249008
rect 1360 248968 1952 248996
rect 1360 248956 1366 248968
rect 1946 248956 1952 248968
rect 2004 248956 2010 249008
rect 569954 247256 569960 247308
rect 570012 247296 570018 247308
rect 570325 247299 570383 247305
rect 570325 247296 570337 247299
rect 570012 247268 570337 247296
rect 570012 247256 570018 247268
rect 570325 247265 570337 247268
rect 570371 247265 570383 247299
rect 570325 247259 570383 247265
rect 570046 246684 570052 246696
rect 570007 246656 570052 246684
rect 570046 246644 570052 246656
rect 570104 246644 570110 246696
rect 570046 246508 570052 246560
rect 570104 246548 570110 246560
rect 570233 246551 570291 246557
rect 570233 246548 570245 246551
rect 570104 246520 570245 246548
rect 570104 246508 570110 246520
rect 570233 246517 570245 246520
rect 570279 246517 570291 246551
rect 570233 246511 570291 246517
rect 569957 246007 570015 246013
rect 569957 245973 569969 246007
rect 570003 246004 570015 246007
rect 570233 246007 570291 246013
rect 570233 246004 570245 246007
rect 570003 245976 570245 246004
rect 570003 245973 570015 245976
rect 569957 245967 570015 245973
rect 570233 245973 570245 245976
rect 570279 245973 570291 246007
rect 570233 245967 570291 245973
rect 569865 245735 569923 245741
rect 569865 245701 569877 245735
rect 569911 245732 569923 245735
rect 569957 245735 570015 245741
rect 569957 245732 569969 245735
rect 569911 245704 569969 245732
rect 569911 245701 569923 245704
rect 569865 245695 569923 245701
rect 569957 245701 569969 245704
rect 570003 245701 570015 245735
rect 569957 245695 570015 245701
rect 569865 245395 569923 245401
rect 569865 245361 569877 245395
rect 569911 245392 569923 245395
rect 570509 245395 570567 245401
rect 570509 245392 570521 245395
rect 569911 245364 570521 245392
rect 569911 245361 569923 245364
rect 569865 245355 569923 245361
rect 570509 245361 570521 245364
rect 570555 245361 570567 245395
rect 570509 245355 570567 245361
rect 569954 243652 569960 243704
rect 570012 243692 570018 243704
rect 570233 243695 570291 243701
rect 570233 243692 570245 243695
rect 570012 243664 570245 243692
rect 570012 243652 570018 243664
rect 570233 243661 570245 243664
rect 570279 243661 570291 243695
rect 570233 243655 570291 243661
rect 569954 243516 569960 243568
rect 570012 243556 570018 243568
rect 570049 243559 570107 243565
rect 570049 243556 570061 243559
rect 570012 243528 570061 243556
rect 570012 243516 570018 243528
rect 570049 243525 570061 243528
rect 570095 243525 570107 243559
rect 570049 243519 570107 243525
rect 1946 243080 1952 243092
rect 1907 243052 1952 243080
rect 1946 243040 1952 243052
rect 2004 243040 2010 243092
rect 1946 242904 1952 242956
rect 2004 242944 2010 242956
rect 2004 242916 2049 242944
rect 2004 242904 2010 242916
rect 1946 242536 1952 242548
rect 1907 242508 1952 242536
rect 1946 242496 1952 242508
rect 2004 242496 2010 242548
rect 1673 242267 1731 242273
rect 1673 242233 1685 242267
rect 1719 242264 1731 242267
rect 1854 242264 1860 242276
rect 1719 242236 1860 242264
rect 1719 242233 1731 242236
rect 1673 242227 1731 242233
rect 1854 242224 1860 242236
rect 1912 242224 1918 242276
rect 1946 242224 1952 242276
rect 2004 242224 2010 242276
rect 1762 242196 1768 242208
rect 1723 242168 1768 242196
rect 1762 242156 1768 242168
rect 1820 242156 1826 242208
rect 1581 242131 1639 242137
rect 1581 242097 1593 242131
rect 1627 242128 1639 242131
rect 1857 242131 1915 242137
rect 1857 242128 1869 242131
rect 1627 242100 1869 242128
rect 1627 242097 1639 242100
rect 1581 242091 1639 242097
rect 1857 242097 1869 242100
rect 1903 242097 1915 242131
rect 1857 242091 1915 242097
rect 1121 242063 1179 242069
rect 1121 242029 1133 242063
rect 1167 242060 1179 242063
rect 1762 242060 1768 242072
rect 1167 242032 1768 242060
rect 1167 242029 1179 242032
rect 1121 242023 1179 242029
rect 1762 242020 1768 242032
rect 1820 242020 1826 242072
rect 1857 241995 1915 242001
rect 1857 241961 1869 241995
rect 1903 241992 1915 241995
rect 1964 241992 1992 242224
rect 1903 241964 1992 241992
rect 1903 241961 1915 241964
rect 1857 241955 1915 241961
rect 474 241612 480 241664
rect 532 241652 538 241664
rect 1946 241652 1952 241664
rect 532 241624 1952 241652
rect 532 241612 538 241624
rect 1946 241612 1952 241624
rect 2004 241612 2010 241664
rect 570138 239436 570144 239488
rect 570196 239476 570202 239488
rect 570417 239479 570475 239485
rect 570417 239476 570429 239479
rect 570196 239448 570429 239476
rect 570196 239436 570202 239448
rect 570417 239445 570429 239448
rect 570463 239445 570475 239479
rect 570417 239439 570475 239445
rect 1946 238456 1952 238468
rect 1412 238428 1952 238456
rect 1412 238252 1440 238428
rect 1946 238416 1952 238428
rect 2004 238416 2010 238468
rect 1489 238323 1547 238329
rect 1489 238289 1501 238323
rect 1535 238320 1547 238323
rect 1946 238320 1952 238332
rect 1535 238292 1952 238320
rect 1535 238289 1547 238292
rect 1489 238283 1547 238289
rect 1946 238280 1952 238292
rect 2004 238280 2010 238332
rect 1412 238224 1992 238252
rect 1964 238196 1992 238224
rect 1489 238187 1547 238193
rect 1489 238153 1501 238187
rect 1535 238184 1547 238187
rect 1762 238184 1768 238196
rect 1535 238156 1768 238184
rect 1535 238153 1547 238156
rect 1489 238147 1547 238153
rect 1762 238144 1768 238156
rect 1820 238144 1826 238196
rect 1946 238144 1952 238196
rect 2004 238144 2010 238196
rect 1673 237983 1731 237989
rect 1673 237949 1685 237983
rect 1719 237980 1731 237983
rect 1854 237980 1860 237992
rect 1719 237952 1860 237980
rect 1719 237949 1731 237952
rect 1673 237943 1731 237949
rect 1854 237940 1860 237952
rect 1912 237940 1918 237992
rect 569954 236036 569960 236088
rect 570012 236076 570018 236088
rect 570049 236079 570107 236085
rect 570049 236076 570061 236079
rect 570012 236048 570061 236076
rect 570012 236036 570018 236048
rect 570049 236045 570061 236048
rect 570095 236045 570107 236079
rect 570049 236039 570107 236045
rect 474 235424 480 235476
rect 532 235464 538 235476
rect 1762 235464 1768 235476
rect 532 235436 1768 235464
rect 532 235424 538 235436
rect 1762 235424 1768 235436
rect 1820 235424 1826 235476
rect 569954 233656 569960 233708
rect 570012 233696 570018 233708
rect 570509 233699 570567 233705
rect 570509 233696 570521 233699
rect 570012 233668 570521 233696
rect 570012 233656 570018 233668
rect 570509 233665 570521 233668
rect 570555 233665 570567 233699
rect 570509 233659 570567 233665
rect 569954 233520 569960 233572
rect 570012 233560 570018 233572
rect 570138 233560 570144 233572
rect 570012 233532 570144 233560
rect 570012 233520 570018 233532
rect 570138 233520 570144 233532
rect 570196 233520 570202 233572
rect 569954 230228 569960 230240
rect 569915 230200 569960 230228
rect 569954 230188 569960 230200
rect 570012 230188 570018 230240
rect 569954 229984 569960 230036
rect 570012 230024 570018 230036
rect 570138 230024 570144 230036
rect 570012 229996 570144 230024
rect 570012 229984 570018 229996
rect 570138 229984 570144 229996
rect 570196 229984 570202 230036
rect 570141 229891 570199 229897
rect 570141 229857 570153 229891
rect 570187 229888 570199 229891
rect 570414 229888 570420 229900
rect 570187 229860 570420 229888
rect 570187 229857 570199 229860
rect 570141 229851 570199 229857
rect 570414 229848 570420 229860
rect 570472 229848 570478 229900
rect 569954 229780 569960 229832
rect 570012 229820 570018 229832
rect 570322 229820 570328 229832
rect 570012 229792 570328 229820
rect 570012 229780 570018 229792
rect 570322 229780 570328 229792
rect 570380 229780 570386 229832
rect 570138 229712 570144 229764
rect 570196 229752 570202 229764
rect 570233 229755 570291 229761
rect 570233 229752 570245 229755
rect 570196 229724 570245 229752
rect 570196 229712 570202 229724
rect 570233 229721 570245 229724
rect 570279 229721 570291 229755
rect 570233 229715 570291 229721
rect 569957 229687 570015 229693
rect 569957 229653 569969 229687
rect 570003 229684 570015 229687
rect 570046 229684 570052 229696
rect 570003 229656 570052 229684
rect 570003 229653 570015 229656
rect 569957 229647 570015 229653
rect 570046 229644 570052 229656
rect 570104 229644 570110 229696
rect 569954 229236 569960 229288
rect 570012 229276 570018 229288
rect 570509 229279 570567 229285
rect 570509 229276 570521 229279
rect 570012 229248 570521 229276
rect 570012 229236 570018 229248
rect 570509 229245 570521 229248
rect 570555 229245 570567 229279
rect 570509 229239 570567 229245
rect 569957 228735 570015 228741
rect 569957 228701 569969 228735
rect 570003 228732 570015 228735
rect 570325 228735 570383 228741
rect 570325 228732 570337 228735
rect 570003 228704 570337 228732
rect 570003 228701 570015 228704
rect 569957 228695 570015 228701
rect 570325 228701 570337 228704
rect 570371 228701 570383 228735
rect 570325 228695 570383 228701
rect 1762 228392 1768 228404
rect 1723 228364 1768 228392
rect 1762 228352 1768 228364
rect 1820 228352 1826 228404
rect 570046 227032 570052 227044
rect 570007 227004 570052 227032
rect 570046 226992 570052 227004
rect 570104 226992 570110 227044
rect 570049 226899 570107 226905
rect 570049 226865 570061 226899
rect 570095 226896 570107 226899
rect 570230 226896 570236 226908
rect 570095 226868 570236 226896
rect 570095 226865 570107 226868
rect 570049 226859 570107 226865
rect 570230 226856 570236 226868
rect 570288 226856 570294 226908
rect 569954 225972 569960 226024
rect 570012 226012 570018 226024
rect 570230 226012 570236 226024
rect 570012 225984 570236 226012
rect 570012 225972 570018 225984
rect 570230 225972 570236 225984
rect 570288 225972 570294 226024
rect 569954 225768 569960 225820
rect 570012 225808 570018 225820
rect 570325 225811 570383 225817
rect 570325 225808 570337 225811
rect 570012 225780 570337 225808
rect 570012 225768 570018 225780
rect 570325 225777 570337 225780
rect 570371 225777 570383 225811
rect 570325 225771 570383 225777
rect 1581 222615 1639 222621
rect 1581 222581 1593 222615
rect 1627 222612 1639 222615
rect 1857 222615 1915 222621
rect 1857 222612 1869 222615
rect 1627 222584 1869 222612
rect 1627 222581 1639 222584
rect 1581 222575 1639 222581
rect 1857 222581 1869 222584
rect 1903 222581 1915 222615
rect 1857 222575 1915 222581
rect 845 221731 903 221737
rect 845 221697 857 221731
rect 891 221728 903 221731
rect 1946 221728 1952 221740
rect 891 221700 1952 221728
rect 891 221697 903 221700
rect 845 221691 903 221697
rect 1946 221688 1952 221700
rect 2004 221688 2010 221740
rect 750 221620 756 221672
rect 808 221660 814 221672
rect 1394 221660 1400 221672
rect 808 221632 1400 221660
rect 808 221620 814 221632
rect 1394 221620 1400 221632
rect 1452 221620 1458 221672
rect 1302 221524 1308 221536
rect 1263 221496 1308 221524
rect 1302 221484 1308 221496
rect 1360 221484 1366 221536
rect 1394 221484 1400 221536
rect 1452 221524 1458 221536
rect 1489 221527 1547 221533
rect 1489 221524 1501 221527
rect 1452 221496 1501 221524
rect 1452 221484 1458 221496
rect 1489 221493 1501 221496
rect 1535 221493 1547 221527
rect 1489 221487 1547 221493
rect 1673 221527 1731 221533
rect 1673 221493 1685 221527
rect 1719 221524 1731 221527
rect 1949 221527 2007 221533
rect 1949 221524 1961 221527
rect 1719 221496 1961 221524
rect 1719 221493 1731 221496
rect 1673 221487 1731 221493
rect 1949 221493 1961 221496
rect 1995 221493 2007 221527
rect 1949 221487 2007 221493
rect 382 221348 388 221400
rect 440 221388 446 221400
rect 1949 221391 2007 221397
rect 1949 221388 1961 221391
rect 440 221360 1961 221388
rect 440 221348 446 221360
rect 1949 221357 1961 221360
rect 1995 221357 2007 221391
rect 1949 221351 2007 221357
rect 1394 221280 1400 221332
rect 1452 221320 1458 221332
rect 1765 221323 1823 221329
rect 1765 221320 1777 221323
rect 1452 221292 1777 221320
rect 1452 221280 1458 221292
rect 1765 221289 1777 221292
rect 1811 221289 1823 221323
rect 1765 221283 1823 221289
rect 293 221051 351 221057
rect 293 221017 305 221051
rect 339 221048 351 221051
rect 1946 221048 1952 221060
rect 339 221020 1952 221048
rect 339 221017 351 221020
rect 293 221011 351 221017
rect 1946 221008 1952 221020
rect 2004 221008 2010 221060
rect 1581 219963 1639 219969
rect 1581 219929 1593 219963
rect 1627 219960 1639 219963
rect 1946 219960 1952 219972
rect 1627 219932 1952 219960
rect 1627 219929 1639 219932
rect 1581 219923 1639 219929
rect 1946 219920 1952 219932
rect 2004 219920 2010 219972
rect 1765 218331 1823 218337
rect 1765 218297 1777 218331
rect 1811 218328 1823 218331
rect 1946 218328 1952 218340
rect 1811 218300 1952 218328
rect 1811 218297 1823 218300
rect 1765 218291 1823 218297
rect 1946 218288 1952 218300
rect 2004 218288 2010 218340
rect 1765 217719 1823 217725
rect 1765 217685 1777 217719
rect 1811 217716 1823 217719
rect 1946 217716 1952 217728
rect 1811 217688 1952 217716
rect 1811 217685 1823 217688
rect 1765 217679 1823 217685
rect 1946 217676 1952 217688
rect 2004 217676 2010 217728
rect 1394 217404 1400 217456
rect 1452 217444 1458 217456
rect 1765 217447 1823 217453
rect 1765 217444 1777 217447
rect 1452 217416 1777 217444
rect 1452 217404 1458 217416
rect 1765 217413 1777 217416
rect 1811 217413 1823 217447
rect 1765 217407 1823 217413
rect 106 216792 112 216844
rect 164 216832 170 216844
rect 1397 216835 1455 216841
rect 1397 216832 1409 216835
rect 164 216804 1409 216832
rect 164 216792 170 216804
rect 1397 216801 1409 216804
rect 1443 216801 1455 216835
rect 1397 216795 1455 216801
rect 569954 215676 569960 215688
rect 569880 215648 569960 215676
rect 569880 215404 569908 215648
rect 569954 215636 569960 215648
rect 570012 215636 570018 215688
rect 569954 215404 569960 215416
rect 569880 215376 569960 215404
rect 569954 215364 569960 215376
rect 570012 215364 570018 215416
rect 569954 214616 569960 214668
rect 570012 214656 570018 214668
rect 570325 214659 570383 214665
rect 570325 214656 570337 214659
rect 570012 214628 570337 214656
rect 570012 214616 570018 214628
rect 570325 214625 570337 214628
rect 570371 214625 570383 214659
rect 570325 214619 570383 214625
rect 570138 214588 570144 214600
rect 570099 214560 570144 214588
rect 570138 214548 570144 214560
rect 570196 214548 570202 214600
rect 1394 214276 1400 214328
rect 1452 214316 1458 214328
rect 1946 214316 1952 214328
rect 1452 214288 1952 214316
rect 1452 214276 1458 214288
rect 1946 214276 1952 214288
rect 2004 214276 2010 214328
rect 566 214140 572 214192
rect 624 214180 630 214192
rect 1946 214180 1952 214192
rect 624 214152 1952 214180
rect 624 214140 630 214152
rect 1946 214140 1952 214152
rect 2004 214140 2010 214192
rect 569954 214004 569960 214056
rect 570012 214044 570018 214056
rect 570230 214044 570236 214056
rect 570012 214016 570236 214044
rect 570012 214004 570018 214016
rect 570230 214004 570236 214016
rect 570288 214004 570294 214056
rect 1305 212891 1363 212897
rect 1305 212857 1317 212891
rect 1351 212888 1363 212891
rect 1946 212888 1952 212900
rect 1351 212860 1952 212888
rect 1351 212857 1363 212860
rect 1305 212851 1363 212857
rect 1946 212848 1952 212860
rect 2004 212848 2010 212900
rect 842 209924 848 209976
rect 900 209964 906 209976
rect 1305 209967 1363 209973
rect 1305 209964 1317 209967
rect 900 209936 1317 209964
rect 900 209924 906 209936
rect 1305 209933 1317 209936
rect 1351 209933 1363 209967
rect 1305 209927 1363 209933
rect 570138 208360 570144 208412
rect 570196 208400 570202 208412
rect 570414 208400 570420 208412
rect 570196 208372 570420 208400
rect 570196 208360 570202 208372
rect 570414 208360 570420 208372
rect 570472 208360 570478 208412
rect 1121 207791 1179 207797
rect 1121 207757 1133 207791
rect 1167 207788 1179 207791
rect 1581 207791 1639 207797
rect 1581 207788 1593 207791
rect 1167 207760 1593 207788
rect 1167 207757 1179 207760
rect 1121 207751 1179 207757
rect 1581 207757 1593 207760
rect 1627 207757 1639 207791
rect 1581 207751 1639 207757
rect 1210 207720 1216 207732
rect 1171 207692 1216 207720
rect 1210 207680 1216 207692
rect 1268 207680 1274 207732
rect 1857 205819 1915 205825
rect 1857 205816 1869 205819
rect 1780 205788 1869 205816
rect 1780 205689 1808 205788
rect 1857 205785 1869 205788
rect 1903 205785 1915 205819
rect 1857 205779 1915 205785
rect 1765 205683 1823 205689
rect 1765 205649 1777 205683
rect 1811 205649 1823 205683
rect 1765 205643 1823 205649
rect 570049 205479 570107 205485
rect 570049 205445 570061 205479
rect 570095 205476 570107 205479
rect 570233 205479 570291 205485
rect 570233 205476 570245 205479
rect 570095 205448 570245 205476
rect 570095 205445 570107 205448
rect 570049 205439 570107 205445
rect 570233 205445 570245 205448
rect 570279 205445 570291 205479
rect 570233 205439 570291 205445
rect 569957 205207 570015 205213
rect 569957 205204 569969 205207
rect 569880 205176 569969 205204
rect 566 205028 572 205080
rect 624 205068 630 205080
rect 1210 205068 1216 205080
rect 624 205040 1216 205068
rect 624 205028 630 205040
rect 1210 205028 1216 205040
rect 1268 205028 1274 205080
rect 1029 204935 1087 204941
rect 1029 204901 1041 204935
rect 1075 204932 1087 204935
rect 1394 204932 1400 204944
rect 1075 204904 1400 204932
rect 1075 204901 1087 204904
rect 1029 204895 1087 204901
rect 1394 204892 1400 204904
rect 1452 204892 1458 204944
rect 569880 204932 569908 205176
rect 569957 205173 569969 205176
rect 570003 205173 570015 205207
rect 569957 205167 570015 205173
rect 569954 205028 569960 205080
rect 570012 205068 570018 205080
rect 570230 205068 570236 205080
rect 570012 205040 570236 205068
rect 570012 205028 570018 205040
rect 570230 205028 570236 205040
rect 570288 205028 570294 205080
rect 569957 204935 570015 204941
rect 569957 204932 569969 204935
rect 569880 204904 569969 204932
rect 569957 204901 569969 204904
rect 570003 204901 570015 204935
rect 569957 204895 570015 204901
rect 1946 204864 1952 204876
rect 1412 204836 1952 204864
rect 1412 204808 1440 204836
rect 1946 204824 1952 204836
rect 2004 204824 2010 204876
rect 1394 204756 1400 204808
rect 1452 204756 1458 204808
rect 569954 204756 569960 204808
rect 570012 204796 570018 204808
rect 570049 204799 570107 204805
rect 570049 204796 570061 204799
rect 570012 204768 570061 204796
rect 570012 204756 570018 204768
rect 570049 204765 570061 204768
rect 570095 204765 570107 204799
rect 570049 204759 570107 204765
rect 1489 204731 1547 204737
rect 1489 204697 1501 204731
rect 1535 204728 1547 204731
rect 1946 204728 1952 204740
rect 1535 204700 1952 204728
rect 1535 204697 1547 204700
rect 1489 204691 1547 204697
rect 1946 204688 1952 204700
rect 2004 204688 2010 204740
rect 570046 204416 570052 204468
rect 570104 204456 570110 204468
rect 570233 204459 570291 204465
rect 570233 204456 570245 204459
rect 570104 204428 570245 204456
rect 570104 204416 570110 204428
rect 570233 204425 570245 204428
rect 570279 204425 570291 204459
rect 570233 204419 570291 204425
rect 574830 204280 574836 204332
rect 574888 204320 574894 204332
rect 580166 204320 580172 204332
rect 574888 204292 580172 204320
rect 574888 204280 574894 204292
rect 580166 204280 580172 204292
rect 580224 204280 580230 204332
rect 569954 203668 569960 203720
rect 570012 203708 570018 203720
rect 570049 203711 570107 203717
rect 570049 203708 570061 203711
rect 570012 203680 570061 203708
rect 570012 203668 570018 203680
rect 570049 203677 570061 203680
rect 570095 203677 570107 203711
rect 570049 203671 570107 203677
rect 569954 203532 569960 203584
rect 570012 203572 570018 203584
rect 570325 203575 570383 203581
rect 570325 203572 570337 203575
rect 570012 203544 570337 203572
rect 570012 203532 570018 203544
rect 570325 203541 570337 203544
rect 570371 203541 570383 203575
rect 570325 203535 570383 203541
rect 569954 203396 569960 203448
rect 570012 203436 570018 203448
rect 570230 203436 570236 203448
rect 570012 203408 570236 203436
rect 570012 203396 570018 203408
rect 570230 203396 570236 203408
rect 570288 203396 570294 203448
rect 569954 203124 569960 203176
rect 570012 203164 570018 203176
rect 570049 203167 570107 203173
rect 570049 203164 570061 203167
rect 570012 203136 570061 203164
rect 570012 203124 570018 203136
rect 570049 203133 570061 203136
rect 570095 203133 570107 203167
rect 570049 203127 570107 203133
rect 569954 202988 569960 203040
rect 570012 203028 570018 203040
rect 570141 203031 570199 203037
rect 570141 203028 570153 203031
rect 570012 203000 570153 203028
rect 570012 202988 570018 203000
rect 570141 202997 570153 203000
rect 570187 202997 570199 203031
rect 570141 202991 570199 202997
rect 569954 202620 569960 202632
rect 569915 202592 569960 202620
rect 569954 202580 569960 202592
rect 570012 202580 570018 202632
rect 661 201875 719 201881
rect 661 201841 673 201875
rect 707 201872 719 201875
rect 1946 201872 1952 201884
rect 707 201844 1952 201872
rect 707 201841 719 201844
rect 661 201835 719 201841
rect 1946 201832 1952 201844
rect 2004 201832 2010 201884
rect 1029 200855 1087 200861
rect 1029 200821 1041 200855
rect 1075 200852 1087 200855
rect 1489 200855 1547 200861
rect 1489 200852 1501 200855
rect 1075 200824 1501 200852
rect 1075 200821 1087 200824
rect 1029 200815 1087 200821
rect 1489 200821 1501 200824
rect 1535 200821 1547 200855
rect 1489 200815 1547 200821
rect 1489 200719 1547 200725
rect 1489 200685 1501 200719
rect 1535 200716 1547 200719
rect 1857 200719 1915 200725
rect 1857 200716 1869 200719
rect 1535 200688 1869 200716
rect 1535 200685 1547 200688
rect 1489 200679 1547 200685
rect 1857 200685 1869 200688
rect 1903 200685 1915 200719
rect 1857 200679 1915 200685
rect 566 200200 572 200252
rect 624 200240 630 200252
rect 1394 200240 1400 200252
rect 624 200212 1400 200240
rect 624 200200 630 200212
rect 1394 200200 1400 200212
rect 1452 200200 1458 200252
rect 290 199492 296 199504
rect 251 199464 296 199492
rect 290 199452 296 199464
rect 348 199452 354 199504
rect 842 199492 848 199504
rect 803 199464 848 199492
rect 842 199452 848 199464
rect 900 199452 906 199504
rect 1029 198883 1087 198889
rect 1029 198849 1041 198883
rect 1075 198880 1087 198883
rect 1075 198852 1164 198880
rect 1075 198849 1087 198852
rect 1029 198843 1087 198849
rect 1136 198744 1164 198852
rect 1581 198747 1639 198753
rect 1581 198744 1593 198747
rect 1136 198716 1593 198744
rect 1581 198713 1593 198716
rect 1627 198713 1639 198747
rect 1581 198707 1639 198713
rect 1394 198228 1400 198280
rect 1452 198268 1458 198280
rect 1452 198240 1992 198268
rect 1452 198228 1458 198240
rect 1964 198212 1992 198240
rect 1581 198203 1639 198209
rect 1581 198169 1593 198203
rect 1627 198200 1639 198203
rect 1857 198203 1915 198209
rect 1857 198200 1869 198203
rect 1627 198172 1869 198200
rect 1627 198169 1639 198172
rect 1581 198163 1639 198169
rect 1857 198169 1869 198172
rect 1903 198169 1915 198203
rect 1857 198163 1915 198169
rect 1946 198160 1952 198212
rect 2004 198160 2010 198212
rect 1394 198024 1400 198076
rect 1452 198064 1458 198076
rect 1581 198067 1639 198073
rect 1452 198036 1497 198064
rect 1452 198024 1458 198036
rect 1581 198033 1593 198067
rect 1627 198064 1639 198067
rect 1949 198067 2007 198073
rect 1949 198064 1961 198067
rect 1627 198036 1961 198064
rect 1627 198033 1639 198036
rect 1581 198027 1639 198033
rect 1949 198033 1961 198036
rect 1995 198033 2007 198067
rect 1949 198027 2007 198033
rect 1121 197931 1179 197937
rect 1121 197897 1133 197931
rect 1167 197928 1179 197931
rect 1305 197931 1363 197937
rect 1305 197928 1317 197931
rect 1167 197900 1317 197928
rect 1167 197897 1179 197900
rect 1121 197891 1179 197897
rect 1305 197897 1317 197900
rect 1351 197897 1363 197931
rect 1305 197891 1363 197897
rect 1121 197795 1179 197801
rect 1121 197761 1133 197795
rect 1167 197792 1179 197795
rect 1946 197792 1952 197804
rect 1167 197764 1952 197792
rect 1167 197761 1179 197764
rect 1121 197755 1179 197761
rect 1946 197752 1952 197764
rect 2004 197752 2010 197804
rect 934 197656 940 197668
rect 895 197628 940 197656
rect 934 197616 940 197628
rect 992 197616 998 197668
rect 1946 197656 1952 197668
rect 1907 197628 1952 197656
rect 1946 197616 1952 197628
rect 2004 197616 2010 197668
rect 934 197480 940 197532
rect 992 197520 998 197532
rect 1673 197523 1731 197529
rect 1673 197520 1685 197523
rect 992 197492 1685 197520
rect 992 197480 998 197492
rect 1673 197489 1685 197492
rect 1719 197489 1731 197523
rect 1673 197483 1731 197489
rect 1946 196364 1952 196376
rect 1907 196336 1952 196364
rect 1946 196324 1952 196336
rect 2004 196324 2010 196376
rect 845 196231 903 196237
rect 845 196197 857 196231
rect 891 196228 903 196231
rect 1946 196228 1952 196240
rect 891 196200 1952 196228
rect 891 196197 903 196200
rect 845 196191 903 196197
rect 1946 196188 1952 196200
rect 2004 196188 2010 196240
rect 1857 196095 1915 196101
rect 1857 196061 1869 196095
rect 1903 196092 1915 196095
rect 1946 196092 1952 196104
rect 1903 196064 1952 196092
rect 1903 196061 1915 196064
rect 1857 196055 1915 196061
rect 1946 196052 1952 196064
rect 2004 196052 2010 196104
rect 937 195959 995 195965
rect 937 195925 949 195959
rect 983 195956 995 195959
rect 1946 195956 1952 195968
rect 983 195928 1952 195956
rect 983 195925 995 195928
rect 937 195919 995 195925
rect 1946 195916 1952 195928
rect 2004 195916 2010 195968
rect 1305 195823 1363 195829
rect 1305 195789 1317 195823
rect 1351 195820 1363 195823
rect 1946 195820 1952 195832
rect 1351 195792 1952 195820
rect 1351 195789 1363 195792
rect 1305 195783 1363 195789
rect 1946 195780 1952 195792
rect 2004 195780 2010 195832
rect 1486 195644 1492 195696
rect 1544 195684 1550 195696
rect 1673 195687 1731 195693
rect 1673 195684 1685 195687
rect 1544 195656 1685 195684
rect 1544 195644 1550 195656
rect 1673 195653 1685 195656
rect 1719 195653 1731 195687
rect 1673 195647 1731 195653
rect 1302 195508 1308 195560
rect 1360 195548 1366 195560
rect 1486 195548 1492 195560
rect 1360 195520 1492 195548
rect 1360 195508 1366 195520
rect 1486 195508 1492 195520
rect 1544 195508 1550 195560
rect 1489 195211 1547 195217
rect 1489 195177 1501 195211
rect 1535 195208 1547 195211
rect 1765 195211 1823 195217
rect 1765 195208 1777 195211
rect 1535 195180 1777 195208
rect 1535 195177 1547 195180
rect 1489 195171 1547 195177
rect 1765 195177 1777 195180
rect 1811 195177 1823 195211
rect 1765 195171 1823 195177
rect 658 195100 664 195152
rect 716 195140 722 195152
rect 1857 195143 1915 195149
rect 1857 195140 1869 195143
rect 716 195112 1869 195140
rect 716 195100 722 195112
rect 1857 195109 1869 195112
rect 1903 195109 1915 195143
rect 1857 195103 1915 195109
rect 1213 195075 1271 195081
rect 1213 195041 1225 195075
rect 1259 195072 1271 195075
rect 1946 195072 1952 195084
rect 1259 195044 1952 195072
rect 1259 195041 1271 195044
rect 1213 195035 1271 195041
rect 1946 195032 1952 195044
rect 2004 195032 2010 195084
rect 1210 194896 1216 194948
rect 1268 194936 1274 194948
rect 1946 194936 1952 194948
rect 1268 194908 1952 194936
rect 1268 194896 1274 194908
rect 1946 194896 1952 194908
rect 2004 194896 2010 194948
rect 1121 194735 1179 194741
rect 1121 194701 1133 194735
rect 1167 194732 1179 194735
rect 1946 194732 1952 194744
rect 1167 194704 1952 194732
rect 1167 194701 1179 194704
rect 1121 194695 1179 194701
rect 1946 194692 1952 194704
rect 2004 194692 2010 194744
rect 658 193984 664 193996
rect 619 193956 664 193984
rect 658 193944 664 193956
rect 716 193944 722 193996
rect 1397 193987 1455 193993
rect 1397 193953 1409 193987
rect 1443 193984 1455 193987
rect 1946 193984 1952 193996
rect 1443 193956 1952 193984
rect 1443 193953 1455 193956
rect 1397 193947 1455 193953
rect 1946 193944 1952 193956
rect 2004 193944 2010 193996
rect 569954 193876 569960 193928
rect 570012 193916 570018 193928
rect 570141 193919 570199 193925
rect 570141 193916 570153 193919
rect 570012 193888 570153 193916
rect 570012 193876 570018 193888
rect 570141 193885 570153 193888
rect 570187 193885 570199 193919
rect 570141 193879 570199 193885
rect 569954 192720 569960 192772
rect 570012 192760 570018 192772
rect 570417 192763 570475 192769
rect 570417 192760 570429 192763
rect 570012 192732 570429 192760
rect 570012 192720 570018 192732
rect 570417 192729 570429 192732
rect 570463 192729 570475 192763
rect 570417 192723 570475 192729
rect 569954 192448 569960 192500
rect 570012 192488 570018 192500
rect 570012 192460 570057 192488
rect 570012 192448 570018 192460
rect 569954 192176 569960 192228
rect 570012 192216 570018 192228
rect 570049 192219 570107 192225
rect 570049 192216 570061 192219
rect 570012 192188 570061 192216
rect 570012 192176 570018 192188
rect 570049 192185 570061 192188
rect 570095 192185 570107 192219
rect 570049 192179 570107 192185
rect 569954 192040 569960 192092
rect 570012 192080 570018 192092
rect 570325 192083 570383 192089
rect 570325 192080 570337 192083
rect 570012 192052 570337 192080
rect 570012 192040 570018 192052
rect 570325 192049 570337 192052
rect 570371 192049 570383 192083
rect 570325 192043 570383 192049
rect 570046 192012 570052 192024
rect 569880 191984 570052 192012
rect 569880 191876 569908 191984
rect 570046 191972 570052 191984
rect 570104 191972 570110 192024
rect 569954 191904 569960 191956
rect 570012 191944 570018 191956
rect 570233 191947 570291 191953
rect 570233 191944 570245 191947
rect 570012 191916 570245 191944
rect 570012 191904 570018 191916
rect 570233 191913 570245 191916
rect 570279 191913 570291 191947
rect 570233 191907 570291 191913
rect 569880 191848 570092 191876
rect 570064 191752 570092 191848
rect 569954 191740 569960 191752
rect 569880 191712 569960 191740
rect 569880 191468 569908 191712
rect 569954 191700 569960 191712
rect 570012 191700 570018 191752
rect 570046 191700 570052 191752
rect 570104 191700 570110 191752
rect 569954 191564 569960 191616
rect 570012 191604 570018 191616
rect 570322 191604 570328 191616
rect 570012 191576 570328 191604
rect 570012 191564 570018 191576
rect 570322 191564 570328 191576
rect 570380 191564 570386 191616
rect 570138 191496 570144 191548
rect 570196 191536 570202 191548
rect 570417 191539 570475 191545
rect 570417 191536 570429 191539
rect 570196 191508 570429 191536
rect 570196 191496 570202 191508
rect 570417 191505 570429 191508
rect 570463 191505 570475 191539
rect 570417 191499 570475 191505
rect 569954 191468 569960 191480
rect 569880 191440 569960 191468
rect 569954 191428 569960 191440
rect 570012 191428 570018 191480
rect 1397 189771 1455 189777
rect 1397 189737 1409 189771
rect 1443 189768 1455 189771
rect 1946 189768 1952 189780
rect 1443 189740 1952 189768
rect 1443 189737 1455 189740
rect 1397 189731 1455 189737
rect 1946 189728 1952 189740
rect 2004 189728 2010 189780
rect 1489 189635 1547 189641
rect 1489 189601 1501 189635
rect 1535 189632 1547 189635
rect 1946 189632 1952 189644
rect 1535 189604 1952 189632
rect 1535 189601 1547 189604
rect 1489 189595 1547 189601
rect 1946 189592 1952 189604
rect 2004 189592 2010 189644
rect 1305 189227 1363 189233
rect 1305 189193 1317 189227
rect 1351 189224 1363 189227
rect 1946 189224 1952 189236
rect 1351 189196 1952 189224
rect 1351 189193 1363 189196
rect 1305 189187 1363 189193
rect 1946 189184 1952 189196
rect 2004 189184 2010 189236
rect 1213 188955 1271 188961
rect 1213 188921 1225 188955
rect 1259 188952 1271 188955
rect 1946 188952 1952 188964
rect 1259 188924 1952 188952
rect 1259 188921 1271 188924
rect 1213 188915 1271 188921
rect 1946 188912 1952 188924
rect 2004 188912 2010 188964
rect 1946 188680 1952 188692
rect 1412 188652 1952 188680
rect 1412 188408 1440 188652
rect 1946 188640 1952 188652
rect 2004 188640 2010 188692
rect 569954 188572 569960 188624
rect 570012 188612 570018 188624
rect 570230 188612 570236 188624
rect 570012 188584 570236 188612
rect 570012 188572 570018 188584
rect 570230 188572 570236 188584
rect 570288 188572 570294 188624
rect 1489 188547 1547 188553
rect 1489 188513 1501 188547
rect 1535 188544 1547 188547
rect 1946 188544 1952 188556
rect 1535 188516 1952 188544
rect 1535 188513 1547 188516
rect 1489 188507 1547 188513
rect 1946 188504 1952 188516
rect 2004 188504 2010 188556
rect 1489 188411 1547 188417
rect 1489 188408 1501 188411
rect 1412 188380 1501 188408
rect 1489 188377 1501 188380
rect 1535 188377 1547 188411
rect 1489 188371 1547 188377
rect 569954 188368 569960 188420
rect 570012 188408 570018 188420
rect 570049 188411 570107 188417
rect 570049 188408 570061 188411
rect 570012 188380 570061 188408
rect 570012 188368 570018 188380
rect 570049 188377 570061 188380
rect 570095 188377 570107 188411
rect 570049 188371 570107 188377
rect 1857 186507 1915 186513
rect 1857 186473 1869 186507
rect 1903 186504 1915 186507
rect 1946 186504 1952 186516
rect 1903 186476 1952 186504
rect 1903 186473 1915 186476
rect 1857 186467 1915 186473
rect 1946 186464 1952 186476
rect 2004 186464 2010 186516
rect 1210 182860 1216 182912
rect 1268 182900 1274 182912
rect 1673 182903 1731 182909
rect 1673 182900 1685 182903
rect 1268 182872 1685 182900
rect 1268 182860 1274 182872
rect 1673 182869 1685 182872
rect 1719 182869 1731 182903
rect 1673 182863 1731 182869
rect 290 182832 296 182844
rect 251 182804 296 182832
rect 290 182792 296 182804
rect 348 182792 354 182844
rect 569954 180412 569960 180464
rect 570012 180452 570018 180464
rect 570049 180455 570107 180461
rect 570049 180452 570061 180455
rect 570012 180424 570061 180452
rect 570012 180412 570018 180424
rect 570049 180421 570061 180424
rect 570095 180421 570107 180455
rect 570049 180415 570107 180421
rect 569954 179800 569960 179852
rect 570012 179840 570018 179852
rect 570141 179843 570199 179849
rect 570141 179840 570153 179843
rect 570012 179812 570153 179840
rect 570012 179800 570018 179812
rect 570141 179809 570153 179812
rect 570187 179809 570199 179843
rect 570141 179803 570199 179809
rect 1854 179636 1860 179648
rect 1815 179608 1860 179636
rect 1854 179596 1860 179608
rect 1912 179596 1918 179648
rect 477 179231 535 179237
rect 477 179197 489 179231
rect 523 179228 535 179231
rect 1949 179231 2007 179237
rect 1949 179228 1961 179231
rect 523 179200 1961 179228
rect 523 179197 535 179200
rect 477 179191 535 179197
rect 1949 179197 1961 179200
rect 1995 179197 2007 179231
rect 1949 179191 2007 179197
rect 1765 179095 1823 179101
rect 1765 179061 1777 179095
rect 1811 179092 1823 179095
rect 1854 179092 1860 179104
rect 1811 179064 1860 179092
rect 1811 179061 1823 179064
rect 1765 179055 1823 179061
rect 1854 179052 1860 179064
rect 1912 179052 1918 179104
rect 1762 178412 1768 178424
rect 1723 178384 1768 178412
rect 1762 178372 1768 178384
rect 1820 178372 1826 178424
rect 570141 178075 570199 178081
rect 570141 178041 570153 178075
rect 570187 178072 570199 178075
rect 570325 178075 570383 178081
rect 570325 178072 570337 178075
rect 570187 178044 570337 178072
rect 570187 178041 570199 178044
rect 570141 178035 570199 178041
rect 570325 178041 570337 178044
rect 570371 178041 570383 178075
rect 570325 178035 570383 178041
rect 569954 177692 569960 177744
rect 570012 177732 570018 177744
rect 570322 177732 570328 177744
rect 570012 177704 570328 177732
rect 570012 177692 570018 177704
rect 570322 177692 570328 177704
rect 570380 177692 570386 177744
rect 1946 177664 1952 177676
rect 1907 177636 1952 177664
rect 1946 177624 1952 177636
rect 2004 177624 2010 177676
rect 569957 177463 570015 177469
rect 569957 177429 569969 177463
rect 570003 177460 570015 177463
rect 570509 177463 570567 177469
rect 570509 177460 570521 177463
rect 570003 177432 570521 177460
rect 570003 177429 570015 177432
rect 569957 177423 570015 177429
rect 570509 177429 570521 177432
rect 570555 177429 570567 177463
rect 570509 177423 570567 177429
rect 569957 177327 570015 177333
rect 569957 177293 569969 177327
rect 570003 177324 570015 177327
rect 570138 177324 570144 177336
rect 570003 177296 570144 177324
rect 570003 177293 570015 177296
rect 569957 177287 570015 177293
rect 570138 177284 570144 177296
rect 570196 177284 570202 177336
rect 1673 176987 1731 176993
rect 1673 176953 1685 176987
rect 1719 176984 1731 176987
rect 1854 176984 1860 176996
rect 1719 176956 1860 176984
rect 1719 176953 1731 176956
rect 1673 176947 1731 176953
rect 1854 176944 1860 176956
rect 1912 176944 1918 176996
rect 569954 176808 569960 176860
rect 570012 176848 570018 176860
rect 570049 176851 570107 176857
rect 570049 176848 570061 176851
rect 570012 176820 570061 176848
rect 570012 176808 570018 176820
rect 570049 176817 570061 176820
rect 570095 176817 570107 176851
rect 570049 176811 570107 176817
rect 1489 176783 1547 176789
rect 1489 176749 1501 176783
rect 1535 176780 1547 176783
rect 1946 176780 1952 176792
rect 1535 176752 1952 176780
rect 1535 176749 1547 176752
rect 1489 176743 1547 176749
rect 1946 176740 1952 176752
rect 2004 176740 2010 176792
rect 1213 176647 1271 176653
rect 1213 176613 1225 176647
rect 1259 176644 1271 176647
rect 1946 176644 1952 176656
rect 1259 176616 1952 176644
rect 1259 176613 1271 176616
rect 1213 176607 1271 176613
rect 1946 176604 1952 176616
rect 2004 176604 2010 176656
rect 1305 176511 1363 176517
rect 1305 176477 1317 176511
rect 1351 176508 1363 176511
rect 1946 176508 1952 176520
rect 1351 176480 1952 176508
rect 1351 176477 1363 176480
rect 1305 176471 1363 176477
rect 1946 176468 1952 176480
rect 2004 176468 2010 176520
rect 1397 176375 1455 176381
rect 1397 176341 1409 176375
rect 1443 176372 1455 176375
rect 1946 176372 1952 176384
rect 1443 176344 1952 176372
rect 1443 176341 1455 176344
rect 1397 176335 1455 176341
rect 1946 176332 1952 176344
rect 2004 176332 2010 176384
rect 1762 176236 1768 176248
rect 1723 176208 1768 176236
rect 1762 176196 1768 176208
rect 1820 176196 1826 176248
rect 1946 176236 1952 176248
rect 1907 176208 1952 176236
rect 1946 176196 1952 176208
rect 2004 176196 2010 176248
rect 382 176060 388 176112
rect 440 176100 446 176112
rect 1857 176103 1915 176109
rect 1857 176100 1869 176103
rect 440 176072 1869 176100
rect 440 176060 446 176072
rect 1857 176069 1869 176072
rect 1903 176069 1915 176103
rect 1857 176063 1915 176069
rect 1581 175967 1639 175973
rect 1581 175933 1593 175967
rect 1627 175964 1639 175967
rect 1946 175964 1952 175976
rect 1627 175936 1952 175964
rect 1627 175933 1639 175936
rect 1581 175927 1639 175933
rect 1946 175924 1952 175936
rect 2004 175924 2010 175976
rect 1210 175584 1216 175636
rect 1268 175624 1274 175636
rect 1489 175627 1547 175633
rect 1489 175624 1501 175627
rect 1268 175596 1501 175624
rect 1268 175584 1274 175596
rect 1489 175593 1501 175596
rect 1535 175593 1547 175627
rect 1489 175587 1547 175593
rect 569954 175176 569960 175228
rect 570012 175216 570018 175228
rect 570233 175219 570291 175225
rect 570233 175216 570245 175219
rect 570012 175188 570245 175216
rect 570012 175176 570018 175188
rect 570233 175185 570245 175188
rect 570279 175185 570291 175219
rect 570233 175179 570291 175185
rect 569954 174944 569960 174956
rect 569915 174916 569960 174944
rect 569954 174904 569960 174916
rect 570012 174904 570018 174956
rect 198 174604 204 174616
rect 159 174576 204 174604
rect 198 174564 204 174576
rect 256 174564 262 174616
rect 198 174428 204 174480
rect 256 174468 262 174480
rect 1486 174468 1492 174480
rect 256 174440 1492 174468
rect 256 174428 262 174440
rect 1486 174428 1492 174440
rect 1544 174428 1550 174480
rect 569954 173612 569960 173664
rect 570012 173652 570018 173664
rect 570138 173652 570144 173664
rect 570012 173624 570144 173652
rect 570012 173612 570018 173624
rect 570138 173612 570144 173624
rect 570196 173612 570202 173664
rect 1486 173136 1492 173188
rect 1544 173176 1550 173188
rect 1854 173176 1860 173188
rect 1544 173148 1860 173176
rect 1544 173136 1550 173148
rect 1854 173136 1860 173148
rect 1912 173136 1918 173188
rect 1673 173043 1731 173049
rect 1673 173009 1685 173043
rect 1719 173040 1731 173043
rect 1854 173040 1860 173052
rect 1719 173012 1860 173040
rect 1719 173009 1731 173012
rect 1673 173003 1731 173009
rect 1854 173000 1860 173012
rect 1912 173000 1918 173052
rect 1210 171912 1216 171964
rect 1268 171952 1274 171964
rect 1394 171952 1400 171964
rect 1268 171924 1400 171952
rect 1268 171912 1274 171924
rect 1394 171912 1400 171924
rect 1452 171912 1458 171964
rect 570046 171912 570052 171964
rect 570104 171952 570110 171964
rect 570417 171955 570475 171961
rect 570417 171952 570429 171955
rect 570104 171924 570429 171952
rect 570104 171912 570110 171924
rect 570417 171921 570429 171924
rect 570463 171921 570475 171955
rect 570417 171915 570475 171921
rect 106 170960 112 171012
rect 164 171000 170 171012
rect 293 171003 351 171009
rect 293 171000 305 171003
rect 164 170972 305 171000
rect 164 170960 170 170972
rect 293 170969 305 170972
rect 339 170969 351 171003
rect 293 170963 351 170969
rect 474 170320 480 170332
rect 435 170292 480 170320
rect 474 170280 480 170292
rect 532 170280 538 170332
rect 569954 169328 569960 169380
rect 570012 169328 570018 169380
rect 569972 169176 570000 169328
rect 569954 169124 569960 169176
rect 570012 169124 570018 169176
rect 1946 169056 1952 169108
rect 2004 169096 2010 169108
rect 570049 169099 570107 169105
rect 2004 169068 2049 169096
rect 2004 169056 2010 169068
rect 570049 169065 570061 169099
rect 570095 169096 570107 169099
rect 570509 169099 570567 169105
rect 570509 169096 570521 169099
rect 570095 169068 570521 169096
rect 570095 169065 570107 169068
rect 570049 169059 570107 169065
rect 570509 169065 570521 169068
rect 570555 169065 570567 169099
rect 570509 169059 570567 169065
rect 569954 168988 569960 169040
rect 570012 169028 570018 169040
rect 570138 169028 570144 169040
rect 570012 169000 570144 169028
rect 570012 168988 570018 169000
rect 570138 168988 570144 169000
rect 570196 168988 570202 169040
rect 1581 168011 1639 168017
rect 1581 167977 1593 168011
rect 1627 168008 1639 168011
rect 1946 168008 1952 168020
rect 1627 167980 1952 168008
rect 1627 167977 1639 167980
rect 1581 167971 1639 167977
rect 1946 167968 1952 167980
rect 2004 167968 2010 168020
rect 293 167807 351 167813
rect 293 167773 305 167807
rect 339 167804 351 167807
rect 1946 167804 1952 167816
rect 339 167776 1952 167804
rect 339 167773 351 167776
rect 293 167767 351 167773
rect 1946 167764 1952 167776
rect 2004 167764 2010 167816
rect 382 167628 388 167680
rect 440 167668 446 167680
rect 937 167671 995 167677
rect 937 167668 949 167671
rect 440 167640 949 167668
rect 440 167628 446 167640
rect 937 167637 949 167640
rect 983 167637 995 167671
rect 937 167631 995 167637
rect 1213 167671 1271 167677
rect 1213 167637 1225 167671
rect 1259 167668 1271 167671
rect 1946 167668 1952 167680
rect 1259 167640 1952 167668
rect 1259 167637 1271 167640
rect 1213 167631 1271 167637
rect 1946 167628 1952 167640
rect 2004 167628 2010 167680
rect 1029 167399 1087 167405
rect 1029 167365 1041 167399
rect 1075 167396 1087 167399
rect 1946 167396 1952 167408
rect 1075 167368 1952 167396
rect 1075 167365 1087 167368
rect 1029 167359 1087 167365
rect 1946 167356 1952 167368
rect 2004 167356 2010 167408
rect 1026 167220 1032 167272
rect 1084 167260 1090 167272
rect 1305 167263 1363 167269
rect 1305 167260 1317 167263
rect 1084 167232 1317 167260
rect 1084 167220 1090 167232
rect 1305 167229 1317 167232
rect 1351 167229 1363 167263
rect 1305 167223 1363 167229
rect 1673 167263 1731 167269
rect 1673 167229 1685 167263
rect 1719 167260 1731 167263
rect 1946 167260 1952 167272
rect 1719 167232 1952 167260
rect 1719 167229 1731 167232
rect 1673 167223 1731 167229
rect 1946 167220 1952 167232
rect 2004 167220 2010 167272
rect 845 166923 903 166929
rect 845 166889 857 166923
rect 891 166920 903 166923
rect 1946 166920 1952 166932
rect 891 166892 1952 166920
rect 891 166889 903 166892
rect 845 166883 903 166889
rect 1946 166880 1952 166892
rect 2004 166880 2010 166932
rect 1026 166744 1032 166796
rect 1084 166784 1090 166796
rect 1946 166784 1952 166796
rect 1084 166756 1952 166784
rect 1084 166744 1090 166756
rect 1946 166744 1952 166756
rect 2004 166744 2010 166796
rect 1397 166447 1455 166453
rect 1397 166413 1409 166447
rect 1443 166444 1455 166447
rect 1946 166444 1952 166456
rect 1443 166416 1952 166444
rect 1443 166413 1455 166416
rect 1397 166407 1455 166413
rect 1946 166404 1952 166416
rect 2004 166404 2010 166456
rect 1946 166308 1952 166320
rect 1320 166280 1952 166308
rect 474 166132 480 166184
rect 532 166172 538 166184
rect 1121 166175 1179 166181
rect 1121 166172 1133 166175
rect 532 166144 1133 166172
rect 532 166132 538 166144
rect 1121 166141 1133 166144
rect 1167 166141 1179 166175
rect 1121 166135 1179 166141
rect 201 165903 259 165909
rect 201 165869 213 165903
rect 247 165900 259 165903
rect 382 165900 388 165912
rect 247 165872 388 165900
rect 247 165869 259 165872
rect 201 165863 259 165869
rect 382 165860 388 165872
rect 440 165860 446 165912
rect 1320 165900 1348 166280
rect 1946 166268 1952 166280
rect 2004 166268 2010 166320
rect 1394 165996 1400 166048
rect 1452 166036 1458 166048
rect 1946 166036 1952 166048
rect 1452 166008 1952 166036
rect 1452 165996 1458 166008
rect 1946 165996 1952 166008
rect 2004 165996 2010 166048
rect 1946 165900 1952 165912
rect 1320 165872 1952 165900
rect 1946 165860 1952 165872
rect 2004 165860 2010 165912
rect 1397 165495 1455 165501
rect 1397 165461 1409 165495
rect 1443 165492 1455 165495
rect 1946 165492 1952 165504
rect 1443 165464 1952 165492
rect 1443 165461 1455 165464
rect 1397 165455 1455 165461
rect 1946 165452 1952 165464
rect 2004 165452 2010 165504
rect 474 163888 480 163940
rect 532 163928 538 163940
rect 1486 163928 1492 163940
rect 532 163900 1492 163928
rect 532 163888 538 163900
rect 1486 163888 1492 163900
rect 1544 163888 1550 163940
rect 1026 163752 1032 163804
rect 1084 163792 1090 163804
rect 1486 163792 1492 163804
rect 1084 163764 1492 163792
rect 1084 163752 1090 163764
rect 1486 163752 1492 163764
rect 1544 163752 1550 163804
rect 569954 163724 569960 163736
rect 569915 163696 569960 163724
rect 569954 163684 569960 163696
rect 570012 163684 570018 163736
rect 1489 163591 1547 163597
rect 1489 163557 1501 163591
rect 1535 163588 1547 163591
rect 1857 163591 1915 163597
rect 1857 163588 1869 163591
rect 1535 163560 1869 163588
rect 1535 163557 1547 163560
rect 1489 163551 1547 163557
rect 1857 163557 1869 163560
rect 1903 163557 1915 163591
rect 1857 163551 1915 163557
rect 569954 163520 569960 163532
rect 569915 163492 569960 163520
rect 569954 163480 569960 163492
rect 570012 163480 570018 163532
rect 1581 163455 1639 163461
rect 1581 163421 1593 163455
rect 1627 163452 1639 163455
rect 1949 163455 2007 163461
rect 1949 163452 1961 163455
rect 1627 163424 1961 163452
rect 1627 163421 1639 163424
rect 1581 163415 1639 163421
rect 1949 163421 1961 163424
rect 1995 163421 2007 163455
rect 1949 163415 2007 163421
rect 750 163276 756 163328
rect 808 163316 814 163328
rect 1581 163319 1639 163325
rect 1581 163316 1593 163319
rect 808 163288 1593 163316
rect 808 163276 814 163288
rect 1581 163285 1593 163288
rect 1627 163285 1639 163319
rect 1581 163279 1639 163285
rect 570414 162228 570420 162240
rect 570375 162200 570420 162228
rect 570414 162188 570420 162200
rect 570472 162188 570478 162240
rect 570046 161984 570052 162036
rect 570104 162024 570110 162036
rect 570233 162027 570291 162033
rect 570233 162024 570245 162027
rect 570104 161996 570245 162024
rect 570104 161984 570110 161996
rect 570233 161993 570245 161996
rect 570279 161993 570291 162027
rect 570233 161987 570291 161993
rect 750 161576 756 161628
rect 808 161616 814 161628
rect 1302 161616 1308 161628
rect 808 161588 1308 161616
rect 808 161576 814 161588
rect 1302 161576 1308 161588
rect 1360 161576 1366 161628
rect 1486 160120 1492 160132
rect 1412 160092 1492 160120
rect 1412 159916 1440 160092
rect 1486 160080 1492 160092
rect 1544 160080 1550 160132
rect 1486 159944 1492 159996
rect 1544 159984 1550 159996
rect 1946 159984 1952 159996
rect 1544 159956 1952 159984
rect 1544 159944 1550 159956
rect 1946 159944 1952 159956
rect 2004 159944 2010 159996
rect 1412 159888 1992 159916
rect 1964 159860 1992 159888
rect 1946 159808 1952 159860
rect 2004 159808 2010 159860
rect 1486 159672 1492 159724
rect 1544 159712 1550 159724
rect 1946 159712 1952 159724
rect 1544 159684 1952 159712
rect 1544 159672 1550 159684
rect 1946 159672 1952 159684
rect 2004 159672 2010 159724
rect 753 159647 811 159653
rect 753 159613 765 159647
rect 799 159644 811 159647
rect 1673 159647 1731 159653
rect 1673 159644 1685 159647
rect 799 159616 1685 159644
rect 799 159613 811 159616
rect 753 159607 811 159613
rect 1673 159613 1685 159616
rect 1719 159613 1731 159647
rect 1673 159607 1731 159613
rect 1026 159536 1032 159588
rect 1084 159576 1090 159588
rect 1765 159579 1823 159585
rect 1765 159576 1777 159579
rect 1084 159548 1777 159576
rect 1084 159536 1090 159548
rect 1765 159545 1777 159548
rect 1811 159545 1823 159579
rect 1765 159539 1823 159545
rect 1489 159511 1547 159517
rect 1489 159477 1501 159511
rect 1535 159508 1547 159511
rect 1673 159511 1731 159517
rect 1673 159508 1685 159511
rect 1535 159480 1685 159508
rect 1535 159477 1547 159480
rect 1489 159471 1547 159477
rect 1673 159477 1685 159480
rect 1719 159477 1731 159511
rect 1673 159471 1731 159477
rect 1305 159443 1363 159449
rect 1305 159409 1317 159443
rect 1351 159440 1363 159443
rect 1765 159443 1823 159449
rect 1765 159440 1777 159443
rect 1351 159412 1777 159440
rect 1351 159409 1363 159412
rect 1305 159403 1363 159409
rect 1765 159409 1777 159412
rect 1811 159409 1823 159443
rect 1765 159403 1823 159409
rect 1397 159375 1455 159381
rect 1397 159341 1409 159375
rect 1443 159372 1455 159375
rect 1486 159372 1492 159384
rect 1443 159344 1492 159372
rect 1443 159341 1455 159344
rect 1397 159335 1455 159341
rect 1486 159332 1492 159344
rect 1544 159332 1550 159384
rect 845 159307 903 159313
rect 845 159273 857 159307
rect 891 159304 903 159307
rect 1946 159304 1952 159316
rect 891 159276 1952 159304
rect 891 159273 903 159276
rect 845 159267 903 159273
rect 1946 159264 1952 159276
rect 2004 159264 2010 159316
rect 1397 159239 1455 159245
rect 1397 159205 1409 159239
rect 1443 159236 1455 159239
rect 1857 159239 1915 159245
rect 1857 159236 1869 159239
rect 1443 159208 1869 159236
rect 1443 159205 1455 159208
rect 1397 159199 1455 159205
rect 1857 159205 1869 159208
rect 1903 159205 1915 159239
rect 1857 159199 1915 159205
rect 1029 159171 1087 159177
rect 1029 159137 1041 159171
rect 1075 159168 1087 159171
rect 1946 159168 1952 159180
rect 1075 159140 1952 159168
rect 1075 159137 1087 159140
rect 1029 159131 1087 159137
rect 1946 159128 1952 159140
rect 2004 159128 2010 159180
rect 750 159060 756 159112
rect 808 159100 814 159112
rect 1857 159103 1915 159109
rect 1857 159100 1869 159103
rect 808 159072 1869 159100
rect 808 159060 814 159072
rect 1857 159069 1869 159072
rect 1903 159069 1915 159103
rect 1857 159063 1915 159069
rect 569957 158763 570015 158769
rect 569957 158729 569969 158763
rect 570003 158760 570015 158763
rect 570325 158763 570383 158769
rect 570325 158760 570337 158763
rect 570003 158732 570337 158760
rect 570003 158729 570015 158732
rect 569957 158723 570015 158729
rect 570325 158729 570337 158732
rect 570371 158729 570383 158763
rect 570325 158723 570383 158729
rect 569957 158015 570015 158021
rect 569957 157981 569969 158015
rect 570003 158012 570015 158015
rect 570141 158015 570199 158021
rect 570141 158012 570153 158015
rect 570003 157984 570153 158012
rect 570003 157981 570015 157984
rect 569957 157975 570015 157981
rect 570141 157981 570153 157984
rect 570187 157981 570199 158015
rect 570141 157975 570199 157981
rect 569954 157836 569960 157888
rect 570012 157876 570018 157888
rect 570012 157848 570057 157876
rect 570012 157836 570018 157848
rect 570138 157632 570144 157684
rect 570196 157672 570202 157684
rect 570509 157675 570567 157681
rect 570509 157672 570521 157675
rect 570196 157644 570521 157672
rect 570196 157632 570202 157644
rect 570509 157641 570521 157644
rect 570555 157641 570567 157675
rect 570509 157635 570567 157641
rect 569954 157496 569960 157548
rect 570012 157536 570018 157548
rect 570138 157536 570144 157548
rect 570012 157508 570144 157536
rect 570012 157496 570018 157508
rect 570138 157496 570144 157508
rect 570196 157496 570202 157548
rect 569954 157360 569960 157412
rect 570012 157400 570018 157412
rect 570325 157403 570383 157409
rect 570325 157400 570337 157403
rect 570012 157372 570337 157400
rect 570012 157360 570018 157372
rect 570325 157369 570337 157372
rect 570371 157369 570383 157403
rect 570325 157363 570383 157369
rect 574922 157360 574928 157412
rect 574980 157400 574986 157412
rect 580166 157400 580172 157412
rect 574980 157372 580172 157400
rect 574980 157360 574986 157372
rect 580166 157360 580172 157372
rect 580224 157360 580230 157412
rect 1489 156383 1547 156389
rect 1489 156349 1501 156383
rect 1535 156380 1547 156383
rect 1578 156380 1584 156392
rect 1535 156352 1584 156380
rect 1535 156349 1547 156352
rect 1489 156343 1547 156349
rect 1578 156340 1584 156352
rect 1636 156340 1642 156392
rect 1394 156204 1400 156256
rect 1452 156244 1458 156256
rect 1578 156244 1584 156256
rect 1452 156216 1584 156244
rect 1452 156204 1458 156216
rect 1578 156204 1584 156216
rect 1636 156204 1642 156256
rect 569954 155864 569960 155916
rect 570012 155864 570018 155916
rect 569972 155768 570000 155864
rect 570230 155768 570236 155780
rect 569972 155740 570236 155768
rect 570230 155728 570236 155740
rect 570288 155728 570294 155780
rect 570046 155592 570052 155644
rect 570104 155632 570110 155644
rect 570325 155635 570383 155641
rect 570325 155632 570337 155635
rect 570104 155604 570337 155632
rect 570104 155592 570110 155604
rect 570325 155601 570337 155604
rect 570371 155601 570383 155635
rect 570325 155595 570383 155601
rect 474 155388 480 155440
rect 532 155428 538 155440
rect 1302 155428 1308 155440
rect 532 155400 1308 155428
rect 532 155388 538 155400
rect 1302 155388 1308 155400
rect 1360 155388 1366 155440
rect 569954 155184 569960 155236
rect 570012 155184 570018 155236
rect 569862 155116 569868 155168
rect 569920 155116 569926 155168
rect 569880 154884 569908 155116
rect 569972 155088 570000 155184
rect 570046 155088 570052 155100
rect 569972 155060 570052 155088
rect 570046 155048 570052 155060
rect 570104 155048 570110 155100
rect 569954 154980 569960 155032
rect 570012 155020 570018 155032
rect 570509 155023 570567 155029
rect 570509 155020 570521 155023
rect 570012 154992 570521 155020
rect 570012 154980 570018 154992
rect 570509 154989 570521 154992
rect 570555 154989 570567 155023
rect 570509 154983 570567 154989
rect 569954 154884 569960 154896
rect 569880 154856 569960 154884
rect 569954 154844 569960 154856
rect 570012 154844 570018 154896
rect 937 154819 995 154825
rect 937 154785 949 154819
rect 983 154816 995 154819
rect 1394 154816 1400 154828
rect 983 154788 1400 154816
rect 983 154785 995 154788
rect 937 154779 995 154785
rect 1394 154776 1400 154788
rect 1452 154776 1458 154828
rect 937 154071 995 154077
rect 937 154037 949 154071
rect 983 154068 995 154071
rect 1946 154068 1952 154080
rect 983 154040 1952 154068
rect 983 154037 995 154040
rect 937 154031 995 154037
rect 1946 154028 1952 154040
rect 2004 154028 2010 154080
rect 661 153935 719 153941
rect 661 153901 673 153935
rect 707 153932 719 153935
rect 1213 153935 1271 153941
rect 1213 153932 1225 153935
rect 707 153904 1225 153932
rect 707 153901 719 153904
rect 661 153895 719 153901
rect 1213 153901 1225 153904
rect 1259 153901 1271 153935
rect 1213 153895 1271 153901
rect 570046 153892 570052 153944
rect 570104 153932 570110 153944
rect 570325 153935 570383 153941
rect 570325 153932 570337 153935
rect 570104 153904 570337 153932
rect 570104 153892 570110 153904
rect 570325 153901 570337 153904
rect 570371 153901 570383 153935
rect 570325 153895 570383 153901
rect 382 153864 388 153876
rect 343 153836 388 153864
rect 382 153824 388 153836
rect 440 153824 446 153876
rect 569954 153824 569960 153876
rect 570012 153864 570018 153876
rect 570230 153864 570236 153876
rect 570012 153836 570236 153864
rect 570012 153824 570018 153836
rect 570230 153824 570236 153836
rect 570288 153824 570294 153876
rect 1213 153799 1271 153805
rect 1213 153765 1225 153799
rect 1259 153796 1271 153799
rect 1854 153796 1860 153808
rect 1259 153768 1860 153796
rect 1259 153765 1271 153768
rect 1213 153759 1271 153765
rect 1854 153756 1860 153768
rect 1912 153756 1918 153808
rect 570230 153456 570236 153468
rect 570191 153428 570236 153456
rect 570230 153416 570236 153428
rect 570288 153416 570294 153468
rect 106 151988 112 152040
rect 164 152028 170 152040
rect 382 152028 388 152040
rect 164 152000 388 152028
rect 164 151988 170 152000
rect 382 151988 388 152000
rect 440 151988 446 152040
rect 1029 150263 1087 150269
rect 1029 150229 1041 150263
rect 1075 150260 1087 150263
rect 1489 150263 1547 150269
rect 1489 150260 1501 150263
rect 1075 150232 1501 150260
rect 1075 150229 1087 150232
rect 1029 150223 1087 150229
rect 1489 150229 1501 150232
rect 1535 150229 1547 150263
rect 1489 150223 1547 150229
rect 937 150127 995 150133
rect 937 150093 949 150127
rect 983 150124 995 150127
rect 1489 150127 1547 150133
rect 1489 150124 1501 150127
rect 983 150096 1501 150124
rect 983 150093 995 150096
rect 937 150087 995 150093
rect 1489 150093 1501 150096
rect 1535 150093 1547 150127
rect 1489 150087 1547 150093
rect 570046 149540 570052 149592
rect 570104 149580 570110 149592
rect 570509 149583 570567 149589
rect 570509 149580 570521 149583
rect 570104 149552 570521 149580
rect 570104 149540 570110 149552
rect 570509 149549 570521 149552
rect 570555 149549 570567 149583
rect 570509 149543 570567 149549
rect 570046 149404 570052 149456
rect 570104 149444 570110 149456
rect 570322 149444 570328 149456
rect 570104 149416 570328 149444
rect 570104 149404 570110 149416
rect 570322 149404 570328 149416
rect 570380 149404 570386 149456
rect 569954 149268 569960 149320
rect 570012 149308 570018 149320
rect 570012 149280 570057 149308
rect 570012 149268 570018 149280
rect 570230 149064 570236 149116
rect 570288 149104 570294 149116
rect 570414 149104 570420 149116
rect 570288 149076 570420 149104
rect 570288 149064 570294 149076
rect 570414 149064 570420 149076
rect 570472 149064 570478 149116
rect 474 148724 480 148776
rect 532 148764 538 148776
rect 1581 148767 1639 148773
rect 1581 148764 1593 148767
rect 532 148736 1593 148764
rect 532 148724 538 148736
rect 1581 148733 1593 148736
rect 1627 148733 1639 148767
rect 1581 148727 1639 148733
rect 1394 148588 1400 148640
rect 1452 148628 1458 148640
rect 1673 148631 1731 148637
rect 1673 148628 1685 148631
rect 1452 148600 1685 148628
rect 1452 148588 1458 148600
rect 1673 148597 1685 148600
rect 1719 148597 1731 148631
rect 1673 148591 1731 148597
rect 569954 148452 569960 148504
rect 570012 148492 570018 148504
rect 570325 148495 570383 148501
rect 570325 148492 570337 148495
rect 570012 148464 570337 148492
rect 570012 148452 570018 148464
rect 570325 148461 570337 148464
rect 570371 148461 570383 148495
rect 570325 148455 570383 148461
rect 569957 148359 570015 148365
rect 569957 148325 569969 148359
rect 570003 148356 570015 148359
rect 570046 148356 570052 148368
rect 570003 148328 570052 148356
rect 570003 148325 570015 148328
rect 569957 148319 570015 148325
rect 570046 148316 570052 148328
rect 570104 148316 570110 148368
rect 569954 147908 569960 147960
rect 570012 147948 570018 147960
rect 570233 147951 570291 147957
rect 570233 147948 570245 147951
rect 570012 147920 570245 147948
rect 570012 147908 570018 147920
rect 570233 147917 570245 147920
rect 570279 147917 570291 147951
rect 570233 147911 570291 147917
rect 569954 147772 569960 147824
rect 570012 147812 570018 147824
rect 570138 147812 570144 147824
rect 570012 147784 570144 147812
rect 570012 147772 570018 147784
rect 570138 147772 570144 147784
rect 570196 147772 570202 147824
rect 569954 147636 569960 147688
rect 570012 147676 570018 147688
rect 570141 147679 570199 147685
rect 570141 147676 570153 147679
rect 570012 147648 570153 147676
rect 570012 147636 570018 147648
rect 570141 147645 570153 147648
rect 570187 147645 570199 147679
rect 570141 147639 570199 147645
rect 106 147092 112 147144
rect 164 147132 170 147144
rect 382 147132 388 147144
rect 164 147104 388 147132
rect 164 147092 170 147104
rect 382 147092 388 147104
rect 440 147092 446 147144
rect 1578 147092 1584 147144
rect 1636 147132 1642 147144
rect 1946 147132 1952 147144
rect 1636 147104 1952 147132
rect 1636 147092 1642 147104
rect 1946 147092 1952 147104
rect 2004 147092 2010 147144
rect 382 146996 388 147008
rect 343 146968 388 146996
rect 382 146956 388 146968
rect 440 146956 446 147008
rect 750 146996 756 147008
rect 711 146968 756 146996
rect 750 146956 756 146968
rect 808 146956 814 147008
rect 937 146999 995 147005
rect 937 146965 949 146999
rect 983 146996 995 146999
rect 1213 146999 1271 147005
rect 1213 146996 1225 146999
rect 983 146968 1225 146996
rect 983 146965 995 146968
rect 937 146959 995 146965
rect 1213 146965 1225 146968
rect 1259 146965 1271 146999
rect 1946 146996 1952 147008
rect 1907 146968 1952 146996
rect 1213 146959 1271 146965
rect 1946 146956 1952 146968
rect 2004 146956 2010 147008
rect 569954 146956 569960 147008
rect 570012 146996 570018 147008
rect 570509 146999 570567 147005
rect 570509 146996 570521 146999
rect 570012 146968 570521 146996
rect 570012 146956 570018 146968
rect 570509 146965 570521 146968
rect 570555 146965 570567 146999
rect 570509 146959 570567 146965
rect 1578 146344 1584 146396
rect 1636 146384 1642 146396
rect 1765 146387 1823 146393
rect 1765 146384 1777 146387
rect 1636 146356 1777 146384
rect 1636 146344 1642 146356
rect 1765 146353 1777 146356
rect 1811 146353 1823 146387
rect 1765 146347 1823 146353
rect 845 146319 903 146325
rect 845 146285 857 146319
rect 891 146316 903 146319
rect 1305 146319 1363 146325
rect 1305 146316 1317 146319
rect 891 146288 1317 146316
rect 891 146285 903 146288
rect 845 146279 903 146285
rect 1305 146285 1317 146288
rect 1351 146285 1363 146319
rect 1305 146279 1363 146285
rect 566 146208 572 146260
rect 624 146248 630 146260
rect 1765 146251 1823 146257
rect 1765 146248 1777 146251
rect 624 146220 1777 146248
rect 624 146208 630 146220
rect 1765 146217 1777 146220
rect 1811 146217 1823 146251
rect 1765 146211 1823 146217
rect 661 146183 719 146189
rect 661 146149 673 146183
rect 707 146180 719 146183
rect 1305 146183 1363 146189
rect 1305 146180 1317 146183
rect 707 146152 1317 146180
rect 707 146149 719 146152
rect 661 146143 719 146149
rect 1305 146149 1317 146152
rect 1351 146149 1363 146183
rect 1305 146143 1363 146149
rect 1210 145936 1216 145988
rect 1268 145976 1274 145988
rect 1581 145979 1639 145985
rect 1581 145976 1593 145979
rect 1268 145948 1593 145976
rect 1268 145936 1274 145948
rect 1581 145945 1593 145948
rect 1627 145945 1639 145979
rect 1581 145939 1639 145945
rect 1854 145908 1860 145920
rect 1815 145880 1860 145908
rect 1854 145868 1860 145880
rect 1912 145868 1918 145920
rect 1946 145800 1952 145852
rect 2004 145800 2010 145852
rect 1121 145707 1179 145713
rect 1121 145673 1133 145707
rect 1167 145704 1179 145707
rect 1854 145704 1860 145716
rect 1167 145676 1860 145704
rect 1167 145673 1179 145676
rect 1121 145667 1179 145673
rect 1854 145664 1860 145676
rect 1912 145664 1918 145716
rect 1964 145648 1992 145800
rect 290 145636 296 145648
rect 251 145608 296 145636
rect 290 145596 296 145608
rect 348 145596 354 145648
rect 1946 145596 1952 145648
rect 2004 145596 2010 145648
rect 569954 144236 569960 144288
rect 570012 144276 570018 144288
rect 570322 144276 570328 144288
rect 570012 144248 570328 144276
rect 570012 144236 570018 144248
rect 570322 144236 570328 144248
rect 570380 144236 570386 144288
rect 2774 143624 2780 143676
rect 2832 143664 2838 143676
rect 3142 143664 3148 143676
rect 2832 143636 3148 143664
rect 2832 143624 2838 143636
rect 3142 143624 3148 143636
rect 3200 143624 3206 143676
rect 1854 143120 1860 143132
rect 1815 143092 1860 143120
rect 1854 143080 1860 143092
rect 1912 143080 1918 143132
rect 569 142987 627 142993
rect 569 142953 581 142987
rect 615 142984 627 142987
rect 1026 142984 1032 142996
rect 615 142956 1032 142984
rect 615 142953 627 142956
rect 569 142947 627 142953
rect 1026 142944 1032 142956
rect 1084 142944 1090 142996
rect 1578 142944 1584 142996
rect 1636 142984 1642 142996
rect 1857 142987 1915 142993
rect 1857 142984 1869 142987
rect 1636 142956 1869 142984
rect 1636 142944 1642 142956
rect 1857 142953 1869 142956
rect 1903 142953 1915 142987
rect 1857 142947 1915 142953
rect 937 142851 995 142857
rect 937 142817 949 142851
rect 983 142848 995 142851
rect 1026 142848 1032 142860
rect 983 142820 1032 142848
rect 983 142817 995 142820
rect 937 142811 995 142817
rect 1026 142808 1032 142820
rect 1084 142808 1090 142860
rect 658 141856 664 141908
rect 716 141896 722 141908
rect 842 141896 848 141908
rect 716 141868 848 141896
rect 716 141856 722 141868
rect 842 141856 848 141868
rect 900 141856 906 141908
rect 566 141720 572 141772
rect 624 141760 630 141772
rect 842 141760 848 141772
rect 624 141732 848 141760
rect 624 141720 630 141732
rect 842 141720 848 141732
rect 900 141720 906 141772
rect 566 141624 572 141636
rect 527 141596 572 141624
rect 566 141584 572 141596
rect 624 141584 630 141636
rect 1486 141488 1492 141500
rect 1447 141460 1492 141488
rect 1486 141448 1492 141460
rect 1544 141448 1550 141500
rect 1489 141355 1547 141361
rect 1489 141321 1501 141355
rect 1535 141352 1547 141355
rect 1946 141352 1952 141364
rect 1535 141324 1952 141352
rect 1535 141321 1547 141324
rect 1489 141315 1547 141321
rect 1946 141312 1952 141324
rect 2004 141312 2010 141364
rect 1397 141287 1455 141293
rect 1397 141253 1409 141287
rect 1443 141284 1455 141287
rect 1854 141284 1860 141296
rect 1443 141256 1860 141284
rect 1443 141253 1455 141256
rect 1397 141247 1455 141253
rect 1854 141244 1860 141256
rect 1912 141244 1918 141296
rect 753 141219 811 141225
rect 753 141185 765 141219
rect 799 141216 811 141219
rect 1946 141216 1952 141228
rect 799 141188 1952 141216
rect 799 141185 811 141188
rect 753 141179 811 141185
rect 1946 141176 1952 141188
rect 2004 141176 2010 141228
rect 1029 141151 1087 141157
rect 1029 141117 1041 141151
rect 1075 141148 1087 141151
rect 1854 141148 1860 141160
rect 1075 141120 1860 141148
rect 1075 141117 1087 141120
rect 1029 141111 1087 141117
rect 1854 141108 1860 141120
rect 1912 141108 1918 141160
rect 1765 140743 1823 140749
rect 1765 140740 1777 140743
rect 860 140712 1777 140740
rect 860 140681 888 140712
rect 1765 140709 1777 140712
rect 1811 140709 1823 140743
rect 1765 140703 1823 140709
rect 845 140675 903 140681
rect 845 140641 857 140675
rect 891 140641 903 140675
rect 845 140635 903 140641
rect 1765 139995 1823 140001
rect 1765 139961 1777 139995
rect 1811 139992 1823 139995
rect 1946 139992 1952 140004
rect 1811 139964 1952 139992
rect 1811 139961 1823 139964
rect 1765 139955 1823 139961
rect 1946 139952 1952 139964
rect 2004 139952 2010 140004
rect 937 139111 995 139117
rect 937 139077 949 139111
rect 983 139108 995 139111
rect 1946 139108 1952 139120
rect 983 139080 1952 139108
rect 983 139077 995 139080
rect 937 139071 995 139077
rect 1946 139068 1952 139080
rect 2004 139068 2010 139120
rect 293 138975 351 138981
rect 293 138941 305 138975
rect 339 138972 351 138975
rect 1765 138975 1823 138981
rect 1765 138972 1777 138975
rect 339 138944 1777 138972
rect 339 138941 351 138944
rect 293 138935 351 138941
rect 1765 138941 1777 138944
rect 1811 138941 1823 138975
rect 1765 138935 1823 138941
rect 1121 138907 1179 138913
rect 1121 138873 1133 138907
rect 1167 138904 1179 138907
rect 1946 138904 1952 138916
rect 1167 138876 1952 138904
rect 1167 138873 1179 138876
rect 1121 138867 1179 138873
rect 1946 138864 1952 138876
rect 2004 138864 2010 138916
rect 1486 138796 1492 138848
rect 1544 138836 1550 138848
rect 1765 138839 1823 138845
rect 1765 138836 1777 138839
rect 1544 138808 1777 138836
rect 1544 138796 1550 138808
rect 1765 138805 1777 138808
rect 1811 138805 1823 138839
rect 1765 138799 1823 138805
rect 750 138728 756 138780
rect 808 138728 814 138780
rect 937 138771 995 138777
rect 937 138737 949 138771
rect 983 138768 995 138771
rect 1397 138771 1455 138777
rect 1397 138768 1409 138771
rect 983 138740 1409 138768
rect 983 138737 995 138740
rect 937 138731 995 138737
rect 1397 138737 1409 138740
rect 1443 138737 1455 138771
rect 1397 138731 1455 138737
rect 768 138632 796 138728
rect 1121 138703 1179 138709
rect 1121 138669 1133 138703
rect 1167 138700 1179 138703
rect 1302 138700 1308 138712
rect 1167 138672 1308 138700
rect 1167 138669 1179 138672
rect 1121 138663 1179 138669
rect 1302 138660 1308 138672
rect 1360 138660 1366 138712
rect 1397 138635 1455 138641
rect 1397 138632 1409 138635
rect 768 138604 1409 138632
rect 1397 138601 1409 138604
rect 1443 138601 1455 138635
rect 1397 138595 1455 138601
rect 1486 138592 1492 138644
rect 1544 138632 1550 138644
rect 1946 138632 1952 138644
rect 1544 138604 1952 138632
rect 1544 138592 1550 138604
rect 1946 138592 1952 138604
rect 2004 138592 2010 138644
rect 198 138524 204 138576
rect 256 138564 262 138576
rect 658 138564 664 138576
rect 256 138536 664 138564
rect 256 138524 262 138536
rect 658 138524 664 138536
rect 716 138524 722 138576
rect 1765 138295 1823 138301
rect 1765 138261 1777 138295
rect 1811 138292 1823 138295
rect 1946 138292 1952 138304
rect 1811 138264 1952 138292
rect 1811 138261 1823 138264
rect 1765 138255 1823 138261
rect 1946 138252 1952 138264
rect 2004 138252 2010 138304
rect 1489 137955 1547 137961
rect 1489 137921 1501 137955
rect 1535 137952 1547 137955
rect 1946 137952 1952 137964
rect 1535 137924 1952 137952
rect 1535 137921 1547 137924
rect 1489 137915 1547 137921
rect 1946 137912 1952 137924
rect 2004 137912 2010 137964
rect 569954 134920 569960 134972
rect 570012 134920 570018 134972
rect 569972 134768 570000 134920
rect 569954 134716 569960 134768
rect 570012 134716 570018 134768
rect 934 134648 940 134700
rect 992 134688 998 134700
rect 1394 134688 1400 134700
rect 992 134660 1400 134688
rect 992 134648 998 134660
rect 1394 134648 1400 134660
rect 1452 134648 1458 134700
rect 1489 134623 1547 134629
rect 1489 134589 1501 134623
rect 1535 134620 1547 134623
rect 1854 134620 1860 134632
rect 1535 134592 1860 134620
rect 1535 134589 1547 134592
rect 1489 134583 1547 134589
rect 1854 134580 1860 134592
rect 1912 134580 1918 134632
rect 937 134555 995 134561
rect 937 134521 949 134555
rect 983 134552 995 134555
rect 1026 134552 1032 134564
rect 983 134524 1032 134552
rect 983 134521 995 134524
rect 937 134515 995 134521
rect 1026 134512 1032 134524
rect 1084 134512 1090 134564
rect 1670 134552 1676 134564
rect 1631 134524 1676 134552
rect 1670 134512 1676 134524
rect 1728 134512 1734 134564
rect 569957 134555 570015 134561
rect 569957 134521 569969 134555
rect 570003 134552 570015 134555
rect 570046 134552 570052 134564
rect 570003 134524 570052 134552
rect 570003 134521 570015 134524
rect 569957 134515 570015 134521
rect 570046 134512 570052 134524
rect 570104 134512 570110 134564
rect 1213 134487 1271 134493
rect 1213 134453 1225 134487
rect 1259 134484 1271 134487
rect 1946 134484 1952 134496
rect 1259 134456 1952 134484
rect 1259 134453 1271 134456
rect 1213 134447 1271 134453
rect 1946 134444 1952 134456
rect 2004 134444 2010 134496
rect 934 134376 940 134428
rect 992 134416 998 134428
rect 1765 134419 1823 134425
rect 1765 134416 1777 134419
rect 992 134388 1777 134416
rect 992 134376 998 134388
rect 1765 134385 1777 134388
rect 1811 134385 1823 134419
rect 1765 134379 1823 134385
rect 569954 134308 569960 134360
rect 570012 134348 570018 134360
rect 570230 134348 570236 134360
rect 570012 134320 570236 134348
rect 570012 134308 570018 134320
rect 570230 134308 570236 134320
rect 570288 134308 570294 134360
rect 569954 134172 569960 134224
rect 570012 134212 570018 134224
rect 570049 134215 570107 134221
rect 570049 134212 570061 134215
rect 570012 134184 570061 134212
rect 570012 134172 570018 134184
rect 570049 134181 570061 134184
rect 570095 134181 570107 134215
rect 570049 134175 570107 134181
rect 1762 133464 1768 133476
rect 1723 133436 1768 133464
rect 1762 133424 1768 133436
rect 1820 133424 1826 133476
rect 1026 133288 1032 133340
rect 1084 133328 1090 133340
rect 1857 133331 1915 133337
rect 1857 133328 1869 133331
rect 1084 133300 1869 133328
rect 1084 133288 1090 133300
rect 1857 133297 1869 133300
rect 1903 133297 1915 133331
rect 1857 133291 1915 133297
rect 569954 133084 569960 133136
rect 570012 133124 570018 133136
rect 570325 133127 570383 133133
rect 570325 133124 570337 133127
rect 570012 133096 570337 133124
rect 570012 133084 570018 133096
rect 570325 133093 570337 133096
rect 570371 133093 570383 133127
rect 570325 133087 570383 133093
rect 661 132107 719 132113
rect 661 132073 673 132107
rect 707 132104 719 132107
rect 1946 132104 1952 132116
rect 707 132076 1952 132104
rect 707 132073 719 132076
rect 661 132067 719 132073
rect 1946 132064 1952 132076
rect 2004 132064 2010 132116
rect 1581 131155 1639 131161
rect 1581 131121 1593 131155
rect 1627 131152 1639 131155
rect 1627 131124 1900 131152
rect 1627 131121 1639 131124
rect 1581 131115 1639 131121
rect 1872 131084 1900 131124
rect 1949 131087 2007 131093
rect 1949 131084 1961 131087
rect 1872 131056 1961 131084
rect 1949 131053 1961 131056
rect 1995 131053 2007 131087
rect 1949 131047 2007 131053
rect 1581 130883 1639 130889
rect 1581 130849 1593 130883
rect 1627 130880 1639 130883
rect 1946 130880 1952 130892
rect 1627 130852 1952 130880
rect 1627 130849 1639 130852
rect 1581 130843 1639 130849
rect 1946 130840 1952 130852
rect 2004 130840 2010 130892
rect 569 130611 627 130617
rect 569 130577 581 130611
rect 615 130608 627 130611
rect 1946 130608 1952 130620
rect 615 130580 1952 130608
rect 615 130577 627 130580
rect 569 130571 627 130577
rect 1946 130568 1952 130580
rect 2004 130568 2010 130620
rect 477 130407 535 130413
rect 477 130373 489 130407
rect 523 130404 535 130407
rect 753 130407 811 130413
rect 753 130404 765 130407
rect 523 130376 765 130404
rect 523 130373 535 130376
rect 477 130367 535 130373
rect 753 130373 765 130376
rect 799 130373 811 130407
rect 753 130367 811 130373
rect 293 130271 351 130277
rect 293 130237 305 130271
rect 339 130268 351 130271
rect 753 130271 811 130277
rect 753 130268 765 130271
rect 339 130240 765 130268
rect 339 130237 351 130240
rect 293 130231 351 130237
rect 753 130237 765 130240
rect 799 130237 811 130271
rect 753 130231 811 130237
rect 477 129455 535 129461
rect 477 129421 489 129455
rect 523 129452 535 129455
rect 1946 129452 1952 129464
rect 523 129424 1952 129452
rect 523 129421 535 129424
rect 477 129415 535 129421
rect 1946 129412 1952 129424
rect 2004 129412 2010 129464
rect 1581 129183 1639 129189
rect 1581 129149 1593 129183
rect 1627 129180 1639 129183
rect 1946 129180 1952 129192
rect 1627 129152 1952 129180
rect 1627 129149 1639 129152
rect 1581 129143 1639 129149
rect 1946 129140 1952 129152
rect 2004 129140 2010 129192
rect 842 128868 848 128920
rect 900 128908 906 128920
rect 1581 128911 1639 128917
rect 1581 128908 1593 128911
rect 900 128880 1593 128908
rect 900 128868 906 128880
rect 1581 128877 1593 128880
rect 1627 128877 1639 128911
rect 1581 128871 1639 128877
rect 937 128367 995 128373
rect 937 128333 949 128367
rect 983 128364 995 128367
rect 1854 128364 1860 128376
rect 983 128336 1860 128364
rect 983 128333 995 128336
rect 937 128327 995 128333
rect 1854 128324 1860 128336
rect 1912 128324 1918 128376
rect 1029 126667 1087 126673
rect 1029 126633 1041 126667
rect 1075 126664 1087 126667
rect 1762 126664 1768 126676
rect 1075 126636 1768 126664
rect 1075 126633 1087 126636
rect 1029 126627 1087 126633
rect 1762 126624 1768 126636
rect 1820 126624 1826 126676
rect 1029 126531 1087 126537
rect 1029 126497 1041 126531
rect 1075 126528 1087 126531
rect 1581 126531 1639 126537
rect 1581 126528 1593 126531
rect 1075 126500 1593 126528
rect 1075 126497 1087 126500
rect 1029 126491 1087 126497
rect 1581 126497 1593 126500
rect 1627 126497 1639 126531
rect 1581 126491 1639 126497
rect 1581 126395 1639 126401
rect 1581 126361 1593 126395
rect 1627 126392 1639 126395
rect 1854 126392 1860 126404
rect 1627 126364 1860 126392
rect 1627 126361 1639 126364
rect 1581 126355 1639 126361
rect 1854 126352 1860 126364
rect 1912 126352 1918 126404
rect 382 126284 388 126336
rect 440 126324 446 126336
rect 842 126324 848 126336
rect 440 126296 848 126324
rect 440 126284 446 126296
rect 842 126284 848 126296
rect 900 126284 906 126336
rect 661 126259 719 126265
rect 661 126225 673 126259
rect 707 126256 719 126259
rect 937 126259 995 126265
rect 937 126256 949 126259
rect 707 126228 949 126256
rect 707 126225 719 126228
rect 661 126219 719 126225
rect 937 126225 949 126228
rect 983 126225 995 126259
rect 937 126219 995 126225
rect 1489 126259 1547 126265
rect 1489 126225 1501 126259
rect 1535 126256 1547 126259
rect 1578 126256 1584 126268
rect 1535 126228 1584 126256
rect 1535 126225 1547 126228
rect 1489 126219 1547 126225
rect 1578 126216 1584 126228
rect 1636 126216 1642 126268
rect 382 126080 388 126132
rect 440 126120 446 126132
rect 845 126123 903 126129
rect 845 126120 857 126123
rect 440 126092 857 126120
rect 440 126080 446 126092
rect 845 126089 857 126092
rect 891 126089 903 126123
rect 845 126083 903 126089
rect 1489 126123 1547 126129
rect 1489 126089 1501 126123
rect 1535 126120 1547 126123
rect 1946 126120 1952 126132
rect 1535 126092 1952 126120
rect 1535 126089 1547 126092
rect 1489 126083 1547 126089
rect 1946 126080 1952 126092
rect 2004 126080 2010 126132
rect 661 126055 719 126061
rect 661 126021 673 126055
rect 707 126052 719 126055
rect 1670 126052 1676 126064
rect 707 126024 1676 126052
rect 707 126021 719 126024
rect 661 126015 719 126021
rect 1670 126012 1676 126024
rect 1728 126012 1734 126064
rect 1854 124964 1860 124976
rect 1815 124936 1860 124964
rect 1854 124924 1860 124936
rect 1912 124924 1918 124976
rect 1946 124924 1952 124976
rect 2004 124964 2010 124976
rect 2004 124936 2049 124964
rect 2004 124924 2010 124936
rect 1670 124896 1676 124908
rect 1631 124868 1676 124896
rect 1670 124856 1676 124868
rect 1728 124856 1734 124908
rect 1394 124720 1400 124772
rect 1452 124760 1458 124772
rect 1673 124763 1731 124769
rect 1673 124760 1685 124763
rect 1452 124732 1685 124760
rect 1452 124720 1458 124732
rect 1673 124729 1685 124732
rect 1719 124729 1731 124763
rect 1673 124723 1731 124729
rect 1762 124720 1768 124772
rect 1820 124760 1826 124772
rect 1820 124732 1865 124760
rect 1820 124720 1826 124732
rect 750 124584 756 124636
rect 808 124624 814 124636
rect 1394 124624 1400 124636
rect 808 124596 1400 124624
rect 808 124584 814 124596
rect 1394 124584 1400 124596
rect 1452 124584 1458 124636
rect 572714 124040 572720 124092
rect 572772 124080 572778 124092
rect 574830 124080 574836 124092
rect 572772 124052 574836 124080
rect 572772 124040 572778 124052
rect 574830 124040 574836 124052
rect 574888 124040 574894 124092
rect 750 121184 756 121236
rect 808 121224 814 121236
rect 934 121224 940 121236
rect 808 121196 940 121224
rect 808 121184 814 121196
rect 934 121184 940 121196
rect 992 121184 998 121236
rect 934 121048 940 121100
rect 992 121088 998 121100
rect 1210 121088 1216 121100
rect 992 121060 1216 121088
rect 992 121048 998 121060
rect 1210 121048 1216 121060
rect 1268 121048 1274 121100
rect 1029 119595 1087 119601
rect 1029 119561 1041 119595
rect 1075 119592 1087 119595
rect 1765 119595 1823 119601
rect 1765 119592 1777 119595
rect 1075 119564 1777 119592
rect 1075 119561 1087 119564
rect 1029 119555 1087 119561
rect 1765 119561 1777 119564
rect 1811 119561 1823 119595
rect 1765 119555 1823 119561
rect 1946 118028 1952 118040
rect 1907 118000 1952 118028
rect 1946 117988 1952 118000
rect 2004 117988 2010 118040
rect 1857 117827 1915 117833
rect 1857 117793 1869 117827
rect 1903 117824 1915 117827
rect 1946 117824 1952 117836
rect 1903 117796 1952 117824
rect 1903 117793 1915 117796
rect 1857 117787 1915 117793
rect 1946 117784 1952 117796
rect 2004 117784 2010 117836
rect 1210 117512 1216 117564
rect 1268 117552 1274 117564
rect 1946 117552 1952 117564
rect 1268 117524 1952 117552
rect 1268 117512 1274 117524
rect 1946 117512 1952 117524
rect 2004 117512 2010 117564
rect 753 117487 811 117493
rect 753 117453 765 117487
rect 799 117484 811 117487
rect 1029 117487 1087 117493
rect 1029 117484 1041 117487
rect 799 117456 1041 117484
rect 799 117453 811 117456
rect 753 117447 811 117453
rect 1029 117453 1041 117456
rect 1075 117453 1087 117487
rect 1029 117447 1087 117453
rect 937 117419 995 117425
rect 937 117385 949 117419
rect 983 117416 995 117419
rect 1946 117416 1952 117428
rect 983 117388 1952 117416
rect 983 117385 995 117388
rect 937 117379 995 117385
rect 1946 117376 1952 117388
rect 2004 117376 2010 117428
rect 1302 116424 1308 116476
rect 1360 116464 1366 116476
rect 1489 116467 1547 116473
rect 1489 116464 1501 116467
rect 1360 116436 1501 116464
rect 1360 116424 1366 116436
rect 1489 116433 1501 116436
rect 1535 116433 1547 116467
rect 1489 116427 1547 116433
rect 1029 115243 1087 115249
rect 1029 115209 1041 115243
rect 1075 115240 1087 115243
rect 1489 115243 1547 115249
rect 1489 115240 1501 115243
rect 1075 115212 1501 115240
rect 1075 115209 1087 115212
rect 1029 115203 1087 115209
rect 1489 115209 1501 115212
rect 1535 115209 1547 115243
rect 1489 115203 1547 115209
rect 937 115107 995 115113
rect 937 115073 949 115107
rect 983 115104 995 115107
rect 1210 115104 1216 115116
rect 983 115076 1216 115104
rect 983 115073 995 115076
rect 937 115067 995 115073
rect 1210 115064 1216 115076
rect 1268 115064 1274 115116
rect 1029 111027 1087 111033
rect 1029 110993 1041 111027
rect 1075 111024 1087 111027
rect 1946 111024 1952 111036
rect 1075 110996 1952 111024
rect 1075 110993 1087 110996
rect 1029 110987 1087 110993
rect 1946 110984 1952 110996
rect 2004 110984 2010 111036
rect 574738 110440 574744 110492
rect 574796 110480 574802 110492
rect 580166 110480 580172 110492
rect 574796 110452 580172 110480
rect 574796 110440 574802 110452
rect 580166 110440 580172 110452
rect 580224 110440 580230 110492
rect 1210 110032 1216 110084
rect 1268 110072 1274 110084
rect 1946 110072 1952 110084
rect 1268 110044 1952 110072
rect 1268 110032 1274 110044
rect 1946 110032 1952 110044
rect 2004 110032 2010 110084
rect 753 109735 811 109741
rect 753 109701 765 109735
rect 799 109732 811 109735
rect 1946 109732 1952 109744
rect 799 109704 1952 109732
rect 799 109701 811 109704
rect 753 109695 811 109701
rect 1946 109692 1952 109704
rect 2004 109692 2010 109744
rect 661 109463 719 109469
rect 661 109429 673 109463
rect 707 109460 719 109463
rect 1946 109460 1952 109472
rect 707 109432 1952 109460
rect 707 109429 719 109432
rect 661 109423 719 109429
rect 1946 109420 1952 109432
rect 2004 109420 2010 109472
rect 569 109327 627 109333
rect 569 109293 581 109327
rect 615 109324 627 109327
rect 1946 109324 1952 109336
rect 615 109296 1952 109324
rect 615 109293 627 109296
rect 569 109287 627 109293
rect 1946 109284 1952 109296
rect 2004 109284 2010 109336
rect 661 109191 719 109197
rect 661 109157 673 109191
rect 707 109188 719 109191
rect 1946 109188 1952 109200
rect 707 109160 1952 109188
rect 707 109157 719 109160
rect 661 109151 719 109157
rect 1946 109148 1952 109160
rect 2004 109148 2010 109200
rect 937 108919 995 108925
rect 937 108885 949 108919
rect 983 108916 995 108919
rect 1946 108916 1952 108928
rect 983 108888 1952 108916
rect 983 108885 995 108888
rect 937 108879 995 108885
rect 1946 108876 1952 108888
rect 2004 108876 2010 108928
rect 753 108783 811 108789
rect 753 108749 765 108783
rect 799 108780 811 108783
rect 1946 108780 1952 108792
rect 799 108752 1952 108780
rect 799 108749 811 108752
rect 753 108743 811 108749
rect 1946 108740 1952 108752
rect 2004 108740 2010 108792
rect 1581 108647 1639 108653
rect 1581 108613 1593 108647
rect 1627 108644 1639 108647
rect 1946 108644 1952 108656
rect 1627 108616 1952 108644
rect 1627 108613 1639 108616
rect 1581 108607 1639 108613
rect 1946 108604 1952 108616
rect 2004 108604 2010 108656
rect 1489 108511 1547 108517
rect 1489 108477 1501 108511
rect 1535 108508 1547 108511
rect 1946 108508 1952 108520
rect 1535 108480 1952 108508
rect 1535 108477 1547 108480
rect 1489 108471 1547 108477
rect 1946 108468 1952 108480
rect 2004 108468 2010 108520
rect 1213 108375 1271 108381
rect 1213 108341 1225 108375
rect 1259 108372 1271 108375
rect 1946 108372 1952 108384
rect 1259 108344 1952 108372
rect 1259 108341 1271 108344
rect 1213 108335 1271 108341
rect 1946 108332 1952 108344
rect 2004 108332 2010 108384
rect 1029 108103 1087 108109
rect 1029 108069 1041 108103
rect 1075 108100 1087 108103
rect 1210 108100 1216 108112
rect 1075 108072 1216 108100
rect 1075 108069 1087 108072
rect 1029 108063 1087 108069
rect 1210 108060 1216 108072
rect 1268 108060 1274 108112
rect 1673 108103 1731 108109
rect 1673 108069 1685 108103
rect 1719 108100 1731 108103
rect 1946 108100 1952 108112
rect 1719 108072 1952 108100
rect 1719 108069 1731 108072
rect 1673 108063 1731 108069
rect 1946 108060 1952 108072
rect 2004 108060 2010 108112
rect 845 107695 903 107701
rect 845 107661 857 107695
rect 891 107692 903 107695
rect 1946 107692 1952 107704
rect 891 107664 1952 107692
rect 891 107661 903 107664
rect 845 107655 903 107661
rect 1946 107652 1952 107664
rect 2004 107652 2010 107704
rect 1302 107312 1308 107364
rect 1360 107352 1366 107364
rect 1946 107352 1952 107364
rect 1360 107324 1952 107352
rect 1360 107312 1366 107324
rect 1946 107312 1952 107324
rect 2004 107312 2010 107364
rect 1305 107219 1363 107225
rect 1305 107185 1317 107219
rect 1351 107216 1363 107219
rect 1946 107216 1952 107228
rect 1351 107188 1952 107216
rect 1351 107185 1363 107188
rect 1305 107179 1363 107185
rect 1946 107176 1952 107188
rect 2004 107176 2010 107228
rect 1946 107080 1952 107092
rect 1907 107052 1952 107080
rect 1946 107040 1952 107052
rect 2004 107040 2010 107092
rect 1210 102552 1216 102604
rect 1268 102592 1274 102604
rect 1765 102595 1823 102601
rect 1765 102592 1777 102595
rect 1268 102564 1777 102592
rect 1268 102552 1274 102564
rect 1765 102561 1777 102564
rect 1811 102561 1823 102595
rect 1765 102555 1823 102561
rect 1765 98447 1823 98453
rect 1765 98413 1777 98447
rect 1811 98444 1823 98447
rect 1946 98444 1952 98456
rect 1811 98416 1952 98444
rect 1811 98413 1823 98416
rect 1765 98407 1823 98413
rect 1946 98404 1952 98416
rect 2004 98404 2010 98456
rect 1302 98308 1308 98320
rect 1263 98280 1308 98308
rect 1302 98268 1308 98280
rect 1360 98268 1366 98320
rect 1673 98311 1731 98317
rect 1673 98277 1685 98311
rect 1719 98308 1731 98311
rect 1946 98308 1952 98320
rect 1719 98280 1952 98308
rect 1719 98277 1731 98280
rect 1673 98271 1731 98277
rect 1946 98268 1952 98280
rect 2004 98268 2010 98320
rect 382 98132 388 98184
rect 440 98172 446 98184
rect 1302 98172 1308 98184
rect 440 98144 1308 98172
rect 440 98132 446 98144
rect 1302 98132 1308 98144
rect 1360 98132 1366 98184
rect 1946 98172 1952 98184
rect 1907 98144 1952 98172
rect 1946 98132 1952 98144
rect 2004 98132 2010 98184
rect 572714 96500 572720 96552
rect 572772 96540 572778 96552
rect 574922 96540 574928 96552
rect 572772 96512 574928 96540
rect 572772 96500 572778 96512
rect 574922 96500 574928 96512
rect 574980 96500 574986 96552
rect 474 96228 480 96280
rect 532 96268 538 96280
rect 1857 96271 1915 96277
rect 1857 96268 1869 96271
rect 532 96240 1869 96268
rect 532 96228 538 96240
rect 1857 96237 1869 96240
rect 1903 96237 1915 96271
rect 1857 96231 1915 96237
rect 1121 96067 1179 96073
rect 1121 96033 1133 96067
rect 1167 96064 1179 96067
rect 1581 96067 1639 96073
rect 1581 96064 1593 96067
rect 1167 96036 1593 96064
rect 1167 96033 1179 96036
rect 1121 96027 1179 96033
rect 1581 96033 1593 96036
rect 1627 96033 1639 96067
rect 1581 96027 1639 96033
rect 1854 94772 1860 94784
rect 1815 94744 1860 94772
rect 1854 94732 1860 94744
rect 1912 94732 1918 94784
rect 1029 94707 1087 94713
rect 1029 94673 1041 94707
rect 1075 94704 1087 94707
rect 1946 94704 1952 94716
rect 1075 94676 1952 94704
rect 1075 94673 1087 94676
rect 1029 94667 1087 94673
rect 1946 94664 1952 94676
rect 2004 94664 2010 94716
rect 1121 94027 1179 94033
rect 1121 93993 1133 94027
rect 1167 94024 1179 94027
rect 1946 94024 1952 94036
rect 1167 93996 1952 94024
rect 1167 93993 1179 93996
rect 1121 93987 1179 93993
rect 1946 93984 1952 93996
rect 2004 93984 2010 94036
rect 1213 93619 1271 93625
rect 1213 93585 1225 93619
rect 1259 93616 1271 93619
rect 1946 93616 1952 93628
rect 1259 93588 1952 93616
rect 1259 93585 1271 93588
rect 1213 93579 1271 93585
rect 1946 93576 1952 93588
rect 2004 93576 2010 93628
rect 1305 93551 1363 93557
rect 1305 93517 1317 93551
rect 1351 93548 1363 93551
rect 1489 93551 1547 93557
rect 1489 93548 1501 93551
rect 1351 93520 1501 93548
rect 1351 93517 1363 93520
rect 1305 93511 1363 93517
rect 1489 93517 1501 93520
rect 1535 93517 1547 93551
rect 1489 93511 1547 93517
rect 1854 93480 1860 93492
rect 1228 93452 1860 93480
rect 1228 93344 1256 93452
rect 1854 93440 1860 93452
rect 1912 93440 1918 93492
rect 1305 93415 1363 93421
rect 1305 93381 1317 93415
rect 1351 93412 1363 93415
rect 1946 93412 1952 93424
rect 1351 93384 1952 93412
rect 1351 93381 1363 93384
rect 1305 93375 1363 93381
rect 1946 93372 1952 93384
rect 2004 93372 2010 93424
rect 1228 93316 1992 93344
rect 1964 93288 1992 93316
rect 1854 93276 1860 93288
rect 1815 93248 1860 93276
rect 1854 93236 1860 93248
rect 1912 93236 1918 93288
rect 1946 93236 1952 93288
rect 2004 93236 2010 93288
rect 566 93100 572 93152
rect 624 93140 630 93152
rect 1857 93143 1915 93149
rect 1857 93140 1869 93143
rect 624 93112 1869 93140
rect 624 93100 630 93112
rect 1857 93109 1869 93112
rect 1903 93109 1915 93143
rect 1857 93103 1915 93109
rect 1946 92188 1952 92200
rect 860 92160 1952 92188
rect 860 91916 888 92160
rect 1946 92148 1952 92160
rect 2004 92148 2010 92200
rect 937 92055 995 92061
rect 937 92021 949 92055
rect 983 92052 995 92055
rect 1946 92052 1952 92064
rect 983 92024 1952 92052
rect 983 92021 995 92024
rect 937 92015 995 92021
rect 1946 92012 1952 92024
rect 2004 92012 2010 92064
rect 1946 91916 1952 91928
rect 860 91888 1952 91916
rect 1946 91876 1952 91888
rect 2004 91876 2010 91928
rect 1213 91783 1271 91789
rect 1213 91749 1225 91783
rect 1259 91780 1271 91783
rect 1946 91780 1952 91792
rect 1259 91752 1952 91780
rect 1259 91749 1271 91752
rect 1213 91743 1271 91749
rect 1946 91740 1952 91752
rect 2004 91740 2010 91792
rect 1121 91647 1179 91653
rect 1121 91613 1133 91647
rect 1167 91644 1179 91647
rect 1946 91644 1952 91656
rect 1167 91616 1952 91644
rect 1167 91613 1179 91616
rect 1121 91607 1179 91613
rect 1946 91604 1952 91616
rect 2004 91604 2010 91656
rect 1305 91511 1363 91517
rect 1305 91477 1317 91511
rect 1351 91508 1363 91511
rect 1946 91508 1952 91520
rect 1351 91480 1952 91508
rect 1351 91477 1363 91480
rect 1305 91471 1363 91477
rect 1946 91468 1952 91480
rect 2004 91468 2010 91520
rect 1397 91375 1455 91381
rect 1397 91341 1409 91375
rect 1443 91372 1455 91375
rect 1946 91372 1952 91384
rect 1443 91344 1952 91372
rect 1443 91341 1455 91344
rect 1397 91335 1455 91341
rect 1946 91332 1952 91344
rect 2004 91332 2010 91384
rect 1765 91239 1823 91245
rect 1765 91205 1777 91239
rect 1811 91236 1823 91239
rect 1946 91236 1952 91248
rect 1811 91208 1952 91236
rect 1811 91205 1823 91208
rect 1765 91199 1823 91205
rect 1946 91196 1952 91208
rect 2004 91196 2010 91248
rect 1029 90423 1087 90429
rect 1029 90389 1041 90423
rect 1075 90420 1087 90423
rect 1397 90423 1455 90429
rect 1397 90420 1409 90423
rect 1075 90392 1409 90420
rect 1075 90389 1087 90392
rect 1029 90383 1087 90389
rect 1397 90389 1409 90392
rect 1443 90389 1455 90423
rect 1397 90383 1455 90389
rect 1213 88791 1271 88797
rect 1213 88757 1225 88791
rect 1259 88788 1271 88791
rect 1949 88791 2007 88797
rect 1949 88788 1961 88791
rect 1259 88760 1961 88788
rect 1259 88757 1271 88760
rect 1213 88751 1271 88757
rect 1949 88757 1961 88760
rect 1995 88757 2007 88791
rect 1949 88751 2007 88757
rect 1029 87635 1087 87641
rect 1029 87601 1041 87635
rect 1075 87632 1087 87635
rect 1489 87635 1547 87641
rect 1489 87632 1501 87635
rect 1075 87604 1501 87632
rect 1075 87601 1087 87604
rect 1029 87595 1087 87601
rect 1489 87601 1501 87604
rect 1535 87601 1547 87635
rect 1489 87595 1547 87601
rect 1489 87363 1547 87369
rect 1489 87329 1501 87363
rect 1535 87360 1547 87363
rect 1673 87363 1731 87369
rect 1673 87360 1685 87363
rect 1535 87332 1685 87360
rect 1535 87329 1547 87332
rect 1489 87323 1547 87329
rect 1673 87329 1685 87332
rect 1719 87329 1731 87363
rect 1673 87323 1731 87329
rect 1946 86408 1952 86420
rect 1907 86380 1952 86408
rect 1946 86368 1952 86380
rect 2004 86368 2010 86420
rect 1673 86343 1731 86349
rect 1673 86309 1685 86343
rect 1719 86340 1731 86343
rect 1854 86340 1860 86352
rect 1719 86312 1860 86340
rect 1719 86309 1731 86312
rect 1673 86303 1731 86309
rect 1854 86300 1860 86312
rect 1912 86300 1918 86352
rect 1765 86207 1823 86213
rect 1765 86173 1777 86207
rect 1811 86204 1823 86207
rect 1946 86204 1952 86216
rect 1811 86176 1952 86204
rect 1811 86173 1823 86176
rect 1765 86167 1823 86173
rect 1946 86164 1952 86176
rect 2004 86164 2010 86216
rect 937 86139 995 86145
rect 937 86105 949 86139
rect 983 86136 995 86139
rect 1854 86136 1860 86148
rect 983 86108 1860 86136
rect 983 86105 995 86108
rect 937 86099 995 86105
rect 1854 86096 1860 86108
rect 1912 86096 1918 86148
rect 937 84779 995 84785
rect 937 84745 949 84779
rect 983 84776 995 84779
rect 1946 84776 1952 84788
rect 983 84748 1952 84776
rect 983 84745 995 84748
rect 937 84739 995 84745
rect 1946 84736 1952 84748
rect 2004 84736 2010 84788
rect 1121 84643 1179 84649
rect 1121 84609 1133 84643
rect 1167 84640 1179 84643
rect 1946 84640 1952 84652
rect 1167 84612 1952 84640
rect 1167 84609 1179 84612
rect 1121 84603 1179 84609
rect 1946 84600 1952 84612
rect 2004 84600 2010 84652
rect 1305 83827 1363 83833
rect 1305 83793 1317 83827
rect 1351 83824 1363 83827
rect 1946 83824 1952 83836
rect 1351 83796 1952 83824
rect 1351 83793 1363 83796
rect 1305 83787 1363 83793
rect 1946 83784 1952 83796
rect 2004 83784 2010 83836
rect 1029 83623 1087 83629
rect 1029 83589 1041 83623
rect 1075 83620 1087 83623
rect 1946 83620 1952 83632
rect 1075 83592 1952 83620
rect 1075 83589 1087 83592
rect 1029 83583 1087 83589
rect 1946 83580 1952 83592
rect 2004 83580 2010 83632
rect 1302 83444 1308 83496
rect 1360 83484 1366 83496
rect 1854 83484 1860 83496
rect 1360 83456 1860 83484
rect 1360 83444 1366 83456
rect 1854 83444 1860 83456
rect 1912 83444 1918 83496
rect 937 82127 995 82133
rect 937 82093 949 82127
rect 983 82124 995 82127
rect 1946 82124 1952 82136
rect 983 82096 1952 82124
rect 983 82093 995 82096
rect 937 82087 995 82093
rect 1946 82084 1952 82096
rect 2004 82084 2010 82136
rect 566 80928 572 80980
rect 624 80968 630 80980
rect 1673 80971 1731 80977
rect 1673 80968 1685 80971
rect 624 80940 1685 80968
rect 624 80928 630 80940
rect 1673 80937 1685 80940
rect 1719 80937 1731 80971
rect 1673 80931 1731 80937
rect 1489 80835 1547 80841
rect 1489 80801 1501 80835
rect 1535 80832 1547 80835
rect 1673 80835 1731 80841
rect 1673 80832 1685 80835
rect 1535 80804 1685 80832
rect 1535 80801 1547 80804
rect 1489 80795 1547 80801
rect 1673 80801 1685 80804
rect 1719 80801 1731 80835
rect 1673 80795 1731 80801
rect 1305 80767 1363 80773
rect 1305 80733 1317 80767
rect 1351 80764 1363 80767
rect 1946 80764 1952 80776
rect 1351 80736 1952 80764
rect 1351 80733 1363 80736
rect 1305 80727 1363 80733
rect 1946 80724 1952 80736
rect 2004 80724 2010 80776
rect 1213 80699 1271 80705
rect 1213 80665 1225 80699
rect 1259 80696 1271 80699
rect 1489 80699 1547 80705
rect 1489 80696 1501 80699
rect 1259 80668 1501 80696
rect 1259 80665 1271 80668
rect 1213 80659 1271 80665
rect 1489 80665 1501 80668
rect 1535 80665 1547 80699
rect 1489 80659 1547 80665
rect 569954 77256 569960 77308
rect 570012 77296 570018 77308
rect 570049 77299 570107 77305
rect 570049 77296 570061 77299
rect 570012 77268 570061 77296
rect 570012 77256 570018 77268
rect 570049 77265 570061 77268
rect 570095 77265 570107 77299
rect 570049 77259 570107 77265
rect 569954 76712 569960 76764
rect 570012 76752 570018 76764
rect 570141 76755 570199 76761
rect 570141 76752 570153 76755
rect 570012 76724 570153 76752
rect 570012 76712 570018 76724
rect 570141 76721 570153 76724
rect 570187 76721 570199 76755
rect 570141 76715 570199 76721
rect 569954 76576 569960 76628
rect 570012 76616 570018 76628
rect 570233 76619 570291 76625
rect 570233 76616 570245 76619
rect 570012 76588 570245 76616
rect 570012 76576 570018 76588
rect 570233 76585 570245 76588
rect 570279 76585 570291 76619
rect 570233 76579 570291 76585
rect 569954 76440 569960 76492
rect 570012 76480 570018 76492
rect 570138 76480 570144 76492
rect 570012 76452 570144 76480
rect 570012 76440 570018 76452
rect 570138 76440 570144 76452
rect 570196 76440 570202 76492
rect 569954 76344 569960 76356
rect 569915 76316 569960 76344
rect 569954 76304 569960 76316
rect 570012 76304 570018 76356
rect 569954 76168 569960 76220
rect 570012 76208 570018 76220
rect 570325 76211 570383 76217
rect 570325 76208 570337 76211
rect 570012 76180 570337 76208
rect 570012 76168 570018 76180
rect 570325 76177 570337 76180
rect 570371 76177 570383 76211
rect 570325 76171 570383 76177
rect 569957 75939 570015 75945
rect 569957 75905 569969 75939
rect 570003 75936 570015 75939
rect 570233 75939 570291 75945
rect 570233 75936 570245 75939
rect 570003 75908 570245 75936
rect 570003 75905 570015 75908
rect 569957 75899 570015 75905
rect 570233 75905 570245 75908
rect 570279 75905 570291 75939
rect 570233 75899 570291 75905
rect 569954 74808 569960 74860
rect 570012 74848 570018 74860
rect 570325 74851 570383 74857
rect 570325 74848 570337 74851
rect 570012 74820 570337 74848
rect 570012 74808 570018 74820
rect 570325 74817 570337 74820
rect 570371 74817 570383 74851
rect 570325 74811 570383 74817
rect 569954 74672 569960 74724
rect 570012 74712 570018 74724
rect 570230 74712 570236 74724
rect 570012 74684 570236 74712
rect 570012 74672 570018 74684
rect 570230 74672 570236 74684
rect 570288 74672 570294 74724
rect 569954 73760 569960 73772
rect 569880 73732 569960 73760
rect 569880 73148 569908 73732
rect 569954 73720 569960 73732
rect 570012 73720 570018 73772
rect 569954 73584 569960 73636
rect 570012 73624 570018 73636
rect 570417 73627 570475 73633
rect 570417 73624 570429 73627
rect 570012 73596 570429 73624
rect 570012 73584 570018 73596
rect 570417 73593 570429 73596
rect 570463 73593 570475 73627
rect 570417 73587 570475 73593
rect 569954 73380 569960 73432
rect 570012 73420 570018 73432
rect 570509 73423 570567 73429
rect 570509 73420 570521 73423
rect 570012 73392 570521 73420
rect 570012 73380 570018 73392
rect 570509 73389 570521 73392
rect 570555 73389 570567 73423
rect 570509 73383 570567 73389
rect 569954 73244 569960 73296
rect 570012 73284 570018 73296
rect 570230 73284 570236 73296
rect 570012 73256 570236 73284
rect 570012 73244 570018 73256
rect 570230 73244 570236 73256
rect 570288 73244 570294 73296
rect 569954 73148 569960 73160
rect 569880 73120 569960 73148
rect 569954 73108 569960 73120
rect 570012 73108 570018 73160
rect 569954 72972 569960 73024
rect 570012 73012 570018 73024
rect 570417 73015 570475 73021
rect 570417 73012 570429 73015
rect 570012 72984 570429 73012
rect 570012 72972 570018 72984
rect 570417 72981 570429 72984
rect 570463 72981 570475 73015
rect 570417 72975 570475 72981
rect 566 72564 572 72616
rect 624 72604 630 72616
rect 1854 72604 1860 72616
rect 624 72576 1860 72604
rect 624 72564 630 72576
rect 1854 72564 1860 72576
rect 1912 72564 1918 72616
rect 1854 72468 1860 72480
rect 1815 72440 1860 72468
rect 1854 72428 1860 72440
rect 1912 72428 1918 72480
rect 569954 72428 569960 72480
rect 570012 72468 570018 72480
rect 570325 72471 570383 72477
rect 570325 72468 570337 72471
rect 570012 72440 570337 72468
rect 570012 72428 570018 72440
rect 570325 72437 570337 72440
rect 570371 72437 570383 72471
rect 570325 72431 570383 72437
rect 1581 72335 1639 72341
rect 1581 72301 1593 72335
rect 1627 72332 1639 72335
rect 1765 72335 1823 72341
rect 1765 72332 1777 72335
rect 1627 72304 1777 72332
rect 1627 72301 1639 72304
rect 1581 72295 1639 72301
rect 1765 72301 1777 72304
rect 1811 72301 1823 72335
rect 1765 72295 1823 72301
rect 1302 72156 1308 72208
rect 1360 72196 1366 72208
rect 1946 72196 1952 72208
rect 1360 72168 1952 72196
rect 1360 72156 1366 72168
rect 1946 72156 1952 72168
rect 2004 72156 2010 72208
rect 1581 71995 1639 72001
rect 1581 71961 1593 71995
rect 1627 71992 1639 71995
rect 1946 71992 1952 72004
rect 1627 71964 1952 71992
rect 1627 71961 1639 71964
rect 1581 71955 1639 71961
rect 1946 71952 1952 71964
rect 2004 71952 2010 72004
rect 1210 71000 1216 71052
rect 1268 71040 1274 71052
rect 1946 71040 1952 71052
rect 1268 71012 1952 71040
rect 1268 71000 1274 71012
rect 1946 71000 1952 71012
rect 2004 71000 2010 71052
rect 1121 70431 1179 70437
rect 1121 70397 1133 70431
rect 1167 70397 1179 70431
rect 1121 70391 1179 70397
rect 1136 70292 1164 70391
rect 1305 70295 1363 70301
rect 1305 70292 1317 70295
rect 1136 70264 1317 70292
rect 1305 70261 1317 70264
rect 1351 70261 1363 70295
rect 1305 70255 1363 70261
rect 1213 69615 1271 69621
rect 1213 69581 1225 69615
rect 1259 69612 1271 69615
rect 1673 69615 1731 69621
rect 1673 69612 1685 69615
rect 1259 69584 1685 69612
rect 1259 69581 1271 69584
rect 1213 69575 1271 69581
rect 1673 69581 1685 69584
rect 1719 69581 1731 69615
rect 1673 69575 1731 69581
rect 1397 69479 1455 69485
rect 1397 69445 1409 69479
rect 1443 69476 1455 69479
rect 1673 69479 1731 69485
rect 1673 69476 1685 69479
rect 1443 69448 1685 69476
rect 1443 69445 1455 69448
rect 1397 69439 1455 69445
rect 1673 69445 1685 69448
rect 1719 69445 1731 69479
rect 1673 69439 1731 69445
rect 1302 69300 1308 69352
rect 1360 69340 1366 69352
rect 1397 69343 1455 69349
rect 1397 69340 1409 69343
rect 1360 69312 1409 69340
rect 1360 69300 1366 69312
rect 1397 69309 1409 69312
rect 1443 69309 1455 69343
rect 1397 69303 1455 69309
rect 569954 68348 569960 68400
rect 570012 68388 570018 68400
rect 570230 68388 570236 68400
rect 570012 68360 570236 68388
rect 570012 68348 570018 68360
rect 570230 68348 570236 68360
rect 570288 68348 570294 68400
rect 569954 68008 569960 68060
rect 570012 68048 570018 68060
rect 570325 68051 570383 68057
rect 570325 68048 570337 68051
rect 570012 68020 570337 68048
rect 570012 68008 570018 68020
rect 570325 68017 570337 68020
rect 570371 68017 570383 68051
rect 570325 68011 570383 68017
rect 569954 67872 569960 67924
rect 570012 67912 570018 67924
rect 570138 67912 570144 67924
rect 570012 67884 570144 67912
rect 570012 67872 570018 67884
rect 570138 67872 570144 67884
rect 570196 67872 570202 67924
rect 1029 67507 1087 67513
rect 1029 67473 1041 67507
rect 1075 67504 1087 67507
rect 1946 67504 1952 67516
rect 1075 67476 1952 67504
rect 1075 67473 1087 67476
rect 1029 67467 1087 67473
rect 1946 67464 1952 67476
rect 2004 67464 2010 67516
rect 1302 67328 1308 67380
rect 1360 67368 1366 67380
rect 1946 67368 1952 67380
rect 1360 67340 1952 67368
rect 1360 67328 1366 67340
rect 1946 67328 1952 67340
rect 2004 67328 2010 67380
rect 937 67235 995 67241
rect 937 67201 949 67235
rect 983 67232 995 67235
rect 1946 67232 1952 67244
rect 983 67204 1952 67232
rect 983 67201 995 67204
rect 937 67195 995 67201
rect 1946 67192 1952 67204
rect 2004 67192 2010 67244
rect 198 66920 204 66972
rect 256 66960 262 66972
rect 1489 66963 1547 66969
rect 1489 66960 1501 66963
rect 256 66932 1501 66960
rect 256 66920 262 66932
rect 1489 66929 1501 66932
rect 1535 66929 1547 66963
rect 1489 66923 1547 66929
rect 753 66759 811 66765
rect 753 66725 765 66759
rect 799 66756 811 66759
rect 1946 66756 1952 66768
rect 799 66728 1952 66756
rect 799 66725 811 66728
rect 753 66719 811 66725
rect 1946 66716 1952 66728
rect 2004 66716 2010 66768
rect 845 66623 903 66629
rect 845 66589 857 66623
rect 891 66620 903 66623
rect 1946 66620 1952 66632
rect 891 66592 1952 66620
rect 891 66589 903 66592
rect 845 66583 903 66589
rect 1946 66580 1952 66592
rect 2004 66580 2010 66632
rect 1946 66484 1952 66496
rect 1907 66456 1952 66484
rect 1946 66444 1952 66456
rect 2004 66444 2010 66496
rect 1673 66351 1731 66357
rect 1673 66317 1685 66351
rect 1719 66348 1731 66351
rect 1949 66351 2007 66357
rect 1949 66348 1961 66351
rect 1719 66320 1961 66348
rect 1719 66317 1731 66320
rect 1673 66311 1731 66317
rect 1949 66317 1961 66320
rect 1995 66317 2007 66351
rect 1949 66311 2007 66317
rect 570138 66104 570144 66156
rect 570196 66144 570202 66156
rect 570509 66147 570567 66153
rect 570509 66144 570521 66147
rect 570196 66116 570521 66144
rect 570196 66104 570202 66116
rect 570509 66113 570521 66116
rect 570555 66113 570567 66147
rect 570509 66107 570567 66113
rect 570046 65968 570052 66020
rect 570104 66008 570110 66020
rect 570509 66011 570567 66017
rect 570509 66008 570521 66011
rect 570104 65980 570521 66008
rect 570104 65968 570110 65980
rect 570509 65977 570521 65980
rect 570555 65977 570567 66011
rect 570509 65971 570567 65977
rect 1670 65872 1676 65884
rect 1631 65844 1676 65872
rect 1670 65832 1676 65844
rect 1728 65832 1734 65884
rect 1121 65467 1179 65473
rect 1121 65433 1133 65467
rect 1167 65464 1179 65467
rect 1210 65464 1216 65476
rect 1167 65436 1216 65464
rect 1167 65433 1179 65436
rect 1121 65427 1179 65433
rect 1210 65424 1216 65436
rect 1268 65424 1274 65476
rect 1581 65467 1639 65473
rect 1581 65433 1593 65467
rect 1627 65464 1639 65467
rect 1857 65467 1915 65473
rect 1857 65464 1869 65467
rect 1627 65436 1869 65464
rect 1627 65433 1639 65436
rect 1581 65427 1639 65433
rect 1857 65433 1869 65436
rect 1903 65433 1915 65467
rect 2038 65464 2044 65476
rect 1857 65427 1915 65433
rect 1964 65436 2044 65464
rect 1964 65396 1992 65436
rect 2038 65424 2044 65436
rect 2096 65424 2102 65476
rect 1320 65368 1992 65396
rect 1320 65272 1348 65368
rect 1302 65220 1308 65272
rect 1360 65220 1366 65272
rect 569954 64948 569960 65000
rect 570012 64988 570018 65000
rect 570417 64991 570475 64997
rect 570417 64988 570429 64991
rect 570012 64960 570429 64988
rect 570012 64948 570018 64960
rect 570417 64957 570429 64960
rect 570463 64957 570475 64991
rect 570417 64951 570475 64957
rect 1670 64784 1676 64796
rect 1631 64756 1676 64784
rect 1670 64744 1676 64756
rect 1728 64744 1734 64796
rect 1857 64787 1915 64793
rect 1857 64753 1869 64787
rect 1903 64784 1915 64787
rect 1946 64784 1952 64796
rect 1903 64756 1952 64784
rect 1903 64753 1915 64756
rect 1857 64747 1915 64753
rect 1946 64744 1952 64756
rect 2004 64744 2010 64796
rect 753 64651 811 64657
rect 753 64617 765 64651
rect 799 64648 811 64651
rect 1946 64648 1952 64660
rect 799 64620 1952 64648
rect 799 64617 811 64620
rect 753 64611 811 64617
rect 1946 64608 1952 64620
rect 2004 64608 2010 64660
rect 574738 63520 574744 63572
rect 574796 63560 574802 63572
rect 580166 63560 580172 63572
rect 574796 63532 580172 63560
rect 574796 63520 574802 63532
rect 580166 63520 580172 63532
rect 580224 63520 580230 63572
rect 1210 63316 1216 63368
rect 1268 63356 1274 63368
rect 1946 63356 1952 63368
rect 1268 63328 1952 63356
rect 1268 63316 1274 63328
rect 1946 63316 1952 63328
rect 2004 63316 2010 63368
rect 937 63155 995 63161
rect 937 63121 949 63155
rect 983 63152 995 63155
rect 1946 63152 1952 63164
rect 983 63124 1952 63152
rect 983 63121 995 63124
rect 937 63115 995 63121
rect 1946 63112 1952 63124
rect 2004 63112 2010 63164
rect 1397 63019 1455 63025
rect 1397 62985 1409 63019
rect 1443 63016 1455 63019
rect 1946 63016 1952 63028
rect 1443 62988 1952 63016
rect 1443 62985 1455 62988
rect 1397 62979 1455 62985
rect 1946 62976 1952 62988
rect 2004 62976 2010 63028
rect 1029 62883 1087 62889
rect 1029 62849 1041 62883
rect 1075 62880 1087 62883
rect 1946 62880 1952 62892
rect 1075 62852 1952 62880
rect 1075 62849 1087 62852
rect 1029 62843 1087 62849
rect 1946 62840 1952 62852
rect 2004 62840 2010 62892
rect 1213 62747 1271 62753
rect 1213 62713 1225 62747
rect 1259 62744 1271 62747
rect 1581 62747 1639 62753
rect 1581 62744 1593 62747
rect 1259 62716 1593 62744
rect 1259 62713 1271 62716
rect 1213 62707 1271 62713
rect 1581 62713 1593 62716
rect 1627 62713 1639 62747
rect 1581 62707 1639 62713
rect 1121 62271 1179 62277
rect 1121 62237 1133 62271
rect 1167 62268 1179 62271
rect 1946 62268 1952 62280
rect 1167 62240 1952 62268
rect 1167 62237 1179 62240
rect 1121 62231 1179 62237
rect 1946 62228 1952 62240
rect 2004 62228 2010 62280
rect 569954 61724 569960 61736
rect 569880 61696 569960 61724
rect 569880 61316 569908 61696
rect 569954 61684 569960 61696
rect 570012 61684 570018 61736
rect 569954 61548 569960 61600
rect 570012 61588 570018 61600
rect 570138 61588 570144 61600
rect 570012 61560 570144 61588
rect 570012 61548 570018 61560
rect 570138 61548 570144 61560
rect 570196 61548 570202 61600
rect 570046 61316 570052 61328
rect 569880 61288 570052 61316
rect 570046 61276 570052 61288
rect 570104 61276 570110 61328
rect 569954 60732 569960 60784
rect 570012 60772 570018 60784
rect 570325 60775 570383 60781
rect 570325 60772 570337 60775
rect 570012 60744 570337 60772
rect 570012 60732 570018 60744
rect 570325 60741 570337 60744
rect 570371 60741 570383 60775
rect 570325 60735 570383 60741
rect 569954 59916 569960 59968
rect 570012 59956 570018 59968
rect 570233 59959 570291 59965
rect 570233 59956 570245 59959
rect 570012 59928 570245 59956
rect 570012 59916 570018 59928
rect 570233 59925 570245 59928
rect 570279 59925 570291 59959
rect 570233 59919 570291 59925
rect 569865 58871 569923 58877
rect 569865 58837 569877 58871
rect 569911 58868 569923 58871
rect 569954 58868 569960 58880
rect 569911 58840 569960 58868
rect 569911 58837 569923 58840
rect 569865 58831 569923 58837
rect 569954 58828 569960 58840
rect 570012 58828 570018 58880
rect 569954 58692 569960 58744
rect 570012 58732 570018 58744
rect 570417 58735 570475 58741
rect 570417 58732 570429 58735
rect 570012 58704 570429 58732
rect 570012 58692 570018 58704
rect 570417 58701 570429 58704
rect 570463 58701 570475 58735
rect 570417 58695 570475 58701
rect 845 57919 903 57925
rect 845 57885 857 57919
rect 891 57916 903 57919
rect 1302 57916 1308 57928
rect 891 57888 1308 57916
rect 891 57885 903 57888
rect 845 57879 903 57885
rect 1302 57876 1308 57888
rect 1360 57876 1366 57928
rect 1213 57103 1271 57109
rect 1213 57069 1225 57103
rect 1259 57100 1271 57103
rect 1946 57100 1952 57112
rect 1259 57072 1952 57100
rect 1259 57069 1271 57072
rect 1213 57063 1271 57069
rect 1946 57060 1952 57072
rect 2004 57060 2010 57112
rect 569954 56964 569960 56976
rect 569915 56936 569960 56964
rect 569954 56924 569960 56936
rect 570012 56924 570018 56976
rect 1946 56896 1952 56908
rect 1320 56868 1952 56896
rect 1320 56624 1348 56868
rect 1946 56856 1952 56868
rect 2004 56856 2010 56908
rect 1397 56763 1455 56769
rect 1397 56729 1409 56763
rect 1443 56760 1455 56763
rect 1946 56760 1952 56772
rect 1443 56732 1952 56760
rect 1443 56729 1455 56732
rect 1397 56723 1455 56729
rect 1946 56720 1952 56732
rect 2004 56720 2010 56772
rect 569954 56652 569960 56704
rect 570012 56692 570018 56704
rect 570141 56695 570199 56701
rect 570141 56692 570153 56695
rect 570012 56664 570153 56692
rect 570012 56652 570018 56664
rect 570141 56661 570153 56664
rect 570187 56661 570199 56695
rect 570141 56655 570199 56661
rect 1946 56624 1952 56636
rect 1320 56596 1952 56624
rect 1946 56584 1952 56596
rect 2004 56584 2010 56636
rect 570509 56627 570567 56633
rect 570509 56593 570521 56627
rect 570555 56593 570567 56627
rect 570509 56587 570567 56593
rect 569954 56516 569960 56568
rect 570012 56556 570018 56568
rect 570524 56556 570552 56587
rect 570012 56528 570552 56556
rect 570012 56516 570018 56528
rect 1213 55879 1271 55885
rect 1213 55845 1225 55879
rect 1259 55876 1271 55879
rect 1946 55876 1952 55888
rect 1259 55848 1952 55876
rect 1259 55845 1271 55848
rect 1213 55839 1271 55845
rect 1946 55836 1952 55848
rect 2004 55836 2010 55888
rect 1397 55199 1455 55205
rect 1397 55165 1409 55199
rect 1443 55196 1455 55199
rect 1946 55196 1952 55208
rect 1443 55168 1952 55196
rect 1443 55165 1455 55168
rect 1397 55159 1455 55165
rect 1946 55156 1952 55168
rect 2004 55156 2010 55208
rect 569954 53728 569960 53780
rect 570012 53768 570018 53780
rect 570049 53771 570107 53777
rect 570049 53768 570061 53771
rect 570012 53740 570061 53768
rect 570012 53728 570018 53740
rect 570049 53737 570061 53740
rect 570095 53737 570107 53771
rect 570049 53731 570107 53737
rect 1305 52751 1363 52757
rect 1305 52717 1317 52751
rect 1351 52748 1363 52751
rect 1946 52748 1952 52760
rect 1351 52720 1952 52748
rect 1351 52717 1363 52720
rect 1305 52711 1363 52717
rect 1946 52708 1952 52720
rect 2004 52708 2010 52760
rect 1489 52615 1547 52621
rect 1489 52581 1501 52615
rect 1535 52612 1547 52615
rect 1946 52612 1952 52624
rect 1535 52584 1952 52612
rect 1535 52581 1547 52584
rect 1489 52575 1547 52581
rect 1946 52572 1952 52584
rect 2004 52572 2010 52624
rect 17 50439 75 50445
rect 17 50405 29 50439
rect 63 50436 75 50439
rect 1857 50439 1915 50445
rect 1857 50436 1869 50439
rect 63 50408 1869 50436
rect 63 50405 75 50408
rect 17 50399 75 50405
rect 1857 50405 1869 50408
rect 1903 50405 1915 50439
rect 1857 50399 1915 50405
rect 1026 50368 1032 50380
rect 987 50340 1032 50368
rect 1026 50328 1032 50340
rect 1084 50328 1090 50380
rect 1765 47651 1823 47657
rect 1765 47617 1777 47651
rect 1811 47648 1823 47651
rect 1949 47651 2007 47657
rect 1949 47648 1961 47651
rect 1811 47620 1961 47648
rect 1811 47617 1823 47620
rect 1765 47611 1823 47617
rect 1949 47617 1961 47620
rect 1995 47617 2007 47651
rect 1949 47611 2007 47617
rect 106 47472 112 47524
rect 164 47512 170 47524
rect 1765 47515 1823 47521
rect 1765 47512 1777 47515
rect 164 47484 1777 47512
rect 164 47472 170 47484
rect 1765 47481 1777 47484
rect 1811 47481 1823 47515
rect 1765 47475 1823 47481
rect 1397 45543 1455 45549
rect 1397 45509 1409 45543
rect 1443 45540 1455 45543
rect 1581 45543 1639 45549
rect 1581 45540 1593 45543
rect 1443 45512 1593 45540
rect 1443 45509 1455 45512
rect 1397 45503 1455 45509
rect 1581 45509 1593 45512
rect 1627 45509 1639 45543
rect 1581 45503 1639 45509
rect 569954 45500 569960 45552
rect 570012 45540 570018 45552
rect 570322 45540 570328 45552
rect 570012 45512 570328 45540
rect 570012 45500 570018 45512
rect 570322 45500 570328 45512
rect 570380 45500 570386 45552
rect 1673 43503 1731 43509
rect 1673 43469 1685 43503
rect 1719 43500 1731 43503
rect 1949 43503 2007 43509
rect 1949 43500 1961 43503
rect 1719 43472 1961 43500
rect 1719 43469 1731 43472
rect 1673 43463 1731 43469
rect 1949 43469 1961 43472
rect 1995 43469 2007 43503
rect 1949 43463 2007 43469
rect 569954 43256 569960 43308
rect 570012 43296 570018 43308
rect 570509 43299 570567 43305
rect 570509 43296 570521 43299
rect 570012 43268 570521 43296
rect 570012 43256 570018 43268
rect 570509 43265 570521 43268
rect 570555 43265 570567 43299
rect 570509 43259 570567 43265
rect 1397 43095 1455 43101
rect 1397 43061 1409 43095
rect 1443 43092 1455 43095
rect 1946 43092 1952 43104
rect 1443 43064 1952 43092
rect 1443 43061 1455 43064
rect 1397 43055 1455 43061
rect 1946 43052 1952 43064
rect 2004 43052 2010 43104
rect 1581 42823 1639 42829
rect 1581 42789 1593 42823
rect 1627 42820 1639 42823
rect 1946 42820 1952 42832
rect 1627 42792 1952 42820
rect 1627 42789 1639 42792
rect 1581 42783 1639 42789
rect 1946 42780 1952 42792
rect 2004 42780 2010 42832
rect 569954 42344 569960 42356
rect 569915 42316 569960 42344
rect 569954 42304 569960 42316
rect 570012 42304 570018 42356
rect 569954 42168 569960 42220
rect 570012 42208 570018 42220
rect 570233 42211 570291 42217
rect 570233 42208 570245 42211
rect 570012 42180 570245 42208
rect 570012 42168 570018 42180
rect 570233 42177 570245 42180
rect 570279 42177 570291 42211
rect 570233 42171 570291 42177
rect 569954 41760 569960 41812
rect 570012 41800 570018 41812
rect 570325 41803 570383 41809
rect 570325 41800 570337 41803
rect 570012 41772 570337 41800
rect 570012 41760 570018 41772
rect 570325 41769 570337 41772
rect 570371 41769 570383 41803
rect 570325 41763 570383 41769
rect 569954 41624 569960 41676
rect 570012 41664 570018 41676
rect 570049 41667 570107 41673
rect 570049 41664 570061 41667
rect 570012 41636 570061 41664
rect 570012 41624 570018 41636
rect 570049 41633 570061 41636
rect 570095 41633 570107 41667
rect 570049 41627 570107 41633
rect 569954 41080 569960 41132
rect 570012 41120 570018 41132
rect 570141 41123 570199 41129
rect 570141 41120 570153 41123
rect 570012 41092 570153 41120
rect 570012 41080 570018 41092
rect 570141 41089 570153 41092
rect 570187 41089 570199 41123
rect 570141 41083 570199 41089
rect 569954 40984 569960 40996
rect 569915 40956 569960 40984
rect 569954 40944 569960 40956
rect 570012 40944 570018 40996
rect 569954 40712 569960 40724
rect 569880 40684 569960 40712
rect 569880 40168 569908 40684
rect 569954 40672 569960 40684
rect 570012 40672 570018 40724
rect 569954 40400 569960 40452
rect 570012 40440 570018 40452
rect 570417 40443 570475 40449
rect 570417 40440 570429 40443
rect 570012 40412 570429 40440
rect 570012 40400 570018 40412
rect 570417 40409 570429 40412
rect 570463 40409 570475 40443
rect 570417 40403 570475 40409
rect 569954 40264 569960 40316
rect 570012 40304 570018 40316
rect 570601 40307 570659 40313
rect 570601 40304 570613 40307
rect 570012 40276 570613 40304
rect 570012 40264 570018 40276
rect 570601 40273 570613 40276
rect 570647 40273 570659 40307
rect 570601 40267 570659 40273
rect 569954 40168 569960 40180
rect 569880 40140 569960 40168
rect 569954 40128 569960 40140
rect 570012 40128 570018 40180
rect 569954 39992 569960 40044
rect 570012 40032 570018 40044
rect 570417 40035 570475 40041
rect 570417 40032 570429 40035
rect 570012 40004 570429 40032
rect 570012 39992 570018 40004
rect 570417 40001 570429 40004
rect 570463 40001 570475 40035
rect 570417 39995 570475 40001
rect 569954 39856 569960 39908
rect 570012 39896 570018 39908
rect 570141 39899 570199 39905
rect 570141 39896 570153 39899
rect 570012 39868 570153 39896
rect 570012 39856 570018 39868
rect 570141 39865 570153 39868
rect 570187 39865 570199 39899
rect 570141 39859 570199 39865
rect 570141 39763 570199 39769
rect 570141 39729 570153 39763
rect 570187 39760 570199 39763
rect 570325 39763 570383 39769
rect 570325 39760 570337 39763
rect 570187 39732 570337 39760
rect 570187 39729 570199 39732
rect 570141 39723 570199 39729
rect 570325 39729 570337 39732
rect 570371 39729 570383 39763
rect 570325 39723 570383 39729
rect 569954 39692 569960 39704
rect 569915 39664 569960 39692
rect 569954 39652 569960 39664
rect 570012 39652 570018 39704
rect 1121 39491 1179 39497
rect 1121 39457 1133 39491
rect 1167 39488 1179 39491
rect 1946 39488 1952 39500
rect 1167 39460 1952 39488
rect 1167 39457 1179 39460
rect 1121 39451 1179 39457
rect 1946 39448 1952 39460
rect 2004 39448 2010 39500
rect 569954 39380 569960 39432
rect 570012 39420 570018 39432
rect 570049 39423 570107 39429
rect 570049 39420 570061 39423
rect 570012 39392 570061 39420
rect 570012 39380 570018 39392
rect 570049 39389 570061 39392
rect 570095 39389 570107 39423
rect 570049 39383 570107 39389
rect 1397 39355 1455 39361
rect 1397 39321 1409 39355
rect 1443 39352 1455 39355
rect 1486 39352 1492 39364
rect 1443 39324 1492 39352
rect 1443 39321 1455 39324
rect 1397 39315 1455 39321
rect 1486 39312 1492 39324
rect 1544 39312 1550 39364
rect 1857 39355 1915 39361
rect 1857 39321 1869 39355
rect 1903 39352 1915 39355
rect 1946 39352 1952 39364
rect 1903 39324 1952 39352
rect 1903 39321 1915 39324
rect 1857 39315 1915 39321
rect 1946 39312 1952 39324
rect 2004 39312 2010 39364
rect 1765 39219 1823 39225
rect 1765 39185 1777 39219
rect 1811 39216 1823 39219
rect 1946 39216 1952 39228
rect 1811 39188 1952 39216
rect 1811 39185 1823 39188
rect 1765 39179 1823 39185
rect 1946 39176 1952 39188
rect 2004 39176 2010 39228
rect 570230 39040 570236 39092
rect 570288 39080 570294 39092
rect 570509 39083 570567 39089
rect 570509 39080 570521 39083
rect 570288 39052 570521 39080
rect 570288 39040 570294 39052
rect 570509 39049 570521 39052
rect 570555 39049 570567 39083
rect 570509 39043 570567 39049
rect 1302 38496 1308 38548
rect 1360 38536 1366 38548
rect 1854 38536 1860 38548
rect 1360 38508 1860 38536
rect 1360 38496 1366 38508
rect 1854 38496 1860 38508
rect 1912 38496 1918 38548
rect 1026 37040 1032 37052
rect 987 37012 1032 37040
rect 1026 37000 1032 37012
rect 1084 37000 1090 37052
rect 1305 35683 1363 35689
rect 1305 35649 1317 35683
rect 1351 35680 1363 35683
rect 1946 35680 1952 35692
rect 1351 35652 1952 35680
rect 1351 35649 1363 35652
rect 1305 35643 1363 35649
rect 1946 35640 1952 35652
rect 2004 35640 2010 35692
rect 1213 35547 1271 35553
rect 1213 35513 1225 35547
rect 1259 35544 1271 35547
rect 1946 35544 1952 35556
rect 1259 35516 1952 35544
rect 1259 35513 1271 35516
rect 1213 35507 1271 35513
rect 1946 35504 1952 35516
rect 2004 35504 2010 35556
rect 1029 35411 1087 35417
rect 1029 35377 1041 35411
rect 1075 35408 1087 35411
rect 1946 35408 1952 35420
rect 1075 35380 1952 35408
rect 1075 35377 1087 35380
rect 1029 35371 1087 35377
rect 1946 35368 1952 35380
rect 2004 35368 2010 35420
rect 382 35232 388 35284
rect 440 35272 446 35284
rect 1946 35272 1952 35284
rect 440 35244 1952 35272
rect 440 35232 446 35244
rect 1946 35232 1952 35244
rect 2004 35232 2010 35284
rect 14 34960 20 35012
rect 72 35000 78 35012
rect 72 34972 117 35000
rect 72 34960 78 34972
rect 570322 34756 570328 34808
rect 570380 34796 570386 34808
rect 570601 34799 570659 34805
rect 570601 34796 570613 34799
rect 570380 34768 570613 34796
rect 570380 34756 570386 34768
rect 570601 34765 570613 34768
rect 570647 34765 570659 34799
rect 570601 34759 570659 34765
rect 658 33572 664 33584
rect 619 33544 664 33572
rect 658 33532 664 33544
rect 716 33532 722 33584
rect 570138 31016 570144 31068
rect 570196 31056 570202 31068
rect 570325 31059 570383 31065
rect 570325 31056 570337 31059
rect 570196 31028 570337 31056
rect 570196 31016 570202 31028
rect 570325 31025 570337 31028
rect 570371 31025 570383 31059
rect 570325 31019 570383 31025
rect 106 29860 112 29912
rect 164 29900 170 29912
rect 1949 29903 2007 29909
rect 1949 29900 1961 29903
rect 164 29872 1961 29900
rect 164 29860 170 29872
rect 1949 29869 1961 29872
rect 1995 29869 2007 29903
rect 1949 29863 2007 29869
rect 1854 29724 1860 29776
rect 1912 29764 1918 29776
rect 1949 29767 2007 29773
rect 1949 29764 1961 29767
rect 1912 29736 1961 29764
rect 1912 29724 1918 29736
rect 1949 29733 1961 29736
rect 1995 29733 2007 29767
rect 1949 29727 2007 29733
rect 1581 29699 1639 29705
rect 1581 29665 1593 29699
rect 1627 29696 1639 29699
rect 1762 29696 1768 29708
rect 1627 29668 1768 29696
rect 1627 29665 1639 29668
rect 1581 29659 1639 29665
rect 1762 29656 1768 29668
rect 1820 29656 1826 29708
rect 1121 29631 1179 29637
rect 1121 29597 1133 29631
rect 1167 29628 1179 29631
rect 1857 29631 1915 29637
rect 1857 29628 1869 29631
rect 1167 29600 1869 29628
rect 1167 29597 1179 29600
rect 1121 29591 1179 29597
rect 1857 29597 1869 29600
rect 1903 29597 1915 29631
rect 1857 29591 1915 29597
rect 1029 29563 1087 29569
rect 1029 29529 1041 29563
rect 1075 29560 1087 29563
rect 1762 29560 1768 29572
rect 1075 29532 1768 29560
rect 1075 29529 1087 29532
rect 1029 29523 1087 29529
rect 1762 29520 1768 29532
rect 1820 29520 1826 29572
rect 1486 29492 1492 29504
rect 1447 29464 1492 29492
rect 1486 29452 1492 29464
rect 1544 29452 1550 29504
rect 1397 29019 1455 29025
rect 1397 28985 1409 29019
rect 1443 29016 1455 29019
rect 1443 28988 1532 29016
rect 1443 28985 1455 28988
rect 1397 28979 1455 28985
rect 937 28883 995 28889
rect 937 28849 949 28883
rect 983 28880 995 28883
rect 1504 28880 1532 28988
rect 983 28852 1532 28880
rect 983 28849 995 28852
rect 937 28843 995 28849
rect 1397 28339 1455 28345
rect 1397 28305 1409 28339
rect 1443 28336 1455 28339
rect 1946 28336 1952 28348
rect 1443 28308 1952 28336
rect 1443 28305 1455 28308
rect 1397 28299 1455 28305
rect 1946 28296 1952 28308
rect 2004 28296 2010 28348
rect 1486 27956 1492 28008
rect 1544 27996 1550 28008
rect 1946 27996 1952 28008
rect 1544 27968 1952 27996
rect 1544 27956 1550 27968
rect 1946 27956 1952 27968
rect 2004 27956 2010 28008
rect 569957 27931 570015 27937
rect 569957 27897 569969 27931
rect 570003 27928 570015 27931
rect 570233 27931 570291 27937
rect 570233 27928 570245 27931
rect 570003 27900 570245 27928
rect 570003 27897 570015 27900
rect 569957 27891 570015 27897
rect 570233 27897 570245 27900
rect 570279 27897 570291 27931
rect 570233 27891 570291 27897
rect 1213 27251 1271 27257
rect 1213 27217 1225 27251
rect 1259 27248 1271 27251
rect 1946 27248 1952 27260
rect 1259 27220 1952 27248
rect 1259 27217 1271 27220
rect 1213 27211 1271 27217
rect 1946 27208 1952 27220
rect 2004 27208 2010 27260
rect 1029 27115 1087 27121
rect 1029 27081 1041 27115
rect 1075 27112 1087 27115
rect 1210 27112 1216 27124
rect 1075 27084 1216 27112
rect 1075 27081 1087 27084
rect 1029 27075 1087 27081
rect 1210 27072 1216 27084
rect 1268 27072 1274 27124
rect 1489 27115 1547 27121
rect 1489 27081 1501 27115
rect 1535 27112 1547 27115
rect 1946 27112 1952 27124
rect 1535 27084 1952 27112
rect 1535 27081 1547 27084
rect 1489 27075 1547 27081
rect 1946 27072 1952 27084
rect 2004 27072 2010 27124
rect 1210 26936 1216 26988
rect 1268 26976 1274 26988
rect 1946 26976 1952 26988
rect 1268 26948 1952 26976
rect 1268 26936 1274 26948
rect 1946 26936 1952 26948
rect 2004 26936 2010 26988
rect 1486 26800 1492 26852
rect 1544 26840 1550 26852
rect 1946 26840 1952 26852
rect 1544 26812 1952 26840
rect 1544 26800 1550 26812
rect 1946 26800 1952 26812
rect 2004 26800 2010 26852
rect 569954 26460 569960 26512
rect 570012 26500 570018 26512
rect 570233 26503 570291 26509
rect 570233 26500 570245 26503
rect 570012 26472 570245 26500
rect 570012 26460 570018 26472
rect 570233 26469 570245 26472
rect 570279 26469 570291 26503
rect 570233 26463 570291 26469
rect 569954 25712 569960 25764
rect 570012 25752 570018 25764
rect 570049 25755 570107 25761
rect 570049 25752 570061 25755
rect 570012 25724 570061 25752
rect 570012 25712 570018 25724
rect 570049 25721 570061 25724
rect 570095 25721 570107 25755
rect 570049 25715 570107 25721
rect 569954 25508 569960 25560
rect 570012 25548 570018 25560
rect 570417 25551 570475 25557
rect 570417 25548 570429 25551
rect 570012 25520 570429 25548
rect 570012 25508 570018 25520
rect 570417 25517 570429 25520
rect 570463 25517 570475 25551
rect 570417 25511 570475 25517
rect 569954 25100 569960 25152
rect 570012 25140 570018 25152
rect 570230 25140 570236 25152
rect 570012 25112 570236 25140
rect 570012 25100 570018 25112
rect 570230 25100 570236 25112
rect 570288 25100 570294 25152
rect 569954 24284 569960 24336
rect 570012 24324 570018 24336
rect 570322 24324 570328 24336
rect 570012 24296 570328 24324
rect 570012 24284 570018 24296
rect 570322 24284 570328 24296
rect 570380 24284 570386 24336
rect 106 24256 112 24268
rect 67 24228 112 24256
rect 106 24216 112 24228
rect 164 24216 170 24268
rect 569954 24148 569960 24200
rect 570012 24188 570018 24200
rect 570417 24191 570475 24197
rect 570417 24188 570429 24191
rect 570012 24160 570429 24188
rect 570012 24148 570018 24160
rect 570417 24157 570429 24160
rect 570463 24157 570475 24191
rect 570417 24151 570475 24157
rect 569 24055 627 24061
rect 569 24021 581 24055
rect 615 24052 627 24055
rect 1486 24052 1492 24064
rect 615 24024 1492 24052
rect 615 24021 627 24024
rect 569 24015 627 24021
rect 1486 24012 1492 24024
rect 1544 24012 1550 24064
rect 937 23783 995 23789
rect 937 23749 949 23783
rect 983 23780 995 23783
rect 1486 23780 1492 23792
rect 983 23752 1492 23780
rect 983 23749 995 23752
rect 937 23743 995 23749
rect 1486 23740 1492 23752
rect 1544 23740 1550 23792
rect 569954 23740 569960 23792
rect 570012 23780 570018 23792
rect 570233 23783 570291 23789
rect 570233 23780 570245 23783
rect 570012 23752 570245 23780
rect 570012 23740 570018 23752
rect 570233 23749 570245 23752
rect 570279 23749 570291 23783
rect 570233 23743 570291 23749
rect 569954 23536 569960 23588
rect 570012 23576 570018 23588
rect 570230 23576 570236 23588
rect 570012 23548 570236 23576
rect 570012 23536 570018 23548
rect 570230 23536 570236 23548
rect 570288 23536 570294 23588
rect 569954 23196 569960 23248
rect 570012 23236 570018 23248
rect 570141 23239 570199 23245
rect 570141 23236 570153 23239
rect 570012 23208 570153 23236
rect 570012 23196 570018 23208
rect 570141 23205 570153 23208
rect 570187 23205 570199 23239
rect 570141 23199 570199 23205
rect 569957 23103 570015 23109
rect 569957 23069 569969 23103
rect 570003 23100 570015 23103
rect 570141 23103 570199 23109
rect 570141 23100 570153 23103
rect 570003 23072 570153 23100
rect 570003 23069 570015 23072
rect 569957 23063 570015 23069
rect 570141 23069 570153 23072
rect 570187 23069 570199 23103
rect 570141 23063 570199 23069
rect 1397 22219 1455 22225
rect 1397 22185 1409 22219
rect 1443 22216 1455 22219
rect 1946 22216 1952 22228
rect 1443 22188 1952 22216
rect 1443 22185 1455 22188
rect 1397 22179 1455 22185
rect 1946 22176 1952 22188
rect 2004 22176 2010 22228
rect 661 22083 719 22089
rect 661 22049 673 22083
rect 707 22080 719 22083
rect 1946 22080 1952 22092
rect 707 22052 1952 22080
rect 707 22049 719 22052
rect 661 22043 719 22049
rect 1946 22040 1952 22052
rect 2004 22040 2010 22092
rect 1302 21564 1308 21616
rect 1360 21604 1366 21616
rect 1489 21607 1547 21613
rect 1489 21604 1501 21607
rect 1360 21576 1501 21604
rect 1360 21564 1366 21576
rect 1489 21573 1501 21576
rect 1535 21573 1547 21607
rect 1489 21567 1547 21573
rect 106 20136 112 20188
rect 164 20176 170 20188
rect 1394 20176 1400 20188
rect 164 20148 1400 20176
rect 164 20136 170 20148
rect 1394 20136 1400 20148
rect 1452 20136 1458 20188
rect 1857 20111 1915 20117
rect 1857 20108 1869 20111
rect 768 20080 1869 20108
rect 768 19848 796 20080
rect 1857 20077 1869 20080
rect 1903 20077 1915 20111
rect 1857 20071 1915 20077
rect 937 20043 995 20049
rect 937 20009 949 20043
rect 983 20040 995 20043
rect 1026 20040 1032 20052
rect 983 20012 1032 20040
rect 983 20009 995 20012
rect 937 20003 995 20009
rect 1026 20000 1032 20012
rect 1084 20000 1090 20052
rect 1394 19932 1400 19984
rect 1452 19972 1458 19984
rect 1765 19975 1823 19981
rect 1765 19972 1777 19975
rect 1452 19944 1777 19972
rect 1452 19932 1458 19944
rect 1765 19941 1777 19944
rect 1811 19941 1823 19975
rect 1765 19935 1823 19941
rect 750 19796 756 19848
rect 808 19796 814 19848
rect 1302 18844 1308 18896
rect 1360 18884 1366 18896
rect 1949 18887 2007 18893
rect 1949 18884 1961 18887
rect 1360 18856 1961 18884
rect 1360 18844 1366 18856
rect 1949 18853 1961 18856
rect 1995 18853 2007 18887
rect 1949 18847 2007 18853
rect 1394 18708 1400 18760
rect 1452 18748 1458 18760
rect 1949 18751 2007 18757
rect 1949 18748 1961 18751
rect 1452 18720 1961 18748
rect 1452 18708 1458 18720
rect 1949 18717 1961 18720
rect 1995 18717 2007 18751
rect 1949 18711 2007 18717
rect 1029 18615 1087 18621
rect 1029 18581 1041 18615
rect 1075 18612 1087 18615
rect 1394 18612 1400 18624
rect 1075 18584 1400 18612
rect 1075 18581 1087 18584
rect 1029 18575 1087 18581
rect 1394 18572 1400 18584
rect 1452 18572 1458 18624
rect 753 18479 811 18485
rect 753 18445 765 18479
rect 799 18476 811 18479
rect 1946 18476 1952 18488
rect 799 18448 1952 18476
rect 799 18445 811 18448
rect 753 18439 811 18445
rect 1946 18436 1952 18448
rect 2004 18436 2010 18488
rect 1026 18368 1032 18420
rect 1084 18408 1090 18420
rect 1581 18411 1639 18417
rect 1581 18408 1593 18411
rect 1084 18380 1593 18408
rect 1084 18368 1090 18380
rect 1581 18377 1593 18380
rect 1627 18377 1639 18411
rect 1581 18371 1639 18377
rect 474 18232 480 18284
rect 532 18272 538 18284
rect 1581 18275 1639 18281
rect 1581 18272 1593 18275
rect 532 18244 1593 18272
rect 532 18232 538 18244
rect 1581 18241 1593 18244
rect 1627 18241 1639 18275
rect 1581 18235 1639 18241
rect 1029 17935 1087 17941
rect 1029 17901 1041 17935
rect 1075 17932 1087 17935
rect 1854 17932 1860 17944
rect 1075 17904 1860 17932
rect 1075 17901 1087 17904
rect 1029 17895 1087 17901
rect 1854 17892 1860 17904
rect 1912 17892 1918 17944
rect 569954 17620 569960 17672
rect 570012 17660 570018 17672
rect 570141 17663 570199 17669
rect 570141 17660 570153 17663
rect 570012 17632 570153 17660
rect 570012 17620 570018 17632
rect 570141 17629 570153 17632
rect 570187 17629 570199 17663
rect 570141 17623 570199 17629
rect 845 17119 903 17125
rect 845 17085 857 17119
rect 891 17116 903 17119
rect 1673 17119 1731 17125
rect 1673 17116 1685 17119
rect 891 17088 1685 17116
rect 891 17085 903 17088
rect 845 17079 903 17085
rect 1673 17085 1685 17088
rect 1719 17085 1731 17119
rect 1673 17079 1731 17085
rect 109 16983 167 16989
rect 109 16949 121 16983
rect 155 16980 167 16983
rect 1673 16983 1731 16989
rect 1673 16980 1685 16983
rect 155 16952 1685 16980
rect 155 16949 167 16952
rect 109 16943 167 16949
rect 1673 16949 1685 16952
rect 1719 16949 1731 16983
rect 1673 16943 1731 16949
rect 1118 16668 1124 16720
rect 1176 16708 1182 16720
rect 1176 16680 1992 16708
rect 1176 16668 1182 16680
rect 661 16575 719 16581
rect 661 16541 673 16575
rect 707 16572 719 16575
rect 1854 16572 1860 16584
rect 707 16544 1860 16572
rect 707 16541 719 16544
rect 661 16535 719 16541
rect 1854 16532 1860 16544
rect 1912 16532 1918 16584
rect 1305 16439 1363 16445
rect 1305 16405 1317 16439
rect 1351 16436 1363 16439
rect 1854 16436 1860 16448
rect 1351 16408 1860 16436
rect 1351 16405 1363 16408
rect 1305 16399 1363 16405
rect 1854 16396 1860 16408
rect 1912 16396 1918 16448
rect 1964 16312 1992 16680
rect 1946 16260 1952 16312
rect 2004 16260 2010 16312
rect 1489 16099 1547 16105
rect 1489 16065 1501 16099
rect 1535 16096 1547 16099
rect 1854 16096 1860 16108
rect 1535 16068 1860 16096
rect 1535 16065 1547 16068
rect 1489 16059 1547 16065
rect 1854 16056 1860 16068
rect 1912 16056 1918 16108
rect 1394 15920 1400 15972
rect 1452 15960 1458 15972
rect 1489 15963 1547 15969
rect 1489 15960 1501 15963
rect 1452 15932 1501 15960
rect 1452 15920 1458 15932
rect 1489 15929 1501 15932
rect 1535 15929 1547 15963
rect 1489 15923 1547 15929
rect 1486 15716 1492 15768
rect 1544 15756 1550 15768
rect 1946 15756 1952 15768
rect 1544 15728 1952 15756
rect 1544 15716 1550 15728
rect 1946 15716 1952 15728
rect 2004 15716 2010 15768
rect 1118 15580 1124 15632
rect 1176 15620 1182 15632
rect 1946 15620 1952 15632
rect 1176 15592 1952 15620
rect 1176 15580 1182 15592
rect 1946 15580 1952 15592
rect 2004 15580 2010 15632
rect 569 15487 627 15493
rect 569 15453 581 15487
rect 615 15484 627 15487
rect 1946 15484 1952 15496
rect 615 15456 1952 15484
rect 615 15453 627 15456
rect 569 15447 627 15453
rect 1946 15444 1952 15456
rect 2004 15444 2010 15496
rect 1213 15351 1271 15357
rect 1213 15317 1225 15351
rect 1259 15348 1271 15351
rect 1946 15348 1952 15360
rect 1259 15320 1952 15348
rect 1259 15317 1271 15320
rect 1213 15311 1271 15317
rect 1946 15308 1952 15320
rect 2004 15308 2010 15360
rect 1121 15215 1179 15221
rect 1121 15181 1133 15215
rect 1167 15212 1179 15215
rect 1167 15184 1992 15212
rect 1167 15181 1179 15184
rect 1121 15175 1179 15181
rect 1964 15156 1992 15184
rect 1486 15104 1492 15156
rect 1544 15144 1550 15156
rect 1544 15116 1900 15144
rect 1544 15104 1550 15116
rect 1486 14968 1492 15020
rect 1544 15008 1550 15020
rect 1762 15008 1768 15020
rect 1544 14980 1768 15008
rect 1544 14968 1550 14980
rect 1762 14968 1768 14980
rect 1820 14968 1826 15020
rect 1872 14816 1900 15116
rect 1946 15104 1952 15156
rect 2004 15104 2010 15156
rect 571610 15104 571616 15156
rect 571668 15144 571674 15156
rect 580166 15144 580172 15156
rect 571668 15116 580172 15144
rect 571668 15104 571674 15116
rect 580166 15104 580172 15116
rect 580224 15104 580230 15156
rect 1118 14804 1124 14816
rect 1079 14776 1124 14804
rect 1118 14764 1124 14776
rect 1176 14764 1182 14816
rect 1854 14764 1860 14816
rect 1912 14764 1918 14816
rect 570049 14739 570107 14745
rect 570049 14705 570061 14739
rect 570095 14736 570107 14739
rect 570322 14736 570328 14748
rect 570095 14708 570328 14736
rect 570095 14705 570107 14708
rect 570049 14699 570107 14705
rect 570322 14696 570328 14708
rect 570380 14696 570386 14748
rect 1118 14628 1124 14680
rect 1176 14668 1182 14680
rect 1489 14671 1547 14677
rect 1489 14668 1501 14671
rect 1176 14640 1501 14668
rect 1176 14628 1182 14640
rect 1489 14637 1501 14640
rect 1535 14637 1547 14671
rect 1489 14631 1547 14637
rect 1029 14603 1087 14609
rect 1029 14569 1041 14603
rect 1075 14600 1087 14603
rect 1075 14572 1164 14600
rect 1075 14569 1087 14572
rect 1029 14563 1087 14569
rect 1136 14473 1164 14572
rect 1121 14467 1179 14473
rect 1121 14433 1133 14467
rect 1167 14433 1179 14467
rect 1121 14427 1179 14433
rect 1213 13515 1271 13521
rect 1213 13481 1225 13515
rect 1259 13512 1271 13515
rect 1946 13512 1952 13524
rect 1259 13484 1952 13512
rect 1259 13481 1271 13484
rect 1213 13475 1271 13481
rect 1946 13472 1952 13484
rect 2004 13472 2010 13524
rect 1029 13379 1087 13385
rect 1029 13345 1041 13379
rect 1075 13376 1087 13379
rect 1946 13376 1952 13388
rect 1075 13348 1952 13376
rect 1075 13345 1087 13348
rect 1029 13339 1087 13345
rect 1946 13336 1952 13348
rect 2004 13336 2010 13388
rect 1118 12996 1124 13048
rect 1176 13036 1182 13048
rect 1946 13036 1952 13048
rect 1176 13008 1952 13036
rect 1176 12996 1182 13008
rect 1946 12996 1952 13008
rect 2004 12996 2010 13048
rect 1118 12792 1124 12844
rect 1176 12832 1182 12844
rect 1946 12832 1952 12844
rect 1176 12804 1952 12832
rect 1176 12792 1182 12804
rect 1946 12792 1952 12804
rect 2004 12792 2010 12844
rect 1486 12452 1492 12504
rect 1544 12492 1550 12504
rect 1946 12492 1952 12504
rect 1544 12464 1952 12492
rect 1544 12452 1550 12464
rect 1946 12452 1952 12464
rect 2004 12452 2010 12504
rect 1118 12316 1124 12368
rect 1176 12356 1182 12368
rect 1305 12359 1363 12365
rect 1305 12356 1317 12359
rect 1176 12328 1317 12356
rect 1176 12316 1182 12328
rect 1305 12325 1317 12328
rect 1351 12325 1363 12359
rect 1305 12319 1363 12325
rect 1397 12359 1455 12365
rect 1397 12325 1409 12359
rect 1443 12356 1455 12359
rect 1765 12359 1823 12365
rect 1765 12356 1777 12359
rect 1443 12328 1777 12356
rect 1443 12325 1455 12328
rect 1397 12319 1455 12325
rect 1765 12325 1777 12328
rect 1811 12325 1823 12359
rect 1765 12319 1823 12325
rect 1302 12180 1308 12232
rect 1360 12220 1366 12232
rect 1765 12223 1823 12229
rect 1765 12220 1777 12223
rect 1360 12192 1777 12220
rect 1360 12180 1366 12192
rect 1765 12189 1777 12192
rect 1811 12189 1823 12223
rect 1765 12183 1823 12189
rect 753 12087 811 12093
rect 753 12053 765 12087
rect 799 12084 811 12087
rect 1302 12084 1308 12096
rect 799 12056 1308 12084
rect 799 12053 811 12056
rect 753 12047 811 12053
rect 1302 12044 1308 12056
rect 1360 12044 1366 12096
rect 842 11840 848 11892
rect 900 11880 906 11892
rect 1305 11883 1363 11889
rect 1305 11880 1317 11883
rect 900 11852 1317 11880
rect 900 11840 906 11852
rect 1305 11849 1317 11852
rect 1351 11849 1363 11883
rect 1305 11843 1363 11849
rect 842 10480 848 10532
rect 900 10520 906 10532
rect 1397 10523 1455 10529
rect 1397 10520 1409 10523
rect 900 10492 1409 10520
rect 900 10480 906 10492
rect 1397 10489 1409 10492
rect 1443 10489 1455 10523
rect 1397 10483 1455 10489
rect 753 10455 811 10461
rect 753 10421 765 10455
rect 799 10452 811 10455
rect 1581 10455 1639 10461
rect 1581 10452 1593 10455
rect 799 10424 1593 10452
rect 799 10421 811 10424
rect 753 10415 811 10421
rect 1581 10421 1593 10424
rect 1627 10421 1639 10455
rect 1581 10415 1639 10421
rect 566 10384 572 10396
rect 527 10356 572 10384
rect 566 10344 572 10356
rect 624 10344 630 10396
rect 658 10344 664 10396
rect 716 10344 722 10396
rect 1026 10384 1032 10396
rect 987 10356 1032 10384
rect 1026 10344 1032 10356
rect 1084 10344 1090 10396
rect 1397 10387 1455 10393
rect 1397 10353 1409 10387
rect 1443 10384 1455 10387
rect 1673 10387 1731 10393
rect 1673 10384 1685 10387
rect 1443 10356 1685 10384
rect 1443 10353 1455 10356
rect 1397 10347 1455 10353
rect 1673 10353 1685 10356
rect 1719 10353 1731 10387
rect 1673 10347 1731 10353
rect 474 10140 480 10192
rect 532 10180 538 10192
rect 676 10180 704 10344
rect 845 10319 903 10325
rect 845 10285 857 10319
rect 891 10316 903 10319
rect 1581 10319 1639 10325
rect 1581 10316 1593 10319
rect 891 10288 1593 10316
rect 891 10285 903 10288
rect 845 10279 903 10285
rect 1581 10285 1593 10288
rect 1627 10285 1639 10319
rect 1581 10279 1639 10285
rect 934 10208 940 10260
rect 992 10248 998 10260
rect 1673 10251 1731 10257
rect 1673 10248 1685 10251
rect 992 10220 1685 10248
rect 992 10208 998 10220
rect 1673 10217 1685 10220
rect 1719 10217 1731 10251
rect 1673 10211 1731 10217
rect 532 10152 704 10180
rect 532 10140 538 10152
rect 661 10115 719 10121
rect 661 10081 673 10115
rect 707 10112 719 10115
rect 1026 10112 1032 10124
rect 707 10084 1032 10112
rect 707 10081 719 10084
rect 661 10075 719 10081
rect 1026 10072 1032 10084
rect 1084 10072 1090 10124
rect 1302 9392 1308 9444
rect 1360 9432 1366 9444
rect 1949 9435 2007 9441
rect 1949 9432 1961 9435
rect 1360 9404 1961 9432
rect 1360 9392 1366 9404
rect 1949 9401 1961 9404
rect 1995 9401 2007 9435
rect 1949 9395 2007 9401
rect 1578 8712 1584 8764
rect 1636 8752 1642 8764
rect 1949 8755 2007 8761
rect 1949 8752 1961 8755
rect 1636 8724 1961 8752
rect 1636 8712 1642 8724
rect 1949 8721 1961 8724
rect 1995 8721 2007 8755
rect 1949 8715 2007 8721
rect 474 8684 480 8696
rect 435 8656 480 8684
rect 474 8644 480 8656
rect 532 8644 538 8696
rect 569954 8576 569960 8628
rect 570012 8616 570018 8628
rect 570322 8616 570328 8628
rect 570012 8588 570328 8616
rect 570012 8576 570018 8588
rect 570322 8576 570328 8588
rect 570380 8576 570386 8628
rect 569954 8140 569960 8152
rect 569915 8112 569960 8140
rect 569954 8100 569960 8112
rect 570012 8100 570018 8152
rect 569954 7828 569960 7880
rect 570012 7868 570018 7880
rect 570325 7871 570383 7877
rect 570325 7868 570337 7871
rect 570012 7840 570337 7868
rect 570012 7828 570018 7840
rect 570325 7837 570337 7840
rect 570371 7837 570383 7871
rect 570325 7831 570383 7837
rect 842 7488 848 7540
rect 900 7528 906 7540
rect 937 7531 995 7537
rect 937 7528 949 7531
rect 900 7500 949 7528
rect 900 7488 906 7500
rect 937 7497 949 7500
rect 983 7497 995 7531
rect 937 7491 995 7497
rect 750 4700 756 4752
rect 808 4740 814 4752
rect 1946 4740 1952 4752
rect 808 4712 1952 4740
rect 808 4700 814 4712
rect 1946 4700 1952 4712
rect 2004 4700 2010 4752
rect 750 3720 756 3732
rect 711 3692 756 3720
rect 750 3680 756 3692
rect 808 3680 814 3732
rect 1854 3720 1860 3732
rect 1815 3692 1860 3720
rect 1854 3680 1860 3692
rect 1912 3680 1918 3732
rect 1210 3312 1216 3324
rect 1171 3284 1216 3312
rect 1210 3272 1216 3284
rect 1268 3272 1274 3324
rect 124306 3068 124312 3120
rect 124364 3108 124370 3120
rect 177942 3108 177948 3120
rect 124364 3080 124409 3108
rect 177903 3080 177948 3108
rect 124364 3068 124370 3080
rect 177942 3068 177948 3080
rect 178000 3068 178006 3120
rect 268378 3068 268384 3120
rect 268436 3108 268442 3120
rect 268436 3080 268481 3108
rect 268436 3068 268442 3080
rect 1486 1776 1492 1828
rect 1544 1816 1550 1828
rect 5537 1819 5595 1825
rect 5537 1816 5549 1819
rect 1544 1788 5549 1816
rect 1544 1776 1550 1788
rect 5537 1785 5549 1788
rect 5583 1785 5595 1819
rect 5537 1779 5595 1785
rect 5629 1819 5687 1825
rect 5629 1785 5641 1819
rect 5675 1816 5687 1819
rect 26973 1819 27031 1825
rect 5675 1788 26924 1816
rect 5675 1785 5687 1788
rect 5629 1779 5687 1785
rect 569 1751 627 1757
rect 569 1717 581 1751
rect 615 1748 627 1751
rect 1670 1748 1676 1760
rect 615 1720 1676 1748
rect 615 1717 627 1720
rect 569 1711 627 1717
rect 1670 1708 1676 1720
rect 1728 1708 1734 1760
rect 3697 1751 3755 1757
rect 3697 1748 3709 1751
rect 1780 1720 3709 1748
rect 1029 1683 1087 1689
rect 1029 1649 1041 1683
rect 1075 1680 1087 1683
rect 1486 1680 1492 1692
rect 1075 1652 1492 1680
rect 1075 1649 1087 1652
rect 1029 1643 1087 1649
rect 1486 1640 1492 1652
rect 1544 1640 1550 1692
rect 14 1572 20 1624
rect 72 1612 78 1624
rect 1780 1612 1808 1720
rect 3697 1717 3709 1720
rect 3743 1717 3755 1751
rect 3697 1711 3755 1717
rect 3786 1708 3792 1760
rect 3844 1748 3850 1760
rect 7650 1748 7656 1760
rect 3844 1720 7656 1748
rect 3844 1708 3850 1720
rect 7650 1708 7656 1720
rect 7708 1708 7714 1760
rect 22094 1748 22100 1760
rect 10244 1720 22100 1748
rect 2958 1640 2964 1692
rect 3016 1680 3022 1692
rect 4062 1680 4068 1692
rect 3016 1652 4068 1680
rect 3016 1640 3022 1652
rect 4062 1640 4068 1652
rect 4120 1640 4126 1692
rect 4157 1683 4215 1689
rect 4157 1649 4169 1683
rect 4203 1680 4215 1683
rect 5261 1683 5319 1689
rect 5261 1680 5273 1683
rect 4203 1652 5273 1680
rect 4203 1649 4215 1652
rect 4157 1643 4215 1649
rect 5261 1649 5273 1652
rect 5307 1649 5319 1683
rect 5442 1680 5448 1692
rect 5403 1652 5448 1680
rect 5261 1643 5319 1649
rect 5442 1640 5448 1652
rect 5500 1640 5506 1692
rect 5537 1683 5595 1689
rect 5537 1649 5549 1683
rect 5583 1680 5595 1683
rect 10137 1683 10195 1689
rect 10137 1680 10149 1683
rect 5583 1652 10149 1680
rect 5583 1649 5595 1652
rect 5537 1643 5595 1649
rect 10137 1649 10149 1652
rect 10183 1649 10195 1683
rect 10137 1643 10195 1649
rect 72 1584 1808 1612
rect 1949 1615 2007 1621
rect 72 1572 78 1584
rect 1949 1581 1961 1615
rect 1995 1612 2007 1615
rect 10244 1612 10272 1720
rect 22094 1708 22100 1720
rect 22152 1708 22158 1760
rect 22186 1708 22192 1760
rect 22244 1748 22250 1760
rect 26237 1751 26295 1757
rect 26237 1748 26249 1751
rect 22244 1720 26249 1748
rect 22244 1708 22250 1720
rect 26237 1717 26249 1720
rect 26283 1717 26295 1751
rect 26237 1711 26295 1717
rect 26418 1708 26424 1760
rect 26476 1748 26482 1760
rect 26896 1748 26924 1788
rect 26973 1785 26985 1819
rect 27019 1816 27031 1819
rect 35253 1819 35311 1825
rect 27019 1788 35204 1816
rect 27019 1785 27031 1788
rect 26973 1779 27031 1785
rect 34977 1751 35035 1757
rect 34977 1748 34989 1751
rect 26476 1720 26740 1748
rect 26896 1720 34989 1748
rect 26476 1708 26482 1720
rect 18322 1680 18328 1692
rect 1995 1584 10272 1612
rect 10336 1652 18328 1680
rect 1995 1581 2007 1584
rect 1949 1575 2007 1581
rect 1305 1547 1363 1553
rect 1305 1513 1317 1547
rect 1351 1544 1363 1547
rect 5077 1547 5135 1553
rect 5077 1544 5089 1547
rect 1351 1516 5089 1544
rect 1351 1513 1363 1516
rect 1305 1507 1363 1513
rect 5077 1513 5089 1516
rect 5123 1513 5135 1547
rect 5077 1507 5135 1513
rect 5169 1547 5227 1553
rect 5169 1513 5181 1547
rect 5215 1544 5227 1547
rect 10336 1544 10364 1652
rect 18322 1640 18328 1652
rect 18380 1640 18386 1692
rect 19334 1640 19340 1692
rect 19392 1680 19398 1692
rect 25133 1683 25191 1689
rect 25133 1680 25145 1683
rect 19392 1652 25145 1680
rect 19392 1640 19398 1652
rect 25133 1649 25145 1652
rect 25179 1649 25191 1683
rect 25133 1643 25191 1649
rect 25777 1683 25835 1689
rect 25777 1649 25789 1683
rect 25823 1680 25835 1683
rect 26602 1680 26608 1692
rect 25823 1652 26608 1680
rect 25823 1649 25835 1652
rect 25777 1643 25835 1649
rect 26602 1640 26608 1652
rect 26660 1640 26666 1692
rect 26712 1680 26740 1720
rect 34977 1717 34989 1720
rect 35023 1717 35035 1751
rect 34977 1711 35035 1717
rect 26973 1683 27031 1689
rect 26973 1680 26985 1683
rect 26712 1652 26985 1680
rect 26973 1649 26985 1652
rect 27019 1649 27031 1683
rect 26973 1643 27031 1649
rect 27065 1683 27123 1689
rect 27065 1649 27077 1683
rect 27111 1680 27123 1683
rect 35069 1683 35127 1689
rect 35069 1680 35081 1683
rect 27111 1652 35081 1680
rect 27111 1649 27123 1652
rect 27065 1643 27123 1649
rect 35069 1649 35081 1652
rect 35115 1649 35127 1683
rect 35176 1680 35204 1788
rect 35253 1785 35265 1819
rect 35299 1816 35311 1819
rect 39577 1819 39635 1825
rect 39577 1816 39589 1819
rect 35299 1788 39589 1816
rect 35299 1785 35311 1788
rect 35253 1779 35311 1785
rect 39577 1785 39589 1788
rect 39623 1785 39635 1819
rect 39577 1779 39635 1785
rect 39669 1819 39727 1825
rect 39669 1785 39681 1819
rect 39715 1816 39727 1819
rect 48961 1819 49019 1825
rect 39715 1788 48912 1816
rect 39715 1785 39727 1788
rect 39669 1779 39727 1785
rect 48884 1760 48912 1788
rect 48961 1785 48973 1819
rect 49007 1816 49019 1819
rect 56781 1819 56839 1825
rect 49007 1788 56456 1816
rect 49007 1785 49019 1788
rect 48961 1779 49019 1785
rect 56428 1760 56456 1788
rect 56781 1785 56793 1819
rect 56827 1816 56839 1819
rect 65429 1819 65487 1825
rect 65429 1816 65441 1819
rect 56827 1788 65441 1816
rect 56827 1785 56839 1788
rect 56781 1779 56839 1785
rect 65429 1785 65441 1788
rect 65475 1785 65487 1819
rect 65429 1779 65487 1785
rect 65521 1819 65579 1825
rect 65521 1785 65533 1819
rect 65567 1816 65579 1819
rect 106001 1819 106059 1825
rect 106001 1816 106013 1819
rect 65567 1788 106013 1816
rect 65567 1785 65579 1788
rect 65521 1779 65579 1785
rect 106001 1785 106013 1788
rect 106047 1785 106059 1819
rect 106001 1779 106059 1785
rect 106093 1819 106151 1825
rect 106093 1785 106105 1819
rect 106139 1816 106151 1819
rect 106829 1819 106887 1825
rect 106829 1816 106841 1819
rect 106139 1788 106841 1816
rect 106139 1785 106151 1788
rect 106093 1779 106151 1785
rect 106829 1785 106841 1788
rect 106875 1785 106887 1819
rect 116121 1819 116179 1825
rect 116121 1816 116133 1819
rect 106829 1779 106887 1785
rect 106936 1788 116133 1816
rect 35345 1751 35403 1757
rect 35345 1717 35357 1751
rect 35391 1748 35403 1751
rect 35391 1720 45692 1748
rect 35391 1717 35403 1720
rect 35345 1711 35403 1717
rect 37734 1680 37740 1692
rect 35176 1652 37740 1680
rect 35069 1643 35127 1649
rect 37734 1640 37740 1652
rect 37792 1640 37798 1692
rect 38013 1683 38071 1689
rect 38013 1649 38025 1683
rect 38059 1680 38071 1683
rect 39022 1680 39028 1692
rect 38059 1652 39028 1680
rect 38059 1649 38071 1652
rect 38013 1643 38071 1649
rect 39022 1640 39028 1652
rect 39080 1640 39086 1692
rect 39117 1683 39175 1689
rect 39117 1649 39129 1683
rect 39163 1680 39175 1683
rect 42702 1680 42708 1692
rect 39163 1652 42708 1680
rect 39163 1649 39175 1652
rect 39117 1643 39175 1649
rect 42702 1640 42708 1652
rect 42760 1640 42766 1692
rect 45554 1680 45560 1692
rect 42812 1652 45560 1680
rect 10410 1572 10416 1624
rect 10468 1612 10474 1624
rect 11149 1615 11207 1621
rect 11149 1612 11161 1615
rect 10468 1584 11161 1612
rect 10468 1572 10474 1584
rect 11149 1581 11161 1584
rect 11195 1581 11207 1615
rect 11149 1575 11207 1581
rect 11241 1615 11299 1621
rect 11241 1581 11253 1615
rect 11287 1612 11299 1615
rect 42429 1615 42487 1621
rect 42429 1612 42441 1615
rect 11287 1584 42441 1612
rect 11287 1581 11299 1584
rect 11241 1575 11299 1581
rect 42429 1581 42441 1584
rect 42475 1581 42487 1615
rect 42429 1575 42487 1581
rect 42518 1572 42524 1624
rect 42576 1612 42582 1624
rect 42812 1612 42840 1652
rect 45554 1640 45560 1652
rect 45612 1640 45618 1692
rect 45664 1680 45692 1720
rect 48682 1708 48688 1760
rect 48740 1748 48746 1760
rect 48740 1720 48785 1748
rect 48740 1708 48746 1720
rect 48866 1708 48872 1760
rect 48924 1708 48930 1760
rect 49053 1751 49111 1757
rect 49053 1717 49065 1751
rect 49099 1748 49111 1751
rect 50614 1748 50620 1760
rect 49099 1720 50620 1748
rect 49099 1717 49111 1720
rect 49053 1711 49111 1717
rect 50614 1708 50620 1720
rect 50672 1708 50678 1760
rect 50798 1748 50804 1760
rect 50759 1720 50804 1748
rect 50798 1708 50804 1720
rect 50856 1708 50862 1760
rect 50985 1751 51043 1757
rect 50985 1717 50997 1751
rect 51031 1748 51043 1751
rect 51031 1720 56364 1748
rect 51031 1717 51043 1720
rect 50985 1711 51043 1717
rect 55769 1683 55827 1689
rect 55769 1680 55781 1683
rect 45664 1652 55781 1680
rect 55769 1649 55781 1652
rect 55815 1649 55827 1683
rect 56336 1680 56364 1720
rect 56410 1708 56416 1760
rect 56468 1708 56474 1760
rect 56686 1708 56692 1760
rect 56744 1748 56750 1760
rect 106936 1748 106964 1788
rect 116121 1785 116133 1788
rect 116167 1785 116179 1819
rect 116121 1779 116179 1785
rect 116213 1819 116271 1825
rect 116213 1785 116225 1819
rect 116259 1816 116271 1819
rect 125597 1819 125655 1825
rect 125597 1816 125609 1819
rect 116259 1788 125609 1816
rect 116259 1785 116271 1788
rect 116213 1779 116271 1785
rect 125597 1785 125609 1788
rect 125643 1785 125655 1819
rect 125597 1779 125655 1785
rect 125689 1819 125747 1825
rect 125689 1785 125701 1819
rect 125735 1816 125747 1819
rect 128449 1819 128507 1825
rect 128449 1816 128461 1819
rect 125735 1788 128461 1816
rect 125735 1785 125747 1788
rect 125689 1779 125747 1785
rect 128449 1785 128461 1788
rect 128495 1785 128507 1819
rect 130473 1819 130531 1825
rect 128449 1779 128507 1785
rect 128556 1788 130424 1816
rect 56744 1720 106964 1748
rect 107013 1751 107071 1757
rect 56744 1708 56750 1720
rect 107013 1717 107025 1751
rect 107059 1748 107071 1751
rect 111613 1751 111671 1757
rect 111613 1748 111625 1751
rect 107059 1720 111625 1748
rect 107059 1717 107071 1720
rect 107013 1711 107071 1717
rect 111613 1717 111625 1720
rect 111659 1717 111671 1751
rect 111613 1711 111671 1717
rect 111978 1708 111984 1760
rect 112036 1748 112042 1760
rect 121549 1751 121607 1757
rect 112036 1720 121500 1748
rect 112036 1708 112042 1720
rect 56597 1683 56655 1689
rect 56597 1680 56609 1683
rect 56336 1652 56609 1680
rect 55769 1643 55827 1649
rect 56597 1649 56609 1652
rect 56643 1649 56655 1683
rect 56597 1643 56655 1649
rect 56778 1640 56784 1692
rect 56836 1680 56842 1692
rect 56836 1652 56881 1680
rect 56836 1640 56842 1652
rect 57882 1640 57888 1692
rect 57940 1680 57946 1692
rect 63221 1683 63279 1689
rect 63221 1680 63233 1683
rect 57940 1652 63233 1680
rect 57940 1640 57946 1652
rect 63221 1649 63233 1652
rect 63267 1649 63279 1683
rect 63221 1643 63279 1649
rect 63313 1683 63371 1689
rect 63313 1649 63325 1683
rect 63359 1680 63371 1683
rect 71774 1680 71780 1692
rect 63359 1652 71780 1680
rect 63359 1649 63371 1652
rect 63313 1643 63371 1649
rect 71774 1640 71780 1652
rect 71832 1640 71838 1692
rect 71869 1683 71927 1689
rect 71869 1649 71881 1683
rect 71915 1680 71927 1683
rect 121365 1683 121423 1689
rect 121365 1680 121377 1683
rect 71915 1652 121377 1680
rect 71915 1649 71927 1652
rect 71869 1643 71927 1649
rect 121365 1649 121377 1652
rect 121411 1649 121423 1683
rect 121472 1680 121500 1720
rect 121549 1717 121561 1751
rect 121595 1748 121607 1751
rect 128081 1751 128139 1757
rect 128081 1748 128093 1751
rect 121595 1720 128093 1748
rect 121595 1717 121607 1720
rect 121549 1711 121607 1717
rect 128081 1717 128093 1720
rect 128127 1717 128139 1751
rect 128262 1748 128268 1760
rect 128223 1720 128268 1748
rect 128081 1711 128139 1717
rect 128262 1708 128268 1720
rect 128320 1708 128326 1760
rect 124582 1680 124588 1692
rect 121472 1652 124588 1680
rect 121365 1643 121423 1649
rect 124582 1640 124588 1652
rect 124640 1640 124646 1692
rect 124677 1683 124735 1689
rect 124677 1649 124689 1683
rect 124723 1680 124735 1683
rect 125597 1683 125655 1689
rect 124723 1652 125456 1680
rect 124723 1649 124735 1652
rect 124677 1643 124735 1649
rect 42576 1584 42840 1612
rect 42889 1615 42947 1621
rect 42576 1572 42582 1584
rect 42889 1581 42901 1615
rect 42935 1612 42947 1615
rect 48961 1615 49019 1621
rect 48961 1612 48973 1615
rect 42935 1584 48973 1612
rect 42935 1581 42947 1584
rect 42889 1575 42947 1581
rect 48961 1581 48973 1584
rect 49007 1581 49019 1615
rect 48961 1575 49019 1581
rect 49053 1615 49111 1621
rect 49053 1581 49065 1615
rect 49099 1612 49111 1615
rect 111245 1615 111303 1621
rect 111245 1612 111257 1615
rect 49099 1584 111257 1612
rect 49099 1581 49111 1584
rect 49053 1575 49111 1581
rect 111245 1581 111257 1584
rect 111291 1581 111303 1615
rect 111245 1575 111303 1581
rect 111334 1572 111340 1624
rect 111392 1612 111398 1624
rect 111429 1615 111487 1621
rect 111429 1612 111441 1615
rect 111392 1584 111441 1612
rect 111392 1572 111398 1584
rect 111429 1581 111441 1584
rect 111475 1581 111487 1615
rect 111429 1575 111487 1581
rect 111797 1615 111855 1621
rect 111797 1581 111809 1615
rect 111843 1612 111855 1615
rect 112162 1612 112168 1624
rect 111843 1584 112168 1612
rect 111843 1581 111855 1584
rect 111797 1575 111855 1581
rect 112162 1572 112168 1584
rect 112220 1572 112226 1624
rect 112349 1615 112407 1621
rect 112349 1581 112361 1615
rect 112395 1612 112407 1615
rect 115109 1615 115167 1621
rect 115109 1612 115121 1615
rect 112395 1584 115121 1612
rect 112395 1581 112407 1584
rect 112349 1575 112407 1581
rect 115109 1581 115121 1584
rect 115155 1581 115167 1615
rect 115109 1575 115167 1581
rect 115198 1572 115204 1624
rect 115256 1612 115262 1624
rect 116489 1615 116547 1621
rect 116489 1612 116501 1615
rect 115256 1584 116501 1612
rect 115256 1572 115262 1584
rect 116489 1581 116501 1584
rect 116535 1581 116547 1615
rect 116489 1575 116547 1581
rect 116581 1615 116639 1621
rect 116581 1581 116593 1615
rect 116627 1612 116639 1615
rect 125321 1615 125379 1621
rect 125321 1612 125333 1615
rect 116627 1584 125333 1612
rect 116627 1581 116639 1584
rect 116581 1575 116639 1581
rect 125321 1581 125333 1584
rect 125367 1581 125379 1615
rect 125428 1612 125456 1652
rect 125597 1649 125609 1683
rect 125643 1680 125655 1683
rect 128556 1680 128584 1788
rect 129553 1751 129611 1757
rect 128648 1720 129504 1748
rect 128648 1689 128676 1720
rect 125643 1652 128584 1680
rect 128633 1683 128691 1689
rect 125643 1649 125655 1652
rect 125597 1643 125655 1649
rect 128633 1649 128645 1683
rect 128679 1649 128691 1683
rect 129369 1683 129427 1689
rect 129369 1680 129381 1683
rect 128633 1643 128691 1649
rect 128740 1652 129381 1680
rect 125689 1615 125747 1621
rect 125689 1612 125701 1615
rect 125428 1584 125701 1612
rect 125321 1575 125379 1581
rect 125689 1581 125701 1584
rect 125735 1581 125747 1615
rect 125689 1575 125747 1581
rect 125778 1572 125784 1624
rect 125836 1612 125842 1624
rect 125965 1615 126023 1621
rect 125965 1612 125977 1615
rect 125836 1584 125977 1612
rect 125836 1572 125842 1584
rect 125965 1581 125977 1584
rect 126011 1581 126023 1615
rect 125965 1575 126023 1581
rect 126057 1615 126115 1621
rect 126057 1581 126069 1615
rect 126103 1612 126115 1615
rect 127345 1615 127403 1621
rect 127345 1612 127357 1615
rect 126103 1584 127357 1612
rect 126103 1581 126115 1584
rect 126057 1575 126115 1581
rect 127345 1581 127357 1584
rect 127391 1581 127403 1615
rect 127345 1575 127403 1581
rect 127437 1615 127495 1621
rect 127437 1581 127449 1615
rect 127483 1612 127495 1615
rect 128081 1615 128139 1621
rect 128081 1612 128093 1615
rect 127483 1584 128093 1612
rect 127483 1581 127495 1584
rect 127437 1575 127495 1581
rect 128081 1581 128093 1584
rect 128127 1581 128139 1615
rect 128081 1575 128139 1581
rect 128173 1615 128231 1621
rect 128173 1581 128185 1615
rect 128219 1612 128231 1615
rect 128740 1612 128768 1652
rect 129369 1649 129381 1652
rect 129415 1649 129427 1683
rect 129476 1680 129504 1720
rect 129553 1717 129565 1751
rect 129599 1748 129611 1751
rect 130289 1751 130347 1757
rect 130289 1748 130301 1751
rect 129599 1720 130301 1748
rect 129599 1717 129611 1720
rect 129553 1711 129611 1717
rect 130289 1717 130301 1720
rect 130335 1717 130347 1751
rect 130396 1748 130424 1788
rect 130473 1785 130485 1819
rect 130519 1816 130531 1819
rect 134245 1819 134303 1825
rect 134245 1816 134257 1819
rect 130519 1788 134257 1816
rect 130519 1785 130531 1788
rect 130473 1779 130531 1785
rect 134245 1785 134257 1788
rect 134291 1785 134303 1819
rect 134245 1779 134303 1785
rect 134337 1819 134395 1825
rect 134337 1785 134349 1819
rect 134383 1816 134395 1819
rect 134613 1819 134671 1825
rect 134383 1788 134564 1816
rect 134383 1785 134395 1788
rect 134337 1779 134395 1785
rect 134429 1751 134487 1757
rect 134429 1748 134441 1751
rect 130396 1720 134441 1748
rect 130289 1711 130347 1717
rect 134429 1717 134441 1720
rect 134475 1717 134487 1751
rect 134536 1748 134564 1788
rect 134613 1785 134625 1819
rect 134659 1816 134671 1819
rect 146849 1819 146907 1825
rect 146849 1816 146861 1819
rect 134659 1788 146861 1816
rect 134659 1785 134671 1788
rect 134613 1779 134671 1785
rect 146849 1785 146861 1788
rect 146895 1785 146907 1819
rect 146849 1779 146907 1785
rect 147125 1819 147183 1825
rect 147125 1785 147137 1819
rect 147171 1785 147183 1819
rect 147125 1779 147183 1785
rect 147217 1819 147275 1825
rect 147217 1785 147229 1819
rect 147263 1816 147275 1819
rect 147861 1819 147919 1825
rect 147861 1816 147873 1819
rect 147263 1788 147873 1816
rect 147263 1785 147275 1788
rect 147217 1779 147275 1785
rect 147861 1785 147873 1788
rect 147907 1785 147919 1819
rect 147861 1779 147919 1785
rect 147953 1819 148011 1825
rect 147953 1785 147965 1819
rect 147999 1785 148011 1819
rect 147953 1779 148011 1785
rect 148045 1819 148103 1825
rect 148045 1785 148057 1819
rect 148091 1816 148103 1819
rect 148505 1819 148563 1825
rect 148505 1816 148517 1819
rect 148091 1788 148517 1816
rect 148091 1785 148103 1788
rect 148045 1779 148103 1785
rect 148505 1785 148517 1788
rect 148551 1785 148563 1819
rect 149057 1819 149115 1825
rect 149057 1816 149069 1819
rect 148505 1779 148563 1785
rect 148612 1788 149069 1816
rect 134536 1720 138888 1748
rect 134429 1711 134487 1717
rect 134518 1680 134524 1692
rect 129476 1652 134524 1680
rect 129369 1643 129427 1649
rect 134518 1640 134524 1652
rect 134576 1640 134582 1692
rect 134613 1683 134671 1689
rect 134613 1649 134625 1683
rect 134659 1680 134671 1683
rect 135073 1683 135131 1689
rect 135073 1680 135085 1683
rect 134659 1652 135085 1680
rect 134659 1649 134671 1652
rect 134613 1643 134671 1649
rect 135073 1649 135085 1652
rect 135119 1649 135131 1683
rect 135073 1643 135131 1649
rect 135162 1640 135168 1692
rect 135220 1680 135226 1692
rect 137186 1680 137192 1692
rect 135220 1652 137192 1680
rect 135220 1640 135226 1652
rect 137186 1640 137192 1652
rect 137244 1640 137250 1692
rect 137281 1683 137339 1689
rect 137281 1649 137293 1683
rect 137327 1680 137339 1683
rect 138290 1680 138296 1692
rect 137327 1652 138296 1680
rect 137327 1649 137339 1652
rect 137281 1643 137339 1649
rect 138290 1640 138296 1652
rect 138348 1640 138354 1692
rect 138382 1640 138388 1692
rect 138440 1680 138446 1692
rect 138477 1683 138535 1689
rect 138477 1680 138489 1683
rect 138440 1652 138489 1680
rect 138440 1640 138446 1652
rect 138477 1649 138489 1652
rect 138523 1649 138535 1683
rect 138477 1643 138535 1649
rect 138569 1683 138627 1689
rect 138569 1649 138581 1683
rect 138615 1680 138627 1683
rect 138750 1680 138756 1692
rect 138615 1652 138756 1680
rect 138615 1649 138627 1652
rect 138569 1643 138627 1649
rect 138750 1640 138756 1652
rect 138808 1640 138814 1692
rect 138860 1680 138888 1720
rect 138934 1708 138940 1760
rect 138992 1748 138998 1760
rect 140501 1751 140559 1757
rect 138992 1720 140452 1748
rect 138992 1708 138998 1720
rect 140317 1683 140375 1689
rect 140317 1680 140329 1683
rect 138860 1652 140329 1680
rect 140317 1649 140329 1652
rect 140363 1649 140375 1683
rect 140424 1680 140452 1720
rect 140501 1717 140513 1751
rect 140547 1748 140559 1751
rect 141605 1751 141663 1757
rect 141605 1748 141617 1751
rect 140547 1720 141617 1748
rect 140547 1717 140559 1720
rect 140501 1711 140559 1717
rect 141605 1717 141617 1720
rect 141651 1717 141663 1751
rect 141605 1711 141663 1717
rect 141697 1751 141755 1757
rect 141697 1717 141709 1751
rect 141743 1748 141755 1751
rect 144825 1751 144883 1757
rect 144825 1748 144837 1751
rect 141743 1720 144837 1748
rect 141743 1717 141755 1720
rect 141697 1711 141755 1717
rect 144825 1717 144837 1720
rect 144871 1717 144883 1751
rect 144825 1711 144883 1717
rect 145558 1708 145564 1760
rect 145616 1748 145622 1760
rect 145834 1748 145840 1760
rect 145616 1720 145840 1748
rect 145616 1708 145622 1720
rect 145834 1708 145840 1720
rect 145892 1708 145898 1760
rect 146202 1708 146208 1760
rect 146260 1748 146266 1760
rect 147030 1748 147036 1760
rect 146260 1720 147036 1748
rect 146260 1708 146266 1720
rect 147030 1708 147036 1720
rect 147088 1708 147094 1760
rect 147140 1748 147168 1779
rect 147968 1748 147996 1779
rect 148612 1760 148640 1788
rect 149057 1785 149069 1788
rect 149103 1785 149115 1819
rect 149057 1779 149115 1785
rect 149149 1819 149207 1825
rect 149149 1785 149161 1819
rect 149195 1785 149207 1819
rect 150253 1819 150311 1825
rect 150253 1816 150265 1819
rect 149149 1779 149207 1785
rect 149256 1788 150265 1816
rect 147140 1720 147996 1748
rect 148318 1708 148324 1760
rect 148376 1748 148382 1760
rect 148413 1751 148471 1757
rect 148413 1748 148425 1751
rect 148376 1720 148425 1748
rect 148376 1708 148382 1720
rect 148413 1717 148425 1720
rect 148459 1717 148471 1751
rect 148413 1711 148471 1717
rect 148594 1708 148600 1760
rect 148652 1708 148658 1760
rect 148965 1751 149023 1757
rect 148965 1717 148977 1751
rect 149011 1748 149023 1751
rect 149164 1748 149192 1779
rect 149256 1760 149284 1788
rect 150253 1785 150265 1788
rect 150299 1785 150311 1819
rect 150253 1779 150311 1785
rect 150345 1819 150403 1825
rect 150345 1785 150357 1819
rect 150391 1816 150403 1819
rect 151449 1819 151507 1825
rect 151449 1816 151461 1819
rect 150391 1788 151461 1816
rect 150391 1785 150403 1788
rect 150345 1779 150403 1785
rect 151449 1785 151461 1788
rect 151495 1785 151507 1819
rect 151449 1779 151507 1785
rect 151633 1819 151691 1825
rect 151633 1785 151645 1819
rect 151679 1816 151691 1819
rect 152277 1819 152335 1825
rect 152277 1816 152289 1819
rect 151679 1788 152289 1816
rect 151679 1785 151691 1788
rect 151633 1779 151691 1785
rect 152277 1785 152289 1788
rect 152323 1785 152335 1819
rect 152277 1779 152335 1785
rect 152369 1819 152427 1825
rect 152369 1785 152381 1819
rect 152415 1816 152427 1819
rect 153289 1819 153347 1825
rect 153289 1816 153301 1819
rect 152415 1788 153301 1816
rect 152415 1785 152427 1788
rect 152369 1779 152427 1785
rect 153289 1785 153301 1788
rect 153335 1785 153347 1819
rect 153289 1779 153347 1785
rect 153381 1819 153439 1825
rect 153381 1785 153393 1819
rect 153427 1816 153439 1819
rect 154209 1819 154267 1825
rect 154209 1816 154221 1819
rect 153427 1788 154221 1816
rect 153427 1785 153439 1788
rect 153381 1779 153439 1785
rect 154209 1785 154221 1788
rect 154255 1785 154267 1819
rect 154209 1779 154267 1785
rect 154485 1819 154543 1825
rect 154485 1785 154497 1819
rect 154531 1816 154543 1819
rect 156141 1819 156199 1825
rect 156141 1816 156153 1819
rect 154531 1788 156153 1816
rect 154531 1785 154543 1788
rect 154485 1779 154543 1785
rect 156141 1785 156153 1788
rect 156187 1785 156199 1819
rect 156509 1819 156567 1825
rect 156509 1816 156521 1819
rect 156141 1779 156199 1785
rect 156248 1788 156521 1816
rect 149011 1720 149192 1748
rect 149011 1717 149023 1720
rect 148965 1711 149023 1717
rect 149238 1708 149244 1760
rect 149296 1708 149302 1760
rect 149330 1708 149336 1760
rect 149388 1748 149394 1760
rect 149974 1748 149980 1760
rect 149388 1720 149980 1748
rect 149388 1708 149394 1720
rect 149974 1708 149980 1720
rect 150032 1708 150038 1760
rect 150069 1751 150127 1757
rect 150069 1717 150081 1751
rect 150115 1748 150127 1751
rect 150437 1751 150495 1757
rect 150115 1720 150296 1748
rect 150115 1717 150127 1720
rect 150069 1711 150127 1717
rect 140869 1683 140927 1689
rect 140869 1680 140881 1683
rect 140424 1652 140881 1680
rect 140317 1643 140375 1649
rect 140869 1649 140881 1652
rect 140915 1649 140927 1683
rect 150158 1680 150164 1692
rect 140869 1643 140927 1649
rect 140976 1652 150164 1680
rect 128219 1584 128768 1612
rect 128219 1581 128231 1584
rect 128173 1575 128231 1581
rect 128814 1572 128820 1624
rect 128872 1612 128878 1624
rect 136545 1615 136603 1621
rect 136545 1612 136557 1615
rect 128872 1584 136557 1612
rect 128872 1572 128878 1584
rect 136545 1581 136557 1584
rect 136591 1581 136603 1615
rect 136545 1575 136603 1581
rect 137005 1615 137063 1621
rect 137005 1581 137017 1615
rect 137051 1612 137063 1615
rect 140976 1612 141004 1652
rect 150158 1640 150164 1652
rect 150216 1640 150222 1692
rect 150268 1680 150296 1720
rect 150437 1717 150449 1751
rect 150483 1748 150495 1751
rect 151265 1751 151323 1757
rect 151265 1748 151277 1751
rect 150483 1720 151277 1748
rect 150483 1717 150495 1720
rect 150437 1711 150495 1717
rect 151265 1717 151277 1720
rect 151311 1717 151323 1751
rect 151265 1711 151323 1717
rect 151357 1751 151415 1757
rect 151357 1717 151369 1751
rect 151403 1748 151415 1751
rect 152001 1751 152059 1757
rect 152001 1748 152013 1751
rect 151403 1720 152013 1748
rect 151403 1717 151415 1720
rect 151357 1711 151415 1717
rect 152001 1717 152013 1720
rect 152047 1717 152059 1751
rect 152001 1711 152059 1717
rect 152093 1751 152151 1757
rect 152093 1717 152105 1751
rect 152139 1748 152151 1751
rect 156248 1748 156276 1788
rect 156509 1785 156521 1788
rect 156555 1785 156567 1819
rect 157245 1819 157303 1825
rect 157245 1816 157257 1819
rect 156509 1779 156567 1785
rect 156616 1788 157257 1816
rect 152139 1720 156276 1748
rect 156325 1751 156383 1757
rect 152139 1717 152151 1720
rect 152093 1711 152151 1717
rect 156325 1717 156337 1751
rect 156371 1748 156383 1751
rect 156616 1748 156644 1788
rect 157245 1785 157257 1788
rect 157291 1785 157303 1819
rect 170033 1819 170091 1825
rect 170033 1816 170045 1819
rect 157245 1779 157303 1785
rect 157352 1788 170045 1816
rect 156371 1720 156644 1748
rect 156371 1717 156383 1720
rect 156325 1711 156383 1717
rect 156782 1708 156788 1760
rect 156840 1748 156846 1760
rect 157352 1748 157380 1788
rect 170033 1785 170045 1788
rect 170079 1785 170091 1819
rect 175553 1819 175611 1825
rect 175553 1816 175565 1819
rect 170033 1779 170091 1785
rect 170140 1788 175565 1816
rect 156840 1720 157380 1748
rect 157429 1751 157487 1757
rect 156840 1708 156846 1720
rect 157429 1717 157441 1751
rect 157475 1748 157487 1751
rect 157797 1751 157855 1757
rect 157475 1720 157748 1748
rect 157475 1717 157487 1720
rect 157429 1711 157487 1717
rect 150268 1652 150572 1680
rect 137051 1584 141004 1612
rect 141053 1615 141111 1621
rect 137051 1581 137063 1584
rect 137005 1575 137063 1581
rect 141053 1581 141065 1615
rect 141099 1612 141111 1615
rect 144730 1612 144736 1624
rect 141099 1584 144736 1612
rect 141099 1581 141111 1584
rect 141053 1575 141111 1581
rect 144730 1572 144736 1584
rect 144788 1572 144794 1624
rect 144825 1615 144883 1621
rect 144825 1581 144837 1615
rect 144871 1612 144883 1615
rect 148873 1615 148931 1621
rect 148873 1612 148885 1615
rect 144871 1584 148885 1612
rect 144871 1581 144883 1584
rect 144825 1575 144883 1581
rect 148873 1581 148885 1584
rect 148919 1581 148931 1615
rect 148873 1575 148931 1581
rect 148962 1572 148968 1624
rect 149020 1612 149026 1624
rect 149057 1615 149115 1621
rect 149057 1612 149069 1615
rect 149020 1584 149069 1612
rect 149020 1572 149026 1584
rect 149057 1581 149069 1584
rect 149103 1581 149115 1615
rect 149057 1575 149115 1581
rect 149149 1615 149207 1621
rect 149149 1581 149161 1615
rect 149195 1612 149207 1615
rect 149517 1615 149575 1621
rect 149517 1612 149529 1615
rect 149195 1584 149529 1612
rect 149195 1581 149207 1584
rect 149149 1575 149207 1581
rect 149517 1581 149529 1584
rect 149563 1581 149575 1615
rect 149517 1575 149575 1581
rect 149609 1615 149667 1621
rect 149609 1581 149621 1615
rect 149655 1612 149667 1615
rect 150437 1615 150495 1621
rect 150437 1612 150449 1615
rect 149655 1584 150449 1612
rect 149655 1581 149667 1584
rect 149609 1575 149667 1581
rect 150437 1581 150449 1584
rect 150483 1581 150495 1615
rect 150544 1612 150572 1652
rect 150618 1640 150624 1692
rect 150676 1680 150682 1692
rect 157720 1680 157748 1720
rect 157797 1717 157809 1751
rect 157843 1748 157855 1751
rect 161566 1748 161572 1760
rect 157843 1720 161572 1748
rect 157843 1717 157855 1720
rect 157797 1711 157855 1717
rect 161566 1708 161572 1720
rect 161624 1708 161630 1760
rect 161661 1751 161719 1757
rect 161661 1717 161673 1751
rect 161707 1748 161719 1751
rect 169478 1748 169484 1760
rect 161707 1720 169484 1748
rect 161707 1717 161719 1720
rect 161661 1711 161719 1717
rect 169478 1708 169484 1720
rect 169536 1708 169542 1760
rect 169665 1751 169723 1757
rect 169665 1717 169677 1751
rect 169711 1748 169723 1751
rect 170140 1748 170168 1788
rect 175553 1785 175565 1788
rect 175599 1785 175611 1819
rect 183557 1819 183615 1825
rect 183557 1816 183569 1819
rect 175553 1779 175611 1785
rect 175660 1788 183569 1816
rect 169711 1720 170168 1748
rect 170217 1751 170275 1757
rect 169711 1717 169723 1720
rect 169665 1711 169723 1717
rect 170217 1717 170229 1751
rect 170263 1748 170275 1751
rect 170950 1748 170956 1760
rect 170263 1720 170956 1748
rect 170263 1717 170275 1720
rect 170217 1711 170275 1717
rect 170950 1708 170956 1720
rect 171008 1708 171014 1760
rect 171042 1708 171048 1760
rect 171100 1748 171106 1760
rect 174173 1751 174231 1757
rect 174173 1748 174185 1751
rect 171100 1720 174185 1748
rect 171100 1708 171106 1720
rect 174173 1717 174185 1720
rect 174219 1717 174231 1751
rect 174173 1711 174231 1717
rect 174262 1708 174268 1760
rect 174320 1748 174326 1760
rect 175274 1748 175280 1760
rect 174320 1720 175280 1748
rect 174320 1708 174326 1720
rect 175274 1708 175280 1720
rect 175332 1708 175338 1760
rect 175369 1751 175427 1757
rect 175369 1717 175381 1751
rect 175415 1748 175427 1751
rect 175660 1748 175688 1788
rect 183557 1785 183569 1788
rect 183603 1785 183615 1819
rect 220265 1819 220323 1825
rect 220265 1816 220277 1819
rect 183557 1779 183615 1785
rect 183664 1788 220277 1816
rect 175415 1720 175688 1748
rect 175737 1751 175795 1757
rect 175415 1717 175427 1720
rect 175369 1711 175427 1717
rect 175737 1717 175749 1751
rect 175783 1748 175795 1751
rect 177761 1751 177819 1757
rect 177761 1748 177773 1751
rect 175783 1720 177773 1748
rect 175783 1717 175795 1720
rect 175737 1711 175795 1717
rect 177761 1717 177773 1720
rect 177807 1717 177819 1751
rect 177761 1711 177819 1717
rect 177850 1708 177856 1760
rect 177908 1748 177914 1760
rect 178865 1751 178923 1757
rect 177908 1720 178724 1748
rect 177908 1708 177914 1720
rect 158898 1680 158904 1692
rect 150676 1652 157564 1680
rect 157720 1652 158904 1680
rect 150676 1640 150682 1652
rect 151173 1615 151231 1621
rect 151173 1612 151185 1615
rect 150544 1584 151185 1612
rect 150437 1575 150495 1581
rect 151173 1581 151185 1584
rect 151219 1581 151231 1615
rect 151541 1615 151599 1621
rect 151541 1612 151553 1615
rect 151173 1575 151231 1581
rect 151372 1584 151553 1612
rect 17954 1544 17960 1556
rect 5215 1516 10364 1544
rect 10428 1516 17960 1544
rect 5215 1513 5227 1516
rect 5169 1507 5227 1513
rect 1578 1436 1584 1488
rect 1636 1476 1642 1488
rect 3421 1479 3479 1485
rect 3421 1476 3433 1479
rect 1636 1448 3433 1476
rect 1636 1436 1642 1448
rect 3421 1445 3433 1448
rect 3467 1445 3479 1479
rect 3421 1439 3479 1445
rect 3510 1436 3516 1488
rect 3568 1476 3574 1488
rect 5353 1479 5411 1485
rect 5353 1476 5365 1479
rect 3568 1448 5365 1476
rect 3568 1436 3574 1448
rect 5353 1445 5365 1448
rect 5399 1445 5411 1479
rect 5353 1439 5411 1445
rect 5445 1479 5503 1485
rect 5445 1445 5457 1479
rect 5491 1476 5503 1479
rect 6822 1476 6828 1488
rect 5491 1448 6828 1476
rect 5491 1445 5503 1448
rect 5445 1439 5503 1445
rect 6822 1436 6828 1448
rect 6880 1436 6886 1488
rect 6917 1479 6975 1485
rect 6917 1445 6929 1479
rect 6963 1476 6975 1479
rect 10428 1476 10456 1516
rect 17954 1504 17960 1516
rect 18012 1504 18018 1556
rect 18046 1504 18052 1556
rect 18104 1544 18110 1556
rect 28261 1547 28319 1553
rect 28261 1544 28273 1547
rect 18104 1516 28273 1544
rect 18104 1504 18110 1516
rect 28261 1513 28273 1516
rect 28307 1513 28319 1547
rect 28261 1507 28319 1513
rect 28350 1504 28356 1556
rect 28408 1544 28414 1556
rect 35253 1547 35311 1553
rect 35253 1544 35265 1547
rect 28408 1516 35265 1544
rect 28408 1504 28414 1516
rect 35253 1513 35265 1516
rect 35299 1513 35311 1547
rect 35253 1507 35311 1513
rect 36170 1504 36176 1556
rect 36228 1544 36234 1556
rect 36228 1516 39528 1544
rect 36228 1504 36234 1516
rect 6963 1448 10456 1476
rect 10597 1479 10655 1485
rect 6963 1445 6975 1448
rect 6917 1439 6975 1445
rect 10597 1445 10609 1479
rect 10643 1476 10655 1479
rect 12897 1479 12955 1485
rect 12897 1476 12909 1479
rect 10643 1448 12909 1476
rect 10643 1445 10655 1448
rect 10597 1439 10655 1445
rect 12897 1445 12909 1448
rect 12943 1445 12955 1479
rect 39500 1476 39528 1516
rect 39574 1504 39580 1556
rect 39632 1544 39638 1556
rect 41138 1544 41144 1556
rect 39632 1516 41144 1544
rect 39632 1504 39638 1516
rect 41138 1504 41144 1516
rect 41196 1504 41202 1556
rect 45462 1504 45468 1556
rect 45520 1544 45526 1556
rect 48777 1547 48835 1553
rect 48777 1544 48789 1547
rect 45520 1516 48789 1544
rect 45520 1504 45526 1516
rect 48777 1513 48789 1516
rect 48823 1513 48835 1547
rect 48777 1507 48835 1513
rect 48869 1547 48927 1553
rect 48869 1513 48881 1547
rect 48915 1513 48927 1547
rect 56594 1544 56600 1556
rect 48869 1507 48927 1513
rect 48976 1516 56600 1544
rect 48884 1476 48912 1507
rect 48976 1488 49004 1516
rect 56594 1504 56600 1516
rect 56652 1504 56658 1556
rect 56689 1547 56747 1553
rect 56689 1513 56701 1547
rect 56735 1544 56747 1547
rect 58066 1544 58072 1556
rect 56735 1516 58072 1544
rect 56735 1513 56747 1516
rect 56689 1507 56747 1513
rect 58066 1504 58072 1516
rect 58124 1504 58130 1556
rect 58253 1547 58311 1553
rect 58253 1513 58265 1547
rect 58299 1544 58311 1547
rect 59262 1544 59268 1556
rect 58299 1516 59268 1544
rect 58299 1513 58311 1516
rect 58253 1507 58311 1513
rect 59262 1504 59268 1516
rect 59320 1504 59326 1556
rect 59354 1504 59360 1556
rect 59412 1544 59418 1556
rect 66898 1544 66904 1556
rect 59412 1516 66904 1544
rect 59412 1504 59418 1516
rect 66898 1504 66904 1516
rect 66956 1504 66962 1556
rect 66993 1547 67051 1553
rect 66993 1513 67005 1547
rect 67039 1544 67051 1547
rect 82817 1547 82875 1553
rect 82817 1544 82829 1547
rect 67039 1516 82829 1544
rect 67039 1513 67051 1516
rect 66993 1507 67051 1513
rect 82817 1513 82829 1516
rect 82863 1513 82875 1547
rect 82817 1507 82875 1513
rect 83461 1547 83519 1553
rect 83461 1513 83473 1547
rect 83507 1544 83519 1547
rect 87509 1547 87567 1553
rect 87509 1544 87521 1547
rect 83507 1516 87521 1544
rect 83507 1513 83519 1516
rect 83461 1507 83519 1513
rect 87509 1513 87521 1516
rect 87555 1513 87567 1547
rect 101401 1547 101459 1553
rect 101401 1544 101413 1547
rect 87509 1507 87567 1513
rect 87616 1516 101413 1544
rect 12897 1439 12955 1445
rect 13004 1448 39344 1476
rect 39500 1448 48912 1476
rect 934 1368 940 1420
rect 992 1408 998 1420
rect 5169 1411 5227 1417
rect 5169 1408 5181 1411
rect 992 1380 5181 1408
rect 992 1368 998 1380
rect 5169 1377 5181 1380
rect 5215 1377 5227 1411
rect 5169 1371 5227 1377
rect 5258 1368 5264 1420
rect 5316 1408 5322 1420
rect 5629 1411 5687 1417
rect 5629 1408 5641 1411
rect 5316 1380 5641 1408
rect 5316 1368 5322 1380
rect 5629 1377 5641 1380
rect 5675 1377 5687 1411
rect 5629 1371 5687 1377
rect 5902 1368 5908 1420
rect 5960 1408 5966 1420
rect 6454 1408 6460 1420
rect 5960 1380 6460 1408
rect 5960 1368 5966 1380
rect 6454 1368 6460 1380
rect 6512 1368 6518 1420
rect 7285 1411 7343 1417
rect 7285 1377 7297 1411
rect 7331 1408 7343 1411
rect 10505 1411 10563 1417
rect 10505 1408 10517 1411
rect 7331 1380 10517 1408
rect 7331 1377 7343 1380
rect 7285 1371 7343 1377
rect 10505 1377 10517 1380
rect 10551 1377 10563 1411
rect 10505 1371 10563 1377
rect 10686 1368 10692 1420
rect 10744 1408 10750 1420
rect 13004 1408 13032 1448
rect 25961 1411 26019 1417
rect 25961 1408 25973 1411
rect 10744 1380 13032 1408
rect 13096 1380 25973 1408
rect 10744 1368 10750 1380
rect 1121 1343 1179 1349
rect 1121 1309 1133 1343
rect 1167 1340 1179 1343
rect 4982 1340 4988 1352
rect 1167 1312 4988 1340
rect 1167 1309 1179 1312
rect 1121 1303 1179 1309
rect 4982 1300 4988 1312
rect 5040 1300 5046 1352
rect 5350 1300 5356 1352
rect 5408 1340 5414 1352
rect 5408 1312 10364 1340
rect 5408 1300 5414 1312
rect 3142 1232 3148 1284
rect 3200 1272 3206 1284
rect 5077 1275 5135 1281
rect 5077 1272 5089 1275
rect 3200 1244 5089 1272
rect 3200 1232 3206 1244
rect 5077 1241 5089 1244
rect 5123 1241 5135 1275
rect 5077 1235 5135 1241
rect 5261 1275 5319 1281
rect 5261 1241 5273 1275
rect 5307 1272 5319 1275
rect 8846 1272 8852 1284
rect 5307 1244 8852 1272
rect 5307 1241 5319 1244
rect 5261 1235 5319 1241
rect 8846 1232 8852 1244
rect 8904 1232 8910 1284
rect 1581 1207 1639 1213
rect 1581 1173 1593 1207
rect 1627 1204 1639 1207
rect 5169 1207 5227 1213
rect 5169 1204 5181 1207
rect 1627 1176 5181 1204
rect 1627 1173 1639 1176
rect 1581 1167 1639 1173
rect 5169 1173 5181 1176
rect 5215 1173 5227 1207
rect 5169 1167 5227 1173
rect 5353 1207 5411 1213
rect 5353 1173 5365 1207
rect 5399 1204 5411 1207
rect 6917 1207 6975 1213
rect 6917 1204 6929 1207
rect 5399 1176 6929 1204
rect 5399 1173 5411 1176
rect 5353 1167 5411 1173
rect 6917 1173 6929 1176
rect 6963 1173 6975 1207
rect 10336 1204 10364 1312
rect 10594 1300 10600 1352
rect 10652 1340 10658 1352
rect 13096 1340 13124 1380
rect 25961 1377 25973 1380
rect 26007 1377 26019 1411
rect 25961 1371 26019 1377
rect 26789 1411 26847 1417
rect 26789 1377 26801 1411
rect 26835 1408 26847 1411
rect 27065 1411 27123 1417
rect 27065 1408 27077 1411
rect 26835 1380 27077 1408
rect 26835 1377 26847 1380
rect 26789 1371 26847 1377
rect 27065 1377 27077 1380
rect 27111 1377 27123 1411
rect 27065 1371 27123 1377
rect 29086 1368 29092 1420
rect 29144 1408 29150 1420
rect 35069 1411 35127 1417
rect 29144 1380 34468 1408
rect 29144 1368 29150 1380
rect 10652 1312 13124 1340
rect 13173 1343 13231 1349
rect 10652 1300 10658 1312
rect 13173 1309 13185 1343
rect 13219 1340 13231 1343
rect 14458 1340 14464 1352
rect 13219 1312 14464 1340
rect 13219 1309 13231 1312
rect 13173 1303 13231 1309
rect 14458 1300 14464 1312
rect 14516 1300 14522 1352
rect 14550 1300 14556 1352
rect 14608 1340 14614 1352
rect 18046 1340 18052 1352
rect 14608 1312 18052 1340
rect 14608 1300 14614 1312
rect 18046 1300 18052 1312
rect 18104 1300 18110 1352
rect 26237 1343 26295 1349
rect 26237 1309 26249 1343
rect 26283 1340 26295 1343
rect 34333 1343 34391 1349
rect 34333 1340 34345 1343
rect 26283 1312 34345 1340
rect 26283 1309 26295 1312
rect 26237 1303 26295 1309
rect 34333 1309 34345 1312
rect 34379 1309 34391 1343
rect 34440 1340 34468 1380
rect 35069 1377 35081 1411
rect 35115 1408 35127 1411
rect 39025 1411 39083 1417
rect 39025 1408 39037 1411
rect 35115 1380 39037 1408
rect 35115 1377 35127 1380
rect 35069 1371 35127 1377
rect 39025 1377 39037 1380
rect 39071 1377 39083 1411
rect 39025 1371 39083 1377
rect 39117 1343 39175 1349
rect 39117 1340 39129 1343
rect 34440 1312 39129 1340
rect 34333 1303 34391 1309
rect 39117 1309 39129 1312
rect 39163 1309 39175 1343
rect 39316 1340 39344 1448
rect 48958 1436 48964 1488
rect 49016 1436 49022 1488
rect 49053 1479 49111 1485
rect 49053 1445 49065 1479
rect 49099 1476 49111 1479
rect 57974 1476 57980 1488
rect 49099 1448 57980 1476
rect 49099 1445 49111 1448
rect 49053 1439 49111 1445
rect 57974 1436 57980 1448
rect 58032 1436 58038 1488
rect 58161 1479 58219 1485
rect 58161 1445 58173 1479
rect 58207 1476 58219 1479
rect 60734 1476 60740 1488
rect 58207 1448 60740 1476
rect 58207 1445 58219 1448
rect 58161 1439 58219 1445
rect 60734 1436 60740 1448
rect 60792 1436 60798 1488
rect 60921 1479 60979 1485
rect 60921 1445 60933 1479
rect 60967 1476 60979 1479
rect 62117 1479 62175 1485
rect 62117 1476 62129 1479
rect 60967 1448 62129 1476
rect 60967 1445 60979 1448
rect 60921 1439 60979 1445
rect 62117 1445 62129 1448
rect 62163 1445 62175 1479
rect 65521 1479 65579 1485
rect 65521 1476 65533 1479
rect 62117 1439 62175 1445
rect 62224 1448 65533 1476
rect 39393 1411 39451 1417
rect 39393 1377 39405 1411
rect 39439 1408 39451 1411
rect 48869 1411 48927 1417
rect 48869 1408 48881 1411
rect 39439 1380 48881 1408
rect 39439 1377 39451 1380
rect 39393 1371 39451 1377
rect 48869 1377 48881 1380
rect 48915 1377 48927 1411
rect 48869 1371 48927 1377
rect 49145 1411 49203 1417
rect 49145 1377 49157 1411
rect 49191 1408 49203 1411
rect 53285 1411 53343 1417
rect 53285 1408 53297 1411
rect 49191 1380 53297 1408
rect 49191 1377 49203 1380
rect 49145 1371 49203 1377
rect 53285 1377 53297 1380
rect 53331 1377 53343 1411
rect 62224 1408 62252 1448
rect 65521 1445 65533 1448
rect 65567 1445 65579 1479
rect 65521 1439 65579 1445
rect 65613 1479 65671 1485
rect 65613 1445 65625 1479
rect 65659 1476 65671 1479
rect 66717 1479 66775 1485
rect 66717 1476 66729 1479
rect 65659 1448 66729 1476
rect 65659 1445 65671 1448
rect 65613 1439 65671 1445
rect 66717 1445 66729 1448
rect 66763 1445 66775 1479
rect 66717 1439 66775 1445
rect 66809 1479 66867 1485
rect 66809 1445 66821 1479
rect 66855 1476 66867 1479
rect 76285 1479 76343 1485
rect 76285 1476 76297 1479
rect 66855 1448 76297 1476
rect 66855 1445 66867 1448
rect 66809 1439 66867 1445
rect 76285 1445 76297 1448
rect 76331 1445 76343 1479
rect 76285 1439 76343 1445
rect 76377 1479 76435 1485
rect 76377 1445 76389 1479
rect 76423 1476 76435 1479
rect 78582 1476 78588 1488
rect 76423 1448 78588 1476
rect 76423 1445 76435 1448
rect 76377 1439 76435 1445
rect 78582 1436 78588 1448
rect 78640 1436 78646 1488
rect 78677 1479 78735 1485
rect 78677 1445 78689 1479
rect 78723 1476 78735 1479
rect 82633 1479 82691 1485
rect 82633 1476 82645 1479
rect 78723 1448 82645 1476
rect 78723 1445 78735 1448
rect 78677 1439 78735 1445
rect 82633 1445 82645 1448
rect 82679 1445 82691 1479
rect 82633 1439 82691 1445
rect 82725 1479 82783 1485
rect 82725 1445 82737 1479
rect 82771 1476 82783 1479
rect 83185 1479 83243 1485
rect 83185 1476 83197 1479
rect 82771 1448 83197 1476
rect 82771 1445 82783 1448
rect 82725 1439 82783 1445
rect 83185 1445 83197 1448
rect 83231 1445 83243 1479
rect 83185 1439 83243 1445
rect 83369 1479 83427 1485
rect 83369 1445 83381 1479
rect 83415 1476 83427 1479
rect 87616 1476 87644 1516
rect 101401 1513 101413 1516
rect 101447 1513 101459 1547
rect 101401 1507 101459 1513
rect 101674 1504 101680 1556
rect 101732 1544 101738 1556
rect 102226 1544 102232 1556
rect 101732 1516 102232 1544
rect 101732 1504 101738 1516
rect 102226 1504 102232 1516
rect 102284 1504 102290 1556
rect 102413 1547 102471 1553
rect 102413 1513 102425 1547
rect 102459 1544 102471 1547
rect 103330 1544 103336 1556
rect 102459 1516 103336 1544
rect 102459 1513 102471 1516
rect 102413 1507 102471 1513
rect 103330 1504 103336 1516
rect 103388 1504 103394 1556
rect 103425 1547 103483 1553
rect 103425 1513 103437 1547
rect 103471 1544 103483 1547
rect 103698 1544 103704 1556
rect 103471 1516 103704 1544
rect 103471 1513 103483 1516
rect 103425 1507 103483 1513
rect 103698 1504 103704 1516
rect 103756 1504 103762 1556
rect 103793 1547 103851 1553
rect 103793 1513 103805 1547
rect 103839 1544 103851 1547
rect 104345 1547 104403 1553
rect 104345 1544 104357 1547
rect 103839 1516 104357 1544
rect 103839 1513 103851 1516
rect 103793 1507 103851 1513
rect 104345 1513 104357 1516
rect 104391 1513 104403 1547
rect 104345 1507 104403 1513
rect 104529 1547 104587 1553
rect 104529 1513 104541 1547
rect 104575 1544 104587 1547
rect 136637 1547 136695 1553
rect 136637 1544 136649 1547
rect 104575 1516 129412 1544
rect 104575 1513 104587 1516
rect 104529 1507 104587 1513
rect 83415 1448 87644 1476
rect 87693 1479 87751 1485
rect 83415 1445 83427 1448
rect 83369 1439 83427 1445
rect 87693 1445 87705 1479
rect 87739 1476 87751 1479
rect 92753 1479 92811 1485
rect 87739 1448 92704 1476
rect 87739 1445 87751 1448
rect 87693 1439 87751 1445
rect 53285 1371 53343 1377
rect 54956 1380 62252 1408
rect 47026 1340 47032 1352
rect 39316 1312 47032 1340
rect 39117 1303 39175 1309
rect 47026 1300 47032 1312
rect 47084 1300 47090 1352
rect 54956 1340 54984 1380
rect 62298 1368 62304 1420
rect 62356 1408 62362 1420
rect 68830 1408 68836 1420
rect 62356 1380 68836 1408
rect 62356 1368 62362 1380
rect 68830 1368 68836 1380
rect 68888 1368 68894 1420
rect 68922 1368 68928 1420
rect 68980 1408 68986 1420
rect 71777 1411 71835 1417
rect 71777 1408 71789 1411
rect 68980 1380 71789 1408
rect 68980 1368 68986 1380
rect 71777 1377 71789 1380
rect 71823 1377 71835 1411
rect 71777 1371 71835 1377
rect 71866 1368 71872 1420
rect 71924 1408 71930 1420
rect 74442 1408 74448 1420
rect 71924 1380 74448 1408
rect 71924 1368 71930 1380
rect 74442 1368 74448 1380
rect 74500 1368 74506 1420
rect 74534 1368 74540 1420
rect 74592 1408 74598 1420
rect 74813 1411 74871 1417
rect 74813 1408 74825 1411
rect 74592 1380 74825 1408
rect 74592 1368 74598 1380
rect 74813 1377 74825 1380
rect 74859 1377 74871 1411
rect 78769 1411 78827 1417
rect 78769 1408 78781 1411
rect 74813 1371 74871 1377
rect 74920 1380 78781 1408
rect 47136 1312 54984 1340
rect 10413 1275 10471 1281
rect 10413 1241 10425 1275
rect 10459 1272 10471 1275
rect 11057 1275 11115 1281
rect 11057 1272 11069 1275
rect 10459 1244 11069 1272
rect 10459 1241 10471 1244
rect 10413 1235 10471 1241
rect 11057 1241 11069 1244
rect 11103 1241 11115 1275
rect 11057 1235 11115 1241
rect 11149 1275 11207 1281
rect 11149 1241 11161 1275
rect 11195 1272 11207 1275
rect 27890 1272 27896 1284
rect 11195 1244 27896 1272
rect 11195 1241 11207 1244
rect 11149 1235 11207 1241
rect 27890 1232 27896 1244
rect 27948 1232 27954 1284
rect 28261 1275 28319 1281
rect 28261 1241 28273 1275
rect 28307 1272 28319 1275
rect 39485 1275 39543 1281
rect 28307 1244 39344 1272
rect 28307 1241 28319 1244
rect 28261 1235 28319 1241
rect 24302 1204 24308 1216
rect 10336 1176 24308 1204
rect 6917 1167 6975 1173
rect 24302 1164 24308 1176
rect 24360 1164 24366 1216
rect 25133 1207 25191 1213
rect 25133 1173 25145 1207
rect 25179 1204 25191 1207
rect 39209 1207 39267 1213
rect 39209 1204 39221 1207
rect 25179 1176 39221 1204
rect 25179 1173 25191 1176
rect 25133 1167 25191 1173
rect 39209 1173 39221 1176
rect 39255 1173 39267 1207
rect 39209 1167 39267 1173
rect 1673 1139 1731 1145
rect 1673 1105 1685 1139
rect 1719 1136 1731 1139
rect 4982 1136 4988 1148
rect 1719 1108 4988 1136
rect 1719 1105 1731 1108
rect 1673 1099 1731 1105
rect 4982 1096 4988 1108
rect 5040 1096 5046 1148
rect 10413 1139 10471 1145
rect 10413 1136 10425 1139
rect 5368 1108 10425 1136
rect 1397 1071 1455 1077
rect 1397 1037 1409 1071
rect 1443 1068 1455 1071
rect 5074 1068 5080 1080
rect 1443 1040 5080 1068
rect 1443 1037 1455 1040
rect 1397 1031 1455 1037
rect 5074 1028 5080 1040
rect 5132 1028 5138 1080
rect 5261 1071 5319 1077
rect 5261 1037 5273 1071
rect 5307 1068 5319 1071
rect 5368 1068 5396 1108
rect 10413 1105 10425 1108
rect 10459 1105 10471 1139
rect 10413 1099 10471 1105
rect 10505 1139 10563 1145
rect 10505 1105 10517 1139
rect 10551 1136 10563 1139
rect 33870 1136 33876 1148
rect 10551 1108 33876 1136
rect 10551 1105 10563 1108
rect 10505 1099 10563 1105
rect 33870 1096 33876 1108
rect 33928 1096 33934 1148
rect 34333 1139 34391 1145
rect 34333 1105 34345 1139
rect 34379 1136 34391 1139
rect 38381 1139 38439 1145
rect 38381 1136 38393 1139
rect 34379 1108 38393 1136
rect 34379 1105 34391 1108
rect 34333 1099 34391 1105
rect 38381 1105 38393 1108
rect 38427 1105 38439 1139
rect 39316 1136 39344 1244
rect 39485 1241 39497 1275
rect 39531 1272 39543 1275
rect 47136 1272 47164 1312
rect 55030 1300 55036 1352
rect 55088 1340 55094 1352
rect 58069 1343 58127 1349
rect 58069 1340 58081 1343
rect 55088 1312 58081 1340
rect 55088 1300 55094 1312
rect 58069 1309 58081 1312
rect 58115 1309 58127 1343
rect 58069 1303 58127 1309
rect 58250 1300 58256 1352
rect 58308 1340 58314 1352
rect 59081 1343 59139 1349
rect 59081 1340 59093 1343
rect 58308 1312 59093 1340
rect 58308 1300 58314 1312
rect 59081 1309 59093 1312
rect 59127 1309 59139 1343
rect 59081 1303 59139 1309
rect 59170 1300 59176 1352
rect 59228 1340 59234 1352
rect 61289 1343 61347 1349
rect 61289 1340 61301 1343
rect 59228 1312 61301 1340
rect 59228 1300 59234 1312
rect 61289 1309 61301 1312
rect 61335 1309 61347 1343
rect 61289 1303 61347 1309
rect 62117 1343 62175 1349
rect 62117 1309 62129 1343
rect 62163 1340 62175 1343
rect 63313 1343 63371 1349
rect 63313 1340 63325 1343
rect 62163 1312 63325 1340
rect 62163 1309 62175 1312
rect 62117 1303 62175 1309
rect 63313 1309 63325 1312
rect 63359 1309 63371 1343
rect 63313 1303 63371 1309
rect 63405 1343 63463 1349
rect 63405 1309 63417 1343
rect 63451 1340 63463 1343
rect 66993 1343 67051 1349
rect 66993 1340 67005 1343
rect 63451 1312 67005 1340
rect 63451 1309 63463 1312
rect 63405 1303 63463 1309
rect 66993 1309 67005 1312
rect 67039 1309 67051 1343
rect 66993 1303 67051 1309
rect 67085 1343 67143 1349
rect 67085 1309 67097 1343
rect 67131 1340 67143 1343
rect 72789 1343 72847 1349
rect 72789 1340 72801 1343
rect 67131 1312 72801 1340
rect 67131 1309 67143 1312
rect 67085 1303 67143 1309
rect 72789 1309 72801 1312
rect 72835 1309 72847 1343
rect 72789 1303 72847 1309
rect 72881 1343 72939 1349
rect 72881 1309 72893 1343
rect 72927 1340 72939 1343
rect 74920 1340 74948 1380
rect 78769 1377 78781 1380
rect 78815 1377 78827 1411
rect 78769 1371 78827 1377
rect 78858 1368 78864 1420
rect 78916 1408 78922 1420
rect 81342 1408 81348 1420
rect 78916 1380 81348 1408
rect 78916 1368 78922 1380
rect 81342 1368 81348 1380
rect 81400 1368 81406 1420
rect 81437 1411 81495 1417
rect 81437 1377 81449 1411
rect 81483 1408 81495 1411
rect 81713 1411 81771 1417
rect 81713 1408 81725 1411
rect 81483 1380 81725 1408
rect 81483 1377 81495 1380
rect 81437 1371 81495 1377
rect 81713 1377 81725 1380
rect 81759 1377 81771 1411
rect 81713 1371 81771 1377
rect 81802 1368 81808 1420
rect 81860 1408 81866 1420
rect 84105 1411 84163 1417
rect 84105 1408 84117 1411
rect 81860 1380 83320 1408
rect 81860 1368 81866 1380
rect 72927 1312 74948 1340
rect 74997 1343 75055 1349
rect 72927 1309 72939 1312
rect 72881 1303 72939 1309
rect 74997 1309 75009 1343
rect 75043 1340 75055 1343
rect 76650 1340 76656 1352
rect 75043 1312 76656 1340
rect 75043 1309 75055 1312
rect 74997 1303 75055 1309
rect 76650 1300 76656 1312
rect 76708 1300 76714 1352
rect 76745 1343 76803 1349
rect 76745 1309 76757 1343
rect 76791 1340 76803 1343
rect 83093 1343 83151 1349
rect 83093 1340 83105 1343
rect 76791 1312 83105 1340
rect 76791 1309 76803 1312
rect 76745 1303 76803 1309
rect 83093 1309 83105 1312
rect 83139 1309 83151 1343
rect 83093 1303 83151 1309
rect 83185 1343 83243 1349
rect 83185 1309 83197 1343
rect 83231 1309 83243 1343
rect 83185 1303 83243 1309
rect 39531 1244 47164 1272
rect 39531 1241 39543 1244
rect 39485 1235 39543 1241
rect 47946 1232 47952 1284
rect 48004 1272 48010 1284
rect 48682 1272 48688 1284
rect 48004 1244 48688 1272
rect 48004 1232 48010 1244
rect 48682 1232 48688 1244
rect 48740 1232 48746 1284
rect 48869 1275 48927 1281
rect 48869 1241 48881 1275
rect 48915 1272 48927 1275
rect 48915 1244 63448 1272
rect 48915 1241 48927 1244
rect 48869 1235 48927 1241
rect 39390 1164 39396 1216
rect 39448 1204 39454 1216
rect 49053 1207 49111 1213
rect 49053 1204 49065 1207
rect 39448 1176 49065 1204
rect 39448 1164 39454 1176
rect 49053 1173 49065 1176
rect 49099 1173 49111 1207
rect 49053 1167 49111 1173
rect 49145 1207 49203 1213
rect 49145 1173 49157 1207
rect 49191 1204 49203 1207
rect 56686 1204 56692 1216
rect 49191 1176 56692 1204
rect 49191 1173 49203 1176
rect 49145 1167 49203 1173
rect 56686 1164 56692 1176
rect 56744 1164 56750 1216
rect 57974 1164 57980 1216
rect 58032 1204 58038 1216
rect 63313 1207 63371 1213
rect 63313 1204 63325 1207
rect 58032 1176 63325 1204
rect 58032 1164 58038 1176
rect 63313 1173 63325 1176
rect 63359 1173 63371 1207
rect 63420 1204 63448 1244
rect 63678 1232 63684 1284
rect 63736 1272 63742 1284
rect 78677 1275 78735 1281
rect 78677 1272 78689 1275
rect 63736 1244 78689 1272
rect 63736 1232 63742 1244
rect 78677 1241 78689 1244
rect 78723 1241 78735 1275
rect 78677 1235 78735 1241
rect 78766 1232 78772 1284
rect 78824 1272 78830 1284
rect 82354 1272 82360 1284
rect 78824 1244 82360 1272
rect 78824 1232 78830 1244
rect 82354 1232 82360 1244
rect 82412 1232 82418 1284
rect 83200 1272 83228 1303
rect 82924 1244 83228 1272
rect 83292 1272 83320 1380
rect 83384 1380 84117 1408
rect 83384 1349 83412 1380
rect 84105 1377 84117 1380
rect 84151 1377 84163 1411
rect 84105 1371 84163 1377
rect 84197 1411 84255 1417
rect 84197 1377 84209 1411
rect 84243 1408 84255 1411
rect 85666 1408 85672 1420
rect 84243 1380 85672 1408
rect 84243 1377 84255 1380
rect 84197 1371 84255 1377
rect 85666 1368 85672 1380
rect 85724 1368 85730 1420
rect 85850 1368 85856 1420
rect 85908 1408 85914 1420
rect 85945 1411 86003 1417
rect 85945 1408 85957 1411
rect 85908 1380 85957 1408
rect 85908 1368 85914 1380
rect 85945 1377 85957 1380
rect 85991 1377 86003 1411
rect 85945 1371 86003 1377
rect 86037 1411 86095 1417
rect 86037 1377 86049 1411
rect 86083 1408 86095 1411
rect 87417 1411 87475 1417
rect 87417 1408 87429 1411
rect 86083 1380 87429 1408
rect 86083 1377 86095 1380
rect 86037 1371 86095 1377
rect 87417 1377 87429 1380
rect 87463 1377 87475 1411
rect 87417 1371 87475 1377
rect 87509 1411 87567 1417
rect 87509 1377 87521 1411
rect 87555 1408 87567 1411
rect 91833 1411 91891 1417
rect 91833 1408 91845 1411
rect 87555 1380 91845 1408
rect 87555 1377 87567 1380
rect 87509 1371 87567 1377
rect 91833 1377 91845 1380
rect 91879 1377 91891 1411
rect 92569 1411 92627 1417
rect 92569 1408 92581 1411
rect 91833 1371 91891 1377
rect 92308 1380 92581 1408
rect 83369 1343 83427 1349
rect 83369 1309 83381 1343
rect 83415 1309 83427 1343
rect 83369 1303 83427 1309
rect 83553 1343 83611 1349
rect 83553 1309 83565 1343
rect 83599 1340 83611 1343
rect 83599 1312 86264 1340
rect 83599 1309 83611 1312
rect 83553 1303 83611 1309
rect 86236 1272 86264 1312
rect 86310 1300 86316 1352
rect 86368 1340 86374 1352
rect 86862 1340 86868 1352
rect 86368 1312 86868 1340
rect 86368 1300 86374 1312
rect 86862 1300 86868 1312
rect 86920 1300 86926 1352
rect 87049 1343 87107 1349
rect 87049 1309 87061 1343
rect 87095 1340 87107 1343
rect 87601 1343 87659 1349
rect 87601 1340 87613 1343
rect 87095 1312 87613 1340
rect 87095 1309 87107 1312
rect 87049 1303 87107 1309
rect 87601 1309 87613 1312
rect 87647 1309 87659 1343
rect 92308 1340 92336 1380
rect 92569 1377 92581 1380
rect 92615 1377 92627 1411
rect 92676 1408 92704 1448
rect 92753 1445 92765 1479
rect 92799 1476 92811 1479
rect 101493 1479 101551 1485
rect 101493 1476 101505 1479
rect 92799 1448 101505 1476
rect 92799 1445 92811 1448
rect 92753 1439 92811 1445
rect 101493 1445 101505 1448
rect 101539 1445 101551 1479
rect 101493 1439 101551 1445
rect 101585 1479 101643 1485
rect 101585 1445 101597 1479
rect 101631 1445 101643 1479
rect 101585 1439 101643 1445
rect 102321 1479 102379 1485
rect 102321 1445 102333 1479
rect 102367 1476 102379 1479
rect 106829 1479 106887 1485
rect 106829 1476 106841 1479
rect 102367 1448 106841 1476
rect 102367 1445 102379 1448
rect 102321 1439 102379 1445
rect 106829 1445 106841 1448
rect 106875 1445 106887 1479
rect 106829 1439 106887 1445
rect 93029 1411 93087 1417
rect 92676 1380 92796 1408
rect 92569 1371 92627 1377
rect 87601 1303 87659 1309
rect 87708 1312 92336 1340
rect 92385 1343 92443 1349
rect 87708 1272 87736 1312
rect 92385 1309 92397 1343
rect 92431 1340 92443 1343
rect 92431 1312 92704 1340
rect 92431 1309 92443 1312
rect 92385 1303 92443 1309
rect 92676 1284 92704 1312
rect 91833 1275 91891 1281
rect 91833 1272 91845 1275
rect 83292 1244 86172 1272
rect 86236 1244 87736 1272
rect 87800 1244 91845 1272
rect 63497 1207 63555 1213
rect 63497 1204 63509 1207
rect 63420 1176 63509 1204
rect 63313 1167 63371 1173
rect 63497 1173 63509 1176
rect 63543 1173 63555 1207
rect 63497 1167 63555 1173
rect 63586 1164 63592 1216
rect 63644 1204 63650 1216
rect 66809 1207 66867 1213
rect 66809 1204 66821 1207
rect 63644 1176 66821 1204
rect 63644 1164 63650 1176
rect 66809 1173 66821 1176
rect 66855 1173 66867 1207
rect 66809 1167 66867 1173
rect 66898 1164 66904 1216
rect 66956 1204 66962 1216
rect 72973 1207 73031 1213
rect 72973 1204 72985 1207
rect 66956 1176 72985 1204
rect 66956 1164 66962 1176
rect 72973 1173 72985 1176
rect 73019 1173 73031 1207
rect 72973 1167 73031 1173
rect 73157 1207 73215 1213
rect 73157 1173 73169 1207
rect 73203 1204 73215 1207
rect 76193 1207 76251 1213
rect 76193 1204 76205 1207
rect 73203 1176 76205 1204
rect 73203 1173 73215 1176
rect 73157 1167 73215 1173
rect 76193 1173 76205 1176
rect 76239 1173 76251 1207
rect 76193 1167 76251 1173
rect 76285 1207 76343 1213
rect 76285 1173 76297 1207
rect 76331 1204 76343 1207
rect 82817 1207 82875 1213
rect 82817 1204 82829 1207
rect 76331 1176 82829 1204
rect 76331 1173 76343 1176
rect 76285 1167 76343 1173
rect 82817 1173 82829 1176
rect 82863 1173 82875 1207
rect 82817 1167 82875 1173
rect 78858 1136 78864 1148
rect 39316 1108 78864 1136
rect 38381 1099 38439 1105
rect 78858 1096 78864 1108
rect 78916 1096 78922 1148
rect 78953 1139 79011 1145
rect 78953 1105 78965 1139
rect 78999 1136 79011 1139
rect 82725 1139 82783 1145
rect 82725 1136 82737 1139
rect 78999 1108 82737 1136
rect 78999 1105 79011 1108
rect 78953 1099 79011 1105
rect 82725 1105 82737 1108
rect 82771 1105 82783 1139
rect 82924 1136 82952 1244
rect 83001 1207 83059 1213
rect 83001 1173 83013 1207
rect 83047 1204 83059 1207
rect 84841 1207 84899 1213
rect 84841 1204 84853 1207
rect 83047 1176 84853 1204
rect 83047 1173 83059 1176
rect 83001 1167 83059 1173
rect 84841 1173 84853 1176
rect 84887 1173 84899 1207
rect 84841 1167 84899 1173
rect 84930 1164 84936 1216
rect 84988 1204 84994 1216
rect 85761 1207 85819 1213
rect 85761 1204 85773 1207
rect 84988 1176 85773 1204
rect 84988 1164 84994 1176
rect 85761 1173 85773 1176
rect 85807 1173 85819 1207
rect 86144 1204 86172 1244
rect 87800 1204 87828 1244
rect 91833 1241 91845 1244
rect 91879 1241 91891 1275
rect 91833 1235 91891 1241
rect 91922 1232 91928 1284
rect 91980 1272 91986 1284
rect 92566 1272 92572 1284
rect 91980 1244 92572 1272
rect 91980 1232 91986 1244
rect 92566 1232 92572 1244
rect 92624 1232 92630 1284
rect 92658 1232 92664 1284
rect 92716 1232 92722 1284
rect 92768 1272 92796 1380
rect 93029 1377 93041 1411
rect 93075 1408 93087 1411
rect 101600 1408 101628 1439
rect 106918 1436 106924 1488
rect 106976 1476 106982 1488
rect 110693 1479 110751 1485
rect 110693 1476 110705 1479
rect 106976 1448 110705 1476
rect 106976 1436 106982 1448
rect 110693 1445 110705 1448
rect 110739 1445 110751 1479
rect 110693 1439 110751 1445
rect 110785 1479 110843 1485
rect 110785 1445 110797 1479
rect 110831 1476 110843 1479
rect 111061 1479 111119 1485
rect 111061 1476 111073 1479
rect 110831 1448 111073 1476
rect 110831 1445 110843 1448
rect 110785 1439 110843 1445
rect 111061 1445 111073 1448
rect 111107 1445 111119 1479
rect 111061 1439 111119 1445
rect 111242 1436 111248 1488
rect 111300 1476 111306 1488
rect 114833 1479 114891 1485
rect 114833 1476 114845 1479
rect 111300 1448 114845 1476
rect 111300 1436 111306 1448
rect 114833 1445 114845 1448
rect 114879 1445 114891 1479
rect 114833 1439 114891 1445
rect 114925 1479 114983 1485
rect 114925 1445 114937 1479
rect 114971 1476 114983 1479
rect 122101 1479 122159 1485
rect 122101 1476 122113 1479
rect 114971 1448 122113 1476
rect 114971 1445 114983 1448
rect 114925 1439 114983 1445
rect 122101 1445 122113 1448
rect 122147 1445 122159 1479
rect 122653 1479 122711 1485
rect 122653 1476 122665 1479
rect 122101 1439 122159 1445
rect 122208 1448 122665 1476
rect 93075 1380 101628 1408
rect 102045 1411 102103 1417
rect 93075 1377 93087 1380
rect 93029 1371 93087 1377
rect 102045 1377 102057 1411
rect 102091 1408 102103 1411
rect 105909 1411 105967 1417
rect 105909 1408 105921 1411
rect 102091 1380 105921 1408
rect 102091 1377 102103 1380
rect 102045 1371 102103 1377
rect 105909 1377 105921 1380
rect 105955 1377 105967 1411
rect 105909 1371 105967 1377
rect 106001 1411 106059 1417
rect 106001 1377 106013 1411
rect 106047 1408 106059 1411
rect 109862 1408 109868 1420
rect 106047 1380 109868 1408
rect 106047 1377 106059 1380
rect 106001 1371 106059 1377
rect 109862 1368 109868 1380
rect 109920 1368 109926 1420
rect 109957 1411 110015 1417
rect 109957 1377 109969 1411
rect 110003 1408 110015 1411
rect 111153 1411 111211 1417
rect 111153 1408 111165 1411
rect 110003 1380 111165 1408
rect 110003 1377 110015 1380
rect 109957 1371 110015 1377
rect 111153 1377 111165 1380
rect 111199 1377 111211 1411
rect 111153 1371 111211 1377
rect 111337 1411 111395 1417
rect 111337 1377 111349 1411
rect 111383 1408 111395 1411
rect 111426 1408 111432 1420
rect 111383 1380 111432 1408
rect 111383 1377 111395 1380
rect 111337 1371 111395 1377
rect 111426 1368 111432 1380
rect 111484 1368 111490 1420
rect 111521 1411 111579 1417
rect 111521 1377 111533 1411
rect 111567 1408 111579 1411
rect 115198 1408 115204 1420
rect 111567 1380 115204 1408
rect 111567 1377 111579 1380
rect 111521 1371 111579 1377
rect 115198 1368 115204 1380
rect 115256 1368 115262 1420
rect 115293 1411 115351 1417
rect 115293 1377 115305 1411
rect 115339 1408 115351 1411
rect 116213 1411 116271 1417
rect 116213 1408 116225 1411
rect 115339 1380 116225 1408
rect 115339 1377 115351 1380
rect 115293 1371 115351 1377
rect 116213 1377 116225 1380
rect 116259 1377 116271 1411
rect 116213 1371 116271 1377
rect 116305 1411 116363 1417
rect 116305 1377 116317 1411
rect 116351 1408 116363 1411
rect 119430 1408 119436 1420
rect 116351 1380 119436 1408
rect 116351 1377 116363 1380
rect 116305 1371 116363 1377
rect 119430 1368 119436 1380
rect 119488 1368 119494 1420
rect 119798 1368 119804 1420
rect 119856 1408 119862 1420
rect 120350 1408 120356 1420
rect 119856 1380 120356 1408
rect 119856 1368 119862 1380
rect 120350 1368 120356 1380
rect 120408 1368 120414 1420
rect 120445 1411 120503 1417
rect 120445 1377 120457 1411
rect 120491 1408 120503 1411
rect 120905 1411 120963 1417
rect 120905 1408 120917 1411
rect 120491 1380 120917 1408
rect 120491 1377 120503 1380
rect 120445 1371 120503 1377
rect 120905 1377 120917 1380
rect 120951 1377 120963 1411
rect 120905 1371 120963 1377
rect 120994 1368 121000 1420
rect 121052 1408 121058 1420
rect 121917 1411 121975 1417
rect 121917 1408 121929 1411
rect 121052 1380 121929 1408
rect 121052 1368 121058 1380
rect 121917 1377 121929 1380
rect 121963 1377 121975 1411
rect 121917 1371 121975 1377
rect 122006 1368 122012 1420
rect 122064 1408 122070 1420
rect 122208 1408 122236 1448
rect 122653 1445 122665 1448
rect 122699 1445 122711 1479
rect 122653 1439 122711 1445
rect 122742 1436 122748 1488
rect 122800 1476 122806 1488
rect 125505 1479 125563 1485
rect 125505 1476 125517 1479
rect 122800 1448 125517 1476
rect 122800 1436 122806 1448
rect 125505 1445 125517 1448
rect 125551 1445 125563 1479
rect 125505 1439 125563 1445
rect 125597 1479 125655 1485
rect 125597 1445 125609 1479
rect 125643 1476 125655 1479
rect 125873 1479 125931 1485
rect 125873 1476 125885 1479
rect 125643 1448 125885 1476
rect 125643 1445 125655 1448
rect 125597 1439 125655 1445
rect 125873 1445 125885 1448
rect 125919 1445 125931 1479
rect 125873 1439 125931 1445
rect 125962 1436 125968 1488
rect 126020 1476 126026 1488
rect 127986 1476 127992 1488
rect 126020 1448 127992 1476
rect 126020 1436 126026 1448
rect 127986 1436 127992 1448
rect 128044 1436 128050 1488
rect 128081 1479 128139 1485
rect 128081 1445 128093 1479
rect 128127 1476 128139 1479
rect 128357 1479 128415 1485
rect 128357 1476 128369 1479
rect 128127 1448 128369 1476
rect 128127 1445 128139 1448
rect 128081 1439 128139 1445
rect 128357 1445 128369 1448
rect 128403 1445 128415 1479
rect 128357 1439 128415 1445
rect 128446 1436 128452 1488
rect 128504 1476 128510 1488
rect 128633 1479 128691 1485
rect 128633 1476 128645 1479
rect 128504 1448 128645 1476
rect 128504 1436 128510 1448
rect 128633 1445 128645 1448
rect 128679 1445 128691 1479
rect 128633 1439 128691 1445
rect 128725 1479 128783 1485
rect 128725 1445 128737 1479
rect 128771 1476 128783 1479
rect 129277 1479 129335 1485
rect 129277 1476 129289 1479
rect 128771 1448 129289 1476
rect 128771 1445 128783 1448
rect 128725 1439 128783 1445
rect 129277 1445 129289 1448
rect 129323 1445 129335 1479
rect 129384 1476 129412 1516
rect 129660 1516 136649 1544
rect 129660 1476 129688 1516
rect 136637 1513 136649 1516
rect 136683 1513 136695 1547
rect 136637 1507 136695 1513
rect 136821 1547 136879 1553
rect 136821 1513 136833 1547
rect 136867 1544 136879 1547
rect 142433 1547 142491 1553
rect 142433 1544 142445 1547
rect 136867 1516 142445 1544
rect 136867 1513 136879 1516
rect 136821 1507 136879 1513
rect 142433 1513 142445 1516
rect 142479 1513 142491 1547
rect 142433 1507 142491 1513
rect 142522 1504 142528 1556
rect 142580 1544 142586 1556
rect 142890 1544 142896 1556
rect 142580 1516 142896 1544
rect 142580 1504 142586 1516
rect 142890 1504 142896 1516
rect 142948 1504 142954 1556
rect 142985 1547 143043 1553
rect 142985 1513 142997 1547
rect 143031 1544 143043 1547
rect 144089 1547 144147 1553
rect 144089 1544 144101 1547
rect 143031 1516 144101 1544
rect 143031 1513 143043 1516
rect 142985 1507 143043 1513
rect 144089 1513 144101 1516
rect 144135 1513 144147 1547
rect 144089 1507 144147 1513
rect 144365 1547 144423 1553
rect 144365 1513 144377 1547
rect 144411 1544 144423 1547
rect 145101 1547 145159 1553
rect 145101 1544 145113 1547
rect 144411 1516 145113 1544
rect 144411 1513 144423 1516
rect 144365 1507 144423 1513
rect 145101 1513 145113 1516
rect 145147 1513 145159 1547
rect 145101 1507 145159 1513
rect 145193 1547 145251 1553
rect 145193 1513 145205 1547
rect 145239 1544 145251 1547
rect 151372 1544 151400 1584
rect 151541 1581 151553 1584
rect 151587 1581 151599 1615
rect 151541 1575 151599 1581
rect 151633 1615 151691 1621
rect 151633 1581 151645 1615
rect 151679 1612 151691 1615
rect 152277 1615 152335 1621
rect 151679 1584 152228 1612
rect 151679 1581 151691 1584
rect 151633 1575 151691 1581
rect 145239 1516 151400 1544
rect 151449 1547 151507 1553
rect 145239 1513 145251 1516
rect 145193 1507 145251 1513
rect 151449 1513 151461 1547
rect 151495 1544 151507 1547
rect 151909 1547 151967 1553
rect 151909 1544 151921 1547
rect 151495 1516 151921 1544
rect 151495 1513 151507 1516
rect 151449 1507 151507 1513
rect 151909 1513 151921 1516
rect 151955 1513 151967 1547
rect 151909 1507 151967 1513
rect 151998 1504 152004 1556
rect 152056 1544 152062 1556
rect 152093 1547 152151 1553
rect 152093 1544 152105 1547
rect 152056 1516 152105 1544
rect 152056 1504 152062 1516
rect 152093 1513 152105 1516
rect 152139 1513 152151 1547
rect 152200 1544 152228 1584
rect 152277 1581 152289 1615
rect 152323 1612 152335 1615
rect 152645 1615 152703 1621
rect 152645 1612 152657 1615
rect 152323 1584 152657 1612
rect 152323 1581 152335 1584
rect 152277 1575 152335 1581
rect 152645 1581 152657 1584
rect 152691 1581 152703 1615
rect 152645 1575 152703 1581
rect 152737 1615 152795 1621
rect 152737 1581 152749 1615
rect 152783 1612 152795 1615
rect 153565 1615 153623 1621
rect 153565 1612 153577 1615
rect 152783 1584 153577 1612
rect 152783 1581 152795 1584
rect 152737 1575 152795 1581
rect 153565 1581 153577 1584
rect 153611 1581 153623 1615
rect 156969 1615 157027 1621
rect 156969 1612 156981 1615
rect 153565 1575 153623 1581
rect 153672 1584 156981 1612
rect 153197 1547 153255 1553
rect 153197 1544 153209 1547
rect 152200 1516 153209 1544
rect 152093 1507 152151 1513
rect 153197 1513 153209 1516
rect 153243 1513 153255 1547
rect 153197 1507 153255 1513
rect 153289 1547 153347 1553
rect 153289 1513 153301 1547
rect 153335 1544 153347 1547
rect 153672 1544 153700 1584
rect 156969 1581 156981 1584
rect 157015 1581 157027 1615
rect 156969 1575 157027 1581
rect 157058 1572 157064 1624
rect 157116 1612 157122 1624
rect 157429 1615 157487 1621
rect 157429 1612 157441 1615
rect 157116 1584 157441 1612
rect 157116 1572 157122 1584
rect 157429 1581 157441 1584
rect 157475 1581 157487 1615
rect 157429 1575 157487 1581
rect 153335 1516 153700 1544
rect 153749 1547 153807 1553
rect 153335 1513 153347 1516
rect 153289 1507 153347 1513
rect 153749 1513 153761 1547
rect 153795 1544 153807 1547
rect 156325 1547 156383 1553
rect 156325 1544 156337 1547
rect 153795 1516 156337 1544
rect 153795 1513 153807 1516
rect 153749 1507 153807 1513
rect 156325 1513 156337 1516
rect 156371 1513 156383 1547
rect 156325 1507 156383 1513
rect 156509 1547 156567 1553
rect 156509 1513 156521 1547
rect 156555 1544 156567 1547
rect 156877 1547 156935 1553
rect 156877 1544 156889 1547
rect 156555 1516 156889 1544
rect 156555 1513 156567 1516
rect 156509 1507 156567 1513
rect 156877 1513 156889 1516
rect 156923 1513 156935 1547
rect 157150 1544 157156 1556
rect 157111 1516 157156 1544
rect 156877 1507 156935 1513
rect 157150 1504 157156 1516
rect 157208 1504 157214 1556
rect 157334 1544 157340 1556
rect 157295 1516 157340 1544
rect 157334 1504 157340 1516
rect 157392 1504 157398 1556
rect 157536 1544 157564 1652
rect 158898 1640 158904 1652
rect 158956 1640 158962 1692
rect 158993 1683 159051 1689
rect 158993 1649 159005 1683
rect 159039 1680 159051 1683
rect 160373 1683 160431 1689
rect 160373 1680 160385 1683
rect 159039 1652 160385 1680
rect 159039 1649 159051 1652
rect 158993 1643 159051 1649
rect 160373 1649 160385 1652
rect 160419 1649 160431 1683
rect 160373 1643 160431 1649
rect 160465 1683 160523 1689
rect 160465 1649 160477 1683
rect 160511 1680 160523 1683
rect 161017 1683 161075 1689
rect 160511 1652 160968 1680
rect 160511 1649 160523 1652
rect 160465 1643 160523 1649
rect 157613 1615 157671 1621
rect 157613 1581 157625 1615
rect 157659 1612 157671 1615
rect 158717 1615 158775 1621
rect 158717 1612 158729 1615
rect 157659 1584 158729 1612
rect 157659 1581 157671 1584
rect 157613 1575 157671 1581
rect 158717 1581 158729 1584
rect 158763 1581 158775 1615
rect 158717 1575 158775 1581
rect 158806 1572 158812 1624
rect 158864 1612 158870 1624
rect 159269 1615 159327 1621
rect 159269 1612 159281 1615
rect 158864 1584 159281 1612
rect 158864 1572 158870 1584
rect 159269 1581 159281 1584
rect 159315 1581 159327 1615
rect 159269 1575 159327 1581
rect 159358 1572 159364 1624
rect 159416 1612 159422 1624
rect 160833 1615 160891 1621
rect 160833 1612 160845 1615
rect 159416 1584 160845 1612
rect 159416 1572 159422 1584
rect 160833 1581 160845 1584
rect 160879 1581 160891 1615
rect 160940 1612 160968 1652
rect 161017 1649 161029 1683
rect 161063 1680 161075 1683
rect 169110 1680 169116 1692
rect 161063 1652 169116 1680
rect 161063 1649 161075 1652
rect 161017 1643 161075 1649
rect 169110 1640 169116 1652
rect 169168 1640 169174 1692
rect 169205 1683 169263 1689
rect 169205 1649 169217 1683
rect 169251 1680 169263 1683
rect 169570 1680 169576 1692
rect 169251 1652 169576 1680
rect 169251 1649 169263 1652
rect 169205 1643 169263 1649
rect 169570 1640 169576 1652
rect 169628 1640 169634 1692
rect 178589 1683 178647 1689
rect 178589 1680 178601 1683
rect 169680 1652 178601 1680
rect 161109 1615 161167 1621
rect 160940 1584 161060 1612
rect 160833 1575 160891 1581
rect 157889 1547 157947 1553
rect 157889 1544 157901 1547
rect 157536 1516 157901 1544
rect 157889 1513 157901 1516
rect 157935 1513 157947 1547
rect 157889 1507 157947 1513
rect 157978 1504 157984 1556
rect 158036 1544 158042 1556
rect 158993 1547 159051 1553
rect 158993 1544 159005 1547
rect 158036 1516 159005 1544
rect 158036 1504 158042 1516
rect 158993 1513 159005 1516
rect 159039 1513 159051 1547
rect 158993 1507 159051 1513
rect 159177 1547 159235 1553
rect 159177 1513 159189 1547
rect 159223 1544 159235 1547
rect 160278 1544 160284 1556
rect 159223 1516 160284 1544
rect 159223 1513 159235 1516
rect 159177 1507 159235 1513
rect 160278 1504 160284 1516
rect 160336 1504 160342 1556
rect 160373 1547 160431 1553
rect 160373 1513 160385 1547
rect 160419 1544 160431 1547
rect 160922 1544 160928 1556
rect 160419 1516 160928 1544
rect 160419 1513 160431 1516
rect 160373 1507 160431 1513
rect 160922 1504 160928 1516
rect 160980 1504 160986 1556
rect 161032 1544 161060 1584
rect 161109 1581 161121 1615
rect 161155 1612 161167 1615
rect 169680 1612 169708 1652
rect 178589 1649 178601 1652
rect 178635 1649 178647 1683
rect 178696 1680 178724 1720
rect 178865 1717 178877 1751
rect 178911 1748 178923 1751
rect 179693 1751 179751 1757
rect 178911 1720 179368 1748
rect 178911 1717 178923 1720
rect 178865 1711 178923 1717
rect 179340 1692 179368 1720
rect 179693 1717 179705 1751
rect 179739 1748 179751 1751
rect 180429 1751 180487 1757
rect 180429 1748 180441 1751
rect 179739 1720 180441 1748
rect 179739 1717 179751 1720
rect 179693 1711 179751 1717
rect 180429 1717 180441 1720
rect 180475 1717 180487 1751
rect 180429 1711 180487 1717
rect 180521 1751 180579 1757
rect 180521 1717 180533 1751
rect 180567 1748 180579 1751
rect 183664 1748 183692 1788
rect 220265 1785 220277 1788
rect 220311 1785 220323 1819
rect 220265 1779 220323 1785
rect 220725 1819 220783 1825
rect 220725 1785 220737 1819
rect 220771 1816 220783 1819
rect 231581 1819 231639 1825
rect 231581 1816 231593 1819
rect 220771 1788 231593 1816
rect 220771 1785 220783 1788
rect 220725 1779 220783 1785
rect 231581 1785 231593 1788
rect 231627 1785 231639 1819
rect 231581 1779 231639 1785
rect 231673 1819 231731 1825
rect 231673 1785 231685 1819
rect 231719 1816 231731 1819
rect 232133 1819 232191 1825
rect 232133 1816 232145 1819
rect 231719 1788 232145 1816
rect 231719 1785 231731 1788
rect 231673 1779 231731 1785
rect 232133 1785 232145 1788
rect 232179 1785 232191 1819
rect 232593 1819 232651 1825
rect 232593 1816 232605 1819
rect 232133 1779 232191 1785
rect 232240 1788 232605 1816
rect 180567 1720 183692 1748
rect 180567 1717 180579 1720
rect 180521 1711 180579 1717
rect 183738 1708 183744 1760
rect 183796 1748 183802 1760
rect 190273 1751 190331 1757
rect 190273 1748 190285 1751
rect 183796 1720 190285 1748
rect 183796 1708 183802 1720
rect 190273 1717 190285 1720
rect 190319 1717 190331 1751
rect 190273 1711 190331 1717
rect 190362 1708 190368 1760
rect 190420 1748 190426 1760
rect 191006 1748 191012 1760
rect 190420 1720 191012 1748
rect 190420 1708 190426 1720
rect 191006 1708 191012 1720
rect 191064 1708 191070 1760
rect 191190 1748 191196 1760
rect 191151 1720 191196 1748
rect 191190 1708 191196 1720
rect 191248 1708 191254 1760
rect 191285 1751 191343 1757
rect 191285 1717 191297 1751
rect 191331 1748 191343 1751
rect 191653 1751 191711 1757
rect 191653 1748 191665 1751
rect 191331 1720 191665 1748
rect 191331 1717 191343 1720
rect 191285 1711 191343 1717
rect 191653 1717 191665 1720
rect 191699 1717 191711 1751
rect 191653 1711 191711 1717
rect 191742 1708 191748 1760
rect 191800 1748 191806 1760
rect 196897 1751 196955 1757
rect 191800 1720 196848 1748
rect 191800 1708 191806 1720
rect 179046 1680 179052 1692
rect 178696 1652 179052 1680
rect 178589 1643 178647 1649
rect 179046 1640 179052 1652
rect 179104 1640 179110 1692
rect 179138 1640 179144 1692
rect 179196 1680 179202 1692
rect 179233 1683 179291 1689
rect 179233 1680 179245 1683
rect 179196 1652 179245 1680
rect 179196 1640 179202 1652
rect 179233 1649 179245 1652
rect 179279 1649 179291 1683
rect 179233 1643 179291 1649
rect 179322 1640 179328 1692
rect 179380 1640 179386 1692
rect 179506 1640 179512 1692
rect 179564 1680 179570 1692
rect 196820 1689 196848 1720
rect 196897 1717 196909 1751
rect 196943 1748 196955 1751
rect 197173 1751 197231 1757
rect 197173 1748 197185 1751
rect 196943 1720 197185 1748
rect 196943 1717 196955 1720
rect 196897 1711 196955 1717
rect 197173 1717 197185 1720
rect 197219 1717 197231 1751
rect 197173 1711 197231 1717
rect 197357 1751 197415 1757
rect 197357 1717 197369 1751
rect 197403 1748 197415 1751
rect 231489 1751 231547 1757
rect 231489 1748 231501 1751
rect 197403 1720 231501 1748
rect 197403 1717 197415 1720
rect 197357 1711 197415 1717
rect 231489 1717 231501 1720
rect 231535 1717 231547 1751
rect 232240 1748 232268 1788
rect 232593 1785 232605 1788
rect 232639 1785 232651 1819
rect 236733 1819 236791 1825
rect 232593 1779 232651 1785
rect 232700 1788 236684 1816
rect 231489 1711 231547 1717
rect 231964 1720 232268 1748
rect 232409 1751 232467 1757
rect 196621 1683 196679 1689
rect 196621 1680 196633 1683
rect 179564 1652 196633 1680
rect 179564 1640 179570 1652
rect 196621 1649 196633 1652
rect 196667 1649 196679 1683
rect 196621 1643 196679 1649
rect 196805 1683 196863 1689
rect 196805 1649 196817 1683
rect 196851 1649 196863 1683
rect 196805 1643 196863 1649
rect 196989 1683 197047 1689
rect 196989 1649 197001 1683
rect 197035 1680 197047 1683
rect 197035 1652 216720 1680
rect 197035 1649 197047 1652
rect 196989 1643 197047 1649
rect 177853 1615 177911 1621
rect 177853 1612 177865 1615
rect 161155 1584 169708 1612
rect 169772 1584 177865 1612
rect 161155 1581 161167 1584
rect 161109 1575 161167 1581
rect 169772 1544 169800 1584
rect 177853 1581 177865 1584
rect 177899 1581 177911 1615
rect 177853 1575 177911 1581
rect 177945 1615 178003 1621
rect 177945 1581 177957 1615
rect 177991 1612 178003 1615
rect 178678 1612 178684 1624
rect 177991 1584 178684 1612
rect 177991 1581 178003 1584
rect 177945 1575 178003 1581
rect 178678 1572 178684 1584
rect 178736 1572 178742 1624
rect 178770 1572 178776 1624
rect 178828 1612 178834 1624
rect 178957 1615 179015 1621
rect 178828 1584 178873 1612
rect 178828 1572 178834 1584
rect 178957 1581 178969 1615
rect 179003 1612 179015 1615
rect 183922 1612 183928 1624
rect 179003 1584 183928 1612
rect 179003 1581 179015 1584
rect 178957 1575 179015 1581
rect 183922 1572 183928 1584
rect 183980 1572 183986 1624
rect 184017 1615 184075 1621
rect 184017 1581 184029 1615
rect 184063 1581 184075 1615
rect 184017 1575 184075 1581
rect 161032 1516 169800 1544
rect 169846 1504 169852 1556
rect 169904 1544 169910 1556
rect 175737 1547 175795 1553
rect 175737 1544 175749 1547
rect 169904 1516 175749 1544
rect 169904 1504 169910 1516
rect 175737 1513 175749 1516
rect 175783 1513 175795 1547
rect 175737 1507 175795 1513
rect 175829 1547 175887 1553
rect 175829 1513 175841 1547
rect 175875 1544 175887 1547
rect 176565 1547 176623 1553
rect 176565 1544 176577 1547
rect 175875 1516 176577 1544
rect 175875 1513 175887 1516
rect 175829 1507 175887 1513
rect 176565 1513 176577 1516
rect 176611 1513 176623 1547
rect 179877 1547 179935 1553
rect 179877 1544 179889 1547
rect 176565 1507 176623 1513
rect 176672 1516 179889 1544
rect 129384 1448 129688 1476
rect 129737 1479 129795 1485
rect 129277 1439 129335 1445
rect 129737 1445 129749 1479
rect 129783 1476 129795 1479
rect 134153 1479 134211 1485
rect 134153 1476 134165 1479
rect 129783 1448 134165 1476
rect 129783 1445 129795 1448
rect 129737 1439 129795 1445
rect 134153 1445 134165 1448
rect 134199 1445 134211 1479
rect 143997 1479 144055 1485
rect 143997 1476 144009 1479
rect 134153 1439 134211 1445
rect 134352 1448 144009 1476
rect 122064 1380 122236 1408
rect 122285 1411 122343 1417
rect 122064 1368 122070 1380
rect 122285 1377 122297 1411
rect 122331 1408 122343 1411
rect 131761 1411 131819 1417
rect 131761 1408 131773 1411
rect 122331 1380 131773 1408
rect 122331 1377 122343 1380
rect 122285 1371 122343 1377
rect 131761 1377 131773 1380
rect 131807 1377 131819 1411
rect 132589 1411 132647 1417
rect 132589 1408 132601 1411
rect 131761 1371 131819 1377
rect 131868 1380 132601 1408
rect 93121 1343 93179 1349
rect 93121 1309 93133 1343
rect 93167 1340 93179 1343
rect 101861 1343 101919 1349
rect 101861 1340 101873 1343
rect 93167 1312 101873 1340
rect 93167 1309 93179 1312
rect 93121 1303 93179 1309
rect 101861 1309 101873 1312
rect 101907 1309 101919 1343
rect 102226 1340 102232 1352
rect 102187 1312 102232 1340
rect 101861 1303 101919 1309
rect 102226 1300 102232 1312
rect 102284 1300 102290 1352
rect 128173 1343 128231 1349
rect 102336 1312 121592 1340
rect 100294 1272 100300 1284
rect 92768 1244 100300 1272
rect 100294 1232 100300 1244
rect 100352 1232 100358 1284
rect 100389 1275 100447 1281
rect 100389 1241 100401 1275
rect 100435 1272 100447 1275
rect 100665 1275 100723 1281
rect 100665 1272 100677 1275
rect 100435 1244 100677 1272
rect 100435 1241 100447 1244
rect 100389 1235 100447 1241
rect 100665 1241 100677 1244
rect 100711 1241 100723 1275
rect 100665 1235 100723 1241
rect 100757 1275 100815 1281
rect 100757 1241 100769 1275
rect 100803 1272 100815 1275
rect 101950 1272 101956 1284
rect 100803 1244 101956 1272
rect 100803 1241 100815 1244
rect 100757 1235 100815 1241
rect 101950 1232 101956 1244
rect 102008 1232 102014 1284
rect 102045 1275 102103 1281
rect 102045 1241 102057 1275
rect 102091 1272 102103 1275
rect 102336 1272 102364 1312
rect 102091 1244 102364 1272
rect 102413 1275 102471 1281
rect 102091 1241 102103 1244
rect 102045 1235 102103 1241
rect 102413 1241 102425 1275
rect 102459 1272 102471 1275
rect 102689 1275 102747 1281
rect 102689 1272 102701 1275
rect 102459 1244 102701 1272
rect 102459 1241 102471 1244
rect 102413 1235 102471 1241
rect 102689 1241 102701 1244
rect 102735 1241 102747 1275
rect 102689 1235 102747 1241
rect 102778 1232 102784 1284
rect 102836 1272 102842 1284
rect 103241 1275 103299 1281
rect 103241 1272 103253 1275
rect 102836 1244 103253 1272
rect 102836 1232 102842 1244
rect 103241 1241 103253 1244
rect 103287 1241 103299 1275
rect 103241 1235 103299 1241
rect 103330 1232 103336 1284
rect 103388 1272 103394 1284
rect 106642 1272 106648 1284
rect 103388 1244 106648 1272
rect 103388 1232 103394 1244
rect 106642 1232 106648 1244
rect 106700 1232 106706 1284
rect 106826 1232 106832 1284
rect 106884 1272 106890 1284
rect 110414 1272 110420 1284
rect 106884 1244 110420 1272
rect 106884 1232 106890 1244
rect 110414 1232 110420 1244
rect 110472 1232 110478 1284
rect 110598 1232 110604 1284
rect 110656 1272 110662 1284
rect 111150 1272 111156 1284
rect 110656 1244 111156 1272
rect 110656 1232 110662 1244
rect 111150 1232 111156 1244
rect 111208 1232 111214 1284
rect 111245 1275 111303 1281
rect 111245 1241 111257 1275
rect 111291 1272 111303 1275
rect 111797 1275 111855 1281
rect 111797 1272 111809 1275
rect 111291 1244 111809 1272
rect 111291 1241 111303 1244
rect 111245 1235 111303 1241
rect 111797 1241 111809 1244
rect 111843 1241 111855 1275
rect 111797 1235 111855 1241
rect 111886 1232 111892 1284
rect 111944 1272 111950 1284
rect 114925 1275 114983 1281
rect 114925 1272 114937 1275
rect 111944 1244 114937 1272
rect 111944 1232 111950 1244
rect 114925 1241 114937 1244
rect 114971 1241 114983 1275
rect 114925 1235 114983 1241
rect 115017 1275 115075 1281
rect 115017 1241 115029 1275
rect 115063 1272 115075 1275
rect 116486 1272 116492 1284
rect 115063 1244 116492 1272
rect 115063 1241 115075 1244
rect 115017 1235 115075 1241
rect 116486 1232 116492 1244
rect 116544 1232 116550 1284
rect 116670 1272 116676 1284
rect 116631 1244 116676 1272
rect 116670 1232 116676 1244
rect 116728 1232 116734 1284
rect 116762 1232 116768 1284
rect 116820 1272 116826 1284
rect 120997 1275 121055 1281
rect 120997 1272 121009 1275
rect 116820 1244 121009 1272
rect 116820 1232 116826 1244
rect 120997 1241 121009 1244
rect 121043 1241 121055 1275
rect 120997 1235 121055 1241
rect 121089 1275 121147 1281
rect 121089 1241 121101 1275
rect 121135 1272 121147 1275
rect 121362 1272 121368 1284
rect 121135 1244 121368 1272
rect 121135 1241 121147 1244
rect 121089 1235 121147 1241
rect 121362 1232 121368 1244
rect 121420 1232 121426 1284
rect 121564 1272 121592 1312
rect 121932 1312 128124 1340
rect 121932 1272 121960 1312
rect 121564 1244 121960 1272
rect 122101 1275 122159 1281
rect 122101 1241 122113 1275
rect 122147 1272 122159 1275
rect 125413 1275 125471 1281
rect 125413 1272 125425 1275
rect 122147 1244 125425 1272
rect 122147 1241 122159 1244
rect 122101 1235 122159 1241
rect 125413 1241 125425 1244
rect 125459 1241 125471 1275
rect 125413 1235 125471 1241
rect 125505 1275 125563 1281
rect 125505 1241 125517 1275
rect 125551 1272 125563 1275
rect 126057 1275 126115 1281
rect 126057 1272 126069 1275
rect 125551 1244 126069 1272
rect 125551 1241 125563 1244
rect 125505 1235 125563 1241
rect 126057 1241 126069 1244
rect 126103 1241 126115 1275
rect 126057 1235 126115 1241
rect 126146 1232 126152 1284
rect 126204 1272 126210 1284
rect 128096 1281 128124 1312
rect 128173 1309 128185 1343
rect 128219 1340 128231 1343
rect 128630 1340 128636 1352
rect 128219 1312 128636 1340
rect 128219 1309 128231 1312
rect 128173 1303 128231 1309
rect 128630 1300 128636 1312
rect 128688 1300 128694 1352
rect 128725 1343 128783 1349
rect 128725 1309 128737 1343
rect 128771 1309 128783 1343
rect 128906 1340 128912 1352
rect 128867 1312 128912 1340
rect 128725 1303 128783 1309
rect 127989 1275 128047 1281
rect 127989 1272 128001 1275
rect 126204 1244 128001 1272
rect 126204 1232 126210 1244
rect 127989 1241 128001 1244
rect 128035 1241 128047 1275
rect 127989 1235 128047 1241
rect 128081 1275 128139 1281
rect 128081 1241 128093 1275
rect 128127 1241 128139 1275
rect 128081 1235 128139 1241
rect 128538 1232 128544 1284
rect 128596 1272 128602 1284
rect 128740 1272 128768 1303
rect 128906 1300 128912 1312
rect 128964 1300 128970 1352
rect 129274 1300 129280 1352
rect 129332 1340 129338 1352
rect 131868 1340 131896 1380
rect 132589 1377 132601 1380
rect 132635 1377 132647 1411
rect 132589 1371 132647 1377
rect 132773 1411 132831 1417
rect 132773 1377 132785 1411
rect 132819 1408 132831 1411
rect 134352 1408 134380 1448
rect 143997 1445 144009 1448
rect 144043 1445 144055 1479
rect 143997 1439 144055 1445
rect 144273 1479 144331 1485
rect 144273 1445 144285 1479
rect 144319 1476 144331 1479
rect 145009 1479 145067 1485
rect 145009 1476 145021 1479
rect 144319 1448 145021 1476
rect 144319 1445 144331 1448
rect 144273 1439 144331 1445
rect 145009 1445 145021 1448
rect 145055 1445 145067 1479
rect 145558 1476 145564 1488
rect 145519 1448 145564 1476
rect 145009 1439 145067 1445
rect 145558 1436 145564 1448
rect 145616 1436 145622 1488
rect 145653 1479 145711 1485
rect 145653 1445 145665 1479
rect 145699 1476 145711 1479
rect 147401 1479 147459 1485
rect 147401 1476 147413 1479
rect 145699 1448 147413 1476
rect 145699 1445 145711 1448
rect 145653 1439 145711 1445
rect 147401 1445 147413 1448
rect 147447 1445 147459 1479
rect 149238 1476 149244 1488
rect 147401 1439 147459 1445
rect 147508 1448 149244 1476
rect 132819 1380 134380 1408
rect 134429 1411 134487 1417
rect 132819 1377 132831 1380
rect 132773 1371 132831 1377
rect 134429 1377 134441 1411
rect 134475 1408 134487 1411
rect 134705 1411 134763 1417
rect 134705 1408 134717 1411
rect 134475 1380 134717 1408
rect 134475 1377 134487 1380
rect 134429 1371 134487 1377
rect 134705 1377 134717 1380
rect 134751 1377 134763 1411
rect 134705 1371 134763 1377
rect 134794 1368 134800 1420
rect 134852 1408 134858 1420
rect 135806 1408 135812 1420
rect 134852 1380 135812 1408
rect 134852 1368 134858 1380
rect 135806 1368 135812 1380
rect 135864 1368 135870 1420
rect 135901 1411 135959 1417
rect 135901 1377 135913 1411
rect 135947 1408 135959 1411
rect 138661 1411 138719 1417
rect 138661 1408 138673 1411
rect 135947 1380 138673 1408
rect 135947 1377 135959 1380
rect 135901 1371 135959 1377
rect 138661 1377 138673 1380
rect 138707 1377 138719 1411
rect 138661 1371 138719 1377
rect 138750 1368 138756 1420
rect 138808 1408 138814 1420
rect 139118 1408 139124 1420
rect 138808 1380 139124 1408
rect 138808 1368 138814 1380
rect 139118 1368 139124 1380
rect 139176 1368 139182 1420
rect 139210 1368 139216 1420
rect 139268 1408 139274 1420
rect 140314 1408 140320 1420
rect 139268 1380 140320 1408
rect 139268 1368 139274 1380
rect 140314 1368 140320 1380
rect 140372 1368 140378 1420
rect 140406 1368 140412 1420
rect 140464 1408 140470 1420
rect 141142 1408 141148 1420
rect 140464 1380 141148 1408
rect 140464 1368 140470 1380
rect 141142 1368 141148 1380
rect 141200 1368 141206 1420
rect 141237 1411 141295 1417
rect 141237 1377 141249 1411
rect 141283 1408 141295 1411
rect 143077 1411 143135 1417
rect 143077 1408 143089 1411
rect 141283 1380 143089 1408
rect 141283 1377 141295 1380
rect 141237 1371 141295 1377
rect 143077 1377 143089 1380
rect 143123 1377 143135 1411
rect 143077 1371 143135 1377
rect 143629 1411 143687 1417
rect 143629 1377 143641 1411
rect 143675 1408 143687 1411
rect 144089 1411 144147 1417
rect 144089 1408 144101 1411
rect 143675 1380 144101 1408
rect 143675 1377 143687 1380
rect 143629 1371 143687 1377
rect 144089 1377 144101 1380
rect 144135 1377 144147 1411
rect 144089 1371 144147 1377
rect 144178 1368 144184 1420
rect 144236 1408 144242 1420
rect 145098 1408 145104 1420
rect 144236 1380 145104 1408
rect 144236 1368 144242 1380
rect 145098 1368 145104 1380
rect 145156 1368 145162 1420
rect 145190 1368 145196 1420
rect 145248 1408 145254 1420
rect 147508 1408 147536 1448
rect 149238 1436 149244 1448
rect 149296 1436 149302 1488
rect 149333 1479 149391 1485
rect 149333 1445 149345 1479
rect 149379 1476 149391 1479
rect 149422 1476 149428 1488
rect 149379 1448 149428 1476
rect 149379 1445 149391 1448
rect 149333 1439 149391 1445
rect 149422 1436 149428 1448
rect 149480 1436 149486 1488
rect 149517 1479 149575 1485
rect 149517 1445 149529 1479
rect 149563 1476 149575 1479
rect 150437 1479 150495 1485
rect 150437 1476 150449 1479
rect 149563 1448 150449 1476
rect 149563 1445 149575 1448
rect 149517 1439 149575 1445
rect 150437 1445 150449 1448
rect 150483 1445 150495 1479
rect 150437 1439 150495 1445
rect 150529 1479 150587 1485
rect 150529 1445 150541 1479
rect 150575 1476 150587 1479
rect 152550 1476 152556 1488
rect 150575 1448 152556 1476
rect 150575 1445 150587 1448
rect 150529 1439 150587 1445
rect 152550 1436 152556 1448
rect 152608 1436 152614 1488
rect 152645 1479 152703 1485
rect 152645 1445 152657 1479
rect 152691 1476 152703 1479
rect 164053 1479 164111 1485
rect 164053 1476 164065 1479
rect 152691 1448 164065 1476
rect 152691 1445 152703 1448
rect 152645 1439 152703 1445
rect 164053 1445 164065 1448
rect 164099 1445 164111 1479
rect 164053 1439 164111 1445
rect 164145 1479 164203 1485
rect 164145 1445 164157 1479
rect 164191 1476 164203 1479
rect 164513 1479 164571 1485
rect 164513 1476 164525 1479
rect 164191 1448 164525 1476
rect 164191 1445 164203 1448
rect 164145 1439 164203 1445
rect 164513 1445 164525 1448
rect 164559 1445 164571 1479
rect 164513 1439 164571 1445
rect 164605 1479 164663 1485
rect 164605 1445 164617 1479
rect 164651 1445 164663 1479
rect 169297 1479 169355 1485
rect 169297 1476 169309 1479
rect 164605 1439 164663 1445
rect 164804 1448 169309 1476
rect 145248 1380 147536 1408
rect 147769 1411 147827 1417
rect 145248 1368 145254 1380
rect 147769 1377 147781 1411
rect 147815 1408 147827 1411
rect 148781 1411 148839 1417
rect 148781 1408 148793 1411
rect 147815 1380 148793 1408
rect 147815 1377 147827 1380
rect 147769 1371 147827 1377
rect 148781 1377 148793 1380
rect 148827 1377 148839 1411
rect 148781 1371 148839 1377
rect 148870 1368 148876 1420
rect 148928 1408 148934 1420
rect 151357 1411 151415 1417
rect 151357 1408 151369 1411
rect 148928 1380 151369 1408
rect 148928 1368 148934 1380
rect 151357 1377 151369 1380
rect 151403 1377 151415 1411
rect 151357 1371 151415 1377
rect 151449 1411 151507 1417
rect 151449 1377 151461 1411
rect 151495 1408 151507 1411
rect 152737 1411 152795 1417
rect 152737 1408 152749 1411
rect 151495 1380 152749 1408
rect 151495 1377 151507 1380
rect 151449 1371 151507 1377
rect 152737 1377 152749 1380
rect 152783 1377 152795 1411
rect 152737 1371 152795 1377
rect 152829 1411 152887 1417
rect 152829 1377 152841 1411
rect 152875 1408 152887 1411
rect 156509 1411 156567 1417
rect 156509 1408 156521 1411
rect 152875 1380 156521 1408
rect 152875 1377 152887 1380
rect 152829 1371 152887 1377
rect 156509 1377 156521 1380
rect 156555 1377 156567 1411
rect 156509 1371 156567 1377
rect 156601 1411 156659 1417
rect 156601 1377 156613 1411
rect 156647 1408 156659 1411
rect 161937 1411 161995 1417
rect 161937 1408 161949 1411
rect 156647 1380 161949 1408
rect 156647 1377 156659 1380
rect 156601 1371 156659 1377
rect 161937 1377 161949 1380
rect 161983 1377 161995 1411
rect 161937 1371 161995 1377
rect 162121 1411 162179 1417
rect 162121 1377 162133 1411
rect 162167 1408 162179 1411
rect 162854 1408 162860 1420
rect 162167 1380 162860 1408
rect 162167 1377 162179 1380
rect 162121 1371 162179 1377
rect 162854 1368 162860 1380
rect 162912 1368 162918 1420
rect 162949 1411 163007 1417
rect 162949 1377 162961 1411
rect 162995 1408 163007 1411
rect 164620 1408 164648 1439
rect 164804 1417 164832 1448
rect 169297 1445 169309 1448
rect 169343 1445 169355 1479
rect 169297 1439 169355 1445
rect 169386 1436 169392 1488
rect 169444 1476 169450 1488
rect 171502 1476 171508 1488
rect 169444 1448 171508 1476
rect 169444 1436 169450 1448
rect 171502 1436 171508 1448
rect 171560 1436 171566 1488
rect 171597 1479 171655 1485
rect 171597 1445 171609 1479
rect 171643 1476 171655 1479
rect 173437 1479 173495 1485
rect 173437 1476 173449 1479
rect 171643 1448 173449 1476
rect 171643 1445 171655 1448
rect 171597 1439 171655 1445
rect 173437 1445 173449 1448
rect 173483 1445 173495 1479
rect 173437 1439 173495 1445
rect 173529 1479 173587 1485
rect 173529 1445 173541 1479
rect 173575 1445 173587 1479
rect 173529 1439 173587 1445
rect 173713 1479 173771 1485
rect 173713 1445 173725 1479
rect 173759 1476 173771 1479
rect 176672 1476 176700 1516
rect 179877 1513 179889 1516
rect 179923 1513 179935 1547
rect 184032 1544 184060 1575
rect 184198 1572 184204 1624
rect 184256 1612 184262 1624
rect 190825 1615 190883 1621
rect 184256 1584 190776 1612
rect 184256 1572 184262 1584
rect 179877 1507 179935 1513
rect 179984 1516 184060 1544
rect 184109 1547 184167 1553
rect 177850 1476 177856 1488
rect 173759 1448 176700 1476
rect 176764 1448 177856 1476
rect 173759 1445 173771 1448
rect 173713 1439 173771 1445
rect 162995 1380 164648 1408
rect 164789 1411 164847 1417
rect 162995 1377 163007 1380
rect 162949 1371 163007 1377
rect 164789 1377 164801 1411
rect 164835 1377 164847 1411
rect 164789 1371 164847 1377
rect 164881 1411 164939 1417
rect 164881 1377 164893 1411
rect 164927 1408 164939 1411
rect 166721 1411 166779 1417
rect 166721 1408 166733 1411
rect 164927 1380 166733 1408
rect 164927 1377 164939 1380
rect 164881 1371 164939 1377
rect 166721 1377 166733 1380
rect 166767 1377 166779 1411
rect 166721 1371 166779 1377
rect 166810 1368 166816 1420
rect 166868 1408 166874 1420
rect 167270 1408 167276 1420
rect 166868 1380 167276 1408
rect 166868 1368 166874 1380
rect 167270 1368 167276 1380
rect 167328 1368 167334 1420
rect 167362 1368 167368 1420
rect 167420 1408 167426 1420
rect 169202 1408 169208 1420
rect 167420 1380 169208 1408
rect 167420 1368 167426 1380
rect 169202 1368 169208 1380
rect 169260 1368 169266 1420
rect 169481 1411 169539 1417
rect 169481 1377 169493 1411
rect 169527 1408 169539 1411
rect 173544 1408 173572 1439
rect 169527 1380 173572 1408
rect 169527 1377 169539 1380
rect 169481 1371 169539 1377
rect 173618 1368 173624 1420
rect 173676 1408 173682 1420
rect 176473 1411 176531 1417
rect 176473 1408 176485 1411
rect 173676 1380 176485 1408
rect 173676 1368 173682 1380
rect 176473 1377 176485 1380
rect 176519 1377 176531 1411
rect 176473 1371 176531 1377
rect 176565 1411 176623 1417
rect 176565 1377 176577 1411
rect 176611 1408 176623 1411
rect 176764 1408 176792 1448
rect 177850 1436 177856 1448
rect 177908 1436 177914 1488
rect 178037 1479 178095 1485
rect 178037 1445 178049 1479
rect 178083 1476 178095 1479
rect 178957 1479 179015 1485
rect 178957 1476 178969 1479
rect 178083 1448 178969 1476
rect 178083 1445 178095 1448
rect 178037 1439 178095 1445
rect 178957 1445 178969 1448
rect 179003 1445 179015 1479
rect 178957 1439 179015 1445
rect 179141 1479 179199 1485
rect 179141 1445 179153 1479
rect 179187 1476 179199 1479
rect 179984 1476 180012 1516
rect 184109 1513 184121 1547
rect 184155 1544 184167 1547
rect 189445 1547 189503 1553
rect 189445 1544 189457 1547
rect 184155 1516 189457 1544
rect 184155 1513 184167 1516
rect 184109 1507 184167 1513
rect 189445 1513 189457 1516
rect 189491 1513 189503 1547
rect 189445 1507 189503 1513
rect 189537 1547 189595 1553
rect 189537 1513 189549 1547
rect 189583 1544 189595 1547
rect 189902 1544 189908 1556
rect 189583 1516 189908 1544
rect 189583 1513 189595 1516
rect 189537 1507 189595 1513
rect 189902 1504 189908 1516
rect 189960 1504 189966 1556
rect 189994 1504 190000 1556
rect 190052 1504 190058 1556
rect 190086 1504 190092 1556
rect 190144 1544 190150 1556
rect 190546 1544 190552 1556
rect 190144 1516 190552 1544
rect 190144 1504 190150 1516
rect 190546 1504 190552 1516
rect 190604 1504 190610 1556
rect 190748 1544 190776 1584
rect 190825 1581 190837 1615
rect 190871 1612 190883 1615
rect 214101 1615 214159 1621
rect 214101 1612 214113 1615
rect 190871 1584 214113 1612
rect 190871 1581 190883 1584
rect 190825 1575 190883 1581
rect 214101 1581 214113 1584
rect 214147 1581 214159 1615
rect 214101 1575 214159 1581
rect 214190 1572 214196 1624
rect 214248 1612 214254 1624
rect 214377 1615 214435 1621
rect 214377 1612 214389 1615
rect 214248 1584 214389 1612
rect 214248 1572 214254 1584
rect 214377 1581 214389 1584
rect 214423 1581 214435 1615
rect 214377 1575 214435 1581
rect 214466 1572 214472 1624
rect 214524 1612 214530 1624
rect 214837 1615 214895 1621
rect 214837 1612 214849 1615
rect 214524 1584 214849 1612
rect 214524 1572 214530 1584
rect 214837 1581 214849 1584
rect 214883 1581 214895 1615
rect 214837 1575 214895 1581
rect 214926 1572 214932 1624
rect 214984 1612 214990 1624
rect 216582 1612 216588 1624
rect 214984 1584 216588 1612
rect 214984 1572 214990 1584
rect 216582 1572 216588 1584
rect 216640 1572 216646 1624
rect 216692 1612 216720 1652
rect 216766 1640 216772 1692
rect 216824 1680 216830 1692
rect 220170 1680 220176 1692
rect 216824 1652 220176 1680
rect 216824 1640 216830 1652
rect 220170 1640 220176 1652
rect 220228 1640 220234 1692
rect 224037 1683 224095 1689
rect 224037 1680 224049 1683
rect 220280 1652 224049 1680
rect 220280 1612 220308 1652
rect 224037 1649 224049 1652
rect 224083 1649 224095 1683
rect 224589 1683 224647 1689
rect 224589 1680 224601 1683
rect 224037 1643 224095 1649
rect 224144 1652 224601 1680
rect 216692 1584 220308 1612
rect 220357 1615 220415 1621
rect 220357 1581 220369 1615
rect 220403 1612 220415 1615
rect 220633 1615 220691 1621
rect 220633 1612 220645 1615
rect 220403 1584 220645 1612
rect 220403 1581 220415 1584
rect 220357 1575 220415 1581
rect 220633 1581 220645 1584
rect 220679 1581 220691 1615
rect 220633 1575 220691 1581
rect 220725 1615 220783 1621
rect 220725 1581 220737 1615
rect 220771 1581 220783 1615
rect 220725 1575 220783 1581
rect 220909 1615 220967 1621
rect 220909 1581 220921 1615
rect 220955 1612 220967 1615
rect 222013 1615 222071 1621
rect 222013 1612 222025 1615
rect 220955 1584 222025 1612
rect 220955 1581 220967 1584
rect 220909 1575 220967 1581
rect 222013 1581 222025 1584
rect 222059 1581 222071 1615
rect 222013 1575 222071 1581
rect 222105 1615 222163 1621
rect 222105 1581 222117 1615
rect 222151 1612 222163 1615
rect 224144 1612 224172 1652
rect 224589 1649 224601 1652
rect 224635 1649 224647 1683
rect 224589 1643 224647 1649
rect 224681 1683 224739 1689
rect 224681 1649 224693 1683
rect 224727 1680 224739 1683
rect 231765 1683 231823 1689
rect 231765 1680 231777 1683
rect 224727 1652 231777 1680
rect 224727 1649 224739 1652
rect 224681 1643 224739 1649
rect 231765 1649 231777 1652
rect 231811 1649 231823 1683
rect 231765 1643 231823 1649
rect 222151 1584 224172 1612
rect 224405 1615 224463 1621
rect 222151 1581 222163 1584
rect 222105 1575 222163 1581
rect 224405 1581 224417 1615
rect 224451 1612 224463 1615
rect 224957 1615 225015 1621
rect 224451 1584 224724 1612
rect 224451 1581 224463 1584
rect 224405 1575 224463 1581
rect 197814 1544 197820 1556
rect 190748 1516 197820 1544
rect 197814 1504 197820 1516
rect 197872 1504 197878 1556
rect 197909 1547 197967 1553
rect 197909 1513 197921 1547
rect 197955 1544 197967 1547
rect 198550 1544 198556 1556
rect 197955 1516 198556 1544
rect 197955 1513 197967 1516
rect 197909 1507 197967 1513
rect 198550 1504 198556 1516
rect 198608 1504 198614 1556
rect 198737 1547 198795 1553
rect 198737 1513 198749 1547
rect 198783 1544 198795 1547
rect 199102 1544 199108 1556
rect 198783 1516 199108 1544
rect 198783 1513 198795 1516
rect 198737 1507 198795 1513
rect 199102 1504 199108 1516
rect 199160 1504 199166 1556
rect 199197 1547 199255 1553
rect 199197 1513 199209 1547
rect 199243 1544 199255 1547
rect 202877 1547 202935 1553
rect 202877 1544 202889 1547
rect 199243 1516 202889 1544
rect 199243 1513 199255 1516
rect 199197 1507 199255 1513
rect 202877 1513 202889 1516
rect 202923 1513 202935 1547
rect 204622 1544 204628 1556
rect 202877 1507 202935 1513
rect 202984 1516 204628 1544
rect 179187 1448 180012 1476
rect 180429 1479 180487 1485
rect 179187 1445 179199 1448
rect 179141 1439 179199 1445
rect 180429 1445 180441 1479
rect 180475 1476 180487 1479
rect 180705 1479 180763 1485
rect 180705 1476 180717 1479
rect 180475 1448 180717 1476
rect 180475 1445 180487 1448
rect 180429 1439 180487 1445
rect 180705 1445 180717 1448
rect 180751 1445 180763 1479
rect 180705 1439 180763 1445
rect 180797 1479 180855 1485
rect 180797 1445 180809 1479
rect 180843 1476 180855 1479
rect 182545 1479 182603 1485
rect 182545 1476 182557 1479
rect 180843 1448 182557 1476
rect 180843 1445 180855 1448
rect 180797 1439 180855 1445
rect 182545 1445 182557 1448
rect 182591 1445 182603 1479
rect 182545 1439 182603 1445
rect 182634 1436 182640 1488
rect 182692 1476 182698 1488
rect 190012 1476 190040 1504
rect 190362 1476 190368 1488
rect 182692 1448 190040 1476
rect 190323 1448 190368 1476
rect 182692 1436 182698 1448
rect 190362 1436 190368 1448
rect 190420 1436 190426 1488
rect 190641 1479 190699 1485
rect 190641 1445 190653 1479
rect 190687 1476 190699 1479
rect 191006 1476 191012 1488
rect 190687 1448 191012 1476
rect 190687 1445 190699 1448
rect 190641 1439 190699 1445
rect 191006 1436 191012 1448
rect 191064 1436 191070 1488
rect 191101 1479 191159 1485
rect 191101 1445 191113 1479
rect 191147 1476 191159 1479
rect 191282 1476 191288 1488
rect 191147 1448 191288 1476
rect 191147 1445 191159 1448
rect 191101 1439 191159 1445
rect 191282 1436 191288 1448
rect 191340 1436 191346 1488
rect 191377 1479 191435 1485
rect 191377 1445 191389 1479
rect 191423 1476 191435 1479
rect 191561 1479 191619 1485
rect 191561 1476 191573 1479
rect 191423 1448 191573 1476
rect 191423 1445 191435 1448
rect 191377 1439 191435 1445
rect 191561 1445 191573 1448
rect 191607 1445 191619 1479
rect 191561 1439 191619 1445
rect 191650 1436 191656 1488
rect 191708 1476 191714 1488
rect 191708 1448 191753 1476
rect 191708 1436 191714 1448
rect 191834 1436 191840 1488
rect 191892 1476 191898 1488
rect 191929 1479 191987 1485
rect 191929 1476 191941 1479
rect 191892 1448 191941 1476
rect 191892 1436 191898 1448
rect 191929 1445 191941 1448
rect 191975 1445 191987 1479
rect 191929 1439 191987 1445
rect 192110 1436 192116 1488
rect 192168 1476 192174 1488
rect 196526 1476 196532 1488
rect 192168 1448 196532 1476
rect 192168 1436 192174 1448
rect 196526 1436 196532 1448
rect 196584 1436 196590 1488
rect 196621 1479 196679 1485
rect 196621 1445 196633 1479
rect 196667 1476 196679 1479
rect 196897 1479 196955 1485
rect 196897 1476 196909 1479
rect 196667 1448 196909 1476
rect 196667 1445 196679 1448
rect 196621 1439 196679 1445
rect 196897 1445 196909 1448
rect 196943 1445 196955 1479
rect 196897 1439 196955 1445
rect 196986 1436 196992 1488
rect 197044 1476 197050 1488
rect 200206 1476 200212 1488
rect 197044 1448 200212 1476
rect 197044 1436 197050 1448
rect 200206 1436 200212 1448
rect 200264 1436 200270 1488
rect 200853 1479 200911 1485
rect 200853 1445 200865 1479
rect 200899 1476 200911 1479
rect 202984 1476 203012 1516
rect 204622 1504 204628 1516
rect 204680 1504 204686 1556
rect 211065 1547 211123 1553
rect 211065 1544 211077 1547
rect 204732 1516 211077 1544
rect 200899 1448 203012 1476
rect 200899 1445 200911 1448
rect 200853 1439 200911 1445
rect 204530 1436 204536 1488
rect 204588 1476 204594 1488
rect 204732 1476 204760 1516
rect 211065 1513 211077 1516
rect 211111 1513 211123 1547
rect 211065 1507 211123 1513
rect 211157 1547 211215 1553
rect 211157 1513 211169 1547
rect 211203 1544 211215 1547
rect 220740 1544 220768 1575
rect 211203 1516 220768 1544
rect 220817 1547 220875 1553
rect 211203 1513 211215 1516
rect 211157 1507 211215 1513
rect 220817 1513 220829 1547
rect 220863 1544 220875 1547
rect 224313 1547 224371 1553
rect 224313 1544 224325 1547
rect 220863 1516 224325 1544
rect 220863 1513 220875 1516
rect 220817 1507 220875 1513
rect 224313 1513 224325 1516
rect 224359 1513 224371 1547
rect 224696 1544 224724 1584
rect 224957 1581 224969 1615
rect 225003 1612 225015 1615
rect 231964 1612 231992 1720
rect 232409 1717 232421 1751
rect 232455 1748 232467 1751
rect 232700 1748 232728 1788
rect 233510 1748 233516 1760
rect 232455 1720 232728 1748
rect 232792 1720 233516 1748
rect 232455 1717 232467 1720
rect 232409 1711 232467 1717
rect 232133 1683 232191 1689
rect 232133 1649 232145 1683
rect 232179 1680 232191 1683
rect 232792 1680 232820 1720
rect 233510 1708 233516 1720
rect 233568 1708 233574 1760
rect 233973 1751 234031 1757
rect 233973 1717 233985 1751
rect 234019 1748 234031 1751
rect 236546 1748 236552 1760
rect 234019 1720 236552 1748
rect 234019 1717 234031 1720
rect 233973 1711 234031 1717
rect 236546 1708 236552 1720
rect 236604 1708 236610 1760
rect 236656 1748 236684 1788
rect 236733 1785 236745 1819
rect 236779 1816 236791 1819
rect 258445 1819 258503 1825
rect 258445 1816 258457 1819
rect 236779 1788 258457 1816
rect 236779 1785 236791 1788
rect 236733 1779 236791 1785
rect 258445 1785 258457 1788
rect 258491 1785 258503 1819
rect 258445 1779 258503 1785
rect 258537 1819 258595 1825
rect 258537 1785 258549 1819
rect 258583 1816 258595 1819
rect 262033 1819 262091 1825
rect 258583 1788 261984 1816
rect 258583 1785 258595 1788
rect 258537 1779 258595 1785
rect 239125 1751 239183 1757
rect 239125 1748 239137 1751
rect 236656 1720 239137 1748
rect 239125 1717 239137 1720
rect 239171 1717 239183 1751
rect 239125 1711 239183 1717
rect 239309 1751 239367 1757
rect 239309 1717 239321 1751
rect 239355 1748 239367 1751
rect 240045 1751 240103 1757
rect 240045 1748 240057 1751
rect 239355 1720 240057 1748
rect 239355 1717 239367 1720
rect 239309 1711 239367 1717
rect 240045 1717 240057 1720
rect 240091 1717 240103 1751
rect 240045 1711 240103 1717
rect 240134 1708 240140 1760
rect 240192 1748 240198 1760
rect 241514 1748 241520 1760
rect 240192 1720 241520 1748
rect 240192 1708 240198 1720
rect 241514 1708 241520 1720
rect 241572 1708 241578 1760
rect 241609 1751 241667 1757
rect 241609 1717 241621 1751
rect 241655 1748 241667 1751
rect 250073 1751 250131 1757
rect 250073 1748 250085 1751
rect 241655 1720 250085 1748
rect 241655 1717 241667 1720
rect 241609 1711 241667 1717
rect 250073 1717 250085 1720
rect 250119 1717 250131 1751
rect 250073 1711 250131 1717
rect 250162 1708 250168 1760
rect 250220 1748 250226 1760
rect 250809 1751 250867 1757
rect 250809 1748 250821 1751
rect 250220 1720 250821 1748
rect 250220 1708 250226 1720
rect 250809 1717 250821 1720
rect 250855 1717 250867 1751
rect 250809 1711 250867 1717
rect 250901 1751 250959 1757
rect 250901 1717 250913 1751
rect 250947 1748 250959 1751
rect 251453 1751 251511 1757
rect 251453 1748 251465 1751
rect 250947 1720 251465 1748
rect 250947 1717 250959 1720
rect 250901 1711 250959 1717
rect 251453 1717 251465 1720
rect 251499 1717 251511 1751
rect 251453 1711 251511 1717
rect 251545 1751 251603 1757
rect 251545 1717 251557 1751
rect 251591 1748 251603 1751
rect 252557 1751 252615 1757
rect 252557 1748 252569 1751
rect 251591 1720 252569 1748
rect 251591 1717 251603 1720
rect 251545 1711 251603 1717
rect 252557 1717 252569 1720
rect 252603 1717 252615 1751
rect 252557 1711 252615 1717
rect 252649 1751 252707 1757
rect 252649 1717 252661 1751
rect 252695 1748 252707 1751
rect 253569 1751 253627 1757
rect 253569 1748 253581 1751
rect 252695 1720 253581 1748
rect 252695 1717 252707 1720
rect 252649 1711 252707 1717
rect 253569 1717 253581 1720
rect 253615 1717 253627 1751
rect 253569 1711 253627 1717
rect 253658 1708 253664 1760
rect 253716 1748 253722 1760
rect 257062 1748 257068 1760
rect 253716 1720 257068 1748
rect 253716 1708 253722 1720
rect 257062 1708 257068 1720
rect 257120 1708 257126 1760
rect 257157 1751 257215 1757
rect 257157 1717 257169 1751
rect 257203 1748 257215 1751
rect 258169 1751 258227 1757
rect 258169 1748 258181 1751
rect 257203 1720 258181 1748
rect 257203 1717 257215 1720
rect 257157 1711 257215 1717
rect 258169 1717 258181 1720
rect 258215 1717 258227 1751
rect 258169 1711 258227 1717
rect 258353 1751 258411 1757
rect 258353 1717 258365 1751
rect 258399 1748 258411 1751
rect 261849 1751 261907 1757
rect 261849 1748 261861 1751
rect 258399 1720 261861 1748
rect 258399 1717 258411 1720
rect 258353 1711 258411 1717
rect 261849 1717 261861 1720
rect 261895 1717 261907 1751
rect 261849 1711 261907 1717
rect 232179 1652 232820 1680
rect 233329 1683 233387 1689
rect 232179 1649 232191 1652
rect 232133 1643 232191 1649
rect 233329 1649 233341 1683
rect 233375 1680 233387 1683
rect 258261 1683 258319 1689
rect 258261 1680 258273 1683
rect 233375 1652 258273 1680
rect 233375 1649 233387 1652
rect 233329 1643 233387 1649
rect 258261 1649 258273 1652
rect 258307 1649 258319 1683
rect 258261 1643 258319 1649
rect 258442 1640 258448 1692
rect 258500 1680 258506 1692
rect 260653 1683 260711 1689
rect 260653 1680 260665 1683
rect 258500 1652 260665 1680
rect 258500 1640 258506 1652
rect 260653 1649 260665 1652
rect 260699 1649 260711 1683
rect 260653 1643 260711 1649
rect 260742 1640 260748 1692
rect 260800 1680 260806 1692
rect 261294 1680 261300 1692
rect 260800 1652 261300 1680
rect 260800 1640 260806 1652
rect 261294 1640 261300 1652
rect 261352 1640 261358 1692
rect 261389 1683 261447 1689
rect 261389 1649 261401 1683
rect 261435 1680 261447 1683
rect 261754 1680 261760 1692
rect 261435 1652 261760 1680
rect 261435 1649 261447 1652
rect 261389 1643 261447 1649
rect 261754 1640 261760 1652
rect 261812 1640 261818 1692
rect 261956 1680 261984 1788
rect 262033 1785 262045 1819
rect 262079 1816 262091 1819
rect 263229 1819 263287 1825
rect 262079 1788 262628 1816
rect 262079 1785 262091 1788
rect 262033 1779 262091 1785
rect 262306 1708 262312 1760
rect 262364 1748 262370 1760
rect 262493 1751 262551 1757
rect 262364 1720 262409 1748
rect 262364 1708 262370 1720
rect 262493 1717 262505 1751
rect 262539 1717 262551 1751
rect 262600 1748 262628 1788
rect 263229 1785 263241 1819
rect 263275 1816 263287 1819
rect 268933 1819 268991 1825
rect 263275 1788 268884 1816
rect 263275 1785 263287 1788
rect 263229 1779 263287 1785
rect 268749 1751 268807 1757
rect 268749 1748 268761 1751
rect 262600 1720 268761 1748
rect 262493 1711 262551 1717
rect 268749 1717 268761 1720
rect 268795 1717 268807 1751
rect 268856 1748 268884 1788
rect 268933 1785 268945 1819
rect 268979 1816 268991 1819
rect 368385 1819 368443 1825
rect 268979 1788 367784 1816
rect 268979 1785 268991 1788
rect 268933 1779 268991 1785
rect 279973 1751 280031 1757
rect 279973 1748 279985 1751
rect 268856 1720 279985 1748
rect 268749 1711 268807 1717
rect 279973 1717 279985 1720
rect 280019 1717 280031 1751
rect 279973 1711 280031 1717
rect 262508 1680 262536 1711
rect 280062 1708 280068 1760
rect 280120 1748 280126 1760
rect 280157 1751 280215 1757
rect 280157 1748 280169 1751
rect 280120 1720 280169 1748
rect 280120 1708 280126 1720
rect 280157 1717 280169 1720
rect 280203 1717 280215 1751
rect 280157 1711 280215 1717
rect 280246 1708 280252 1760
rect 280304 1748 280310 1760
rect 289725 1751 289783 1757
rect 289725 1748 289737 1751
rect 280304 1720 289737 1748
rect 280304 1708 280310 1720
rect 289725 1717 289737 1720
rect 289771 1717 289783 1751
rect 289725 1711 289783 1717
rect 290274 1708 290280 1760
rect 290332 1748 290338 1760
rect 290461 1751 290519 1757
rect 290461 1748 290473 1751
rect 290332 1720 290473 1748
rect 290332 1708 290338 1720
rect 290461 1717 290473 1720
rect 290507 1717 290519 1751
rect 290461 1711 290519 1717
rect 293865 1751 293923 1757
rect 293865 1717 293877 1751
rect 293911 1748 293923 1751
rect 295153 1751 295211 1757
rect 295153 1748 295165 1751
rect 293911 1720 295165 1748
rect 293911 1717 293923 1720
rect 293865 1711 293923 1717
rect 295153 1717 295165 1720
rect 295199 1717 295211 1751
rect 295153 1711 295211 1717
rect 295245 1751 295303 1757
rect 295245 1717 295257 1751
rect 295291 1748 295303 1751
rect 337838 1748 337844 1760
rect 295291 1720 337844 1748
rect 295291 1717 295303 1720
rect 295245 1711 295303 1717
rect 337838 1708 337844 1720
rect 337896 1708 337902 1760
rect 337933 1751 337991 1757
rect 337933 1717 337945 1751
rect 337979 1748 337991 1751
rect 348973 1751 349031 1757
rect 348973 1748 348985 1751
rect 337979 1720 348985 1748
rect 337979 1717 337991 1720
rect 337933 1711 337991 1717
rect 348973 1717 348985 1720
rect 349019 1717 349031 1751
rect 348973 1711 349031 1717
rect 349433 1751 349491 1757
rect 349433 1717 349445 1751
rect 349479 1748 349491 1751
rect 352837 1751 352895 1757
rect 352837 1748 352849 1751
rect 349479 1720 352849 1748
rect 349479 1717 349491 1720
rect 349433 1711 349491 1717
rect 352837 1717 352849 1720
rect 352883 1717 352895 1751
rect 352837 1711 352895 1717
rect 352926 1708 352932 1760
rect 352984 1748 352990 1760
rect 366358 1748 366364 1760
rect 352984 1720 366364 1748
rect 352984 1708 352990 1720
rect 366358 1708 366364 1720
rect 366416 1708 366422 1760
rect 367756 1748 367784 1788
rect 368385 1785 368397 1819
rect 368431 1816 368443 1819
rect 374825 1819 374883 1825
rect 374825 1816 374837 1819
rect 368431 1788 374837 1816
rect 368431 1785 368443 1788
rect 368385 1779 368443 1785
rect 374825 1785 374837 1788
rect 374871 1785 374883 1819
rect 374825 1779 374883 1785
rect 388441 1819 388499 1825
rect 388441 1785 388453 1819
rect 388487 1816 388499 1819
rect 391569 1819 391627 1825
rect 391569 1816 391581 1819
rect 388487 1788 391581 1816
rect 388487 1785 388499 1788
rect 388441 1779 388499 1785
rect 391569 1785 391581 1788
rect 391615 1785 391627 1819
rect 391569 1779 391627 1785
rect 569034 1776 569040 1828
rect 569092 1816 569098 1828
rect 569218 1816 569224 1828
rect 569092 1788 569224 1816
rect 569092 1776 569098 1788
rect 569218 1776 569224 1788
rect 569276 1776 569282 1828
rect 375926 1748 375932 1760
rect 367756 1720 375932 1748
rect 375926 1708 375932 1720
rect 375984 1708 375990 1760
rect 376021 1751 376079 1757
rect 376021 1717 376033 1751
rect 376067 1748 376079 1751
rect 404446 1748 404452 1760
rect 376067 1720 404452 1748
rect 376067 1717 376079 1720
rect 376021 1711 376079 1717
rect 404446 1708 404452 1720
rect 404504 1708 404510 1760
rect 474918 1708 474924 1760
rect 474976 1748 474982 1760
rect 481266 1748 481272 1760
rect 474976 1720 481272 1748
rect 474976 1708 474982 1720
rect 481266 1708 481272 1720
rect 481324 1708 481330 1760
rect 488994 1708 489000 1760
rect 489052 1748 489058 1760
rect 501782 1748 501788 1760
rect 489052 1720 501788 1748
rect 489052 1708 489058 1720
rect 501782 1708 501788 1720
rect 501840 1708 501846 1760
rect 512362 1708 512368 1760
rect 512420 1748 512426 1760
rect 529382 1748 529388 1760
rect 512420 1720 529388 1748
rect 512420 1708 512426 1720
rect 529382 1708 529388 1720
rect 529440 1708 529446 1760
rect 559098 1708 559104 1760
rect 559156 1748 559162 1760
rect 567286 1748 567292 1760
rect 559156 1720 567292 1748
rect 559156 1708 559162 1720
rect 567286 1708 567292 1720
rect 567344 1708 567350 1760
rect 568298 1748 568304 1760
rect 568259 1720 568304 1748
rect 568298 1708 568304 1720
rect 568356 1708 568362 1760
rect 261956 1652 262536 1680
rect 262861 1683 262919 1689
rect 262861 1649 262873 1683
rect 262907 1680 262919 1683
rect 296806 1680 296812 1692
rect 262907 1652 296812 1680
rect 262907 1649 262919 1652
rect 262861 1643 262919 1649
rect 296806 1640 296812 1652
rect 296864 1640 296870 1692
rect 296901 1683 296959 1689
rect 296901 1649 296913 1683
rect 296947 1680 296959 1683
rect 298373 1683 298431 1689
rect 298373 1680 298385 1683
rect 296947 1652 298385 1680
rect 296947 1649 296959 1652
rect 296901 1643 296959 1649
rect 298373 1649 298385 1652
rect 298419 1649 298431 1683
rect 298373 1643 298431 1649
rect 298465 1683 298523 1689
rect 298465 1649 298477 1683
rect 298511 1680 298523 1683
rect 299934 1680 299940 1692
rect 298511 1652 299940 1680
rect 298511 1649 298523 1652
rect 298465 1643 298523 1649
rect 299934 1640 299940 1652
rect 299992 1640 299998 1692
rect 300029 1683 300087 1689
rect 300029 1649 300041 1683
rect 300075 1680 300087 1683
rect 304077 1683 304135 1689
rect 304077 1680 304089 1683
rect 300075 1652 304089 1680
rect 300075 1649 300087 1652
rect 300029 1643 300087 1649
rect 304077 1649 304089 1652
rect 304123 1649 304135 1683
rect 304077 1643 304135 1649
rect 304169 1683 304227 1689
rect 304169 1649 304181 1683
rect 304215 1680 304227 1683
rect 314657 1683 314715 1689
rect 314657 1680 314669 1683
rect 304215 1652 314669 1680
rect 304215 1649 304227 1652
rect 304169 1643 304227 1649
rect 314657 1649 314669 1652
rect 314703 1649 314715 1683
rect 314657 1643 314715 1649
rect 314746 1640 314752 1692
rect 314804 1680 314810 1692
rect 319714 1680 319720 1692
rect 314804 1652 319720 1680
rect 314804 1640 314810 1652
rect 319714 1640 319720 1652
rect 319772 1640 319778 1692
rect 319809 1683 319867 1689
rect 319809 1649 319821 1683
rect 319855 1680 319867 1683
rect 345753 1683 345811 1689
rect 345753 1680 345765 1683
rect 319855 1652 345765 1680
rect 319855 1649 319867 1652
rect 319809 1643 319867 1649
rect 345753 1649 345765 1652
rect 345799 1649 345811 1683
rect 345753 1643 345811 1649
rect 348694 1640 348700 1692
rect 348752 1680 348758 1692
rect 358081 1683 358139 1689
rect 358081 1680 358093 1683
rect 348752 1652 358093 1680
rect 348752 1640 348758 1652
rect 358081 1649 358093 1652
rect 358127 1649 358139 1683
rect 358081 1643 358139 1649
rect 358170 1640 358176 1692
rect 358228 1680 358234 1692
rect 413830 1680 413836 1692
rect 358228 1652 413836 1680
rect 358228 1640 358234 1652
rect 413830 1640 413836 1652
rect 413888 1640 413894 1692
rect 415670 1640 415676 1692
rect 415728 1680 415734 1692
rect 418798 1680 418804 1692
rect 415728 1652 418804 1680
rect 415728 1640 415734 1652
rect 418798 1640 418804 1652
rect 418856 1640 418862 1692
rect 432322 1640 432328 1692
rect 432380 1680 432386 1692
rect 443638 1680 443644 1692
rect 432380 1652 443644 1680
rect 432380 1640 432386 1652
rect 443638 1640 443644 1652
rect 443696 1640 443702 1692
rect 453298 1640 453304 1692
rect 453356 1680 453362 1692
rect 462866 1680 462872 1692
rect 453356 1652 462872 1680
rect 453356 1640 453362 1652
rect 462866 1640 462872 1652
rect 462924 1640 462930 1692
rect 509050 1640 509056 1692
rect 509108 1680 509114 1692
rect 528189 1683 528247 1689
rect 528189 1680 528201 1683
rect 509108 1652 528201 1680
rect 509108 1640 509114 1652
rect 528189 1649 528201 1652
rect 528235 1649 528247 1683
rect 528189 1643 528247 1649
rect 557994 1640 558000 1692
rect 558052 1680 558058 1692
rect 569770 1680 569776 1692
rect 558052 1652 569776 1680
rect 558052 1640 558058 1652
rect 569770 1640 569776 1652
rect 569828 1640 569834 1692
rect 225003 1584 231992 1612
rect 225003 1581 225015 1584
rect 224957 1575 225015 1581
rect 232038 1572 232044 1624
rect 232096 1612 232102 1624
rect 232498 1612 232504 1624
rect 232096 1584 232504 1612
rect 232096 1572 232102 1584
rect 232498 1572 232504 1584
rect 232556 1572 232562 1624
rect 232593 1615 232651 1621
rect 232593 1581 232605 1615
rect 232639 1612 232651 1615
rect 233973 1615 234031 1621
rect 233973 1612 233985 1615
rect 232639 1584 233985 1612
rect 232639 1581 232651 1584
rect 232593 1575 232651 1581
rect 233973 1581 233985 1584
rect 234019 1581 234031 1615
rect 233973 1575 234031 1581
rect 234062 1572 234068 1624
rect 234120 1612 234126 1624
rect 237926 1612 237932 1624
rect 234120 1584 237932 1612
rect 234120 1572 234126 1584
rect 237926 1572 237932 1584
rect 237984 1572 237990 1624
rect 238110 1572 238116 1624
rect 238168 1612 238174 1624
rect 238662 1612 238668 1624
rect 238168 1584 238668 1612
rect 238168 1572 238174 1584
rect 238662 1572 238668 1584
rect 238720 1572 238726 1624
rect 238754 1572 238760 1624
rect 238812 1612 238818 1624
rect 260285 1615 260343 1621
rect 260285 1612 260297 1615
rect 238812 1584 260297 1612
rect 238812 1572 238818 1584
rect 260285 1581 260297 1584
rect 260331 1581 260343 1615
rect 260837 1615 260895 1621
rect 260285 1575 260343 1581
rect 260392 1584 260788 1612
rect 260392 1544 260420 1584
rect 260760 1544 260788 1584
rect 260837 1581 260849 1615
rect 260883 1612 260895 1615
rect 262217 1615 262275 1621
rect 262217 1612 262229 1615
rect 260883 1584 262229 1612
rect 260883 1581 260895 1584
rect 260837 1575 260895 1581
rect 262217 1581 262229 1584
rect 262263 1581 262275 1615
rect 262217 1575 262275 1581
rect 262306 1572 262312 1624
rect 262364 1612 262370 1624
rect 262401 1615 262459 1621
rect 262401 1612 262413 1615
rect 262364 1584 262413 1612
rect 262364 1572 262370 1584
rect 262401 1581 262413 1584
rect 262447 1581 262459 1615
rect 262401 1575 262459 1581
rect 262769 1615 262827 1621
rect 262769 1581 262781 1615
rect 262815 1612 262827 1615
rect 270497 1615 270555 1621
rect 270497 1612 270509 1615
rect 262815 1584 270509 1612
rect 262815 1581 262827 1584
rect 262769 1575 262827 1581
rect 270497 1581 270509 1584
rect 270543 1581 270555 1615
rect 270497 1575 270555 1581
rect 272150 1572 272156 1624
rect 272208 1612 272214 1624
rect 273898 1612 273904 1624
rect 272208 1584 273904 1612
rect 272208 1572 272214 1584
rect 273898 1572 273904 1584
rect 273956 1572 273962 1624
rect 273990 1572 273996 1624
rect 274048 1612 274054 1624
rect 280246 1612 280252 1624
rect 274048 1584 280252 1612
rect 274048 1572 274054 1584
rect 280246 1572 280252 1584
rect 280304 1572 280310 1624
rect 280341 1615 280399 1621
rect 280341 1581 280353 1615
rect 280387 1612 280399 1615
rect 280522 1612 280528 1624
rect 280387 1584 280528 1612
rect 280387 1581 280399 1584
rect 280341 1575 280399 1581
rect 280522 1572 280528 1584
rect 280580 1572 280586 1624
rect 280617 1615 280675 1621
rect 280617 1581 280629 1615
rect 280663 1612 280675 1615
rect 290366 1612 290372 1624
rect 280663 1584 290372 1612
rect 280663 1581 280675 1584
rect 280617 1575 280675 1581
rect 290366 1572 290372 1584
rect 290424 1572 290430 1624
rect 290461 1615 290519 1621
rect 290461 1581 290473 1615
rect 290507 1612 290519 1615
rect 290918 1612 290924 1624
rect 290507 1584 290924 1612
rect 290507 1581 290519 1584
rect 290461 1575 290519 1581
rect 290918 1572 290924 1584
rect 290976 1572 290982 1624
rect 291013 1615 291071 1621
rect 291013 1581 291025 1615
rect 291059 1612 291071 1615
rect 293678 1612 293684 1624
rect 291059 1584 293684 1612
rect 291059 1581 291071 1584
rect 291013 1575 291071 1581
rect 293678 1572 293684 1584
rect 293736 1572 293742 1624
rect 293773 1615 293831 1621
rect 293773 1581 293785 1615
rect 293819 1612 293831 1615
rect 298833 1615 298891 1621
rect 293819 1584 298784 1612
rect 293819 1581 293831 1584
rect 293773 1575 293831 1581
rect 285766 1544 285772 1556
rect 224313 1507 224371 1513
rect 224420 1516 224632 1544
rect 224696 1516 232084 1544
rect 204588 1448 204760 1476
rect 204588 1436 204594 1448
rect 204806 1436 204812 1488
rect 204864 1476 204870 1488
rect 211338 1476 211344 1488
rect 204864 1448 211344 1476
rect 204864 1436 204870 1448
rect 211338 1436 211344 1448
rect 211396 1436 211402 1488
rect 211433 1479 211491 1485
rect 211433 1445 211445 1479
rect 211479 1476 211491 1479
rect 220173 1479 220231 1485
rect 220173 1476 220185 1479
rect 211479 1448 220185 1476
rect 211479 1445 211491 1448
rect 211433 1439 211491 1445
rect 220173 1445 220185 1448
rect 220219 1445 220231 1479
rect 220173 1439 220231 1445
rect 220357 1479 220415 1485
rect 220357 1445 220369 1479
rect 220403 1476 220415 1479
rect 224420 1476 224448 1516
rect 220403 1448 224448 1476
rect 220403 1445 220415 1448
rect 220357 1439 220415 1445
rect 176611 1380 176792 1408
rect 176841 1411 176899 1417
rect 176611 1377 176623 1380
rect 176565 1371 176623 1377
rect 176841 1377 176853 1411
rect 176887 1408 176899 1411
rect 177482 1408 177488 1420
rect 176887 1380 177488 1408
rect 176887 1377 176899 1380
rect 176841 1371 176899 1377
rect 177482 1368 177488 1380
rect 177540 1368 177546 1420
rect 177577 1411 177635 1417
rect 177577 1377 177589 1411
rect 177623 1408 177635 1411
rect 177945 1411 178003 1417
rect 177945 1408 177957 1411
rect 177623 1380 177957 1408
rect 177623 1377 177635 1380
rect 177577 1371 177635 1377
rect 177945 1377 177957 1380
rect 177991 1377 178003 1411
rect 177945 1371 178003 1377
rect 178681 1411 178739 1417
rect 178681 1377 178693 1411
rect 178727 1408 178739 1411
rect 179782 1408 179788 1420
rect 178727 1380 179788 1408
rect 178727 1377 178739 1380
rect 178681 1371 178739 1377
rect 179782 1368 179788 1380
rect 179840 1368 179846 1420
rect 179874 1368 179880 1420
rect 179932 1408 179938 1420
rect 180061 1411 180119 1417
rect 179932 1380 179977 1408
rect 179932 1368 179938 1380
rect 180061 1377 180073 1411
rect 180107 1408 180119 1411
rect 189813 1411 189871 1417
rect 189813 1408 189825 1411
rect 180107 1380 189825 1408
rect 180107 1377 180119 1380
rect 180061 1371 180119 1377
rect 189813 1377 189825 1380
rect 189859 1377 189871 1411
rect 189813 1371 189871 1377
rect 189997 1411 190055 1417
rect 189997 1377 190009 1411
rect 190043 1408 190055 1411
rect 190457 1411 190515 1417
rect 190457 1408 190469 1411
rect 190043 1380 190469 1408
rect 190043 1377 190055 1380
rect 189997 1371 190055 1377
rect 190457 1377 190469 1380
rect 190503 1377 190515 1411
rect 190457 1371 190515 1377
rect 190549 1411 190607 1417
rect 190549 1377 190561 1411
rect 190595 1408 190607 1411
rect 217686 1408 217692 1420
rect 190595 1380 217692 1408
rect 190595 1377 190607 1380
rect 190549 1371 190607 1377
rect 217686 1368 217692 1380
rect 217744 1368 217750 1420
rect 217781 1411 217839 1417
rect 217781 1377 217793 1411
rect 217827 1408 217839 1411
rect 218054 1408 218060 1420
rect 217827 1380 218060 1408
rect 217827 1377 217839 1380
rect 217781 1371 217839 1377
rect 218054 1368 218060 1380
rect 218112 1368 218118 1420
rect 218333 1411 218391 1417
rect 218333 1377 218345 1411
rect 218379 1408 218391 1411
rect 218422 1408 218428 1420
rect 218379 1380 218428 1408
rect 218379 1377 218391 1380
rect 218333 1371 218391 1377
rect 218422 1368 218428 1380
rect 218480 1368 218486 1420
rect 218701 1411 218759 1417
rect 218701 1408 218713 1411
rect 218532 1380 218713 1408
rect 129332 1312 131896 1340
rect 131945 1343 132003 1349
rect 129332 1300 129338 1312
rect 131945 1309 131957 1343
rect 131991 1340 132003 1343
rect 150250 1340 150256 1352
rect 131991 1312 150256 1340
rect 131991 1309 132003 1312
rect 131945 1303 132003 1309
rect 150250 1300 150256 1312
rect 150308 1300 150314 1352
rect 150360 1312 151860 1340
rect 128596 1244 128768 1272
rect 128817 1275 128875 1281
rect 128596 1232 128602 1244
rect 128817 1241 128829 1275
rect 128863 1272 128875 1275
rect 129185 1275 129243 1281
rect 129185 1272 129197 1275
rect 128863 1244 129197 1272
rect 128863 1241 128875 1244
rect 128817 1235 128875 1241
rect 129185 1241 129197 1244
rect 129231 1241 129243 1275
rect 129185 1235 129243 1241
rect 129369 1275 129427 1281
rect 129369 1241 129381 1275
rect 129415 1272 129427 1275
rect 134429 1275 134487 1281
rect 134429 1272 134441 1275
rect 129415 1244 134441 1272
rect 129415 1241 129427 1244
rect 129369 1235 129427 1241
rect 134429 1241 134441 1244
rect 134475 1241 134487 1275
rect 134429 1235 134487 1241
rect 134610 1232 134616 1284
rect 134668 1272 134674 1284
rect 134705 1275 134763 1281
rect 134705 1272 134717 1275
rect 134668 1244 134717 1272
rect 134668 1232 134674 1244
rect 134705 1241 134717 1244
rect 134751 1241 134763 1275
rect 134705 1235 134763 1241
rect 134794 1232 134800 1284
rect 134852 1272 134858 1284
rect 135349 1275 135407 1281
rect 135349 1272 135361 1275
rect 134852 1244 135361 1272
rect 134852 1232 134858 1244
rect 135349 1241 135361 1244
rect 135395 1241 135407 1275
rect 135349 1235 135407 1241
rect 135533 1275 135591 1281
rect 135533 1241 135545 1275
rect 135579 1272 135591 1275
rect 140774 1272 140780 1284
rect 135579 1244 140780 1272
rect 135579 1241 135591 1244
rect 135533 1235 135591 1241
rect 140774 1232 140780 1244
rect 140832 1232 140838 1284
rect 140869 1275 140927 1281
rect 140869 1241 140881 1275
rect 140915 1272 140927 1275
rect 142798 1272 142804 1284
rect 140915 1244 142804 1272
rect 140915 1241 140927 1244
rect 140869 1235 140927 1241
rect 142798 1232 142804 1244
rect 142856 1232 142862 1284
rect 142893 1275 142951 1281
rect 142893 1241 142905 1275
rect 142939 1272 142951 1275
rect 150360 1272 150388 1312
rect 142939 1244 150388 1272
rect 150437 1275 150495 1281
rect 142939 1241 142951 1244
rect 142893 1235 142951 1241
rect 150437 1241 150449 1275
rect 150483 1272 150495 1275
rect 151081 1275 151139 1281
rect 151081 1272 151093 1275
rect 150483 1244 151093 1272
rect 150483 1241 150495 1244
rect 150437 1235 150495 1241
rect 151081 1241 151093 1244
rect 151127 1241 151139 1275
rect 151081 1235 151139 1241
rect 151265 1275 151323 1281
rect 151265 1241 151277 1275
rect 151311 1272 151323 1275
rect 151725 1275 151783 1281
rect 151725 1272 151737 1275
rect 151311 1244 151737 1272
rect 151311 1241 151323 1244
rect 151265 1235 151323 1241
rect 151725 1241 151737 1244
rect 151771 1241 151783 1275
rect 151832 1272 151860 1312
rect 151906 1300 151912 1352
rect 151964 1340 151970 1352
rect 175737 1343 175795 1349
rect 175737 1340 175749 1343
rect 151964 1312 152228 1340
rect 151964 1300 151970 1312
rect 152090 1272 152096 1284
rect 151832 1244 152096 1272
rect 151725 1235 151783 1241
rect 152090 1232 152096 1244
rect 152148 1232 152154 1284
rect 152200 1272 152228 1312
rect 152476 1312 175749 1340
rect 152476 1272 152504 1312
rect 175737 1309 175749 1312
rect 175783 1309 175795 1343
rect 175737 1303 175795 1309
rect 175921 1343 175979 1349
rect 175921 1309 175933 1343
rect 175967 1340 175979 1343
rect 175967 1312 189948 1340
rect 175967 1309 175979 1312
rect 175921 1303 175979 1309
rect 152200 1244 152504 1272
rect 152553 1275 152611 1281
rect 152553 1241 152565 1275
rect 152599 1272 152611 1275
rect 152642 1272 152648 1284
rect 152599 1244 152648 1272
rect 152599 1241 152611 1244
rect 152553 1235 152611 1241
rect 152642 1232 152648 1244
rect 152700 1232 152706 1284
rect 152737 1275 152795 1281
rect 152737 1241 152749 1275
rect 152783 1272 152795 1275
rect 153013 1275 153071 1281
rect 152783 1244 152964 1272
rect 152783 1241 152795 1244
rect 152737 1235 152795 1241
rect 86144 1176 87828 1204
rect 85761 1167 85819 1173
rect 87874 1164 87880 1216
rect 87932 1204 87938 1216
rect 87932 1176 87977 1204
rect 87932 1164 87938 1176
rect 88150 1164 88156 1216
rect 88208 1204 88214 1216
rect 88518 1204 88524 1216
rect 88208 1176 88524 1204
rect 88208 1164 88214 1176
rect 88518 1164 88524 1176
rect 88576 1164 88582 1216
rect 88610 1164 88616 1216
rect 88668 1204 88674 1216
rect 91649 1207 91707 1213
rect 91649 1204 91661 1207
rect 88668 1176 91661 1204
rect 88668 1164 88674 1176
rect 91649 1173 91661 1176
rect 91695 1173 91707 1207
rect 91649 1167 91707 1173
rect 91741 1207 91799 1213
rect 91741 1173 91753 1207
rect 91787 1204 91799 1207
rect 92109 1207 92167 1213
rect 92109 1204 92121 1207
rect 91787 1176 92121 1204
rect 91787 1173 91799 1176
rect 91741 1167 91799 1173
rect 92109 1173 92121 1176
rect 92155 1173 92167 1207
rect 92109 1167 92167 1173
rect 92198 1164 92204 1216
rect 92256 1204 92262 1216
rect 93118 1204 93124 1216
rect 92256 1176 93124 1204
rect 92256 1164 92262 1176
rect 93118 1164 93124 1176
rect 93176 1164 93182 1216
rect 93305 1207 93363 1213
rect 93305 1173 93317 1207
rect 93351 1204 93363 1207
rect 104529 1207 104587 1213
rect 104529 1204 104541 1207
rect 93351 1176 104541 1204
rect 93351 1173 93363 1176
rect 93305 1167 93363 1173
rect 104529 1173 104541 1176
rect 104575 1173 104587 1207
rect 104529 1167 104587 1173
rect 104618 1164 104624 1216
rect 104676 1204 104682 1216
rect 106277 1207 106335 1213
rect 106277 1204 106289 1207
rect 104676 1176 106289 1204
rect 104676 1164 104682 1176
rect 106277 1173 106289 1176
rect 106323 1173 106335 1207
rect 106277 1167 106335 1173
rect 106550 1164 106556 1216
rect 106608 1204 106614 1216
rect 110506 1204 110512 1216
rect 106608 1176 110512 1204
rect 106608 1164 106614 1176
rect 110506 1164 110512 1176
rect 110564 1164 110570 1216
rect 111978 1204 111984 1216
rect 111939 1176 111984 1204
rect 111978 1164 111984 1176
rect 112036 1164 112042 1216
rect 112073 1207 112131 1213
rect 112073 1173 112085 1207
rect 112119 1204 112131 1207
rect 116581 1207 116639 1213
rect 116581 1204 116593 1207
rect 112119 1176 116593 1204
rect 112119 1173 112131 1176
rect 112073 1167 112131 1173
rect 116581 1173 116593 1176
rect 116627 1173 116639 1207
rect 116581 1167 116639 1173
rect 116857 1207 116915 1213
rect 116857 1173 116869 1207
rect 116903 1204 116915 1207
rect 119249 1207 119307 1213
rect 119249 1204 119261 1207
rect 116903 1176 119261 1204
rect 116903 1173 116915 1176
rect 116857 1167 116915 1173
rect 119249 1173 119261 1176
rect 119295 1173 119307 1207
rect 119249 1167 119307 1173
rect 119338 1164 119344 1216
rect 119396 1204 119402 1216
rect 119433 1207 119491 1213
rect 119433 1204 119445 1207
rect 119396 1176 119445 1204
rect 119396 1164 119402 1176
rect 119433 1173 119445 1176
rect 119479 1173 119491 1207
rect 119433 1167 119491 1173
rect 119525 1207 119583 1213
rect 119525 1173 119537 1207
rect 119571 1204 119583 1207
rect 139305 1207 139363 1213
rect 139305 1204 139317 1207
rect 119571 1176 139317 1204
rect 119571 1173 119583 1176
rect 119525 1167 119583 1173
rect 139305 1173 139317 1176
rect 139351 1173 139363 1207
rect 139305 1167 139363 1173
rect 139397 1207 139455 1213
rect 139397 1173 139409 1207
rect 139443 1204 139455 1207
rect 139486 1204 139492 1216
rect 139443 1176 139492 1204
rect 139443 1173 139455 1176
rect 139397 1167 139455 1173
rect 139486 1164 139492 1176
rect 139544 1164 139550 1216
rect 139581 1207 139639 1213
rect 139581 1173 139593 1207
rect 139627 1204 139639 1207
rect 144822 1204 144828 1216
rect 139627 1176 144828 1204
rect 139627 1173 139639 1176
rect 139581 1167 139639 1173
rect 144822 1164 144828 1176
rect 144880 1164 144886 1216
rect 144914 1164 144920 1216
rect 144972 1204 144978 1216
rect 149517 1207 149575 1213
rect 149517 1204 149529 1207
rect 144972 1176 149529 1204
rect 144972 1164 144978 1176
rect 149517 1173 149529 1176
rect 149563 1173 149575 1207
rect 149790 1204 149796 1216
rect 149517 1167 149575 1173
rect 149624 1176 149796 1204
rect 83182 1136 83188 1148
rect 82924 1108 83188 1136
rect 82725 1099 82783 1105
rect 83182 1096 83188 1108
rect 83240 1096 83246 1148
rect 83277 1139 83335 1145
rect 83277 1105 83289 1139
rect 83323 1136 83335 1139
rect 83366 1136 83372 1148
rect 83323 1108 83372 1136
rect 83323 1105 83335 1108
rect 83277 1099 83335 1105
rect 83366 1096 83372 1108
rect 83424 1096 83430 1148
rect 83550 1096 83556 1148
rect 83608 1136 83614 1148
rect 92293 1139 92351 1145
rect 83608 1108 92152 1136
rect 83608 1096 83614 1108
rect 5307 1040 5396 1068
rect 5307 1037 5319 1040
rect 5261 1031 5319 1037
rect 5534 1028 5540 1080
rect 5592 1068 5598 1080
rect 62298 1068 62304 1080
rect 5592 1040 62304 1068
rect 5592 1028 5598 1040
rect 62298 1028 62304 1040
rect 62356 1028 62362 1080
rect 62390 1028 62396 1080
rect 62448 1068 62454 1080
rect 66622 1068 66628 1080
rect 62448 1040 66628 1068
rect 62448 1028 62454 1040
rect 66622 1028 66628 1040
rect 66680 1028 66686 1080
rect 66714 1028 66720 1080
rect 66772 1068 66778 1080
rect 68830 1068 68836 1080
rect 66772 1040 68836 1068
rect 66772 1028 66778 1040
rect 68830 1028 68836 1040
rect 68888 1028 68894 1080
rect 68925 1071 68983 1077
rect 68925 1037 68937 1071
rect 68971 1068 68983 1071
rect 72973 1071 73031 1077
rect 72973 1068 72985 1071
rect 68971 1040 72985 1068
rect 68971 1037 68983 1040
rect 68925 1031 68983 1037
rect 72973 1037 72985 1040
rect 73019 1037 73031 1071
rect 72973 1031 73031 1037
rect 73065 1071 73123 1077
rect 73065 1037 73077 1071
rect 73111 1068 73123 1071
rect 73111 1040 82952 1068
rect 73111 1037 73123 1040
rect 73065 1031 73123 1037
rect 3234 960 3240 1012
rect 3292 1000 3298 1012
rect 25869 1003 25927 1009
rect 25869 1000 25881 1003
rect 3292 972 25881 1000
rect 3292 960 3298 972
rect 25869 969 25881 972
rect 25915 969 25927 1003
rect 25869 963 25927 969
rect 25961 1003 26019 1009
rect 25961 969 25973 1003
rect 26007 1000 26019 1003
rect 35345 1003 35403 1009
rect 35345 1000 35357 1003
rect 26007 972 35357 1000
rect 26007 969 26019 972
rect 25961 963 26019 969
rect 35345 969 35357 972
rect 35391 969 35403 1003
rect 35345 963 35403 969
rect 38289 1003 38347 1009
rect 38289 969 38301 1003
rect 38335 1000 38347 1003
rect 82817 1003 82875 1009
rect 82817 1000 82829 1003
rect 38335 972 82829 1000
rect 38335 969 38347 972
rect 38289 963 38347 969
rect 82817 969 82829 972
rect 82863 969 82875 1003
rect 82924 1000 82952 1040
rect 82998 1028 83004 1080
rect 83056 1068 83062 1080
rect 91833 1071 91891 1077
rect 91833 1068 91845 1071
rect 83056 1040 91845 1068
rect 83056 1028 83062 1040
rect 91833 1037 91845 1040
rect 91879 1037 91891 1071
rect 91833 1031 91891 1037
rect 91925 1071 91983 1077
rect 91925 1037 91937 1071
rect 91971 1068 91983 1071
rect 92014 1068 92020 1080
rect 91971 1040 92020 1068
rect 91971 1037 91983 1040
rect 91925 1031 91983 1037
rect 92014 1028 92020 1040
rect 92072 1028 92078 1080
rect 92124 1068 92152 1108
rect 92293 1105 92305 1139
rect 92339 1136 92351 1139
rect 92661 1139 92719 1145
rect 92661 1136 92673 1139
rect 92339 1108 92673 1136
rect 92339 1105 92351 1108
rect 92293 1099 92351 1105
rect 92661 1105 92673 1108
rect 92707 1105 92719 1139
rect 92661 1099 92719 1105
rect 93213 1139 93271 1145
rect 93213 1105 93225 1139
rect 93259 1136 93271 1139
rect 103517 1139 103575 1145
rect 103517 1136 103529 1139
rect 93259 1108 103529 1136
rect 93259 1105 93271 1108
rect 93213 1099 93271 1105
rect 103517 1105 103529 1108
rect 103563 1105 103575 1139
rect 103517 1099 103575 1105
rect 103701 1139 103759 1145
rect 103701 1105 103713 1139
rect 103747 1136 103759 1139
rect 103974 1136 103980 1148
rect 103747 1108 103980 1136
rect 103747 1105 103759 1108
rect 103701 1099 103759 1105
rect 103974 1096 103980 1108
rect 104032 1096 104038 1148
rect 104069 1139 104127 1145
rect 104069 1105 104081 1139
rect 104115 1136 104127 1139
rect 104802 1136 104808 1148
rect 104115 1108 104808 1136
rect 104115 1105 104127 1108
rect 104069 1099 104127 1105
rect 104802 1096 104808 1108
rect 104860 1096 104866 1148
rect 104897 1139 104955 1145
rect 104897 1105 104909 1139
rect 104943 1136 104955 1139
rect 105814 1136 105820 1148
rect 104943 1108 105820 1136
rect 104943 1105 104955 1108
rect 104897 1099 104955 1105
rect 105814 1096 105820 1108
rect 105872 1096 105878 1148
rect 105909 1139 105967 1145
rect 105909 1105 105921 1139
rect 105955 1136 105967 1139
rect 115845 1139 115903 1145
rect 115845 1136 115857 1139
rect 105955 1108 115857 1136
rect 105955 1105 105967 1108
rect 105909 1099 105967 1105
rect 115845 1105 115857 1108
rect 115891 1105 115903 1139
rect 115845 1099 115903 1105
rect 115934 1096 115940 1148
rect 115992 1136 115998 1148
rect 122834 1136 122840 1148
rect 115992 1108 122840 1136
rect 115992 1096 115998 1108
rect 122834 1096 122840 1108
rect 122892 1096 122898 1148
rect 123202 1096 123208 1148
rect 123260 1136 123266 1148
rect 134794 1136 134800 1148
rect 123260 1108 134800 1136
rect 123260 1096 123266 1108
rect 134794 1096 134800 1108
rect 134852 1096 134858 1148
rect 134889 1139 134947 1145
rect 134889 1105 134901 1139
rect 134935 1136 134947 1139
rect 140222 1136 140228 1148
rect 134935 1108 140228 1136
rect 134935 1105 134947 1108
rect 134889 1099 134947 1105
rect 140222 1096 140228 1108
rect 140280 1096 140286 1148
rect 140685 1139 140743 1145
rect 140685 1105 140697 1139
rect 140731 1136 140743 1139
rect 142249 1139 142307 1145
rect 142249 1136 142261 1139
rect 140731 1108 142261 1136
rect 140731 1105 140743 1108
rect 140685 1099 140743 1105
rect 142249 1105 142261 1108
rect 142295 1105 142307 1139
rect 142249 1099 142307 1105
rect 142338 1096 142344 1148
rect 142396 1136 142402 1148
rect 147582 1136 147588 1148
rect 142396 1108 147588 1136
rect 142396 1096 142402 1108
rect 147582 1096 147588 1108
rect 147640 1096 147646 1148
rect 147953 1139 148011 1145
rect 147953 1136 147965 1139
rect 147692 1108 147965 1136
rect 92750 1068 92756 1080
rect 92124 1040 92756 1068
rect 92750 1028 92756 1040
rect 92808 1028 92814 1080
rect 92842 1028 92848 1080
rect 92900 1068 92906 1080
rect 100849 1071 100907 1077
rect 100849 1068 100861 1071
rect 92900 1040 100861 1068
rect 92900 1028 92906 1040
rect 100849 1037 100861 1040
rect 100895 1037 100907 1071
rect 100849 1031 100907 1037
rect 100941 1071 100999 1077
rect 100941 1037 100953 1071
rect 100987 1068 100999 1071
rect 111797 1071 111855 1077
rect 111797 1068 111809 1071
rect 100987 1040 111809 1068
rect 100987 1037 100999 1040
rect 100941 1031 100999 1037
rect 111797 1037 111809 1040
rect 111843 1037 111855 1071
rect 111797 1031 111855 1037
rect 112073 1071 112131 1077
rect 112073 1037 112085 1071
rect 112119 1068 112131 1071
rect 116397 1071 116455 1077
rect 116397 1068 116409 1071
rect 112119 1040 116409 1068
rect 112119 1037 112131 1040
rect 112073 1031 112131 1037
rect 116397 1037 116409 1040
rect 116443 1037 116455 1071
rect 116397 1031 116455 1037
rect 116489 1071 116547 1077
rect 116489 1037 116501 1071
rect 116535 1068 116547 1071
rect 121178 1068 121184 1080
rect 116535 1040 121184 1068
rect 116535 1037 116547 1040
rect 116489 1031 116547 1037
rect 121178 1028 121184 1040
rect 121236 1028 121242 1080
rect 121273 1071 121331 1077
rect 121273 1037 121285 1071
rect 121319 1068 121331 1071
rect 123021 1071 123079 1077
rect 123021 1068 123033 1071
rect 121319 1040 123033 1068
rect 121319 1037 121331 1040
rect 121273 1031 121331 1037
rect 123021 1037 123033 1040
rect 123067 1037 123079 1071
rect 140041 1071 140099 1077
rect 140041 1068 140053 1071
rect 123021 1031 123079 1037
rect 124232 1040 140053 1068
rect 83461 1003 83519 1009
rect 83461 1000 83473 1003
rect 82924 972 83473 1000
rect 82817 963 82875 969
rect 83461 969 83473 972
rect 83507 969 83519 1003
rect 83461 963 83519 969
rect 83553 1003 83611 1009
rect 83553 969 83565 1003
rect 83599 1000 83611 1003
rect 116121 1003 116179 1009
rect 116121 1000 116133 1003
rect 83599 972 116133 1000
rect 83599 969 83611 972
rect 83553 963 83611 969
rect 116121 969 116133 972
rect 116167 969 116179 1003
rect 116121 963 116179 969
rect 116210 960 116216 1012
rect 116268 1000 116274 1012
rect 120074 1000 120080 1012
rect 116268 972 120080 1000
rect 116268 960 116274 972
rect 120074 960 120080 972
rect 120132 960 120138 1012
rect 120169 1003 120227 1009
rect 120169 969 120181 1003
rect 120215 1000 120227 1003
rect 121365 1003 121423 1009
rect 121365 1000 121377 1003
rect 120215 972 121377 1000
rect 120215 969 120227 972
rect 120169 963 120227 969
rect 121365 969 121377 972
rect 121411 969 121423 1003
rect 121365 963 121423 969
rect 121457 1003 121515 1009
rect 121457 969 121469 1003
rect 121503 1000 121515 1003
rect 121825 1003 121883 1009
rect 121825 1000 121837 1003
rect 121503 972 121837 1000
rect 121503 969 121515 972
rect 121457 963 121515 969
rect 121825 969 121837 972
rect 121871 969 121883 1003
rect 121825 963 121883 969
rect 121917 1003 121975 1009
rect 121917 969 121929 1003
rect 121963 1000 121975 1003
rect 122377 1003 122435 1009
rect 122377 1000 122389 1003
rect 121963 972 122389 1000
rect 121963 969 121975 972
rect 121917 963 121975 969
rect 122377 969 122389 972
rect 122423 969 122435 1003
rect 122377 963 122435 969
rect 122466 960 122472 1012
rect 122524 1000 122530 1012
rect 123938 1000 123944 1012
rect 122524 972 123944 1000
rect 122524 960 122530 972
rect 123938 960 123944 972
rect 123996 960 124002 1012
rect 124033 1003 124091 1009
rect 124033 969 124045 1003
rect 124079 1000 124091 1003
rect 124232 1000 124260 1040
rect 140041 1037 140053 1040
rect 140087 1037 140099 1071
rect 140041 1031 140099 1037
rect 140593 1071 140651 1077
rect 140593 1037 140605 1071
rect 140639 1068 140651 1071
rect 147401 1071 147459 1077
rect 147401 1068 147413 1071
rect 140639 1040 147413 1068
rect 140639 1037 140651 1040
rect 140593 1031 140651 1037
rect 147401 1037 147413 1040
rect 147447 1037 147459 1071
rect 147401 1031 147459 1037
rect 147490 1028 147496 1080
rect 147548 1068 147554 1080
rect 147692 1068 147720 1108
rect 147953 1105 147965 1108
rect 147999 1105 148011 1139
rect 149624 1136 149652 1176
rect 149790 1164 149796 1176
rect 149848 1164 149854 1216
rect 149885 1207 149943 1213
rect 149885 1173 149897 1207
rect 149931 1204 149943 1207
rect 152458 1204 152464 1216
rect 149931 1176 152464 1204
rect 149931 1173 149943 1176
rect 149885 1167 149943 1173
rect 152458 1164 152464 1176
rect 152516 1164 152522 1216
rect 147953 1099 148011 1105
rect 148060 1108 149652 1136
rect 149701 1139 149759 1145
rect 147548 1040 147720 1068
rect 147769 1071 147827 1077
rect 147548 1028 147554 1040
rect 147769 1037 147781 1071
rect 147815 1068 147827 1071
rect 148060 1068 148088 1108
rect 149701 1105 149713 1139
rect 149747 1136 149759 1139
rect 149974 1136 149980 1148
rect 149747 1108 149980 1136
rect 149747 1105 149759 1108
rect 149701 1099 149759 1105
rect 149974 1096 149980 1108
rect 150032 1096 150038 1148
rect 150069 1139 150127 1145
rect 150069 1105 150081 1139
rect 150115 1136 150127 1139
rect 151449 1139 151507 1145
rect 151449 1136 151461 1139
rect 150115 1108 151461 1136
rect 150115 1105 150127 1108
rect 150069 1099 150127 1105
rect 151449 1105 151461 1108
rect 151495 1105 151507 1139
rect 151449 1099 151507 1105
rect 151541 1139 151599 1145
rect 151541 1105 151553 1139
rect 151587 1136 151599 1139
rect 152829 1139 152887 1145
rect 152829 1136 152841 1139
rect 151587 1108 152841 1136
rect 151587 1105 151599 1108
rect 151541 1099 151599 1105
rect 152829 1105 152841 1108
rect 152875 1105 152887 1139
rect 152936 1136 152964 1244
rect 153013 1241 153025 1275
rect 153059 1272 153071 1275
rect 153289 1275 153347 1281
rect 153289 1272 153301 1275
rect 153059 1244 153301 1272
rect 153059 1241 153071 1244
rect 153013 1235 153071 1241
rect 153289 1241 153301 1244
rect 153335 1241 153347 1275
rect 153289 1235 153347 1241
rect 153565 1275 153623 1281
rect 153565 1241 153577 1275
rect 153611 1272 153623 1275
rect 154577 1275 154635 1281
rect 154577 1272 154589 1275
rect 153611 1244 154589 1272
rect 153611 1241 153623 1244
rect 153565 1235 153623 1241
rect 154577 1241 154589 1244
rect 154623 1241 154635 1275
rect 154577 1235 154635 1241
rect 155037 1275 155095 1281
rect 155037 1241 155049 1275
rect 155083 1272 155095 1275
rect 156414 1272 156420 1284
rect 155083 1244 156420 1272
rect 155083 1241 155095 1244
rect 155037 1235 155095 1241
rect 156414 1232 156420 1244
rect 156472 1232 156478 1284
rect 156509 1275 156567 1281
rect 156509 1241 156521 1275
rect 156555 1272 156567 1275
rect 157337 1275 157395 1281
rect 157337 1272 157349 1275
rect 156555 1244 157349 1272
rect 156555 1241 156567 1244
rect 156509 1235 156567 1241
rect 157337 1241 157349 1244
rect 157383 1241 157395 1275
rect 157337 1235 157395 1241
rect 157426 1232 157432 1284
rect 157484 1272 157490 1284
rect 158162 1272 158168 1284
rect 157484 1244 158168 1272
rect 157484 1232 157490 1244
rect 158162 1232 158168 1244
rect 158220 1232 158226 1284
rect 158257 1275 158315 1281
rect 158257 1241 158269 1275
rect 158303 1272 158315 1275
rect 158622 1272 158628 1284
rect 158303 1244 158628 1272
rect 158303 1241 158315 1244
rect 158257 1235 158315 1241
rect 158622 1232 158628 1244
rect 158680 1232 158686 1284
rect 158717 1275 158775 1281
rect 158717 1241 158729 1275
rect 158763 1272 158775 1275
rect 158806 1272 158812 1284
rect 158763 1244 158812 1272
rect 158763 1241 158775 1244
rect 158717 1235 158775 1241
rect 158806 1232 158812 1244
rect 158864 1232 158870 1284
rect 158993 1275 159051 1281
rect 158993 1241 159005 1275
rect 159039 1272 159051 1275
rect 159450 1272 159456 1284
rect 159039 1244 159456 1272
rect 159039 1241 159051 1244
rect 158993 1235 159051 1241
rect 159450 1232 159456 1244
rect 159508 1232 159514 1284
rect 159545 1275 159603 1281
rect 159545 1241 159557 1275
rect 159591 1272 159603 1275
rect 161477 1275 161535 1281
rect 161477 1272 161489 1275
rect 159591 1244 161489 1272
rect 159591 1241 159603 1244
rect 159545 1235 159603 1241
rect 161477 1241 161489 1244
rect 161523 1241 161535 1275
rect 161477 1235 161535 1241
rect 161753 1275 161811 1281
rect 161753 1241 161765 1275
rect 161799 1272 161811 1275
rect 162302 1272 162308 1284
rect 161799 1244 162308 1272
rect 161799 1241 161811 1244
rect 161753 1235 161811 1241
rect 162302 1232 162308 1244
rect 162360 1232 162366 1284
rect 162397 1275 162455 1281
rect 162397 1241 162409 1275
rect 162443 1272 162455 1275
rect 163593 1275 163651 1281
rect 163593 1272 163605 1275
rect 162443 1244 163605 1272
rect 162443 1241 162455 1244
rect 162397 1235 162455 1241
rect 163593 1241 163605 1244
rect 163639 1241 163651 1275
rect 163593 1235 163651 1241
rect 163682 1232 163688 1284
rect 163740 1272 163746 1284
rect 169938 1272 169944 1284
rect 163740 1244 169944 1272
rect 163740 1232 163746 1244
rect 169938 1232 169944 1244
rect 169996 1232 170002 1284
rect 170033 1275 170091 1281
rect 170033 1241 170045 1275
rect 170079 1272 170091 1275
rect 175829 1275 175887 1281
rect 175829 1272 175841 1275
rect 170079 1244 175841 1272
rect 170079 1241 170091 1244
rect 170033 1235 170091 1241
rect 175829 1241 175841 1244
rect 175875 1241 175887 1275
rect 175829 1235 175887 1241
rect 176010 1232 176016 1284
rect 176068 1272 176074 1284
rect 176933 1275 176991 1281
rect 176933 1272 176945 1275
rect 176068 1244 176945 1272
rect 176068 1232 176074 1244
rect 176933 1241 176945 1244
rect 176979 1241 176991 1275
rect 176933 1235 176991 1241
rect 177666 1232 177672 1284
rect 177724 1272 177730 1284
rect 177853 1275 177911 1281
rect 177724 1244 177769 1272
rect 177724 1232 177730 1244
rect 177853 1241 177865 1275
rect 177899 1272 177911 1275
rect 178034 1272 178040 1284
rect 177899 1244 178040 1272
rect 177899 1241 177911 1244
rect 177853 1235 177911 1241
rect 178034 1232 178040 1244
rect 178092 1232 178098 1284
rect 178126 1232 178132 1284
rect 178184 1272 178190 1284
rect 189721 1275 189779 1281
rect 189721 1272 189733 1275
rect 178184 1244 189733 1272
rect 178184 1232 178190 1244
rect 189721 1241 189733 1244
rect 189767 1241 189779 1275
rect 189920 1272 189948 1312
rect 190178 1300 190184 1352
rect 190236 1340 190242 1352
rect 190641 1343 190699 1349
rect 190641 1340 190653 1343
rect 190236 1312 190653 1340
rect 190236 1300 190242 1312
rect 190641 1309 190653 1312
rect 190687 1309 190699 1343
rect 190641 1303 190699 1309
rect 190822 1300 190828 1352
rect 190880 1340 190886 1352
rect 191009 1343 191067 1349
rect 191009 1340 191021 1343
rect 190880 1312 191021 1340
rect 190880 1300 190886 1312
rect 191009 1309 191021 1312
rect 191055 1309 191067 1343
rect 191009 1303 191067 1309
rect 191101 1343 191159 1349
rect 191101 1309 191113 1343
rect 191147 1340 191159 1343
rect 191377 1343 191435 1349
rect 191377 1340 191389 1343
rect 191147 1312 191389 1340
rect 191147 1309 191159 1312
rect 191101 1303 191159 1309
rect 191377 1309 191389 1312
rect 191423 1309 191435 1343
rect 191377 1303 191435 1309
rect 191466 1300 191472 1352
rect 191524 1340 191530 1352
rect 195238 1340 195244 1352
rect 191524 1312 195244 1340
rect 191524 1300 191530 1312
rect 195238 1300 195244 1312
rect 195296 1300 195302 1352
rect 195333 1343 195391 1349
rect 195333 1309 195345 1343
rect 195379 1340 195391 1343
rect 196621 1343 196679 1349
rect 196621 1340 196633 1343
rect 195379 1312 196633 1340
rect 195379 1309 195391 1312
rect 195333 1303 195391 1309
rect 196621 1309 196633 1312
rect 196667 1309 196679 1343
rect 196621 1303 196679 1309
rect 196805 1343 196863 1349
rect 196805 1309 196817 1343
rect 196851 1340 196863 1343
rect 197173 1343 197231 1349
rect 197173 1340 197185 1343
rect 196851 1312 197185 1340
rect 196851 1309 196863 1312
rect 196805 1303 196863 1309
rect 197173 1309 197185 1312
rect 197219 1309 197231 1343
rect 197173 1303 197231 1309
rect 197262 1300 197268 1352
rect 197320 1340 197326 1352
rect 198458 1340 198464 1352
rect 197320 1312 198464 1340
rect 197320 1300 197326 1312
rect 198458 1300 198464 1312
rect 198516 1300 198522 1352
rect 198553 1343 198611 1349
rect 198553 1309 198565 1343
rect 198599 1340 198611 1343
rect 199105 1343 199163 1349
rect 199105 1340 199117 1343
rect 198599 1312 199117 1340
rect 198599 1309 198611 1312
rect 198553 1303 198611 1309
rect 199105 1309 199117 1312
rect 199151 1309 199163 1343
rect 199105 1303 199163 1309
rect 199194 1300 199200 1352
rect 199252 1340 199258 1352
rect 200393 1343 200451 1349
rect 199252 1312 199297 1340
rect 199252 1300 199258 1312
rect 200393 1309 200405 1343
rect 200439 1340 200451 1343
rect 202877 1343 202935 1349
rect 202877 1340 202889 1343
rect 200439 1312 202889 1340
rect 200439 1309 200451 1312
rect 200393 1303 200451 1309
rect 202877 1309 202889 1312
rect 202923 1309 202935 1343
rect 202877 1303 202935 1309
rect 202966 1300 202972 1352
rect 203024 1340 203030 1352
rect 211154 1340 211160 1352
rect 203024 1312 211160 1340
rect 203024 1300 203030 1312
rect 211154 1300 211160 1312
rect 211212 1300 211218 1352
rect 211249 1343 211307 1349
rect 211249 1309 211261 1343
rect 211295 1340 211307 1343
rect 214193 1343 214251 1349
rect 214193 1340 214205 1343
rect 211295 1312 214205 1340
rect 211295 1309 211307 1312
rect 211249 1303 211307 1309
rect 214193 1309 214205 1312
rect 214239 1309 214251 1343
rect 214193 1303 214251 1309
rect 214285 1343 214343 1349
rect 214285 1309 214297 1343
rect 214331 1340 214343 1343
rect 214374 1340 214380 1352
rect 214331 1312 214380 1340
rect 214331 1309 214343 1312
rect 214285 1303 214343 1309
rect 214374 1300 214380 1312
rect 214432 1300 214438 1352
rect 214469 1343 214527 1349
rect 214469 1309 214481 1343
rect 214515 1340 214527 1343
rect 214742 1340 214748 1352
rect 214515 1312 214748 1340
rect 214515 1309 214527 1312
rect 214469 1303 214527 1309
rect 214742 1300 214748 1312
rect 214800 1300 214806 1352
rect 214837 1343 214895 1349
rect 214837 1309 214849 1343
rect 214883 1340 214895 1343
rect 218532 1340 218560 1380
rect 218701 1377 218713 1380
rect 218747 1377 218759 1411
rect 218701 1371 218759 1377
rect 218790 1368 218796 1420
rect 218848 1408 218854 1420
rect 224497 1411 224555 1417
rect 224497 1408 224509 1411
rect 218848 1380 224509 1408
rect 218848 1368 218854 1380
rect 224497 1377 224509 1380
rect 224543 1377 224555 1411
rect 224604 1408 224632 1516
rect 231949 1479 232007 1485
rect 231949 1476 231961 1479
rect 224972 1448 231961 1476
rect 224972 1408 225000 1448
rect 231949 1445 231961 1448
rect 231995 1445 232007 1479
rect 232056 1476 232084 1516
rect 232516 1516 260420 1544
rect 260484 1516 260696 1544
rect 260760 1516 285772 1544
rect 232516 1476 232544 1516
rect 232056 1448 232544 1476
rect 231949 1439 232007 1445
rect 232590 1436 232596 1488
rect 232648 1476 232654 1488
rect 233142 1476 233148 1488
rect 232648 1448 233148 1476
rect 232648 1436 232654 1448
rect 233142 1436 233148 1448
rect 233200 1436 233206 1488
rect 233237 1479 233295 1485
rect 233237 1445 233249 1479
rect 233283 1476 233295 1479
rect 236549 1479 236607 1485
rect 236549 1476 236561 1479
rect 233283 1448 236561 1476
rect 233283 1445 233295 1448
rect 233237 1439 233295 1445
rect 236549 1445 236561 1448
rect 236595 1445 236607 1479
rect 236549 1439 236607 1445
rect 236641 1479 236699 1485
rect 236641 1445 236653 1479
rect 236687 1476 236699 1479
rect 238938 1476 238944 1488
rect 236687 1448 238944 1476
rect 236687 1445 236699 1448
rect 236641 1439 236699 1445
rect 238938 1436 238944 1448
rect 238996 1436 239002 1488
rect 239033 1479 239091 1485
rect 239033 1445 239045 1479
rect 239079 1476 239091 1479
rect 241330 1476 241336 1488
rect 239079 1448 241336 1476
rect 239079 1445 239091 1448
rect 239033 1439 239091 1445
rect 241330 1436 241336 1448
rect 241388 1436 241394 1488
rect 241425 1479 241483 1485
rect 241425 1445 241437 1479
rect 241471 1476 241483 1479
rect 249797 1479 249855 1485
rect 249797 1476 249809 1479
rect 241471 1448 249809 1476
rect 241471 1445 241483 1448
rect 241425 1439 241483 1445
rect 249797 1445 249809 1448
rect 249843 1445 249855 1479
rect 249797 1439 249855 1445
rect 249886 1436 249892 1488
rect 249944 1476 249950 1488
rect 250714 1476 250720 1488
rect 249944 1448 250720 1476
rect 249944 1436 249950 1448
rect 250714 1436 250720 1448
rect 250772 1436 250778 1488
rect 250809 1479 250867 1485
rect 250809 1445 250821 1479
rect 250855 1476 250867 1479
rect 260484 1476 260512 1516
rect 250855 1448 260512 1476
rect 260561 1479 260619 1485
rect 250855 1445 250867 1448
rect 250809 1439 250867 1445
rect 260561 1445 260573 1479
rect 260607 1445 260619 1479
rect 260668 1476 260696 1516
rect 285766 1504 285772 1516
rect 285824 1504 285830 1556
rect 285861 1547 285919 1553
rect 285861 1513 285873 1547
rect 285907 1544 285919 1547
rect 289633 1547 289691 1553
rect 289633 1544 289645 1547
rect 285907 1516 289645 1544
rect 285907 1513 285919 1516
rect 285861 1507 285919 1513
rect 289633 1513 289645 1516
rect 289679 1513 289691 1547
rect 289633 1507 289691 1513
rect 289722 1504 289728 1556
rect 289780 1544 289786 1556
rect 298465 1547 298523 1553
rect 298465 1544 298477 1547
rect 289780 1516 298477 1544
rect 289780 1504 289786 1516
rect 298465 1513 298477 1516
rect 298511 1513 298523 1547
rect 298465 1507 298523 1513
rect 298554 1504 298560 1556
rect 298612 1544 298618 1556
rect 298649 1547 298707 1553
rect 298649 1544 298661 1547
rect 298612 1516 298661 1544
rect 298612 1504 298618 1516
rect 298649 1513 298661 1516
rect 298695 1513 298707 1547
rect 298756 1544 298784 1584
rect 298833 1581 298845 1615
rect 298879 1612 298891 1615
rect 394878 1612 394884 1624
rect 298879 1584 394884 1612
rect 298879 1581 298891 1584
rect 298833 1575 298891 1581
rect 394878 1572 394884 1584
rect 394936 1572 394942 1624
rect 395430 1572 395436 1624
rect 395488 1612 395494 1624
rect 398650 1612 398656 1624
rect 395488 1584 398656 1612
rect 395488 1572 395494 1584
rect 398650 1572 398656 1584
rect 398708 1572 398714 1624
rect 399570 1572 399576 1624
rect 399628 1612 399634 1624
rect 403710 1612 403716 1624
rect 399628 1584 403716 1612
rect 399628 1572 399634 1584
rect 403710 1572 403716 1584
rect 403768 1572 403774 1624
rect 412177 1615 412235 1621
rect 412177 1581 412189 1615
rect 412223 1612 412235 1615
rect 432966 1612 432972 1624
rect 412223 1584 432972 1612
rect 412223 1581 412235 1584
rect 412177 1575 412235 1581
rect 432966 1572 432972 1584
rect 433024 1572 433030 1624
rect 443454 1572 443460 1624
rect 443512 1612 443518 1624
rect 453206 1612 453212 1624
rect 443512 1584 453212 1612
rect 443512 1572 443518 1584
rect 453206 1572 453212 1584
rect 453264 1572 453270 1624
rect 515582 1572 515588 1624
rect 515640 1612 515646 1624
rect 528830 1612 528836 1624
rect 515640 1584 528836 1612
rect 515640 1572 515646 1584
rect 528830 1572 528836 1584
rect 528888 1572 528894 1624
rect 549254 1572 549260 1624
rect 549312 1612 549318 1624
rect 556157 1615 556215 1621
rect 556157 1612 556169 1615
rect 549312 1584 556169 1612
rect 549312 1572 549318 1584
rect 556157 1581 556169 1584
rect 556203 1581 556215 1615
rect 556157 1575 556215 1581
rect 568298 1572 568304 1624
rect 568356 1612 568362 1624
rect 568666 1612 568672 1624
rect 568356 1584 568672 1612
rect 568356 1572 568362 1584
rect 568666 1572 568672 1584
rect 568724 1572 568730 1624
rect 304169 1547 304227 1553
rect 304169 1544 304181 1547
rect 298756 1516 304181 1544
rect 298649 1507 298707 1513
rect 304169 1513 304181 1516
rect 304215 1513 304227 1547
rect 304169 1507 304227 1513
rect 304261 1547 304319 1553
rect 304261 1513 304273 1547
rect 304307 1544 304319 1547
rect 305546 1544 305552 1556
rect 304307 1516 305552 1544
rect 304307 1513 304319 1516
rect 304261 1507 304319 1513
rect 305546 1504 305552 1516
rect 305604 1504 305610 1556
rect 305638 1504 305644 1556
rect 305696 1544 305702 1556
rect 318886 1544 318892 1556
rect 305696 1516 318892 1544
rect 305696 1504 305702 1516
rect 318886 1504 318892 1516
rect 318944 1504 318950 1556
rect 318981 1547 319039 1553
rect 318981 1513 318993 1547
rect 319027 1544 319039 1547
rect 319349 1547 319407 1553
rect 319349 1544 319361 1547
rect 319027 1516 319361 1544
rect 319027 1513 319039 1516
rect 318981 1507 319039 1513
rect 319349 1513 319361 1516
rect 319395 1513 319407 1547
rect 319349 1507 319407 1513
rect 319441 1547 319499 1553
rect 319441 1513 319453 1547
rect 319487 1544 319499 1547
rect 423398 1544 423404 1556
rect 319487 1516 423404 1544
rect 319487 1513 319499 1516
rect 319441 1507 319499 1513
rect 423398 1504 423404 1516
rect 423456 1504 423462 1556
rect 425054 1504 425060 1556
rect 425112 1544 425118 1556
rect 432233 1547 432291 1553
rect 432233 1544 432245 1547
rect 425112 1516 432245 1544
rect 425112 1504 425118 1516
rect 432233 1513 432245 1516
rect 432279 1513 432291 1547
rect 432233 1507 432291 1513
rect 500957 1547 501015 1553
rect 500957 1513 500969 1547
rect 501003 1544 501015 1547
rect 509513 1547 509571 1553
rect 509513 1544 509525 1547
rect 501003 1516 509525 1544
rect 501003 1513 501015 1516
rect 500957 1507 501015 1513
rect 509513 1513 509525 1516
rect 509559 1513 509571 1547
rect 509513 1507 509571 1513
rect 568482 1504 568488 1556
rect 568540 1544 568546 1556
rect 568758 1544 568764 1556
rect 568540 1516 568764 1544
rect 568540 1504 568546 1516
rect 568758 1504 568764 1516
rect 568816 1504 568822 1556
rect 263042 1476 263048 1488
rect 260668 1448 263048 1476
rect 260561 1439 260619 1445
rect 224604 1380 225000 1408
rect 225049 1411 225107 1417
rect 224497 1371 224555 1377
rect 225049 1377 225061 1411
rect 225095 1408 225107 1411
rect 258353 1411 258411 1417
rect 258353 1408 258365 1411
rect 225095 1380 258365 1408
rect 225095 1377 225107 1380
rect 225049 1371 225107 1377
rect 258353 1377 258365 1380
rect 258399 1377 258411 1411
rect 258353 1371 258411 1377
rect 258445 1411 258503 1417
rect 258445 1377 258457 1411
rect 258491 1408 258503 1411
rect 259086 1408 259092 1420
rect 258491 1380 259092 1408
rect 258491 1377 258503 1380
rect 258445 1371 258503 1377
rect 259086 1368 259092 1380
rect 259144 1368 259150 1420
rect 259178 1368 259184 1420
rect 259236 1408 259242 1420
rect 260576 1408 260604 1439
rect 263042 1436 263048 1448
rect 263100 1436 263106 1488
rect 263137 1479 263195 1485
rect 263137 1445 263149 1479
rect 263183 1476 263195 1479
rect 265069 1479 265127 1485
rect 265069 1476 265081 1479
rect 263183 1448 265081 1476
rect 263183 1445 263195 1448
rect 263137 1439 263195 1445
rect 265069 1445 265081 1448
rect 265115 1445 265127 1479
rect 265069 1439 265127 1445
rect 265158 1436 265164 1488
rect 265216 1476 265222 1488
rect 265253 1479 265311 1485
rect 265253 1476 265265 1479
rect 265216 1448 265265 1476
rect 265216 1436 265222 1448
rect 265253 1445 265265 1448
rect 265299 1445 265311 1479
rect 265434 1476 265440 1488
rect 265395 1448 265440 1476
rect 265253 1439 265311 1445
rect 265434 1436 265440 1448
rect 265492 1436 265498 1488
rect 265618 1436 265624 1488
rect 265676 1476 265682 1488
rect 268654 1476 268660 1488
rect 265676 1448 268660 1476
rect 265676 1436 265682 1448
rect 268654 1436 268660 1448
rect 268712 1436 268718 1488
rect 268838 1476 268844 1488
rect 268799 1448 268844 1476
rect 268838 1436 268844 1448
rect 268896 1436 268902 1488
rect 269482 1436 269488 1488
rect 269540 1476 269546 1488
rect 271322 1476 271328 1488
rect 269540 1448 271328 1476
rect 269540 1436 269546 1448
rect 271322 1436 271328 1448
rect 271380 1436 271386 1488
rect 271417 1479 271475 1485
rect 271417 1445 271429 1479
rect 271463 1476 271475 1479
rect 272242 1476 272248 1488
rect 271463 1448 272248 1476
rect 271463 1445 271475 1448
rect 271417 1439 271475 1445
rect 272242 1436 272248 1448
rect 272300 1436 272306 1488
rect 272334 1436 272340 1488
rect 272392 1476 272398 1488
rect 273806 1476 273812 1488
rect 272392 1448 273812 1476
rect 272392 1436 272398 1448
rect 273806 1436 273812 1448
rect 273864 1436 273870 1488
rect 273993 1479 274051 1485
rect 273993 1445 274005 1479
rect 274039 1476 274051 1479
rect 274545 1479 274603 1485
rect 274545 1476 274557 1479
rect 274039 1448 274557 1476
rect 274039 1445 274051 1448
rect 273993 1439 274051 1445
rect 274545 1445 274557 1448
rect 274591 1445 274603 1479
rect 279510 1476 279516 1488
rect 279471 1448 279516 1476
rect 274545 1439 274603 1445
rect 279510 1436 279516 1448
rect 279568 1436 279574 1488
rect 280246 1436 280252 1488
rect 280304 1476 280310 1488
rect 281718 1476 281724 1488
rect 280304 1448 281724 1476
rect 280304 1436 280310 1448
rect 281718 1436 281724 1448
rect 281776 1436 281782 1488
rect 281905 1479 281963 1485
rect 281905 1445 281917 1479
rect 281951 1476 281963 1479
rect 282086 1476 282092 1488
rect 281951 1448 282092 1476
rect 281951 1445 281963 1448
rect 281905 1439 281963 1445
rect 282086 1436 282092 1448
rect 282144 1436 282150 1488
rect 282178 1436 282184 1488
rect 282236 1476 282242 1488
rect 285585 1479 285643 1485
rect 282236 1448 285260 1476
rect 282236 1436 282242 1448
rect 259236 1380 260604 1408
rect 261021 1411 261079 1417
rect 259236 1368 259242 1380
rect 261021 1377 261033 1411
rect 261067 1408 261079 1411
rect 285125 1411 285183 1417
rect 285125 1408 285137 1411
rect 261067 1380 285137 1408
rect 261067 1377 261079 1380
rect 261021 1371 261079 1377
rect 285125 1377 285137 1380
rect 285171 1377 285183 1411
rect 285232 1408 285260 1448
rect 285585 1445 285597 1479
rect 285631 1476 285643 1479
rect 285677 1479 285735 1485
rect 285677 1476 285689 1479
rect 285631 1448 285689 1476
rect 285631 1445 285643 1448
rect 285585 1439 285643 1445
rect 285677 1445 285689 1448
rect 285723 1445 285735 1479
rect 285677 1439 285735 1445
rect 285953 1479 286011 1485
rect 285953 1445 285965 1479
rect 285999 1476 286011 1479
rect 289265 1479 289323 1485
rect 289265 1476 289277 1479
rect 285999 1448 289277 1476
rect 285999 1445 286011 1448
rect 285953 1439 286011 1445
rect 289265 1445 289277 1448
rect 289311 1445 289323 1479
rect 289265 1439 289323 1445
rect 289354 1436 289360 1488
rect 289412 1476 289418 1488
rect 289541 1479 289599 1485
rect 289541 1476 289553 1479
rect 289412 1448 289553 1476
rect 289412 1436 289418 1448
rect 289541 1445 289553 1448
rect 289587 1445 289599 1479
rect 289541 1439 289599 1445
rect 290366 1436 290372 1488
rect 290424 1476 290430 1488
rect 293865 1479 293923 1485
rect 293865 1476 293877 1479
rect 290424 1448 293877 1476
rect 290424 1436 290430 1448
rect 293865 1445 293877 1448
rect 293911 1445 293923 1479
rect 293865 1439 293923 1445
rect 293954 1436 293960 1488
rect 294012 1476 294018 1488
rect 294782 1476 294788 1488
rect 294012 1448 294788 1476
rect 294012 1436 294018 1448
rect 294782 1436 294788 1448
rect 294840 1436 294846 1488
rect 295334 1436 295340 1488
rect 295392 1476 295398 1488
rect 296717 1479 296775 1485
rect 296717 1476 296729 1479
rect 295392 1448 296729 1476
rect 295392 1436 295398 1448
rect 296717 1445 296729 1448
rect 296763 1445 296775 1479
rect 296717 1439 296775 1445
rect 296806 1436 296812 1488
rect 296864 1476 296870 1488
rect 299934 1476 299940 1488
rect 296864 1448 299940 1476
rect 296864 1436 296870 1448
rect 299934 1436 299940 1448
rect 299992 1436 299998 1488
rect 300029 1479 300087 1485
rect 300029 1445 300041 1479
rect 300075 1476 300087 1479
rect 309137 1479 309195 1485
rect 309137 1476 309149 1479
rect 300075 1448 309149 1476
rect 300075 1445 300087 1448
rect 300029 1439 300087 1445
rect 309137 1445 309149 1448
rect 309183 1445 309195 1479
rect 309137 1439 309195 1445
rect 309226 1436 309232 1488
rect 309284 1476 309290 1488
rect 309962 1476 309968 1488
rect 309284 1448 309968 1476
rect 309284 1436 309290 1448
rect 309962 1436 309968 1448
rect 310020 1436 310026 1488
rect 318426 1436 318432 1488
rect 318484 1476 318490 1488
rect 318613 1479 318671 1485
rect 318484 1448 318529 1476
rect 318484 1436 318490 1448
rect 318613 1445 318625 1479
rect 318659 1476 318671 1479
rect 320177 1479 320235 1485
rect 320177 1476 320189 1479
rect 318659 1448 320189 1476
rect 318659 1445 318671 1448
rect 318613 1439 318671 1445
rect 320177 1445 320189 1448
rect 320223 1445 320235 1479
rect 320177 1439 320235 1445
rect 320266 1436 320272 1488
rect 320324 1476 320330 1488
rect 329653 1479 329711 1485
rect 329653 1476 329665 1479
rect 320324 1448 329665 1476
rect 320324 1436 320330 1448
rect 329653 1445 329665 1448
rect 329699 1445 329711 1479
rect 329653 1439 329711 1445
rect 329742 1436 329748 1488
rect 329800 1476 329806 1488
rect 356330 1476 356336 1488
rect 329800 1448 356336 1476
rect 329800 1436 329806 1448
rect 356330 1436 356336 1448
rect 356388 1436 356394 1488
rect 356425 1479 356483 1485
rect 356425 1445 356437 1479
rect 356471 1476 356483 1479
rect 385310 1476 385316 1488
rect 356471 1448 385316 1476
rect 356471 1445 356483 1448
rect 356425 1439 356483 1445
rect 385310 1436 385316 1448
rect 385368 1436 385374 1488
rect 386509 1479 386567 1485
rect 386509 1445 386521 1479
rect 386555 1476 386567 1479
rect 391201 1479 391259 1485
rect 391201 1476 391213 1479
rect 386555 1448 391213 1476
rect 386555 1445 386567 1448
rect 386509 1439 386567 1445
rect 391201 1445 391213 1448
rect 391247 1445 391259 1479
rect 391201 1439 391259 1445
rect 393593 1479 393651 1485
rect 393593 1445 393605 1479
rect 393639 1476 393651 1479
rect 451918 1476 451924 1488
rect 393639 1448 451924 1476
rect 393639 1445 393651 1448
rect 393593 1439 393651 1445
rect 451918 1436 451924 1448
rect 451976 1436 451982 1488
rect 459557 1479 459615 1485
rect 459557 1445 459569 1479
rect 459603 1476 459615 1479
rect 473173 1479 473231 1485
rect 473173 1476 473185 1479
rect 459603 1448 473185 1476
rect 459603 1445 459615 1448
rect 459557 1439 459615 1445
rect 473173 1445 473185 1448
rect 473219 1445 473231 1479
rect 473173 1439 473231 1445
rect 555421 1479 555479 1485
rect 555421 1445 555433 1479
rect 555467 1476 555479 1479
rect 560205 1479 560263 1485
rect 560205 1476 560217 1479
rect 555467 1448 560217 1476
rect 555467 1445 555479 1448
rect 555421 1439 555479 1445
rect 560205 1445 560217 1448
rect 560251 1445 560263 1479
rect 560205 1439 560263 1445
rect 285769 1411 285827 1417
rect 285769 1408 285781 1411
rect 285232 1380 285781 1408
rect 285125 1371 285183 1377
rect 285769 1377 285781 1380
rect 285815 1377 285827 1411
rect 285769 1371 285827 1377
rect 287333 1411 287391 1417
rect 287333 1377 287345 1411
rect 287379 1408 287391 1411
rect 309318 1408 309324 1420
rect 287379 1380 309324 1408
rect 287379 1377 287391 1380
rect 287333 1371 287391 1377
rect 309318 1368 309324 1380
rect 309376 1368 309382 1420
rect 309413 1411 309471 1417
rect 309413 1377 309425 1411
rect 309459 1408 309471 1411
rect 309689 1411 309747 1417
rect 309689 1408 309701 1411
rect 309459 1380 309701 1408
rect 309459 1377 309471 1380
rect 309413 1371 309471 1377
rect 309689 1377 309701 1380
rect 309735 1377 309747 1411
rect 309689 1371 309747 1377
rect 309778 1368 309784 1420
rect 309836 1408 309842 1420
rect 319625 1411 319683 1417
rect 319625 1408 319637 1411
rect 309836 1380 319637 1408
rect 309836 1368 309842 1380
rect 319625 1377 319637 1380
rect 319671 1377 319683 1411
rect 319625 1371 319683 1377
rect 319717 1411 319775 1417
rect 319717 1377 319729 1411
rect 319763 1408 319775 1411
rect 356790 1408 356796 1420
rect 319763 1380 356796 1408
rect 319763 1377 319775 1380
rect 319717 1371 319775 1377
rect 356790 1368 356796 1380
rect 356848 1368 356854 1420
rect 358081 1411 358139 1417
rect 358081 1377 358093 1411
rect 358127 1408 358139 1411
rect 367281 1411 367339 1417
rect 367281 1408 367293 1411
rect 358127 1380 367293 1408
rect 358127 1377 358139 1380
rect 358081 1371 358139 1377
rect 367281 1377 367293 1380
rect 367327 1377 367339 1411
rect 367281 1371 367339 1377
rect 368477 1411 368535 1417
rect 368477 1377 368489 1411
rect 368523 1408 368535 1411
rect 374641 1411 374699 1417
rect 374641 1408 374653 1411
rect 368523 1380 374653 1408
rect 368523 1377 368535 1380
rect 368477 1371 368535 1377
rect 374641 1377 374653 1380
rect 374687 1377 374699 1411
rect 374641 1371 374699 1377
rect 374733 1411 374791 1417
rect 374733 1377 374745 1411
rect 374779 1408 374791 1411
rect 388441 1411 388499 1417
rect 388441 1408 388453 1411
rect 374779 1380 388453 1408
rect 374779 1377 374791 1380
rect 374733 1371 374791 1377
rect 388441 1377 388453 1380
rect 388487 1377 388499 1411
rect 388441 1371 388499 1377
rect 391569 1411 391627 1417
rect 391569 1377 391581 1411
rect 391615 1408 391627 1411
rect 565814 1408 565820 1420
rect 391615 1380 565820 1408
rect 391615 1377 391627 1380
rect 391569 1371 391627 1377
rect 565814 1368 565820 1380
rect 565872 1368 565878 1420
rect 214883 1312 218560 1340
rect 218609 1343 218667 1349
rect 214883 1309 214895 1312
rect 214837 1303 214895 1309
rect 218609 1309 218621 1343
rect 218655 1340 218667 1343
rect 224589 1343 224647 1349
rect 218655 1312 224540 1340
rect 218655 1309 218667 1312
rect 218609 1303 218667 1309
rect 190733 1275 190791 1281
rect 190733 1272 190745 1275
rect 189920 1244 190745 1272
rect 189721 1235 189779 1241
rect 190733 1241 190745 1244
rect 190779 1241 190791 1275
rect 190733 1235 190791 1241
rect 191285 1275 191343 1281
rect 191285 1241 191297 1275
rect 191331 1272 191343 1275
rect 224405 1275 224463 1281
rect 224405 1272 224417 1275
rect 191331 1244 224417 1272
rect 191331 1241 191343 1244
rect 191285 1235 191343 1241
rect 224405 1241 224417 1244
rect 224451 1241 224463 1275
rect 224512 1272 224540 1312
rect 224589 1309 224601 1343
rect 224635 1340 224647 1343
rect 225417 1343 225475 1349
rect 225417 1340 225429 1343
rect 224635 1312 225429 1340
rect 224635 1309 224647 1312
rect 224589 1303 224647 1309
rect 225417 1309 225429 1312
rect 225463 1309 225475 1343
rect 225417 1303 225475 1309
rect 225506 1300 225512 1352
rect 225564 1340 225570 1352
rect 228177 1343 228235 1349
rect 228177 1340 228189 1343
rect 225564 1312 228189 1340
rect 225564 1300 225570 1312
rect 228177 1309 228189 1312
rect 228223 1309 228235 1343
rect 228177 1303 228235 1309
rect 228269 1343 228327 1349
rect 228269 1309 228281 1343
rect 228315 1340 228327 1343
rect 390373 1343 390431 1349
rect 390373 1340 390385 1343
rect 228315 1312 390385 1340
rect 228315 1309 228327 1312
rect 228269 1303 228327 1309
rect 390373 1309 390385 1312
rect 390419 1309 390431 1343
rect 390373 1303 390431 1309
rect 390741 1343 390799 1349
rect 390741 1309 390753 1343
rect 390787 1340 390799 1343
rect 560205 1343 560263 1349
rect 390787 1312 549392 1340
rect 390787 1309 390799 1312
rect 390741 1303 390799 1309
rect 224957 1275 225015 1281
rect 224512 1244 224908 1272
rect 224405 1235 224463 1241
rect 153838 1164 153844 1216
rect 153896 1204 153902 1216
rect 161106 1204 161112 1216
rect 153896 1176 160692 1204
rect 153896 1164 153902 1176
rect 153381 1139 153439 1145
rect 153381 1136 153393 1139
rect 152936 1108 153393 1136
rect 152829 1099 152887 1105
rect 153381 1105 153393 1108
rect 153427 1105 153439 1139
rect 153381 1099 153439 1105
rect 153749 1139 153807 1145
rect 153749 1105 153761 1139
rect 153795 1136 153807 1139
rect 154025 1139 154083 1145
rect 154025 1136 154037 1139
rect 153795 1108 154037 1136
rect 153795 1105 153807 1108
rect 153749 1099 153807 1105
rect 154025 1105 154037 1108
rect 154071 1105 154083 1139
rect 154025 1099 154083 1105
rect 154117 1139 154175 1145
rect 154117 1105 154129 1139
rect 154163 1136 154175 1139
rect 154206 1136 154212 1148
rect 154163 1108 154212 1136
rect 154163 1105 154175 1108
rect 154117 1099 154175 1105
rect 154206 1096 154212 1108
rect 154264 1096 154270 1148
rect 154301 1139 154359 1145
rect 154301 1105 154313 1139
rect 154347 1136 154359 1139
rect 157429 1139 157487 1145
rect 157429 1136 157441 1139
rect 154347 1108 157441 1136
rect 154347 1105 154359 1108
rect 154301 1099 154359 1105
rect 157429 1105 157441 1108
rect 157475 1105 157487 1139
rect 157429 1099 157487 1105
rect 157518 1096 157524 1148
rect 157576 1136 157582 1148
rect 158257 1139 158315 1145
rect 158257 1136 158269 1139
rect 157576 1108 158269 1136
rect 157576 1096 157582 1108
rect 158257 1105 158269 1108
rect 158303 1105 158315 1139
rect 158257 1099 158315 1105
rect 158438 1096 158444 1148
rect 158496 1136 158502 1148
rect 160554 1136 160560 1148
rect 158496 1108 160560 1136
rect 158496 1096 158502 1108
rect 160554 1096 160560 1108
rect 160612 1096 160618 1148
rect 160664 1136 160692 1176
rect 160940 1176 161112 1204
rect 160940 1136 160968 1176
rect 161106 1164 161112 1176
rect 161164 1164 161170 1216
rect 161290 1164 161296 1216
rect 161348 1204 161354 1216
rect 178954 1204 178960 1216
rect 161348 1176 178960 1204
rect 161348 1164 161354 1176
rect 178954 1164 178960 1176
rect 179012 1164 179018 1216
rect 179230 1164 179236 1216
rect 179288 1204 179294 1216
rect 180061 1207 180119 1213
rect 180061 1204 180073 1207
rect 179288 1176 180073 1204
rect 179288 1164 179294 1176
rect 180061 1173 180073 1176
rect 180107 1173 180119 1207
rect 180061 1167 180119 1173
rect 180153 1207 180211 1213
rect 180153 1173 180165 1207
rect 180199 1204 180211 1207
rect 180521 1207 180579 1213
rect 180521 1204 180533 1207
rect 180199 1176 180533 1204
rect 180199 1173 180211 1176
rect 180153 1167 180211 1173
rect 180521 1173 180533 1176
rect 180567 1173 180579 1207
rect 180521 1167 180579 1173
rect 180613 1207 180671 1213
rect 180613 1173 180625 1207
rect 180659 1204 180671 1207
rect 183833 1207 183891 1213
rect 183833 1204 183845 1207
rect 180659 1176 183845 1204
rect 180659 1173 180671 1176
rect 180613 1167 180671 1173
rect 183833 1173 183845 1176
rect 183879 1173 183891 1207
rect 183833 1167 183891 1173
rect 183922 1164 183928 1216
rect 183980 1204 183986 1216
rect 189442 1204 189448 1216
rect 183980 1176 189448 1204
rect 183980 1164 183986 1176
rect 189442 1164 189448 1176
rect 189500 1164 189506 1216
rect 190546 1164 190552 1216
rect 190604 1204 190610 1216
rect 190914 1204 190920 1216
rect 190604 1176 190920 1204
rect 190604 1164 190610 1176
rect 190914 1164 190920 1176
rect 190972 1164 190978 1216
rect 191009 1207 191067 1213
rect 191009 1173 191021 1207
rect 191055 1204 191067 1207
rect 224129 1207 224187 1213
rect 224129 1204 224141 1207
rect 191055 1176 224141 1204
rect 191055 1173 191067 1176
rect 191009 1167 191067 1173
rect 224129 1173 224141 1176
rect 224175 1173 224187 1207
rect 224129 1167 224187 1173
rect 224221 1207 224279 1213
rect 224221 1173 224233 1207
rect 224267 1204 224279 1207
rect 224770 1204 224776 1216
rect 224267 1176 224776 1204
rect 224267 1173 224279 1176
rect 224221 1167 224279 1173
rect 224770 1164 224776 1176
rect 224828 1164 224834 1216
rect 224880 1204 224908 1244
rect 224957 1241 224969 1275
rect 225003 1272 225015 1275
rect 232225 1275 232283 1281
rect 232225 1272 232237 1275
rect 225003 1244 232237 1272
rect 225003 1241 225015 1244
rect 224957 1235 225015 1241
rect 232225 1241 232237 1244
rect 232271 1241 232283 1275
rect 232225 1235 232283 1241
rect 232406 1232 232412 1284
rect 232464 1272 232470 1284
rect 233050 1272 233056 1284
rect 232464 1244 233056 1272
rect 232464 1232 232470 1244
rect 233050 1232 233056 1244
rect 233108 1232 233114 1284
rect 233142 1232 233148 1284
rect 233200 1272 233206 1284
rect 238110 1272 238116 1284
rect 233200 1244 238116 1272
rect 233200 1232 233206 1244
rect 238110 1232 238116 1244
rect 238168 1232 238174 1284
rect 238205 1275 238263 1281
rect 238205 1241 238217 1275
rect 238251 1272 238263 1275
rect 238665 1275 238723 1281
rect 238665 1272 238677 1275
rect 238251 1244 238677 1272
rect 238251 1241 238263 1244
rect 238205 1235 238263 1241
rect 238665 1241 238677 1244
rect 238711 1241 238723 1275
rect 238665 1235 238723 1241
rect 239122 1232 239128 1284
rect 239180 1272 239186 1284
rect 239306 1272 239312 1284
rect 239180 1244 239225 1272
rect 239267 1244 239312 1272
rect 239180 1232 239186 1244
rect 239306 1232 239312 1244
rect 239364 1232 239370 1284
rect 239585 1275 239643 1281
rect 239585 1241 239597 1275
rect 239631 1272 239643 1275
rect 239766 1272 239772 1284
rect 239631 1244 239772 1272
rect 239631 1241 239643 1244
rect 239585 1235 239643 1241
rect 239766 1232 239772 1244
rect 239824 1232 239830 1284
rect 239858 1232 239864 1284
rect 239916 1272 239922 1284
rect 241238 1272 241244 1284
rect 239916 1244 241244 1272
rect 239916 1232 239922 1244
rect 241238 1232 241244 1244
rect 241296 1232 241302 1284
rect 241330 1232 241336 1284
rect 241388 1272 241394 1284
rect 251453 1275 251511 1281
rect 251453 1272 251465 1275
rect 241388 1244 251465 1272
rect 241388 1232 241394 1244
rect 251453 1241 251465 1244
rect 251499 1241 251511 1275
rect 251453 1235 251511 1241
rect 251545 1275 251603 1281
rect 251545 1241 251557 1275
rect 251591 1272 251603 1275
rect 253106 1272 253112 1284
rect 251591 1244 253112 1272
rect 251591 1241 251603 1244
rect 251545 1235 251603 1241
rect 253106 1232 253112 1244
rect 253164 1232 253170 1284
rect 253290 1232 253296 1284
rect 253348 1272 253354 1284
rect 254026 1272 254032 1284
rect 253348 1244 254032 1272
rect 253348 1232 253354 1244
rect 254026 1232 254032 1244
rect 254084 1232 254090 1284
rect 254118 1232 254124 1284
rect 254176 1272 254182 1284
rect 256510 1272 256516 1284
rect 254176 1244 256516 1272
rect 254176 1232 254182 1244
rect 256510 1232 256516 1244
rect 256568 1232 256574 1284
rect 256602 1232 256608 1284
rect 256660 1272 256666 1284
rect 260374 1272 260380 1284
rect 256660 1244 260380 1272
rect 256660 1232 256666 1244
rect 260374 1232 260380 1244
rect 260432 1232 260438 1284
rect 260466 1232 260472 1284
rect 260524 1272 260530 1284
rect 270681 1275 270739 1281
rect 270681 1272 270693 1275
rect 260524 1244 270693 1272
rect 260524 1232 260530 1244
rect 270681 1241 270693 1244
rect 270727 1241 270739 1275
rect 270681 1235 270739 1241
rect 271322 1232 271328 1284
rect 271380 1272 271386 1284
rect 272150 1272 272156 1284
rect 271380 1244 272156 1272
rect 271380 1232 271386 1244
rect 272150 1232 272156 1244
rect 272208 1232 272214 1284
rect 272334 1272 272340 1284
rect 272295 1244 272340 1272
rect 272334 1232 272340 1244
rect 272392 1232 272398 1284
rect 273806 1272 273812 1284
rect 273767 1244 273812 1272
rect 273806 1232 273812 1244
rect 273864 1232 273870 1284
rect 273898 1232 273904 1284
rect 273956 1272 273962 1284
rect 279510 1272 279516 1284
rect 273956 1244 279516 1272
rect 273956 1232 273962 1244
rect 279510 1232 279516 1244
rect 279568 1232 279574 1284
rect 279973 1275 280031 1281
rect 279973 1241 279985 1275
rect 280019 1272 280031 1275
rect 290921 1275 290979 1281
rect 290921 1272 290933 1275
rect 280019 1244 290933 1272
rect 280019 1241 280031 1244
rect 279973 1235 280031 1241
rect 290921 1241 290933 1244
rect 290967 1241 290979 1275
rect 290921 1235 290979 1241
rect 291105 1275 291163 1281
rect 291105 1241 291117 1275
rect 291151 1272 291163 1275
rect 296714 1272 296720 1284
rect 291151 1244 296720 1272
rect 291151 1241 291163 1244
rect 291105 1235 291163 1241
rect 296714 1232 296720 1244
rect 296772 1232 296778 1284
rect 296809 1275 296867 1281
rect 296809 1241 296821 1275
rect 296855 1272 296867 1275
rect 297913 1275 297971 1281
rect 297913 1272 297925 1275
rect 296855 1244 297925 1272
rect 296855 1241 296867 1244
rect 296809 1235 296867 1241
rect 297913 1241 297925 1244
rect 297959 1241 297971 1275
rect 309229 1275 309287 1281
rect 309229 1272 309241 1275
rect 297913 1235 297971 1241
rect 298020 1244 309241 1272
rect 228269 1207 228327 1213
rect 228269 1204 228281 1207
rect 224880 1176 228281 1204
rect 228269 1173 228281 1176
rect 228315 1173 228327 1207
rect 228269 1167 228327 1173
rect 228361 1207 228419 1213
rect 228361 1173 228373 1207
rect 228407 1204 228419 1207
rect 236641 1207 236699 1213
rect 236641 1204 236653 1207
rect 228407 1176 236653 1204
rect 228407 1173 228419 1176
rect 228361 1167 228419 1173
rect 236641 1173 236653 1176
rect 236687 1173 236699 1207
rect 236641 1167 236699 1173
rect 236733 1207 236791 1213
rect 236733 1173 236745 1207
rect 236779 1204 236791 1207
rect 237929 1207 237987 1213
rect 237929 1204 237941 1207
rect 236779 1176 237941 1204
rect 236779 1173 236791 1176
rect 236733 1167 236791 1173
rect 237929 1173 237941 1176
rect 237975 1173 237987 1207
rect 237929 1167 237987 1173
rect 238018 1164 238024 1216
rect 238076 1204 238082 1216
rect 238386 1204 238392 1216
rect 238076 1176 238392 1204
rect 238076 1164 238082 1176
rect 238386 1164 238392 1176
rect 238444 1164 238450 1216
rect 238570 1164 238576 1216
rect 238628 1204 238634 1216
rect 238757 1207 238815 1213
rect 238757 1204 238769 1207
rect 238628 1176 238769 1204
rect 238628 1164 238634 1176
rect 238757 1173 238769 1176
rect 238803 1173 238815 1207
rect 238757 1167 238815 1173
rect 238938 1164 238944 1216
rect 238996 1204 239002 1216
rect 251177 1207 251235 1213
rect 251177 1204 251189 1207
rect 238996 1176 251189 1204
rect 238996 1164 239002 1176
rect 251177 1173 251189 1176
rect 251223 1173 251235 1207
rect 251177 1167 251235 1173
rect 251358 1164 251364 1216
rect 251416 1204 251422 1216
rect 260558 1204 260564 1216
rect 251416 1176 260564 1204
rect 251416 1164 251422 1176
rect 260558 1164 260564 1176
rect 260616 1164 260622 1216
rect 260745 1207 260803 1213
rect 260745 1173 260757 1207
rect 260791 1204 260803 1207
rect 270586 1204 270592 1216
rect 260791 1176 270592 1204
rect 260791 1173 260803 1176
rect 260745 1167 260803 1173
rect 270586 1164 270592 1176
rect 270644 1164 270650 1216
rect 270770 1164 270776 1216
rect 270828 1204 270834 1216
rect 279878 1204 279884 1216
rect 270828 1176 279884 1204
rect 270828 1164 270834 1176
rect 279878 1164 279884 1176
rect 279936 1164 279942 1216
rect 280065 1207 280123 1213
rect 280065 1173 280077 1207
rect 280111 1204 280123 1207
rect 281537 1207 281595 1213
rect 281537 1204 281549 1207
rect 280111 1176 281549 1204
rect 280111 1173 280123 1176
rect 280065 1167 280123 1173
rect 281537 1173 281549 1176
rect 281583 1173 281595 1207
rect 281537 1167 281595 1173
rect 281902 1164 281908 1216
rect 281960 1204 281966 1216
rect 281997 1207 282055 1213
rect 281997 1204 282009 1207
rect 281960 1176 282009 1204
rect 281960 1164 281966 1176
rect 281997 1173 282009 1176
rect 282043 1173 282055 1207
rect 281997 1167 282055 1173
rect 282089 1207 282147 1213
rect 282089 1173 282101 1207
rect 282135 1204 282147 1207
rect 290182 1204 290188 1216
rect 282135 1176 290188 1204
rect 282135 1173 282147 1176
rect 282089 1167 282147 1173
rect 290182 1164 290188 1176
rect 290240 1164 290246 1216
rect 290277 1207 290335 1213
rect 290277 1173 290289 1207
rect 290323 1204 290335 1207
rect 290550 1204 290556 1216
rect 290323 1176 290556 1204
rect 290323 1173 290335 1176
rect 290277 1167 290335 1173
rect 290550 1164 290556 1176
rect 290608 1164 290614 1216
rect 290645 1207 290703 1213
rect 290645 1173 290657 1207
rect 290691 1204 290703 1207
rect 290829 1207 290887 1213
rect 290829 1204 290841 1207
rect 290691 1176 290841 1204
rect 290691 1173 290703 1176
rect 290645 1167 290703 1173
rect 290829 1173 290841 1176
rect 290875 1173 290887 1207
rect 290829 1167 290887 1173
rect 291010 1164 291016 1216
rect 291068 1204 291074 1216
rect 293957 1207 294015 1213
rect 293957 1204 293969 1207
rect 291068 1176 293969 1204
rect 291068 1164 291074 1176
rect 293957 1173 293969 1176
rect 294003 1173 294015 1207
rect 293957 1167 294015 1173
rect 294049 1207 294107 1213
rect 294049 1173 294061 1207
rect 294095 1204 294107 1207
rect 295245 1207 295303 1213
rect 295245 1204 295257 1207
rect 294095 1176 295257 1204
rect 294095 1173 294107 1176
rect 294049 1167 294107 1173
rect 295245 1173 295257 1176
rect 295291 1173 295303 1207
rect 295245 1167 295303 1173
rect 295337 1207 295395 1213
rect 295337 1173 295349 1207
rect 295383 1204 295395 1207
rect 298020 1204 298048 1244
rect 309229 1241 309241 1244
rect 309275 1241 309287 1275
rect 318613 1275 318671 1281
rect 309229 1235 309287 1241
rect 309336 1244 318564 1272
rect 295383 1176 298048 1204
rect 298097 1207 298155 1213
rect 295383 1173 295395 1176
rect 295337 1167 295395 1173
rect 298097 1173 298109 1207
rect 298143 1204 298155 1207
rect 300670 1204 300676 1216
rect 298143 1176 300676 1204
rect 298143 1173 298155 1176
rect 298097 1167 298155 1173
rect 300670 1164 300676 1176
rect 300728 1164 300734 1216
rect 300765 1207 300823 1213
rect 300765 1173 300777 1207
rect 300811 1204 300823 1207
rect 309336 1204 309364 1244
rect 300811 1176 309364 1204
rect 309413 1207 309471 1213
rect 300811 1173 300823 1176
rect 300765 1167 300823 1173
rect 309413 1173 309425 1207
rect 309459 1204 309471 1207
rect 318426 1204 318432 1216
rect 309459 1176 318432 1204
rect 309459 1173 309471 1176
rect 309413 1167 309471 1173
rect 318426 1164 318432 1176
rect 318484 1164 318490 1216
rect 318536 1204 318564 1244
rect 318613 1241 318625 1275
rect 318659 1272 318671 1275
rect 327077 1275 327135 1281
rect 318659 1244 327028 1272
rect 318659 1241 318671 1244
rect 318613 1235 318671 1241
rect 326893 1207 326951 1213
rect 326893 1204 326905 1207
rect 318536 1176 326905 1204
rect 326893 1173 326905 1176
rect 326939 1173 326951 1207
rect 327000 1204 327028 1244
rect 327077 1241 327089 1275
rect 327123 1272 327135 1275
rect 327445 1275 327503 1281
rect 327445 1272 327457 1275
rect 327123 1244 327457 1272
rect 327123 1241 327135 1244
rect 327077 1235 327135 1241
rect 327445 1241 327457 1244
rect 327491 1241 327503 1275
rect 327445 1235 327503 1241
rect 327534 1232 327540 1284
rect 327592 1272 327598 1284
rect 329650 1272 329656 1284
rect 327592 1244 329656 1272
rect 327592 1232 327598 1244
rect 329650 1232 329656 1244
rect 329708 1232 329714 1284
rect 329745 1275 329803 1281
rect 329745 1241 329757 1275
rect 329791 1272 329803 1275
rect 335817 1275 335875 1281
rect 335817 1272 335829 1275
rect 329791 1244 335829 1272
rect 329791 1241 329803 1244
rect 329745 1235 329803 1241
rect 335817 1241 335829 1244
rect 335863 1241 335875 1275
rect 337565 1275 337623 1281
rect 337565 1272 337577 1275
rect 335817 1235 335875 1241
rect 335924 1244 337577 1272
rect 335924 1204 335952 1244
rect 337565 1241 337577 1244
rect 337611 1241 337623 1275
rect 338853 1275 338911 1281
rect 338853 1272 338865 1275
rect 337565 1235 337623 1241
rect 337672 1244 338865 1272
rect 327000 1176 335952 1204
rect 336001 1207 336059 1213
rect 326893 1167 326951 1173
rect 336001 1173 336013 1207
rect 336047 1204 336059 1207
rect 337672 1204 337700 1244
rect 338853 1241 338865 1244
rect 338899 1241 338911 1275
rect 338853 1235 338911 1241
rect 345385 1275 345443 1281
rect 345385 1241 345397 1275
rect 345431 1272 345443 1275
rect 357897 1275 357955 1281
rect 357897 1272 357909 1275
rect 345431 1244 357909 1272
rect 345431 1241 345443 1244
rect 345385 1235 345443 1241
rect 357897 1241 357909 1244
rect 357943 1241 357955 1275
rect 357897 1235 357955 1241
rect 357986 1232 357992 1284
rect 358044 1272 358050 1284
rect 365254 1272 365260 1284
rect 358044 1244 365260 1272
rect 358044 1232 358050 1244
rect 365254 1232 365260 1244
rect 365312 1232 365318 1284
rect 367281 1275 367339 1281
rect 367281 1241 367293 1275
rect 367327 1272 367339 1275
rect 374641 1275 374699 1281
rect 367327 1244 372660 1272
rect 367327 1241 367339 1244
rect 367281 1235 367339 1241
rect 336047 1176 337700 1204
rect 336047 1173 336059 1176
rect 336001 1167 336059 1173
rect 338298 1164 338304 1216
rect 338356 1204 338362 1216
rect 348513 1207 348571 1213
rect 348513 1204 348525 1207
rect 338356 1176 348525 1204
rect 338356 1164 338362 1176
rect 348513 1173 348525 1176
rect 348559 1173 348571 1207
rect 348513 1167 348571 1173
rect 348973 1207 349031 1213
rect 348973 1173 348985 1207
rect 349019 1204 349031 1207
rect 354030 1204 354036 1216
rect 349019 1176 354036 1204
rect 349019 1173 349031 1176
rect 348973 1167 349031 1173
rect 354030 1164 354036 1176
rect 354088 1164 354094 1216
rect 354125 1207 354183 1213
rect 354125 1173 354137 1207
rect 354171 1204 354183 1207
rect 355965 1207 356023 1213
rect 355965 1204 355977 1207
rect 354171 1176 355977 1204
rect 354171 1173 354183 1176
rect 354125 1167 354183 1173
rect 355965 1173 355977 1176
rect 356011 1173 356023 1207
rect 355965 1167 356023 1173
rect 356149 1207 356207 1213
rect 356149 1173 356161 1207
rect 356195 1204 356207 1207
rect 356974 1204 356980 1216
rect 356195 1176 356980 1204
rect 356195 1173 356207 1176
rect 356149 1167 356207 1173
rect 356974 1164 356980 1176
rect 357032 1164 357038 1216
rect 357069 1207 357127 1213
rect 357069 1173 357081 1207
rect 357115 1204 357127 1207
rect 367005 1207 367063 1213
rect 367005 1204 367017 1207
rect 357115 1176 367017 1204
rect 357115 1173 357127 1176
rect 357069 1167 357127 1173
rect 367005 1173 367017 1176
rect 367051 1173 367063 1207
rect 367005 1167 367063 1173
rect 367097 1207 367155 1213
rect 367097 1173 367109 1207
rect 367143 1204 367155 1207
rect 368385 1207 368443 1213
rect 368385 1204 368397 1207
rect 367143 1176 368397 1204
rect 367143 1173 367155 1176
rect 367097 1167 367155 1173
rect 368385 1173 368397 1176
rect 368431 1173 368443 1207
rect 372632 1204 372660 1244
rect 374641 1241 374653 1275
rect 374687 1272 374699 1275
rect 386417 1275 386475 1281
rect 386417 1272 386429 1275
rect 374687 1244 386429 1272
rect 374687 1241 374699 1244
rect 374641 1235 374699 1241
rect 386417 1241 386429 1244
rect 386463 1241 386475 1275
rect 386417 1235 386475 1241
rect 404265 1275 404323 1281
rect 404265 1241 404277 1275
rect 404311 1272 404323 1275
rect 424962 1272 424968 1284
rect 404311 1244 424968 1272
rect 404311 1241 404323 1244
rect 404265 1235 404323 1241
rect 424962 1232 424968 1244
rect 425020 1232 425026 1284
rect 432233 1275 432291 1281
rect 432233 1241 432245 1275
rect 432279 1272 432291 1275
rect 459557 1275 459615 1281
rect 459557 1272 459569 1275
rect 432279 1244 459569 1272
rect 432279 1241 432291 1244
rect 432233 1235 432291 1241
rect 459557 1241 459569 1244
rect 459603 1241 459615 1275
rect 459557 1235 459615 1241
rect 473173 1275 473231 1281
rect 473173 1241 473185 1275
rect 473219 1272 473231 1275
rect 473357 1275 473415 1281
rect 473357 1272 473369 1275
rect 473219 1244 473369 1272
rect 473219 1241 473231 1244
rect 473173 1235 473231 1241
rect 473357 1241 473369 1244
rect 473403 1241 473415 1275
rect 473357 1235 473415 1241
rect 480162 1232 480168 1284
rect 480220 1272 480226 1284
rect 492490 1272 492496 1284
rect 480220 1244 492496 1272
rect 480220 1232 480226 1244
rect 492490 1232 492496 1244
rect 492548 1232 492554 1284
rect 492674 1232 492680 1284
rect 492732 1272 492738 1284
rect 500957 1275 501015 1281
rect 500957 1272 500969 1275
rect 492732 1244 500969 1272
rect 492732 1232 492738 1244
rect 500957 1241 500969 1244
rect 501003 1241 501015 1275
rect 500957 1235 501015 1241
rect 509513 1275 509571 1281
rect 509513 1241 509525 1275
rect 509559 1272 509571 1275
rect 511994 1272 512000 1284
rect 509559 1244 512000 1272
rect 509559 1241 509571 1244
rect 509513 1235 509571 1241
rect 511994 1232 512000 1244
rect 512052 1232 512058 1284
rect 535362 1232 535368 1284
rect 535420 1272 535426 1284
rect 549162 1272 549168 1284
rect 535420 1244 549168 1272
rect 535420 1232 535426 1244
rect 549162 1232 549168 1244
rect 549220 1232 549226 1284
rect 549364 1272 549392 1312
rect 560205 1309 560217 1343
rect 560251 1340 560263 1343
rect 568298 1340 568304 1352
rect 560251 1312 568304 1340
rect 560251 1309 560263 1312
rect 560205 1303 560263 1309
rect 568298 1300 568304 1312
rect 568356 1300 568362 1352
rect 555421 1275 555479 1281
rect 555421 1272 555433 1275
rect 549364 1244 555433 1272
rect 555421 1241 555433 1244
rect 555467 1241 555479 1275
rect 555421 1235 555479 1241
rect 556157 1275 556215 1281
rect 556157 1241 556169 1275
rect 556203 1272 556215 1275
rect 564434 1272 564440 1284
rect 556203 1244 564440 1272
rect 556203 1241 556215 1244
rect 556157 1235 556215 1241
rect 564434 1232 564440 1244
rect 564492 1232 564498 1284
rect 374733 1207 374791 1213
rect 374733 1204 374745 1207
rect 372632 1176 374745 1204
rect 368385 1167 368443 1173
rect 374733 1173 374745 1176
rect 374779 1173 374791 1207
rect 374733 1167 374791 1173
rect 374825 1207 374883 1213
rect 374825 1173 374837 1207
rect 374871 1204 374883 1207
rect 386509 1207 386567 1213
rect 386509 1204 386521 1207
rect 374871 1176 386521 1204
rect 374871 1173 374883 1176
rect 374825 1167 374883 1173
rect 386509 1173 386521 1176
rect 386555 1173 386567 1207
rect 386509 1167 386567 1173
rect 391201 1207 391259 1213
rect 391201 1173 391213 1207
rect 391247 1204 391259 1207
rect 493962 1204 493968 1216
rect 391247 1176 493968 1204
rect 391247 1173 391259 1176
rect 391201 1167 391259 1173
rect 493962 1164 493968 1176
rect 494020 1164 494026 1216
rect 494238 1164 494244 1216
rect 494296 1204 494302 1216
rect 569494 1204 569500 1216
rect 494296 1176 569500 1204
rect 494296 1164 494302 1176
rect 569494 1164 569500 1176
rect 569552 1164 569558 1216
rect 160664 1108 160968 1136
rect 161014 1096 161020 1148
rect 161072 1136 161078 1148
rect 166902 1136 166908 1148
rect 161072 1108 166908 1136
rect 161072 1096 161078 1108
rect 166902 1096 166908 1108
rect 166960 1096 166966 1148
rect 166997 1139 167055 1145
rect 166997 1105 167009 1139
rect 167043 1136 167055 1139
rect 168929 1139 168987 1145
rect 168929 1136 168941 1139
rect 167043 1108 168941 1136
rect 167043 1105 167055 1108
rect 166997 1099 167055 1105
rect 168929 1105 168941 1108
rect 168975 1105 168987 1139
rect 168929 1099 168987 1105
rect 169018 1096 169024 1148
rect 169076 1136 169082 1148
rect 169573 1139 169631 1145
rect 169573 1136 169585 1139
rect 169076 1108 169585 1136
rect 169076 1096 169082 1108
rect 169573 1105 169585 1108
rect 169619 1105 169631 1139
rect 169573 1099 169631 1105
rect 169665 1139 169723 1145
rect 169665 1105 169677 1139
rect 169711 1136 169723 1139
rect 217873 1139 217931 1145
rect 217873 1136 217885 1139
rect 169711 1108 217885 1136
rect 169711 1105 169723 1108
rect 169665 1099 169723 1105
rect 217873 1105 217885 1108
rect 217919 1105 217931 1139
rect 217873 1099 217931 1105
rect 217962 1096 217968 1148
rect 218020 1136 218026 1148
rect 223758 1136 223764 1148
rect 218020 1108 223764 1136
rect 218020 1096 218026 1108
rect 223758 1096 223764 1108
rect 223816 1096 223822 1148
rect 223850 1096 223856 1148
rect 223908 1136 223914 1148
rect 223908 1108 223953 1136
rect 223908 1096 223914 1108
rect 224034 1096 224040 1148
rect 224092 1136 224098 1148
rect 225046 1136 225052 1148
rect 224092 1108 225052 1136
rect 224092 1096 224098 1108
rect 225046 1096 225052 1108
rect 225104 1096 225110 1148
rect 225141 1139 225199 1145
rect 225141 1105 225153 1139
rect 225187 1136 225199 1139
rect 225230 1136 225236 1148
rect 225187 1108 225236 1136
rect 225187 1105 225199 1108
rect 225141 1099 225199 1105
rect 225230 1096 225236 1108
rect 225288 1096 225294 1148
rect 225506 1136 225512 1148
rect 225467 1108 225512 1136
rect 225506 1096 225512 1108
rect 225564 1096 225570 1148
rect 225601 1139 225659 1145
rect 225601 1105 225613 1139
rect 225647 1136 225659 1139
rect 231673 1139 231731 1145
rect 231673 1136 231685 1139
rect 225647 1108 231685 1136
rect 225647 1105 225659 1108
rect 225601 1099 225659 1105
rect 231673 1105 231685 1108
rect 231719 1105 231731 1139
rect 231673 1099 231731 1105
rect 231765 1139 231823 1145
rect 231765 1105 231777 1139
rect 231811 1136 231823 1139
rect 247313 1139 247371 1145
rect 247313 1136 247325 1139
rect 231811 1108 247325 1136
rect 231811 1105 231823 1108
rect 231765 1099 231823 1105
rect 247313 1105 247325 1108
rect 247359 1105 247371 1139
rect 247313 1099 247371 1105
rect 247589 1139 247647 1145
rect 247589 1105 247601 1139
rect 247635 1136 247647 1139
rect 390649 1139 390707 1145
rect 390649 1136 390661 1139
rect 247635 1108 390661 1136
rect 247635 1105 247647 1108
rect 247589 1099 247647 1105
rect 390649 1105 390661 1108
rect 390695 1105 390707 1139
rect 390649 1099 390707 1105
rect 390833 1139 390891 1145
rect 390833 1105 390845 1139
rect 390879 1136 390891 1139
rect 493873 1139 493931 1145
rect 493873 1136 493885 1139
rect 390879 1108 493885 1136
rect 390879 1105 390891 1108
rect 390833 1099 390891 1105
rect 493873 1105 493885 1108
rect 493919 1105 493931 1139
rect 521657 1139 521715 1145
rect 521657 1136 521669 1139
rect 493873 1099 493931 1105
rect 494256 1108 521669 1136
rect 147815 1040 148088 1068
rect 148137 1071 148195 1077
rect 147815 1037 147827 1040
rect 147769 1031 147827 1037
rect 148137 1037 148149 1071
rect 148183 1068 148195 1071
rect 148870 1068 148876 1080
rect 148183 1040 148876 1068
rect 148183 1037 148195 1040
rect 148137 1031 148195 1037
rect 148870 1028 148876 1040
rect 148928 1028 148934 1080
rect 148965 1071 149023 1077
rect 148965 1037 148977 1071
rect 149011 1068 149023 1071
rect 149333 1071 149391 1077
rect 149333 1068 149345 1071
rect 149011 1040 149345 1068
rect 149011 1037 149023 1040
rect 148965 1031 149023 1037
rect 149333 1037 149345 1040
rect 149379 1037 149391 1071
rect 149333 1031 149391 1037
rect 149425 1071 149483 1077
rect 149425 1037 149437 1071
rect 149471 1068 149483 1071
rect 179325 1071 179383 1077
rect 179325 1068 179337 1071
rect 149471 1040 179337 1068
rect 149471 1037 149483 1040
rect 149425 1031 149483 1037
rect 179325 1037 179337 1040
rect 179371 1037 179383 1071
rect 179325 1031 179383 1037
rect 179601 1071 179659 1077
rect 179601 1037 179613 1071
rect 179647 1068 179659 1071
rect 224957 1071 225015 1077
rect 224957 1068 224969 1071
rect 179647 1040 224969 1068
rect 179647 1037 179659 1040
rect 179601 1031 179659 1037
rect 224957 1037 224969 1040
rect 225003 1037 225015 1071
rect 224957 1031 225015 1037
rect 225417 1071 225475 1077
rect 225417 1037 225429 1071
rect 225463 1068 225475 1071
rect 239033 1071 239091 1077
rect 239033 1068 239045 1071
rect 225463 1040 239045 1068
rect 225463 1037 225475 1040
rect 225417 1031 225475 1037
rect 239033 1037 239045 1040
rect 239079 1037 239091 1071
rect 239214 1068 239220 1080
rect 239175 1040 239220 1068
rect 239033 1031 239091 1037
rect 239214 1028 239220 1040
rect 239272 1028 239278 1080
rect 239309 1071 239367 1077
rect 239309 1037 239321 1071
rect 239355 1068 239367 1071
rect 245473 1071 245531 1077
rect 245473 1068 245485 1071
rect 239355 1040 245485 1068
rect 239355 1037 239367 1040
rect 239309 1031 239367 1037
rect 245473 1037 245485 1040
rect 245519 1037 245531 1071
rect 245473 1031 245531 1037
rect 245562 1028 245568 1080
rect 245620 1068 245626 1080
rect 247126 1068 247132 1080
rect 245620 1040 247132 1068
rect 245620 1028 245626 1040
rect 247126 1028 247132 1040
rect 247184 1028 247190 1080
rect 247494 1028 247500 1080
rect 247552 1068 247558 1080
rect 248230 1068 248236 1080
rect 247552 1040 248236 1068
rect 247552 1028 247558 1040
rect 248230 1028 248236 1040
rect 248288 1028 248294 1080
rect 248325 1071 248383 1077
rect 248325 1037 248337 1071
rect 248371 1068 248383 1071
rect 342165 1071 342223 1077
rect 342165 1068 342177 1071
rect 248371 1040 342177 1068
rect 248371 1037 248383 1040
rect 248325 1031 248383 1037
rect 342165 1037 342177 1040
rect 342211 1037 342223 1071
rect 345385 1071 345443 1077
rect 345385 1068 345397 1071
rect 342165 1031 342223 1037
rect 342272 1040 345397 1068
rect 124079 972 124260 1000
rect 124309 1003 124367 1009
rect 124079 969 124091 972
rect 124033 963 124091 969
rect 124309 969 124321 1003
rect 124355 1000 124367 1003
rect 125505 1003 125563 1009
rect 125505 1000 125517 1003
rect 124355 972 125517 1000
rect 124355 969 124367 972
rect 124309 963 124367 969
rect 125505 969 125517 972
rect 125551 969 125563 1003
rect 125505 963 125563 969
rect 125594 960 125600 1012
rect 125652 1000 125658 1012
rect 128909 1003 128967 1009
rect 128909 1000 128921 1003
rect 125652 972 128921 1000
rect 125652 960 125658 972
rect 128909 969 128921 972
rect 128955 969 128967 1003
rect 131666 1000 131672 1012
rect 128909 963 128967 969
rect 129016 972 131672 1000
rect 3326 892 3332 944
rect 3384 932 3390 944
rect 56778 932 56784 944
rect 3384 904 56784 932
rect 3384 892 3390 904
rect 56778 892 56784 904
rect 56836 892 56842 944
rect 56873 935 56931 941
rect 56873 901 56885 935
rect 56919 932 56931 935
rect 57977 935 58035 941
rect 57977 932 57989 935
rect 56919 904 57989 932
rect 56919 901 56931 904
rect 56873 895 56931 901
rect 57977 901 57989 904
rect 58023 901 58035 935
rect 57977 895 58035 901
rect 58066 892 58072 944
rect 58124 932 58130 944
rect 61194 932 61200 944
rect 58124 904 61200 932
rect 58124 892 58130 904
rect 61194 892 61200 904
rect 61252 892 61258 944
rect 61289 935 61347 941
rect 61289 901 61301 935
rect 61335 932 61347 935
rect 62942 932 62948 944
rect 61335 904 62948 932
rect 61335 901 61347 904
rect 61289 895 61347 901
rect 62942 892 62948 904
rect 63000 892 63006 944
rect 63313 935 63371 941
rect 63313 901 63325 935
rect 63359 932 63371 935
rect 64874 932 64880 944
rect 63359 904 64880 932
rect 63359 901 63371 904
rect 63313 895 63371 901
rect 64874 892 64880 904
rect 64932 892 64938 944
rect 64969 935 65027 941
rect 64969 901 64981 935
rect 65015 932 65027 935
rect 68833 935 68891 941
rect 68833 932 68845 935
rect 65015 904 68845 932
rect 65015 901 65027 904
rect 64969 895 65027 901
rect 68833 901 68845 904
rect 68879 901 68891 935
rect 68833 895 68891 901
rect 68922 892 68928 944
rect 68980 932 68986 944
rect 69385 935 69443 941
rect 69385 932 69397 935
rect 68980 904 69397 932
rect 68980 892 68986 904
rect 69385 901 69397 904
rect 69431 901 69443 935
rect 69385 895 69443 901
rect 69477 935 69535 941
rect 69477 901 69489 935
rect 69523 932 69535 935
rect 70581 935 70639 941
rect 70581 932 70593 935
rect 69523 904 70593 932
rect 69523 901 69535 904
rect 69477 895 69535 901
rect 70581 901 70593 904
rect 70627 901 70639 935
rect 70581 895 70639 901
rect 70670 892 70676 944
rect 70728 932 70734 944
rect 72973 935 73031 941
rect 70728 904 72924 932
rect 70728 892 70734 904
rect 1118 824 1124 876
rect 1176 864 1182 876
rect 4982 864 4988 876
rect 1176 836 4988 864
rect 1176 824 1182 836
rect 4982 824 4988 836
rect 5040 824 5046 876
rect 5629 867 5687 873
rect 5629 833 5641 867
rect 5675 864 5687 867
rect 25777 867 25835 873
rect 25777 864 25789 867
rect 5675 836 25789 864
rect 5675 833 5687 836
rect 5629 827 5687 833
rect 25777 833 25789 836
rect 25823 833 25835 867
rect 25777 827 25835 833
rect 25869 867 25927 873
rect 25869 833 25881 867
rect 25915 864 25927 867
rect 28169 867 28227 873
rect 28169 864 28181 867
rect 25915 836 28181 864
rect 25915 833 25927 836
rect 25869 827 25927 833
rect 28169 833 28181 836
rect 28215 833 28227 867
rect 28169 827 28227 833
rect 28258 824 28264 876
rect 28316 864 28322 876
rect 38289 867 38347 873
rect 38289 864 38301 867
rect 28316 836 38301 864
rect 28316 824 28322 836
rect 38289 833 38301 836
rect 38335 833 38347 867
rect 38289 827 38347 833
rect 38381 867 38439 873
rect 38381 833 38393 867
rect 38427 864 38439 867
rect 42150 864 42156 876
rect 38427 836 42156 864
rect 38427 833 38439 836
rect 38381 827 38439 833
rect 42150 824 42156 836
rect 42208 824 42214 876
rect 42429 867 42487 873
rect 42429 833 42441 867
rect 42475 864 42487 867
rect 46658 864 46664 876
rect 42475 836 46664 864
rect 42475 833 42487 836
rect 42429 827 42487 833
rect 46658 824 46664 836
rect 46716 824 46722 876
rect 63497 867 63555 873
rect 63497 864 63509 867
rect 46952 836 63509 864
rect 3050 756 3056 808
rect 3108 796 3114 808
rect 19337 799 19395 805
rect 19337 796 19349 799
rect 3108 768 19349 796
rect 3108 756 3114 768
rect 19337 765 19349 768
rect 19383 765 19395 799
rect 19337 759 19395 765
rect 19426 756 19432 808
rect 19484 796 19490 808
rect 19484 768 19529 796
rect 19484 756 19490 768
rect 29730 756 29736 808
rect 29788 796 29794 808
rect 38105 799 38163 805
rect 38105 796 38117 799
rect 29788 768 38117 796
rect 29788 756 29794 768
rect 38105 765 38117 768
rect 38151 765 38163 799
rect 38105 759 38163 765
rect 38194 756 38200 808
rect 38252 796 38258 808
rect 39485 799 39543 805
rect 39485 796 39497 799
rect 38252 768 39497 796
rect 38252 756 38258 768
rect 39485 765 39497 768
rect 39531 765 39543 799
rect 39485 759 39543 765
rect 42058 756 42064 808
rect 42116 796 42122 808
rect 42889 799 42947 805
rect 42889 796 42901 799
rect 42116 768 42901 796
rect 42116 756 42122 768
rect 42889 765 42901 768
rect 42935 765 42947 799
rect 42889 759 42947 765
rect 43346 756 43352 808
rect 43404 796 43410 808
rect 46952 796 46980 836
rect 63497 833 63509 836
rect 63543 833 63555 867
rect 63497 827 63555 833
rect 63681 867 63739 873
rect 63681 833 63693 867
rect 63727 864 63739 867
rect 63770 864 63776 876
rect 63727 836 63776 864
rect 63727 833 63739 836
rect 63681 827 63739 833
rect 63770 824 63776 836
rect 63828 824 63834 876
rect 63862 824 63868 876
rect 63920 864 63926 876
rect 72789 867 72847 873
rect 72789 864 72801 867
rect 63920 836 72801 864
rect 63920 824 63926 836
rect 72789 833 72801 836
rect 72835 833 72847 867
rect 72896 864 72924 904
rect 72973 901 72985 935
rect 73019 932 73031 935
rect 75457 935 75515 941
rect 75457 932 75469 935
rect 73019 904 75469 932
rect 73019 901 73031 904
rect 72973 895 73031 901
rect 75457 901 75469 904
rect 75503 901 75515 935
rect 75457 895 75515 901
rect 75549 935 75607 941
rect 75549 901 75561 935
rect 75595 932 75607 935
rect 76466 932 76472 944
rect 75595 904 76472 932
rect 75595 901 75607 904
rect 75549 895 75607 901
rect 76466 892 76472 904
rect 76524 892 76530 944
rect 76561 935 76619 941
rect 76561 901 76573 935
rect 76607 932 76619 935
rect 82909 935 82967 941
rect 82909 932 82921 935
rect 76607 904 82921 932
rect 76607 901 76619 904
rect 76561 895 76619 901
rect 82909 901 82921 904
rect 82955 901 82967 935
rect 82909 895 82967 901
rect 83093 935 83151 941
rect 83093 901 83105 935
rect 83139 932 83151 935
rect 97258 932 97264 944
rect 83139 904 97264 932
rect 83139 901 83151 904
rect 83093 895 83151 901
rect 97258 892 97264 904
rect 97316 892 97322 944
rect 97353 935 97411 941
rect 97353 901 97365 935
rect 97399 932 97411 935
rect 101033 935 101091 941
rect 101033 932 101045 935
rect 97399 904 101045 932
rect 97399 901 97411 904
rect 97353 895 97411 901
rect 101033 901 101045 904
rect 101079 901 101091 935
rect 101033 895 101091 901
rect 101309 935 101367 941
rect 101309 901 101321 935
rect 101355 932 101367 935
rect 101355 904 101628 932
rect 101355 901 101367 904
rect 101309 895 101367 901
rect 75917 867 75975 873
rect 75917 864 75929 867
rect 72896 836 75929 864
rect 72789 827 72847 833
rect 75917 833 75929 836
rect 75963 833 75975 867
rect 75917 827 75975 833
rect 76009 867 76067 873
rect 76009 833 76021 867
rect 76055 864 76067 867
rect 76745 867 76803 873
rect 76745 864 76757 867
rect 76055 836 76757 864
rect 76055 833 76067 836
rect 76009 827 76067 833
rect 76745 833 76757 836
rect 76791 833 76803 867
rect 76745 827 76803 833
rect 76834 824 76840 876
rect 76892 864 76898 876
rect 82538 864 82544 876
rect 76892 836 82544 864
rect 76892 824 76898 836
rect 82538 824 82544 836
rect 82596 824 82602 876
rect 82722 824 82728 876
rect 82780 864 82786 876
rect 83369 867 83427 873
rect 82780 836 83136 864
rect 82780 824 82786 836
rect 43404 768 46980 796
rect 43404 756 43410 768
rect 48038 756 48044 808
rect 48096 796 48102 808
rect 49145 799 49203 805
rect 49145 796 49157 799
rect 48096 768 49157 796
rect 48096 756 48102 768
rect 49145 765 49157 768
rect 49191 765 49203 799
rect 49145 759 49203 765
rect 49697 799 49755 805
rect 49697 765 49709 799
rect 49743 796 49755 799
rect 55214 796 55220 808
rect 49743 768 55220 796
rect 49743 765 49755 768
rect 49697 759 49755 765
rect 55214 756 55220 768
rect 55272 756 55278 808
rect 55309 799 55367 805
rect 55309 765 55321 799
rect 55355 796 55367 799
rect 76561 799 76619 805
rect 76561 796 76573 799
rect 55355 768 76573 796
rect 55355 765 55367 768
rect 55309 759 55367 765
rect 76561 765 76573 768
rect 76607 765 76619 799
rect 76561 759 76619 765
rect 76653 799 76711 805
rect 76653 765 76665 799
rect 76699 796 76711 799
rect 78953 799 79011 805
rect 78953 796 78965 799
rect 76699 768 78965 796
rect 76699 765 76711 768
rect 76653 759 76711 765
rect 78953 765 78965 768
rect 78999 765 79011 799
rect 78953 759 79011 765
rect 79042 756 79048 808
rect 79100 796 79106 808
rect 83001 799 83059 805
rect 83001 796 83013 799
rect 79100 768 83013 796
rect 79100 756 79106 768
rect 83001 765 83013 768
rect 83047 765 83059 799
rect 83108 796 83136 836
rect 83369 833 83381 867
rect 83415 864 83427 867
rect 83826 864 83832 876
rect 83415 836 83832 864
rect 83415 833 83427 836
rect 83369 827 83427 833
rect 83826 824 83832 836
rect 83884 824 83890 876
rect 84105 867 84163 873
rect 84105 833 84117 867
rect 84151 864 84163 867
rect 84746 864 84752 876
rect 84151 836 84752 864
rect 84151 833 84163 836
rect 84105 827 84163 833
rect 84746 824 84752 836
rect 84804 824 84810 876
rect 84841 867 84899 873
rect 84841 833 84853 867
rect 84887 864 84899 867
rect 85853 867 85911 873
rect 85853 864 85865 867
rect 84887 836 85865 864
rect 84887 833 84899 836
rect 84841 827 84899 833
rect 85853 833 85865 836
rect 85899 833 85911 867
rect 85853 827 85911 833
rect 86405 867 86463 873
rect 86405 833 86417 867
rect 86451 864 86463 867
rect 87785 867 87843 873
rect 87785 864 87797 867
rect 86451 836 87797 864
rect 86451 833 86463 836
rect 86405 827 86463 833
rect 87785 833 87797 836
rect 87831 833 87843 867
rect 87785 827 87843 833
rect 87874 824 87880 876
rect 87932 864 87938 876
rect 93397 867 93455 873
rect 93397 864 93409 867
rect 87932 836 93409 864
rect 87932 824 87938 836
rect 93397 833 93409 836
rect 93443 833 93455 867
rect 93397 827 93455 833
rect 93486 824 93492 876
rect 93544 864 93550 876
rect 93949 867 94007 873
rect 93949 864 93961 867
rect 93544 836 93961 864
rect 93544 824 93550 836
rect 93949 833 93961 836
rect 93995 833 94007 867
rect 93949 827 94007 833
rect 94038 824 94044 876
rect 94096 864 94102 876
rect 96341 867 96399 873
rect 96341 864 96353 867
rect 94096 836 96353 864
rect 94096 824 94102 836
rect 96341 833 96353 836
rect 96387 833 96399 867
rect 96341 827 96399 833
rect 96433 867 96491 873
rect 96433 833 96445 867
rect 96479 864 96491 867
rect 96985 867 97043 873
rect 96985 864 96997 867
rect 96479 836 96997 864
rect 96479 833 96491 836
rect 96433 827 96491 833
rect 96985 833 96997 836
rect 97031 833 97043 867
rect 96985 827 97043 833
rect 97074 824 97080 876
rect 97132 864 97138 876
rect 101125 867 101183 873
rect 101125 864 101137 867
rect 97132 836 101137 864
rect 97132 824 97138 836
rect 101125 833 101137 836
rect 101171 833 101183 867
rect 101125 827 101183 833
rect 101217 867 101275 873
rect 101217 833 101229 867
rect 101263 864 101275 867
rect 101600 864 101628 904
rect 101674 892 101680 944
rect 101732 932 101738 944
rect 101861 935 101919 941
rect 101861 932 101873 935
rect 101732 904 101873 932
rect 101732 892 101738 904
rect 101861 901 101873 904
rect 101907 901 101919 935
rect 101861 895 101919 901
rect 102873 935 102931 941
rect 102873 901 102885 935
rect 102919 932 102931 935
rect 116578 932 116584 944
rect 102919 904 116584 932
rect 102919 901 102931 904
rect 102873 895 102931 901
rect 116578 892 116584 904
rect 116636 892 116642 944
rect 116673 935 116731 941
rect 116673 901 116685 935
rect 116719 932 116731 935
rect 117041 935 117099 941
rect 117041 932 117053 935
rect 116719 904 117053 932
rect 116719 901 116731 904
rect 116673 895 116731 901
rect 117041 901 117053 904
rect 117087 901 117099 935
rect 117041 895 117099 901
rect 117130 892 117136 944
rect 117188 932 117194 944
rect 122558 932 122564 944
rect 117188 904 122564 932
rect 117188 892 117194 904
rect 122558 892 122564 904
rect 122616 892 122622 944
rect 122653 935 122711 941
rect 122653 901 122665 935
rect 122699 932 122711 935
rect 123478 932 123484 944
rect 122699 904 123484 932
rect 122699 901 122711 904
rect 122653 895 122711 901
rect 123478 892 123484 904
rect 123536 892 123542 944
rect 123570 892 123576 944
rect 123628 932 123634 944
rect 129016 932 129044 972
rect 131666 960 131672 972
rect 131724 960 131730 1012
rect 131761 1003 131819 1009
rect 131761 969 131773 1003
rect 131807 1000 131819 1003
rect 140685 1003 140743 1009
rect 140685 1000 140697 1003
rect 131807 972 140697 1000
rect 131807 969 131819 972
rect 131761 963 131819 969
rect 140685 969 140697 972
rect 140731 969 140743 1003
rect 140685 963 140743 969
rect 140869 1003 140927 1009
rect 140869 969 140881 1003
rect 140915 1000 140927 1003
rect 145561 1003 145619 1009
rect 145561 1000 145573 1003
rect 140915 972 145573 1000
rect 140915 969 140927 972
rect 140869 963 140927 969
rect 145561 969 145573 972
rect 145607 969 145619 1003
rect 146110 1000 146116 1012
rect 145561 963 145619 969
rect 145668 972 146116 1000
rect 123628 904 129044 932
rect 123628 892 123634 904
rect 129090 892 129096 944
rect 129148 932 129154 944
rect 129277 935 129335 941
rect 129148 904 129193 932
rect 129148 892 129154 904
rect 129277 901 129289 935
rect 129323 932 129335 935
rect 129458 932 129464 944
rect 129323 904 129464 932
rect 129323 901 129335 904
rect 129277 895 129335 901
rect 129458 892 129464 904
rect 129516 892 129522 944
rect 129553 935 129611 941
rect 129553 901 129565 935
rect 129599 932 129611 935
rect 134613 935 134671 941
rect 134613 932 134625 935
rect 129599 904 134625 932
rect 129599 901 129611 904
rect 129553 895 129611 901
rect 134613 901 134625 904
rect 134659 901 134671 935
rect 134613 895 134671 901
rect 134797 935 134855 941
rect 134797 901 134809 935
rect 134843 932 134855 935
rect 135257 935 135315 941
rect 135257 932 135269 935
rect 134843 904 135269 932
rect 134843 901 134855 904
rect 134797 895 134855 901
rect 135257 901 135269 904
rect 135303 901 135315 935
rect 135257 895 135315 901
rect 135349 935 135407 941
rect 135349 901 135361 935
rect 135395 932 135407 935
rect 136085 935 136143 941
rect 136085 932 136097 935
rect 135395 904 136097 932
rect 135395 901 135407 904
rect 135349 895 135407 901
rect 136085 901 136097 904
rect 136131 901 136143 935
rect 136085 895 136143 901
rect 136177 935 136235 941
rect 136177 901 136189 935
rect 136223 932 136235 935
rect 140409 935 140467 941
rect 140409 932 140421 935
rect 136223 904 140421 932
rect 136223 901 136235 904
rect 136177 895 136235 901
rect 140409 901 140421 904
rect 140455 901 140467 935
rect 140409 895 140467 901
rect 140498 892 140504 944
rect 140556 932 140562 944
rect 141145 935 141203 941
rect 140556 904 140601 932
rect 140556 892 140562 904
rect 141145 901 141157 935
rect 141191 932 141203 935
rect 142341 935 142399 941
rect 142341 932 142353 935
rect 141191 904 142353 932
rect 141191 901 141203 904
rect 141145 895 141203 901
rect 142341 901 142353 904
rect 142387 901 142399 935
rect 142341 895 142399 901
rect 142430 892 142436 944
rect 142488 932 142494 944
rect 143169 935 143227 941
rect 143169 932 143181 935
rect 142488 904 143181 932
rect 142488 892 142494 904
rect 143169 901 143181 904
rect 143215 901 143227 935
rect 143169 895 143227 901
rect 143261 935 143319 941
rect 143261 901 143273 935
rect 143307 932 143319 935
rect 145668 932 145696 972
rect 146110 960 146116 972
rect 146168 960 146174 1012
rect 152001 1003 152059 1009
rect 152001 1000 152013 1003
rect 146220 972 152013 1000
rect 143307 904 145696 932
rect 145745 935 145803 941
rect 143307 901 143319 904
rect 143261 895 143319 901
rect 145745 901 145757 935
rect 145791 932 145803 935
rect 146220 932 146248 972
rect 152001 969 152013 972
rect 152047 969 152059 1003
rect 152001 963 152059 969
rect 152277 1003 152335 1009
rect 152277 969 152289 1003
rect 152323 1000 152335 1003
rect 179233 1003 179291 1009
rect 179233 1000 179245 1003
rect 152323 972 160968 1000
rect 152323 969 152335 972
rect 152277 963 152335 969
rect 145791 904 146248 932
rect 146297 935 146355 941
rect 145791 901 145803 904
rect 145745 895 145803 901
rect 146297 901 146309 935
rect 146343 932 146355 935
rect 147309 935 147367 941
rect 147309 932 147321 935
rect 146343 904 147321 932
rect 146343 901 146355 904
rect 146297 895 146355 901
rect 147309 901 147321 904
rect 147355 901 147367 935
rect 147309 895 147367 901
rect 147401 935 147459 941
rect 147401 901 147413 935
rect 147447 932 147459 935
rect 149425 935 149483 941
rect 149425 932 149437 935
rect 147447 904 149437 932
rect 147447 901 147459 904
rect 147401 895 147459 901
rect 149425 901 149437 904
rect 149471 901 149483 935
rect 149425 895 149483 901
rect 149514 892 149520 944
rect 149572 932 149578 944
rect 150069 935 150127 941
rect 150069 932 150081 935
rect 149572 904 150081 932
rect 149572 892 149578 904
rect 150069 901 150081 904
rect 150115 901 150127 935
rect 150069 895 150127 901
rect 150161 935 150219 941
rect 150161 901 150173 935
rect 150207 932 150219 935
rect 152366 932 152372 944
rect 150207 904 152372 932
rect 150207 901 150219 904
rect 150161 895 150219 901
rect 152366 892 152372 904
rect 152424 892 152430 944
rect 152461 935 152519 941
rect 152461 901 152473 935
rect 152507 932 152519 935
rect 154114 932 154120 944
rect 152507 904 154120 932
rect 152507 901 152519 904
rect 152461 895 152519 901
rect 154114 892 154120 904
rect 154172 892 154178 944
rect 154390 892 154396 944
rect 154448 932 154454 944
rect 155126 932 155132 944
rect 154448 904 155132 932
rect 154448 892 154454 904
rect 155126 892 155132 904
rect 155184 892 155190 944
rect 155221 935 155279 941
rect 155221 901 155233 935
rect 155267 932 155279 935
rect 157153 935 157211 941
rect 155267 904 157104 932
rect 155267 901 155279 904
rect 155221 895 155279 901
rect 103422 864 103428 876
rect 101263 836 101536 864
rect 101600 836 103428 864
rect 101263 833 101275 836
rect 101217 827 101275 833
rect 83642 796 83648 808
rect 83108 768 83648 796
rect 83001 759 83059 765
rect 83642 756 83648 768
rect 83700 756 83706 808
rect 92569 799 92627 805
rect 92569 796 92581 799
rect 83752 768 92581 796
rect 842 688 848 740
rect 900 728 906 740
rect 5261 731 5319 737
rect 5261 728 5273 731
rect 900 700 5273 728
rect 900 688 906 700
rect 5261 697 5273 700
rect 5307 697 5319 731
rect 5261 691 5319 697
rect 5353 731 5411 737
rect 5353 697 5365 731
rect 5399 728 5411 731
rect 13173 731 13231 737
rect 13173 728 13185 731
rect 5399 700 13185 728
rect 5399 697 5411 700
rect 5353 691 5411 697
rect 13173 697 13185 700
rect 13219 697 13231 731
rect 13173 691 13231 697
rect 13262 688 13268 740
rect 13320 728 13326 740
rect 15194 728 15200 740
rect 13320 700 15200 728
rect 13320 688 13326 700
rect 15194 688 15200 700
rect 15252 688 15258 740
rect 17954 688 17960 740
rect 18012 728 18018 740
rect 83752 728 83780 768
rect 92569 765 92581 768
rect 92615 765 92627 799
rect 92569 759 92627 765
rect 92658 756 92664 808
rect 92716 796 92722 808
rect 92842 796 92848 808
rect 92716 768 92848 796
rect 92716 756 92722 768
rect 92842 756 92848 768
rect 92900 756 92906 808
rect 92937 799 92995 805
rect 92937 765 92949 799
rect 92983 796 92995 799
rect 93026 796 93032 808
rect 92983 768 93032 796
rect 92983 765 92995 768
rect 92937 759 92995 765
rect 93026 756 93032 768
rect 93084 756 93090 808
rect 93121 799 93179 805
rect 93121 765 93133 799
rect 93167 796 93179 799
rect 100573 799 100631 805
rect 100573 796 100585 799
rect 93167 768 100585 796
rect 93167 765 93179 768
rect 93121 759 93179 765
rect 100573 765 100585 768
rect 100619 765 100631 799
rect 100573 759 100631 765
rect 100849 799 100907 805
rect 100849 765 100861 799
rect 100895 796 100907 799
rect 101398 796 101404 808
rect 100895 768 101404 796
rect 100895 765 100907 768
rect 100849 759 100907 765
rect 101398 756 101404 768
rect 101456 756 101462 808
rect 101508 796 101536 836
rect 103422 824 103428 836
rect 103480 824 103486 876
rect 103517 867 103575 873
rect 103517 833 103529 867
rect 103563 864 103575 867
rect 106369 867 106427 873
rect 106369 864 106381 867
rect 103563 836 106381 864
rect 103563 833 103575 836
rect 103517 827 103575 833
rect 106369 833 106381 836
rect 106415 833 106427 867
rect 106369 827 106427 833
rect 106458 824 106464 876
rect 106516 864 106522 876
rect 106553 867 106611 873
rect 106553 864 106565 867
rect 106516 836 106565 864
rect 106516 824 106522 836
rect 106553 833 106565 836
rect 106599 833 106611 867
rect 106553 827 106611 833
rect 107289 867 107347 873
rect 107289 833 107301 867
rect 107335 864 107347 867
rect 108850 864 108856 876
rect 107335 836 108856 864
rect 107335 833 107347 836
rect 107289 827 107347 833
rect 108850 824 108856 836
rect 108908 824 108914 876
rect 109313 867 109371 873
rect 109313 864 109325 867
rect 108960 836 109325 864
rect 101950 796 101956 808
rect 101508 768 101956 796
rect 101950 756 101956 768
rect 102008 756 102014 808
rect 102229 799 102287 805
rect 102229 765 102241 799
rect 102275 796 102287 799
rect 106918 796 106924 808
rect 102275 768 106924 796
rect 102275 765 102287 768
rect 102229 759 102287 765
rect 106918 756 106924 768
rect 106976 756 106982 808
rect 107010 756 107016 808
rect 107068 796 107074 808
rect 107068 768 107976 796
rect 107068 756 107074 768
rect 18012 700 83780 728
rect 18012 688 18018 700
rect 83826 688 83832 740
rect 83884 728 83890 740
rect 91557 731 91615 737
rect 91557 728 91569 731
rect 83884 700 91569 728
rect 83884 688 83890 700
rect 91557 697 91569 700
rect 91603 697 91615 731
rect 91557 691 91615 697
rect 91649 731 91707 737
rect 91649 697 91661 731
rect 91695 728 91707 731
rect 97353 731 97411 737
rect 97353 728 97365 731
rect 91695 700 97365 728
rect 91695 697 91707 700
rect 91649 691 91707 697
rect 97353 697 97365 700
rect 97399 697 97411 731
rect 97353 691 97411 697
rect 97445 731 97503 737
rect 97445 697 97457 731
rect 97491 728 97503 731
rect 100113 731 100171 737
rect 100113 728 100125 731
rect 97491 700 100125 728
rect 97491 697 97503 700
rect 97445 691 97503 697
rect 100113 697 100125 700
rect 100159 697 100171 731
rect 100113 691 100171 697
rect 100481 731 100539 737
rect 100481 697 100493 731
rect 100527 728 100539 731
rect 100665 731 100723 737
rect 100665 728 100677 731
rect 100527 700 100677 728
rect 100527 697 100539 700
rect 100481 691 100539 697
rect 100665 697 100677 700
rect 100711 697 100723 731
rect 100665 691 100723 697
rect 100754 688 100760 740
rect 100812 728 100818 740
rect 102321 731 102379 737
rect 102321 728 102333 731
rect 100812 700 102333 728
rect 100812 688 100818 700
rect 102321 697 102333 700
rect 102367 697 102379 731
rect 102321 691 102379 697
rect 102410 688 102416 740
rect 102468 728 102474 740
rect 102597 731 102655 737
rect 102597 728 102609 731
rect 102468 700 102609 728
rect 102468 688 102474 700
rect 102597 697 102609 700
rect 102643 697 102655 731
rect 102597 691 102655 697
rect 102686 688 102692 740
rect 102744 728 102750 740
rect 107838 728 107844 740
rect 102744 700 107844 728
rect 102744 688 102750 700
rect 107838 688 107844 700
rect 107896 688 107902 740
rect 107948 728 107976 768
rect 108022 756 108028 808
rect 108080 796 108086 808
rect 108960 796 108988 836
rect 109313 833 109325 836
rect 109359 833 109371 867
rect 109313 827 109371 833
rect 109402 824 109408 876
rect 109460 864 109466 876
rect 109954 864 109960 876
rect 109460 836 109960 864
rect 109460 824 109466 836
rect 109954 824 109960 836
rect 110012 824 110018 876
rect 110046 824 110052 876
rect 110104 864 110110 876
rect 110785 867 110843 873
rect 110785 864 110797 867
rect 110104 836 110797 864
rect 110104 824 110110 836
rect 110785 833 110797 836
rect 110831 833 110843 867
rect 110785 827 110843 833
rect 110877 867 110935 873
rect 110877 833 110889 867
rect 110923 864 110935 867
rect 111797 867 111855 873
rect 111797 864 111809 867
rect 110923 836 111809 864
rect 110923 833 110935 836
rect 110877 827 110935 833
rect 111797 833 111809 836
rect 111843 833 111855 867
rect 112533 867 112591 873
rect 111797 827 111855 833
rect 111904 836 112484 864
rect 108080 768 108988 796
rect 109037 799 109095 805
rect 108080 756 108086 768
rect 109037 765 109049 799
rect 109083 796 109095 799
rect 111061 799 111119 805
rect 111061 796 111073 799
rect 109083 768 111073 796
rect 109083 765 109095 768
rect 109037 759 109095 765
rect 111061 765 111073 768
rect 111107 765 111119 799
rect 111061 759 111119 765
rect 111153 799 111211 805
rect 111153 765 111165 799
rect 111199 796 111211 799
rect 111705 799 111763 805
rect 111705 796 111717 799
rect 111199 768 111717 796
rect 111199 765 111211 768
rect 111153 759 111211 765
rect 111705 765 111717 768
rect 111751 765 111763 799
rect 111705 759 111763 765
rect 111518 728 111524 740
rect 107948 700 111524 728
rect 111518 688 111524 700
rect 111576 688 111582 740
rect 111610 688 111616 740
rect 111668 728 111674 740
rect 111904 728 111932 836
rect 111981 799 112039 805
rect 111981 765 111993 799
rect 112027 796 112039 799
rect 112346 796 112352 808
rect 112027 768 112352 796
rect 112027 765 112039 768
rect 111981 759 112039 765
rect 112346 756 112352 768
rect 112404 756 112410 808
rect 112456 796 112484 836
rect 112533 833 112545 867
rect 112579 864 112591 867
rect 114741 867 114799 873
rect 114741 864 114753 867
rect 112579 836 114753 864
rect 112579 833 112591 836
rect 112533 827 112591 833
rect 114741 833 114753 836
rect 114787 833 114799 867
rect 114741 827 114799 833
rect 114833 867 114891 873
rect 114833 833 114845 867
rect 114879 864 114891 867
rect 121365 867 121423 873
rect 114879 836 121316 864
rect 114879 833 114891 836
rect 114833 827 114891 833
rect 112806 796 112812 808
rect 112456 768 112812 796
rect 112806 756 112812 768
rect 112864 756 112870 808
rect 112901 799 112959 805
rect 112901 765 112913 799
rect 112947 796 112959 799
rect 113542 796 113548 808
rect 112947 768 113548 796
rect 112947 765 112959 768
rect 112901 759 112959 765
rect 113542 756 113548 768
rect 113600 756 113606 808
rect 113726 756 113732 808
rect 113784 796 113790 808
rect 120534 796 120540 808
rect 113784 768 120540 796
rect 113784 756 113790 768
rect 120534 756 120540 768
rect 120592 756 120598 808
rect 120718 796 120724 808
rect 120679 768 120724 796
rect 120718 756 120724 768
rect 120776 756 120782 808
rect 121288 805 121316 836
rect 121365 833 121377 867
rect 121411 864 121423 867
rect 153289 867 153347 873
rect 153289 864 153301 867
rect 121411 836 153301 864
rect 121411 833 121423 836
rect 121365 827 121423 833
rect 153289 833 153301 836
rect 153335 833 153347 867
rect 153289 827 153347 833
rect 153396 836 157012 864
rect 121273 799 121331 805
rect 121273 765 121285 799
rect 121319 765 121331 799
rect 121273 759 121331 765
rect 121457 799 121515 805
rect 121457 765 121469 799
rect 121503 796 121515 799
rect 122466 796 122472 808
rect 121503 768 122472 796
rect 121503 765 121515 768
rect 121457 759 121515 765
rect 122466 756 122472 768
rect 122524 756 122530 808
rect 122558 756 122564 808
rect 122616 796 122622 808
rect 152001 799 152059 805
rect 152001 796 152013 799
rect 122616 768 152013 796
rect 122616 756 122622 768
rect 152001 765 152013 768
rect 152047 765 152059 799
rect 152001 759 152059 765
rect 152090 756 152096 808
rect 152148 796 152154 808
rect 153396 805 153424 836
rect 153197 799 153255 805
rect 153197 796 153209 799
rect 152148 768 153209 796
rect 152148 756 152154 768
rect 153197 765 153209 768
rect 153243 765 153255 799
rect 153197 759 153255 765
rect 153381 799 153439 805
rect 153381 765 153393 799
rect 153427 765 153439 799
rect 153381 759 153439 765
rect 153470 756 153476 808
rect 153528 796 153534 808
rect 153841 799 153899 805
rect 153841 796 153853 799
rect 153528 768 153853 796
rect 153528 756 153534 768
rect 153841 765 153853 768
rect 153887 765 153899 799
rect 153841 759 153899 765
rect 153933 799 153991 805
rect 153933 765 153945 799
rect 153979 796 153991 799
rect 154301 799 154359 805
rect 154301 796 154313 799
rect 153979 768 154313 796
rect 153979 765 153991 768
rect 153933 759 153991 765
rect 154301 765 154313 768
rect 154347 765 154359 799
rect 154301 759 154359 765
rect 154393 799 154451 805
rect 154393 765 154405 799
rect 154439 796 154451 799
rect 156877 799 156935 805
rect 156877 796 156889 799
rect 154439 768 156889 796
rect 154439 765 154451 768
rect 154393 759 154451 765
rect 156877 765 156889 768
rect 156923 765 156935 799
rect 156877 759 156935 765
rect 111668 700 111932 728
rect 111668 688 111674 700
rect 112070 688 112076 740
rect 112128 728 112134 740
rect 152182 728 152188 740
rect 112128 700 152188 728
rect 112128 688 112134 700
rect 152182 688 152188 700
rect 152240 688 152246 740
rect 152277 731 152335 737
rect 152277 697 152289 731
rect 152323 728 152335 731
rect 152323 700 153516 728
rect 152323 697 152335 700
rect 152277 691 152335 697
rect 1302 620 1308 672
rect 1360 660 1366 672
rect 5077 663 5135 669
rect 5077 660 5089 663
rect 1360 632 5089 660
rect 1360 620 1366 632
rect 5077 629 5089 632
rect 5123 629 5135 663
rect 7285 663 7343 669
rect 7285 660 7297 663
rect 5077 623 5135 629
rect 5276 632 7297 660
rect 106 552 112 604
rect 164 592 170 604
rect 4890 592 4896 604
rect 164 564 4896 592
rect 164 552 170 564
rect 4890 552 4896 564
rect 4948 552 4954 604
rect 5169 595 5227 601
rect 5169 561 5181 595
rect 5215 592 5227 595
rect 5276 592 5304 632
rect 7285 629 7297 632
rect 7331 629 7343 663
rect 7285 623 7343 629
rect 7374 620 7380 672
rect 7432 660 7438 672
rect 7432 632 26648 660
rect 7432 620 7438 632
rect 5215 564 5304 592
rect 9677 595 9735 601
rect 5215 561 5227 564
rect 5169 555 5227 561
rect 9677 561 9689 595
rect 9723 592 9735 595
rect 10413 595 10471 601
rect 10413 592 10425 595
rect 9723 564 10425 592
rect 9723 561 9735 564
rect 9677 555 9735 561
rect 10413 561 10425 564
rect 10459 561 10471 595
rect 10413 555 10471 561
rect 10502 552 10508 604
rect 10560 592 10566 604
rect 13446 592 13452 604
rect 10560 564 13452 592
rect 10560 552 10566 564
rect 13446 552 13452 564
rect 13504 552 13510 604
rect 14277 595 14335 601
rect 14277 561 14289 595
rect 14323 592 14335 595
rect 22186 592 22192 604
rect 14323 564 22192 592
rect 14323 561 14335 564
rect 14277 555 14335 561
rect 22186 552 22192 564
rect 22244 552 22250 604
rect 26620 592 26648 632
rect 26694 620 26700 672
rect 26752 660 26758 672
rect 39301 663 39359 669
rect 39301 660 39313 663
rect 26752 632 39313 660
rect 26752 620 26758 632
rect 39301 629 39313 632
rect 39347 629 39359 663
rect 39301 623 39359 629
rect 39577 663 39635 669
rect 39577 629 39589 663
rect 39623 660 39635 663
rect 46750 660 46756 672
rect 39623 632 46756 660
rect 39623 629 39635 632
rect 39577 623 39635 629
rect 46750 620 46756 632
rect 46808 620 46814 672
rect 46934 620 46940 672
rect 46992 660 46998 672
rect 49697 663 49755 669
rect 49697 660 49709 663
rect 46992 632 49709 660
rect 46992 620 46998 632
rect 49697 629 49709 632
rect 49743 629 49755 663
rect 49697 623 49755 629
rect 49789 663 49847 669
rect 49789 629 49801 663
rect 49835 660 49847 663
rect 59354 660 59360 672
rect 49835 632 59360 660
rect 49835 629 49847 632
rect 49789 623 49847 629
rect 59354 620 59360 632
rect 59412 620 59418 672
rect 59998 620 60004 672
rect 60056 660 60062 672
rect 73157 663 73215 669
rect 73157 660 73169 663
rect 60056 632 73169 660
rect 60056 620 60062 632
rect 73157 629 73169 632
rect 73203 629 73215 663
rect 73157 623 73215 629
rect 73249 663 73307 669
rect 73249 629 73261 663
rect 73295 660 73307 663
rect 75549 663 75607 669
rect 75549 660 75561 663
rect 73295 632 75561 660
rect 73295 629 73307 632
rect 73249 623 73307 629
rect 75549 629 75561 632
rect 75595 629 75607 663
rect 75549 623 75607 629
rect 75638 620 75644 672
rect 75696 660 75702 672
rect 75825 663 75883 669
rect 75825 660 75837 663
rect 75696 632 75837 660
rect 75696 620 75702 632
rect 75825 629 75837 632
rect 75871 629 75883 663
rect 75825 623 75883 629
rect 75917 663 75975 669
rect 75917 629 75929 663
rect 75963 660 75975 663
rect 82265 663 82323 669
rect 82265 660 82277 663
rect 75963 632 82277 660
rect 75963 629 75975 632
rect 75917 623 75975 629
rect 82265 629 82277 632
rect 82311 629 82323 663
rect 82265 623 82323 629
rect 82725 663 82783 669
rect 82725 629 82737 663
rect 82771 660 82783 663
rect 92109 663 92167 669
rect 92109 660 92121 663
rect 82771 632 92121 660
rect 82771 629 82783 632
rect 82725 623 82783 629
rect 92109 629 92121 632
rect 92155 629 92167 663
rect 92109 623 92167 629
rect 92477 663 92535 669
rect 92477 629 92489 663
rect 92523 660 92535 663
rect 111705 663 111763 669
rect 92523 632 111564 660
rect 92523 629 92535 632
rect 92477 623 92535 629
rect 49237 595 49295 601
rect 49237 592 49249 595
rect 26620 564 49249 592
rect 49237 561 49249 564
rect 49283 561 49295 595
rect 49237 555 49295 561
rect 52822 552 52828 604
rect 52880 592 52886 604
rect 52880 564 93348 592
rect 52880 552 52886 564
rect 3602 484 3608 536
rect 3660 524 3666 536
rect 3660 496 4844 524
rect 3660 484 3666 496
rect 1026 416 1032 468
rect 1084 456 1090 468
rect 4709 459 4767 465
rect 4709 456 4721 459
rect 1084 428 4721 456
rect 1084 416 1090 428
rect 4709 425 4721 428
rect 4755 425 4767 459
rect 4816 456 4844 496
rect 4982 484 4988 536
rect 5040 524 5046 536
rect 5077 527 5135 533
rect 5077 524 5089 527
rect 5040 496 5089 524
rect 5040 484 5046 496
rect 5077 493 5089 496
rect 5123 493 5135 527
rect 5997 527 6055 533
rect 5997 524 6009 527
rect 5077 487 5135 493
rect 5184 496 6009 524
rect 5184 456 5212 496
rect 5997 493 6009 496
rect 6043 493 6055 527
rect 5997 487 6055 493
rect 6089 527 6147 533
rect 6089 493 6101 527
rect 6135 524 6147 527
rect 73246 524 73252 536
rect 6135 496 73252 524
rect 6135 493 6147 496
rect 6089 487 6147 493
rect 73246 484 73252 496
rect 73304 484 73310 536
rect 73341 527 73399 533
rect 73341 493 73353 527
rect 73387 524 73399 527
rect 93213 527 93271 533
rect 93213 524 93225 527
rect 73387 496 93225 524
rect 73387 493 73399 496
rect 73341 487 73399 493
rect 93213 493 93225 496
rect 93259 493 93271 527
rect 93320 524 93348 564
rect 93394 552 93400 604
rect 93452 592 93458 604
rect 93452 564 93497 592
rect 93452 552 93458 564
rect 93854 552 93860 604
rect 93912 592 93918 604
rect 94133 595 94191 601
rect 94133 592 94145 595
rect 93912 564 94145 592
rect 93912 552 93918 564
rect 94133 561 94145 564
rect 94179 561 94191 595
rect 98181 595 98239 601
rect 98181 592 98193 595
rect 94133 555 94191 561
rect 94240 564 98193 592
rect 94240 524 94268 564
rect 98181 561 98193 564
rect 98227 561 98239 595
rect 98181 555 98239 561
rect 98273 595 98331 601
rect 98273 561 98285 595
rect 98319 592 98331 595
rect 102321 595 102379 601
rect 102321 592 102333 595
rect 98319 564 102333 592
rect 98319 561 98331 564
rect 98273 555 98331 561
rect 102321 561 102333 564
rect 102367 561 102379 595
rect 102321 555 102379 561
rect 102413 595 102471 601
rect 102413 561 102425 595
rect 102459 592 102471 595
rect 103054 592 103060 604
rect 102459 564 103060 592
rect 102459 561 102471 564
rect 102413 555 102471 561
rect 103054 552 103060 564
rect 103112 552 103118 604
rect 103149 595 103207 601
rect 103149 561 103161 595
rect 103195 592 103207 595
rect 110877 595 110935 601
rect 110877 592 110889 595
rect 103195 564 110889 592
rect 103195 561 103207 564
rect 103149 555 103207 561
rect 110877 561 110889 564
rect 110923 561 110935 595
rect 110877 555 110935 561
rect 110969 595 111027 601
rect 110969 561 110981 595
rect 111015 592 111027 595
rect 111429 595 111487 601
rect 111429 592 111441 595
rect 111015 564 111441 592
rect 111015 561 111027 564
rect 110969 555 111027 561
rect 111429 561 111441 564
rect 111475 561 111487 595
rect 111536 592 111564 632
rect 111705 629 111717 663
rect 111751 660 111763 663
rect 112165 663 112223 669
rect 112165 660 112177 663
rect 111751 632 112177 660
rect 111751 629 111763 632
rect 111705 623 111763 629
rect 112165 629 112177 632
rect 112211 629 112223 663
rect 121457 663 121515 669
rect 121457 660 121469 663
rect 112165 623 112223 629
rect 112272 632 121469 660
rect 112272 592 112300 632
rect 121457 629 121469 632
rect 121503 629 121515 663
rect 121457 623 121515 629
rect 121549 663 121607 669
rect 121549 629 121561 663
rect 121595 660 121607 663
rect 122101 663 122159 669
rect 122101 660 122113 663
rect 121595 632 122113 660
rect 121595 629 121607 632
rect 121549 623 121607 629
rect 122101 629 122113 632
rect 122147 629 122159 663
rect 122101 623 122159 629
rect 122190 620 122196 672
rect 122248 660 122254 672
rect 124493 663 124551 669
rect 124493 660 124505 663
rect 122248 632 124505 660
rect 122248 620 122254 632
rect 124493 629 124505 632
rect 124539 629 124551 663
rect 124493 623 124551 629
rect 124677 663 124735 669
rect 124677 629 124689 663
rect 124723 660 124735 663
rect 149701 663 149759 669
rect 149701 660 149713 663
rect 124723 632 149713 660
rect 124723 629 124735 632
rect 124677 623 124735 629
rect 149701 629 149713 632
rect 149747 629 149759 663
rect 150069 663 150127 669
rect 150069 660 150081 663
rect 149701 623 149759 629
rect 149808 632 150081 660
rect 111536 564 112300 592
rect 112441 595 112499 601
rect 111429 555 111487 561
rect 112441 561 112453 595
rect 112487 592 112499 595
rect 149808 592 149836 632
rect 150069 629 150081 632
rect 150115 629 150127 663
rect 150250 660 150256 672
rect 150211 632 150256 660
rect 150069 623 150127 629
rect 150250 620 150256 632
rect 150308 620 150314 672
rect 153381 663 153439 669
rect 153381 660 153393 663
rect 150360 632 153393 660
rect 112487 564 149836 592
rect 149885 595 149943 601
rect 112487 561 112499 564
rect 112441 555 112499 561
rect 149885 561 149897 595
rect 149931 592 149943 595
rect 150360 592 150388 632
rect 153381 629 153393 632
rect 153427 629 153439 663
rect 153488 660 153516 700
rect 153562 688 153568 740
rect 153620 728 153626 740
rect 154669 731 154727 737
rect 154669 728 154681 731
rect 153620 700 154681 728
rect 153620 688 153626 700
rect 154669 697 154681 700
rect 154715 697 154727 731
rect 156598 728 156604 740
rect 156559 700 156604 728
rect 154669 691 154727 697
rect 156598 688 156604 700
rect 156656 688 156662 740
rect 156782 728 156788 740
rect 156743 700 156788 728
rect 156782 688 156788 700
rect 156840 688 156846 740
rect 156984 728 157012 836
rect 157076 796 157104 904
rect 157153 901 157165 935
rect 157199 932 157211 935
rect 158349 935 158407 941
rect 158349 932 158361 935
rect 157199 904 158361 932
rect 157199 901 157211 904
rect 157153 895 157211 901
rect 158349 901 158361 904
rect 158395 901 158407 935
rect 158349 895 158407 901
rect 159637 935 159695 941
rect 159637 901 159649 935
rect 159683 932 159695 935
rect 160833 935 160891 941
rect 160833 932 160845 935
rect 159683 904 160845 932
rect 159683 901 159695 904
rect 159637 895 159695 901
rect 160833 901 160845 904
rect 160879 901 160891 935
rect 160940 932 160968 972
rect 161124 972 179245 1000
rect 161124 932 161152 972
rect 179233 969 179245 972
rect 179279 969 179291 1003
rect 179233 963 179291 969
rect 179417 1003 179475 1009
rect 179417 969 179429 1003
rect 179463 1000 179475 1003
rect 218333 1003 218391 1009
rect 218333 1000 218345 1003
rect 179463 972 218345 1000
rect 179463 969 179475 972
rect 179417 963 179475 969
rect 218333 969 218345 972
rect 218379 969 218391 1003
rect 218333 963 218391 969
rect 218517 1003 218575 1009
rect 218517 969 218529 1003
rect 218563 1000 218575 1003
rect 241793 1003 241851 1009
rect 241793 1000 241805 1003
rect 218563 972 241805 1000
rect 218563 969 218575 972
rect 218517 963 218575 969
rect 241793 969 241805 972
rect 241839 969 241851 1003
rect 241793 963 241851 969
rect 241974 960 241980 1012
rect 242032 960 242038 1012
rect 242069 1003 242127 1009
rect 242069 969 242081 1003
rect 242115 1000 242127 1003
rect 296809 1003 296867 1009
rect 296809 1000 296821 1003
rect 242115 972 296821 1000
rect 242115 969 242127 972
rect 242069 963 242127 969
rect 296809 969 296821 972
rect 296855 969 296867 1003
rect 296809 963 296867 969
rect 296898 960 296904 1012
rect 296956 1000 296962 1012
rect 306837 1003 306895 1009
rect 306837 1000 306849 1003
rect 296956 972 306849 1000
rect 296956 960 296962 972
rect 306837 969 306849 972
rect 306883 969 306895 1003
rect 306837 963 306895 969
rect 306926 960 306932 1012
rect 306984 1000 306990 1012
rect 318610 1000 318616 1012
rect 306984 972 318616 1000
rect 306984 960 306990 972
rect 318610 960 318616 972
rect 318668 960 318674 1012
rect 318705 1003 318763 1009
rect 318705 969 318717 1003
rect 318751 1000 318763 1003
rect 319438 1000 319444 1012
rect 318751 972 319444 1000
rect 318751 969 318763 972
rect 318705 963 318763 969
rect 319438 960 319444 972
rect 319496 960 319502 1012
rect 319530 960 319536 1012
rect 319588 1000 319594 1012
rect 327718 1000 327724 1012
rect 319588 972 327724 1000
rect 319588 960 319594 972
rect 327718 960 327724 972
rect 327776 960 327782 1012
rect 327810 960 327816 1012
rect 327868 1000 327874 1012
rect 329558 1000 329564 1012
rect 327868 972 329564 1000
rect 327868 960 327874 972
rect 329558 960 329564 972
rect 329616 960 329622 1012
rect 331674 1000 331680 1012
rect 329668 972 331680 1000
rect 160940 904 161152 932
rect 161201 935 161259 941
rect 160833 895 160891 901
rect 161201 901 161213 935
rect 161247 932 161259 935
rect 162397 935 162455 941
rect 162397 932 162409 935
rect 161247 904 162409 932
rect 161247 901 161259 904
rect 161201 895 161259 901
rect 162397 901 162409 904
rect 162443 901 162455 935
rect 162397 895 162455 901
rect 162489 935 162547 941
rect 162489 901 162501 935
rect 162535 932 162547 935
rect 162578 932 162584 944
rect 162535 904 162584 932
rect 162535 901 162547 904
rect 162489 895 162547 901
rect 162578 892 162584 904
rect 162636 892 162642 944
rect 162673 935 162731 941
rect 162673 901 162685 935
rect 162719 932 162731 935
rect 163041 935 163099 941
rect 163041 932 163053 935
rect 162719 904 163053 932
rect 162719 901 162731 904
rect 162673 895 162731 901
rect 163041 901 163053 904
rect 163087 901 163099 935
rect 163041 895 163099 901
rect 163133 935 163191 941
rect 163133 901 163145 935
rect 163179 932 163191 935
rect 164329 935 164387 941
rect 164329 932 164341 935
rect 163179 904 164341 932
rect 163179 901 163191 904
rect 163133 895 163191 901
rect 164329 901 164341 904
rect 164375 901 164387 935
rect 179325 935 179383 941
rect 179325 932 179337 935
rect 164329 895 164387 901
rect 164436 904 179337 932
rect 157429 867 157487 873
rect 157429 833 157441 867
rect 157475 864 157487 867
rect 161017 867 161075 873
rect 161017 864 161029 867
rect 157475 836 161029 864
rect 157475 833 157487 836
rect 157429 827 157487 833
rect 161017 833 161029 836
rect 161063 833 161075 867
rect 161017 827 161075 833
rect 161293 867 161351 873
rect 161293 833 161305 867
rect 161339 864 161351 867
rect 164436 864 164464 904
rect 179325 901 179337 904
rect 179371 901 179383 935
rect 179325 895 179383 901
rect 179509 935 179567 941
rect 179509 901 179521 935
rect 179555 932 179567 935
rect 218057 935 218115 941
rect 218057 932 218069 935
rect 179555 904 218069 932
rect 179555 901 179567 904
rect 179509 895 179567 901
rect 218057 901 218069 904
rect 218103 901 218115 935
rect 218057 895 218115 901
rect 218425 935 218483 941
rect 218425 901 218437 935
rect 218471 932 218483 935
rect 241885 935 241943 941
rect 241885 932 241897 935
rect 218471 904 241897 932
rect 218471 901 218483 904
rect 218425 895 218483 901
rect 241885 901 241897 904
rect 241931 901 241943 935
rect 241885 895 241943 901
rect 161339 836 164464 864
rect 164513 867 164571 873
rect 161339 833 161351 836
rect 161293 827 161351 833
rect 164513 833 164525 867
rect 164559 864 164571 867
rect 165893 867 165951 873
rect 165893 864 165905 867
rect 164559 836 165905 864
rect 164559 833 164571 836
rect 164513 827 164571 833
rect 165893 833 165905 836
rect 165939 833 165951 867
rect 177574 864 177580 876
rect 165893 827 165951 833
rect 166000 836 175964 864
rect 157797 799 157855 805
rect 157797 796 157809 799
rect 157076 768 157809 796
rect 157797 765 157809 768
rect 157843 765 157855 799
rect 157797 759 157855 765
rect 157981 799 158039 805
rect 157981 765 157993 799
rect 158027 796 158039 799
rect 160557 799 160615 805
rect 160557 796 160569 799
rect 158027 768 160569 796
rect 158027 765 158039 768
rect 157981 759 158039 765
rect 160557 765 160569 768
rect 160603 765 160615 799
rect 160557 759 160615 765
rect 160830 756 160836 808
rect 160888 796 160894 808
rect 161109 799 161167 805
rect 161109 796 161121 799
rect 160888 768 161121 796
rect 160888 756 160894 768
rect 161109 765 161121 768
rect 161155 765 161167 799
rect 161109 759 161167 765
rect 161201 799 161259 805
rect 161201 765 161213 799
rect 161247 796 161259 799
rect 163041 799 163099 805
rect 163041 796 163053 799
rect 161247 768 163053 796
rect 161247 765 161259 768
rect 161201 759 161259 765
rect 163041 765 163053 768
rect 163087 765 163099 799
rect 166000 796 166028 836
rect 163041 759 163099 765
rect 163148 768 166028 796
rect 166077 799 166135 805
rect 157153 731 157211 737
rect 156984 700 157104 728
rect 154485 663 154543 669
rect 154485 660 154497 663
rect 153488 632 154497 660
rect 153381 623 153439 629
rect 154485 629 154497 632
rect 154531 629 154543 663
rect 154485 623 154543 629
rect 154577 663 154635 669
rect 154577 629 154589 663
rect 154623 660 154635 663
rect 156693 663 156751 669
rect 156693 660 156705 663
rect 154623 632 156705 660
rect 154623 629 154635 632
rect 154577 623 154635 629
rect 156693 629 156705 632
rect 156739 629 156751 663
rect 157076 660 157104 700
rect 157153 697 157165 731
rect 157199 728 157211 731
rect 159913 731 159971 737
rect 159913 728 159925 731
rect 157199 700 159925 728
rect 157199 697 157211 700
rect 157153 691 157211 697
rect 159913 697 159925 700
rect 159959 697 159971 731
rect 159913 691 159971 697
rect 160005 731 160063 737
rect 160005 697 160017 731
rect 160051 728 160063 731
rect 160649 731 160707 737
rect 160649 728 160661 731
rect 160051 700 160661 728
rect 160051 697 160063 700
rect 160005 691 160063 697
rect 160649 697 160661 700
rect 160695 697 160707 731
rect 160649 691 160707 697
rect 160738 688 160744 740
rect 160796 728 160802 740
rect 163148 728 163176 768
rect 166077 765 166089 799
rect 166123 796 166135 799
rect 169478 796 169484 808
rect 166123 768 169484 796
rect 166123 765 166135 768
rect 166077 759 166135 765
rect 169478 756 169484 768
rect 169536 756 169542 808
rect 175642 796 175648 808
rect 169588 768 175648 796
rect 160796 700 163176 728
rect 160796 688 160802 700
rect 163222 688 163228 740
rect 163280 728 163286 740
rect 163866 728 163872 740
rect 163280 700 163872 728
rect 163280 688 163286 700
rect 163866 688 163872 700
rect 163924 688 163930 740
rect 163958 688 163964 740
rect 164016 728 164022 740
rect 169113 731 169171 737
rect 164016 700 169064 728
rect 164016 688 164022 700
rect 157334 660 157340 672
rect 156693 623 156751 629
rect 156800 632 157012 660
rect 157076 632 157340 660
rect 149931 564 150388 592
rect 150437 595 150495 601
rect 149931 561 149943 564
rect 149885 555 149943 561
rect 150437 561 150449 595
rect 150483 592 150495 595
rect 151357 595 151415 601
rect 151357 592 151369 595
rect 150483 564 151369 592
rect 150483 561 150495 564
rect 150437 555 150495 561
rect 151357 561 151369 564
rect 151403 561 151415 595
rect 151357 555 151415 561
rect 151449 595 151507 601
rect 151449 561 151461 595
rect 151495 592 151507 595
rect 151495 564 156644 592
rect 151495 561 151507 564
rect 151449 555 151507 561
rect 93320 496 94268 524
rect 94317 527 94375 533
rect 93213 487 93271 493
rect 94317 493 94329 527
rect 94363 524 94375 527
rect 97353 527 97411 533
rect 94363 496 97304 524
rect 94363 493 94375 496
rect 94317 487 94375 493
rect 4816 428 5212 456
rect 5445 459 5503 465
rect 4709 419 4767 425
rect 5445 425 5457 459
rect 5491 456 5503 459
rect 10229 459 10287 465
rect 10229 456 10241 459
rect 5491 428 10241 456
rect 5491 425 5503 428
rect 5445 419 5503 425
rect 10229 425 10241 428
rect 10275 425 10287 459
rect 92566 456 92572 468
rect 10229 419 10287 425
rect 10336 428 74028 456
rect 1489 391 1547 397
rect 1489 357 1501 391
rect 1535 388 1547 391
rect 5353 391 5411 397
rect 5353 388 5365 391
rect 1535 360 5365 388
rect 1535 357 1547 360
rect 1489 351 1547 357
rect 5353 357 5365 360
rect 5399 357 5411 391
rect 5353 351 5411 357
rect 5721 391 5779 397
rect 5721 357 5733 391
rect 5767 357 5779 391
rect 5721 351 5779 357
rect 5813 391 5871 397
rect 5813 357 5825 391
rect 5859 388 5871 391
rect 10336 388 10364 428
rect 5859 360 10364 388
rect 10413 391 10471 397
rect 5859 357 5871 360
rect 5813 351 5871 357
rect 10413 357 10425 391
rect 10459 388 10471 391
rect 14277 391 14335 397
rect 14277 388 14289 391
rect 10459 360 14289 388
rect 10459 357 10471 360
rect 10413 351 10471 357
rect 14277 357 14289 360
rect 14323 357 14335 391
rect 14277 351 14335 357
rect 14461 391 14519 397
rect 14461 357 14473 391
rect 14507 388 14519 391
rect 38657 391 38715 397
rect 38657 388 38669 391
rect 14507 360 38669 388
rect 14507 357 14519 360
rect 14461 351 14519 357
rect 38657 357 38669 360
rect 38703 357 38715 391
rect 39209 391 39267 397
rect 39209 388 39221 391
rect 38657 351 38715 357
rect 38764 360 39221 388
rect 477 323 535 329
rect 477 289 489 323
rect 523 320 535 323
rect 5261 323 5319 329
rect 5261 320 5273 323
rect 523 292 5273 320
rect 523 289 535 292
rect 477 283 535 289
rect 5261 289 5273 292
rect 5307 289 5319 323
rect 5736 320 5764 351
rect 9677 323 9735 329
rect 9677 320 9689 323
rect 5736 292 9689 320
rect 5261 283 5319 289
rect 9677 289 9689 292
rect 9723 289 9735 323
rect 9677 283 9735 289
rect 9769 323 9827 329
rect 9769 289 9781 323
rect 9815 320 9827 323
rect 26789 323 26847 329
rect 26789 320 26801 323
rect 9815 292 26801 320
rect 9815 289 9827 292
rect 9769 283 9827 289
rect 26789 289 26801 292
rect 26835 289 26847 323
rect 26789 283 26847 289
rect 26878 280 26884 332
rect 26936 320 26942 332
rect 35158 320 35164 332
rect 26936 292 35164 320
rect 26936 280 26942 292
rect 35158 280 35164 292
rect 35216 280 35222 332
rect 35253 323 35311 329
rect 35253 289 35265 323
rect 35299 320 35311 323
rect 38764 320 38792 360
rect 39209 357 39221 360
rect 39255 357 39267 391
rect 39209 351 39267 357
rect 39301 391 39359 397
rect 39301 357 39313 391
rect 39347 388 39359 391
rect 73893 391 73951 397
rect 73893 388 73905 391
rect 39347 360 73905 388
rect 39347 357 39359 360
rect 39301 351 39359 357
rect 73893 357 73905 360
rect 73939 357 73951 391
rect 74000 388 74028 428
rect 74276 428 92572 456
rect 74276 388 74304 428
rect 92566 416 92572 428
rect 92624 416 92630 468
rect 92750 416 92756 468
rect 92808 456 92814 468
rect 95697 459 95755 465
rect 95697 456 95709 459
rect 92808 428 95709 456
rect 92808 416 92814 428
rect 95697 425 95709 428
rect 95743 425 95755 459
rect 95697 419 95755 425
rect 96709 459 96767 465
rect 96709 425 96721 459
rect 96755 456 96767 459
rect 97169 459 97227 465
rect 97169 456 97181 459
rect 96755 428 97181 456
rect 96755 425 96767 428
rect 96709 419 96767 425
rect 97169 425 97181 428
rect 97215 425 97227 459
rect 97276 456 97304 496
rect 97353 493 97365 527
rect 97399 524 97411 527
rect 100297 527 100355 533
rect 100297 524 100309 527
rect 97399 496 100309 524
rect 97399 493 97411 496
rect 97353 487 97411 493
rect 100297 493 100309 496
rect 100343 493 100355 527
rect 100297 487 100355 493
rect 100665 527 100723 533
rect 100665 493 100677 527
rect 100711 524 100723 527
rect 111981 527 112039 533
rect 111981 524 111993 527
rect 100711 496 111993 524
rect 100711 493 100723 496
rect 100665 487 100723 493
rect 111981 493 111993 496
rect 112027 493 112039 527
rect 111981 487 112039 493
rect 112165 527 112223 533
rect 112165 493 112177 527
rect 112211 524 112223 527
rect 156509 527 156567 533
rect 156509 524 156521 527
rect 112211 496 156521 524
rect 112211 493 112223 496
rect 112165 487 112223 493
rect 156509 493 156521 496
rect 156555 493 156567 527
rect 156616 524 156644 564
rect 156800 524 156828 632
rect 156984 592 157012 632
rect 157334 620 157340 632
rect 157392 620 157398 672
rect 157610 660 157616 672
rect 157571 632 157616 660
rect 157610 620 157616 632
rect 157668 620 157674 672
rect 157794 620 157800 672
rect 157852 660 157858 672
rect 158993 663 159051 669
rect 158993 660 159005 663
rect 157852 632 159005 660
rect 157852 620 157858 632
rect 158993 629 159005 632
rect 159039 629 159051 663
rect 158993 623 159051 629
rect 159269 663 159327 669
rect 159269 629 159281 663
rect 159315 660 159327 663
rect 159450 660 159456 672
rect 159315 632 159456 660
rect 159315 629 159327 632
rect 159269 623 159327 629
rect 159450 620 159456 632
rect 159508 620 159514 672
rect 159729 663 159787 669
rect 159729 629 159741 663
rect 159775 660 159787 663
rect 160922 660 160928 672
rect 159775 632 160928 660
rect 159775 629 159787 632
rect 159729 623 159787 629
rect 160922 620 160928 632
rect 160980 620 160986 672
rect 161017 663 161075 669
rect 161017 629 161029 663
rect 161063 660 161075 663
rect 162213 663 162271 669
rect 162213 660 162225 663
rect 161063 632 162225 660
rect 161063 629 161075 632
rect 161017 623 161075 629
rect 162213 629 162225 632
rect 162259 629 162271 663
rect 162213 623 162271 629
rect 162305 663 162363 669
rect 162305 629 162317 663
rect 162351 660 162363 663
rect 163041 663 163099 669
rect 163041 660 163053 663
rect 162351 632 163053 660
rect 162351 629 162363 632
rect 162305 623 162363 629
rect 163041 629 163053 632
rect 163087 629 163099 663
rect 163041 623 163099 629
rect 163130 620 163136 672
rect 163188 660 163194 672
rect 166077 663 166135 669
rect 166077 660 166089 663
rect 163188 632 166089 660
rect 163188 620 163194 632
rect 166077 629 166089 632
rect 166123 629 166135 663
rect 166077 623 166135 629
rect 166166 620 166172 672
rect 166224 660 166230 672
rect 166261 663 166319 669
rect 166261 660 166273 663
rect 166224 632 166273 660
rect 166224 620 166230 632
rect 166261 629 166273 632
rect 166307 629 166319 663
rect 166261 623 166319 629
rect 166626 620 166632 672
rect 166684 660 166690 672
rect 167089 663 167147 669
rect 167089 660 167101 663
rect 166684 632 167101 660
rect 166684 620 166690 632
rect 167089 629 167101 632
rect 167135 629 167147 663
rect 167089 623 167147 629
rect 167181 663 167239 669
rect 167181 629 167193 663
rect 167227 660 167239 663
rect 168929 663 168987 669
rect 168929 660 168941 663
rect 167227 632 168941 660
rect 167227 629 167239 632
rect 167181 623 167239 629
rect 168929 629 168941 632
rect 168975 629 168987 663
rect 169036 660 169064 700
rect 169113 697 169125 731
rect 169159 728 169171 731
rect 169588 728 169616 768
rect 175642 756 175648 768
rect 175700 756 175706 808
rect 175936 796 175964 836
rect 176396 836 177580 864
rect 176396 796 176424 836
rect 177574 824 177580 836
rect 177632 824 177638 876
rect 177758 824 177764 876
rect 177816 864 177822 876
rect 179598 864 179604 876
rect 177816 836 179604 864
rect 177816 824 177822 836
rect 179598 824 179604 836
rect 179656 824 179662 876
rect 179690 824 179696 876
rect 179748 864 179754 876
rect 180061 867 180119 873
rect 180061 864 180073 867
rect 179748 836 180073 864
rect 179748 824 179754 836
rect 180061 833 180073 836
rect 180107 833 180119 867
rect 180061 827 180119 833
rect 180245 867 180303 873
rect 180245 833 180257 867
rect 180291 864 180303 867
rect 180610 864 180616 876
rect 180291 836 180616 864
rect 180291 833 180303 836
rect 180245 827 180303 833
rect 180610 824 180616 836
rect 180668 824 180674 876
rect 180702 824 180708 876
rect 180760 864 180766 876
rect 239033 867 239091 873
rect 239033 864 239045 867
rect 180760 836 239045 864
rect 180760 824 180766 836
rect 239033 833 239045 836
rect 239079 833 239091 867
rect 239033 827 239091 833
rect 239401 867 239459 873
rect 239401 833 239413 867
rect 239447 864 239459 867
rect 241701 867 241759 873
rect 241701 864 241713 867
rect 239447 836 241713 864
rect 239447 833 239459 836
rect 239401 827 239459 833
rect 241701 833 241713 836
rect 241747 833 241759 867
rect 241992 864 242020 960
rect 242161 935 242219 941
rect 242161 901 242173 935
rect 242207 932 242219 935
rect 317601 935 317659 941
rect 317601 932 317613 935
rect 242207 904 317613 932
rect 242207 901 242219 904
rect 242161 895 242219 901
rect 317601 901 317613 904
rect 317647 901 317659 935
rect 317601 895 317659 901
rect 317690 892 317696 944
rect 317748 932 317754 944
rect 323397 935 323455 941
rect 323397 932 323409 935
rect 317748 904 323409 932
rect 317748 892 317754 904
rect 323397 901 323409 904
rect 323443 901 323455 935
rect 323397 895 323455 901
rect 323489 935 323547 941
rect 323489 901 323501 935
rect 323535 932 323547 935
rect 328730 932 328736 944
rect 323535 904 328736 932
rect 323535 901 323547 904
rect 323489 895 323547 901
rect 328730 892 328736 904
rect 328788 892 328794 944
rect 328822 892 328828 944
rect 328880 932 328886 944
rect 329668 932 329696 972
rect 331674 960 331680 972
rect 331732 960 331738 1012
rect 331766 960 331772 1012
rect 331824 1000 331830 1012
rect 335722 1000 335728 1012
rect 331824 972 335728 1000
rect 331824 960 331830 972
rect 335722 960 335728 972
rect 335780 960 335786 1012
rect 335814 960 335820 1012
rect 335872 1000 335878 1012
rect 337933 1003 337991 1009
rect 337933 1000 337945 1003
rect 335872 972 337945 1000
rect 335872 960 335878 972
rect 337933 969 337945 972
rect 337979 969 337991 1003
rect 337933 963 337991 969
rect 338761 1003 338819 1009
rect 338761 969 338773 1003
rect 338807 1000 338819 1003
rect 342272 1000 342300 1040
rect 345385 1037 345397 1040
rect 345431 1037 345443 1071
rect 352190 1068 352196 1080
rect 345385 1031 345443 1037
rect 345676 1040 352196 1068
rect 338807 972 342300 1000
rect 338807 969 338819 972
rect 338761 963 338819 969
rect 328880 904 329696 932
rect 328880 892 328886 904
rect 329742 892 329748 944
rect 329800 932 329806 944
rect 343082 932 343088 944
rect 329800 904 343088 932
rect 329800 892 329806 904
rect 343082 892 343088 904
rect 343140 892 343146 944
rect 343177 935 343235 941
rect 343177 901 343189 935
rect 343223 932 343235 935
rect 345676 932 345704 1040
rect 352190 1028 352196 1040
rect 352248 1028 352254 1080
rect 352653 1071 352711 1077
rect 352653 1037 352665 1071
rect 352699 1068 352711 1071
rect 357069 1071 357127 1077
rect 357069 1068 357081 1071
rect 352699 1040 357081 1068
rect 352699 1037 352711 1040
rect 352653 1031 352711 1037
rect 357069 1037 357081 1040
rect 357115 1037 357127 1071
rect 357069 1031 357127 1037
rect 357897 1071 357955 1077
rect 357897 1037 357909 1071
rect 357943 1068 357955 1071
rect 364153 1071 364211 1077
rect 364153 1068 364165 1071
rect 357943 1040 364165 1068
rect 357943 1037 357955 1040
rect 357897 1031 357955 1037
rect 364153 1037 364165 1040
rect 364199 1037 364211 1071
rect 364153 1031 364211 1037
rect 364245 1071 364303 1077
rect 364245 1037 364257 1071
rect 364291 1068 364303 1071
rect 372798 1068 372804 1080
rect 364291 1040 372804 1068
rect 364291 1037 364303 1040
rect 364245 1031 364303 1037
rect 372798 1028 372804 1040
rect 372856 1028 372862 1080
rect 376021 1071 376079 1077
rect 376021 1068 376033 1071
rect 372908 1040 376033 1068
rect 345753 1003 345811 1009
rect 345753 969 345765 1003
rect 345799 1000 345811 1003
rect 372709 1003 372767 1009
rect 372709 1000 372721 1003
rect 345799 972 372721 1000
rect 345799 969 345811 972
rect 345753 963 345811 969
rect 372709 969 372721 972
rect 372755 969 372767 1003
rect 372908 1000 372936 1040
rect 376021 1037 376033 1040
rect 376067 1037 376079 1071
rect 376021 1031 376079 1037
rect 378413 1071 378471 1077
rect 378413 1037 378425 1071
rect 378459 1068 378471 1071
rect 393593 1071 393651 1077
rect 393593 1068 393605 1071
rect 378459 1040 393605 1068
rect 378459 1037 378471 1040
rect 378413 1031 378471 1037
rect 393593 1037 393605 1040
rect 393639 1037 393651 1071
rect 393593 1031 393651 1037
rect 413646 1028 413652 1080
rect 413704 1068 413710 1080
rect 453298 1068 453304 1080
rect 413704 1040 453304 1068
rect 413704 1028 413710 1040
rect 453298 1028 453304 1040
rect 453356 1028 453362 1080
rect 473357 1071 473415 1077
rect 473357 1037 473369 1071
rect 473403 1068 473415 1071
rect 480162 1068 480168 1080
rect 473403 1040 480168 1068
rect 473403 1037 473415 1040
rect 473357 1031 473415 1037
rect 480162 1028 480168 1040
rect 480220 1028 480226 1080
rect 494057 1071 494115 1077
rect 494057 1037 494069 1071
rect 494103 1068 494115 1071
rect 494256 1068 494284 1108
rect 521657 1105 521669 1108
rect 521703 1105 521715 1139
rect 521657 1099 521715 1105
rect 521749 1139 521807 1145
rect 521749 1105 521761 1139
rect 521795 1136 521807 1139
rect 538217 1139 538275 1145
rect 538217 1136 538229 1139
rect 521795 1108 538229 1136
rect 521795 1105 521807 1108
rect 521749 1099 521807 1105
rect 538217 1105 538229 1108
rect 538263 1105 538275 1139
rect 538217 1099 538275 1105
rect 543093 1139 543151 1145
rect 543093 1105 543105 1139
rect 543139 1136 543151 1139
rect 549257 1139 549315 1145
rect 549257 1136 549269 1139
rect 543139 1108 549269 1136
rect 543139 1105 543151 1108
rect 543093 1099 543151 1105
rect 549257 1105 549269 1108
rect 549303 1105 549315 1139
rect 549257 1099 549315 1105
rect 549349 1139 549407 1145
rect 549349 1105 549361 1139
rect 549395 1136 549407 1139
rect 559469 1139 559527 1145
rect 559469 1136 559481 1139
rect 549395 1108 559481 1136
rect 549395 1105 549407 1108
rect 549349 1099 549407 1105
rect 559469 1105 559481 1108
rect 559515 1105 559527 1139
rect 559469 1099 559527 1105
rect 494103 1040 494284 1068
rect 494103 1037 494115 1040
rect 494057 1031 494115 1037
rect 501322 1028 501328 1080
rect 501380 1068 501386 1080
rect 512638 1068 512644 1080
rect 501380 1040 512644 1068
rect 501380 1028 501386 1040
rect 512638 1028 512644 1040
rect 512696 1028 512702 1080
rect 516781 1071 516839 1077
rect 516781 1037 516793 1071
rect 516827 1068 516839 1071
rect 535362 1068 535368 1080
rect 516827 1040 535368 1068
rect 516827 1037 516839 1040
rect 516781 1031 516839 1037
rect 535362 1028 535368 1040
rect 535420 1028 535426 1080
rect 372709 963 372767 969
rect 372816 972 372936 1000
rect 373077 1003 373135 1009
rect 343223 904 345704 932
rect 348237 935 348295 941
rect 343223 901 343235 904
rect 343177 895 343235 901
rect 348237 901 348249 935
rect 348283 932 348295 935
rect 349433 935 349491 941
rect 349433 932 349445 935
rect 348283 904 349445 932
rect 348283 901 348295 904
rect 348237 895 348295 901
rect 349433 901 349445 904
rect 349479 901 349491 935
rect 349433 895 349491 901
rect 349522 892 349528 944
rect 349580 932 349586 944
rect 356149 935 356207 941
rect 356149 932 356161 935
rect 349580 904 356161 932
rect 349580 892 349586 904
rect 356149 901 356161 904
rect 356195 901 356207 935
rect 356149 895 356207 901
rect 356238 892 356244 944
rect 356296 932 356302 944
rect 364245 935 364303 941
rect 364245 932 364257 935
rect 356296 904 364257 932
rect 356296 892 356302 904
rect 364245 901 364257 904
rect 364291 901 364303 935
rect 364245 895 364303 901
rect 364337 935 364395 941
rect 364337 901 364349 935
rect 364383 932 364395 935
rect 368477 935 368535 941
rect 368477 932 368489 935
rect 364383 904 368489 932
rect 364383 901 364395 904
rect 364337 895 364395 901
rect 368477 901 368489 904
rect 368523 901 368535 935
rect 372816 932 372844 972
rect 373077 969 373089 1003
rect 373123 1000 373135 1003
rect 568206 1000 568212 1012
rect 373123 972 568212 1000
rect 373123 969 373135 972
rect 373077 963 373135 969
rect 568206 960 568212 972
rect 568264 960 568270 1012
rect 373902 932 373908 944
rect 368477 895 368535 901
rect 372724 904 372844 932
rect 372908 904 373908 932
rect 241701 827 241759 833
rect 241808 836 242020 864
rect 242069 867 242127 873
rect 183649 799 183707 805
rect 183649 796 183661 799
rect 175936 768 176424 796
rect 176488 768 183661 796
rect 169159 700 169616 728
rect 169159 697 169171 700
rect 169113 691 169171 697
rect 169662 688 169668 740
rect 169720 728 169726 740
rect 169941 731 169999 737
rect 169941 728 169953 731
rect 169720 700 169953 728
rect 169720 688 169726 700
rect 169941 697 169953 700
rect 169987 697 169999 731
rect 169941 691 169999 697
rect 170033 731 170091 737
rect 170033 697 170045 731
rect 170079 697 170091 731
rect 175918 728 175924 740
rect 170033 691 170091 697
rect 170232 700 175924 728
rect 170048 660 170076 691
rect 170232 669 170260 700
rect 175918 688 175924 700
rect 175976 688 175982 740
rect 176010 688 176016 740
rect 176068 728 176074 740
rect 176488 728 176516 768
rect 183649 765 183661 768
rect 183695 765 183707 799
rect 183649 759 183707 765
rect 183738 756 183744 808
rect 183796 796 183802 808
rect 190181 799 190239 805
rect 190181 796 190193 799
rect 183796 768 190193 796
rect 183796 756 183802 768
rect 190181 765 190193 768
rect 190227 765 190239 799
rect 190181 759 190239 765
rect 190273 799 190331 805
rect 190273 765 190285 799
rect 190319 796 190331 799
rect 208029 799 208087 805
rect 208029 796 208041 799
rect 190319 768 208041 796
rect 190319 765 190331 768
rect 190273 759 190331 765
rect 208029 765 208041 768
rect 208075 765 208087 799
rect 208029 759 208087 765
rect 208210 756 208216 808
rect 208268 796 208274 808
rect 213733 799 213791 805
rect 213733 796 213745 799
rect 208268 768 213745 796
rect 208268 756 208274 768
rect 213733 765 213745 768
rect 213779 765 213791 799
rect 213733 759 213791 765
rect 213822 756 213828 808
rect 213880 796 213886 808
rect 219342 796 219348 808
rect 213880 768 219348 796
rect 213880 756 213886 768
rect 219342 756 219348 768
rect 219400 756 219406 808
rect 219434 756 219440 808
rect 219492 796 219498 808
rect 223853 799 223911 805
rect 223853 796 223865 799
rect 219492 768 223865 796
rect 219492 756 219498 768
rect 223853 765 223865 768
rect 223899 765 223911 799
rect 223853 759 223911 765
rect 224221 799 224279 805
rect 224221 765 224233 799
rect 224267 796 224279 799
rect 231949 799 232007 805
rect 231949 796 231961 799
rect 224267 768 231961 796
rect 224267 765 224279 768
rect 224221 759 224279 765
rect 231949 765 231961 768
rect 231995 765 232007 799
rect 231949 759 232007 765
rect 232041 799 232099 805
rect 232041 765 232053 799
rect 232087 796 232099 799
rect 232869 799 232927 805
rect 232869 796 232881 799
rect 232087 768 232881 796
rect 232087 765 232099 768
rect 232041 759 232099 765
rect 232869 765 232881 768
rect 232915 765 232927 799
rect 232869 759 232927 765
rect 232958 756 232964 808
rect 233016 796 233022 808
rect 233421 799 233479 805
rect 233016 768 233372 796
rect 233016 756 233022 768
rect 176068 700 176516 728
rect 176565 731 176623 737
rect 176068 688 176074 700
rect 176565 697 176577 731
rect 176611 728 176623 731
rect 177301 731 177359 737
rect 177301 728 177313 731
rect 176611 700 177313 728
rect 176611 697 176623 700
rect 176565 691 176623 697
rect 177301 697 177313 700
rect 177347 697 177359 731
rect 177301 691 177359 697
rect 178310 688 178316 740
rect 178368 728 178374 740
rect 180150 728 180156 740
rect 178368 700 180156 728
rect 178368 688 178374 700
rect 180150 688 180156 700
rect 180208 688 180214 740
rect 180242 688 180248 740
rect 180300 728 180306 740
rect 183925 731 183983 737
rect 183925 728 183937 731
rect 180300 700 183937 728
rect 180300 688 180306 700
rect 183925 697 183937 700
rect 183971 697 183983 731
rect 183925 691 183983 697
rect 184014 688 184020 740
rect 184072 728 184078 740
rect 204257 731 204315 737
rect 204257 728 204269 731
rect 184072 700 204269 728
rect 184072 688 184078 700
rect 204257 697 204269 700
rect 204303 697 204315 731
rect 204257 691 204315 697
rect 204533 731 204591 737
rect 204533 697 204545 731
rect 204579 728 204591 731
rect 208121 731 208179 737
rect 208121 728 208133 731
rect 204579 700 208133 728
rect 204579 697 204591 700
rect 204533 691 204591 697
rect 208121 697 208133 700
rect 208167 697 208179 731
rect 208121 691 208179 697
rect 208765 731 208823 737
rect 208765 697 208777 731
rect 208811 728 208823 731
rect 213917 731 213975 737
rect 213917 728 213929 731
rect 208811 700 213929 728
rect 208811 697 208823 700
rect 208765 691 208823 697
rect 213917 697 213929 700
rect 213963 697 213975 731
rect 213917 691 213975 697
rect 214285 731 214343 737
rect 214285 697 214297 731
rect 214331 728 214343 731
rect 221366 728 221372 740
rect 214331 700 221372 728
rect 214331 697 214343 700
rect 214285 691 214343 697
rect 221366 688 221372 700
rect 221424 688 221430 740
rect 221461 731 221519 737
rect 221461 697 221473 731
rect 221507 728 221519 731
rect 225049 731 225107 737
rect 225049 728 225061 731
rect 221507 700 225061 728
rect 221507 697 221519 700
rect 221461 691 221519 697
rect 225049 697 225061 700
rect 225095 697 225107 731
rect 225049 691 225107 697
rect 225141 731 225199 737
rect 225141 697 225153 731
rect 225187 728 225199 731
rect 231765 731 231823 737
rect 225187 700 231624 728
rect 225187 697 225199 700
rect 225141 691 225199 697
rect 169036 632 170076 660
rect 170217 663 170275 669
rect 168929 623 168987 629
rect 170217 629 170229 663
rect 170263 629 170275 663
rect 170217 623 170275 629
rect 170309 663 170367 669
rect 170309 629 170321 663
rect 170355 660 170367 663
rect 176102 660 176108 672
rect 170355 632 176108 660
rect 170355 629 170367 632
rect 170309 623 170367 629
rect 176102 620 176108 632
rect 176160 620 176166 672
rect 176197 663 176255 669
rect 176197 629 176209 663
rect 176243 660 176255 663
rect 176243 632 176608 660
rect 176243 629 176255 632
rect 176197 623 176255 629
rect 175645 595 175703 601
rect 175645 592 175657 595
rect 156984 564 175657 592
rect 175645 561 175657 564
rect 175691 561 175703 595
rect 175918 592 175924 604
rect 175879 564 175924 592
rect 175645 555 175703 561
rect 175918 552 175924 564
rect 175976 552 175982 604
rect 176381 595 176439 601
rect 176381 592 176393 595
rect 176028 564 176393 592
rect 156616 496 156828 524
rect 156969 527 157027 533
rect 156509 487 156567 493
rect 156969 493 156981 527
rect 157015 524 157027 527
rect 175734 524 175740 536
rect 157015 496 175740 524
rect 157015 493 157027 496
rect 156969 487 157027 493
rect 175734 484 175740 496
rect 175792 484 175798 536
rect 175829 527 175887 533
rect 175829 493 175841 527
rect 175875 524 175887 527
rect 176028 524 176056 564
rect 176381 561 176393 564
rect 176427 561 176439 595
rect 176580 592 176608 632
rect 176654 620 176660 672
rect 176712 660 176718 672
rect 177025 663 177083 669
rect 177025 660 177037 663
rect 176712 632 177037 660
rect 176712 620 176718 632
rect 177025 629 177037 632
rect 177071 629 177083 663
rect 177025 623 177083 629
rect 177114 620 177120 672
rect 177172 660 177178 672
rect 177393 663 177451 669
rect 177393 660 177405 663
rect 177172 632 177405 660
rect 177172 620 177178 632
rect 177393 629 177405 632
rect 177439 629 177451 663
rect 177393 623 177451 629
rect 177577 663 177635 669
rect 177577 629 177589 663
rect 177623 660 177635 663
rect 177942 660 177948 672
rect 177623 632 177948 660
rect 177623 629 177635 632
rect 177577 623 177635 629
rect 177942 620 177948 632
rect 178000 620 178006 672
rect 178037 663 178095 669
rect 178037 629 178049 663
rect 178083 660 178095 663
rect 183465 663 183523 669
rect 183465 660 183477 663
rect 178083 632 183477 660
rect 178083 629 178095 632
rect 178037 623 178095 629
rect 183465 629 183477 632
rect 183511 629 183523 663
rect 183465 623 183523 629
rect 183554 620 183560 672
rect 183612 660 183618 672
rect 183741 663 183799 669
rect 183741 660 183753 663
rect 183612 632 183753 660
rect 183612 620 183618 632
rect 183741 629 183753 632
rect 183787 629 183799 663
rect 196989 663 197047 669
rect 196989 660 197001 663
rect 183741 623 183799 629
rect 183848 632 197001 660
rect 183848 601 183876 632
rect 196989 629 197001 632
rect 197035 629 197047 663
rect 196989 623 197047 629
rect 197081 663 197139 669
rect 197081 629 197093 663
rect 197127 660 197139 663
rect 199013 663 199071 669
rect 199013 660 199025 663
rect 197127 632 199025 660
rect 197127 629 197139 632
rect 197081 623 197139 629
rect 199013 629 199025 632
rect 199059 629 199071 663
rect 199013 623 199071 629
rect 199105 663 199163 669
rect 199105 629 199117 663
rect 199151 660 199163 663
rect 204346 660 204352 672
rect 199151 632 204352 660
rect 199151 629 199163 632
rect 199105 623 199163 629
rect 204346 620 204352 632
rect 204404 620 204410 672
rect 204441 663 204499 669
rect 204441 629 204453 663
rect 204487 660 204499 663
rect 207750 660 207756 672
rect 204487 632 207756 660
rect 204487 629 204499 632
rect 204441 623 204499 629
rect 207750 620 207756 632
rect 207808 620 207814 672
rect 207842 620 207848 672
rect 207900 660 207906 672
rect 212537 663 212595 669
rect 212537 660 212549 663
rect 207900 632 212549 660
rect 207900 620 207906 632
rect 212537 629 212549 632
rect 212583 629 212595 663
rect 212537 623 212595 629
rect 212721 663 212779 669
rect 212721 629 212733 663
rect 212767 660 212779 663
rect 214009 663 214067 669
rect 214009 660 214021 663
rect 212767 632 214021 660
rect 212767 629 212779 632
rect 212721 623 212779 629
rect 214009 629 214021 632
rect 214055 629 214067 663
rect 214009 623 214067 629
rect 214098 620 214104 672
rect 214156 660 214162 672
rect 214929 663 214987 669
rect 214929 660 214941 663
rect 214156 632 214941 660
rect 214156 620 214162 632
rect 214929 629 214941 632
rect 214975 629 214987 663
rect 214929 623 214987 629
rect 215018 620 215024 672
rect 215076 660 215082 672
rect 217594 660 217600 672
rect 215076 632 217600 660
rect 215076 620 215082 632
rect 217594 620 217600 632
rect 217652 620 217658 672
rect 217689 663 217747 669
rect 217689 629 217701 663
rect 217735 660 217747 663
rect 219434 660 219440 672
rect 217735 632 219440 660
rect 217735 629 217747 632
rect 217689 623 217747 629
rect 219434 620 219440 632
rect 219492 620 219498 672
rect 219618 620 219624 672
rect 219676 660 219682 672
rect 221001 663 221059 669
rect 221001 660 221013 663
rect 219676 632 221013 660
rect 219676 620 219682 632
rect 221001 629 221013 632
rect 221047 629 221059 663
rect 221001 623 221059 629
rect 221090 620 221096 672
rect 221148 660 221154 672
rect 224129 663 224187 669
rect 224129 660 224141 663
rect 221148 632 224141 660
rect 221148 620 221154 632
rect 224129 629 224141 632
rect 224175 629 224187 663
rect 224129 623 224187 629
rect 224218 620 224224 672
rect 224276 660 224282 672
rect 224313 663 224371 669
rect 224313 660 224325 663
rect 224276 632 224325 660
rect 224276 620 224282 632
rect 224313 629 224325 632
rect 224359 629 224371 663
rect 224313 623 224371 629
rect 224402 620 224408 672
rect 224460 660 224466 672
rect 224460 632 224505 660
rect 224460 620 224466 632
rect 224586 620 224592 672
rect 224644 660 224650 672
rect 225322 660 225328 672
rect 224644 632 225328 660
rect 224644 620 224650 632
rect 225322 620 225328 632
rect 225380 620 225386 672
rect 225417 663 225475 669
rect 225417 629 225429 663
rect 225463 660 225475 663
rect 231486 660 231492 672
rect 225463 632 231492 660
rect 225463 629 225475 632
rect 225417 623 225475 629
rect 231486 620 231492 632
rect 231544 620 231550 672
rect 231596 669 231624 700
rect 231765 697 231777 731
rect 231811 728 231823 731
rect 233344 728 233372 768
rect 233421 765 233433 799
rect 233467 796 233479 799
rect 238389 799 238447 805
rect 238389 796 238401 799
rect 233467 768 238401 796
rect 233467 765 233479 768
rect 233421 759 233479 765
rect 238389 765 238401 768
rect 238435 765 238447 799
rect 238389 759 238447 765
rect 238478 756 238484 808
rect 238536 796 238542 808
rect 238757 799 238815 805
rect 238757 796 238769 799
rect 238536 768 238769 796
rect 238536 756 238542 768
rect 238757 765 238769 768
rect 238803 765 238815 799
rect 238757 759 238815 765
rect 239214 756 239220 808
rect 239272 796 239278 808
rect 241808 796 241836 836
rect 242069 833 242081 867
rect 242115 864 242127 867
rect 286137 867 286195 873
rect 286137 864 286149 867
rect 242115 836 286149 864
rect 242115 833 242127 836
rect 242069 827 242127 833
rect 286137 833 286149 836
rect 286183 833 286195 867
rect 286137 827 286195 833
rect 286226 824 286232 876
rect 286284 864 286290 876
rect 287425 867 287483 873
rect 287425 864 287437 867
rect 286284 836 287437 864
rect 286284 824 286290 836
rect 287425 833 287437 836
rect 287471 833 287483 867
rect 287425 827 287483 833
rect 287514 824 287520 876
rect 287572 864 287578 876
rect 289630 864 289636 876
rect 287572 836 289636 864
rect 287572 824 287578 836
rect 289630 824 289636 836
rect 289688 824 289694 876
rect 289725 867 289783 873
rect 289725 833 289737 867
rect 289771 864 289783 867
rect 293770 864 293776 876
rect 289771 836 293776 864
rect 289771 833 289783 836
rect 289725 827 289783 833
rect 293770 824 293776 836
rect 293828 824 293834 876
rect 293865 867 293923 873
rect 293865 833 293877 867
rect 293911 864 293923 867
rect 306742 864 306748 876
rect 293911 836 306748 864
rect 293911 833 293923 836
rect 293865 827 293923 833
rect 306742 824 306748 836
rect 306800 824 306806 876
rect 306837 867 306895 873
rect 306837 833 306849 867
rect 306883 864 306895 867
rect 309962 864 309968 876
rect 306883 836 309968 864
rect 306883 833 306895 836
rect 306837 827 306895 833
rect 309962 824 309968 836
rect 310020 824 310026 876
rect 310054 824 310060 876
rect 310112 864 310118 876
rect 319625 867 319683 873
rect 310112 836 319576 864
rect 310112 824 310118 836
rect 239272 768 241836 796
rect 241885 799 241943 805
rect 239272 756 239278 768
rect 241885 765 241897 799
rect 241931 796 241943 799
rect 314657 799 314715 805
rect 314657 796 314669 799
rect 241931 768 314669 796
rect 241931 765 241943 768
rect 241885 759 241943 765
rect 314657 765 314669 768
rect 314703 765 314715 799
rect 314657 759 314715 765
rect 314749 799 314807 805
rect 314749 765 314761 799
rect 314795 796 314807 799
rect 317509 799 317567 805
rect 317509 796 317521 799
rect 314795 768 317521 796
rect 314795 765 314807 768
rect 314749 759 314807 765
rect 317509 765 317521 768
rect 317555 765 317567 799
rect 317509 759 317567 765
rect 317601 799 317659 805
rect 317601 765 317613 799
rect 317647 796 317659 799
rect 319441 799 319499 805
rect 319441 796 319453 799
rect 317647 768 319453 796
rect 317647 765 317659 768
rect 317601 759 317659 765
rect 319441 765 319453 768
rect 319487 765 319499 799
rect 319441 759 319499 765
rect 261297 731 261355 737
rect 261297 728 261309 731
rect 231811 700 233280 728
rect 233344 700 261309 728
rect 231811 697 231823 700
rect 231765 691 231823 697
rect 231581 663 231639 669
rect 231581 629 231593 663
rect 231627 629 231639 663
rect 231581 623 231639 629
rect 231670 620 231676 672
rect 231728 660 231734 672
rect 233142 660 233148 672
rect 231728 632 233148 660
rect 231728 620 231734 632
rect 233142 620 233148 632
rect 233200 620 233206 672
rect 233252 660 233280 700
rect 261297 697 261309 700
rect 261343 697 261355 731
rect 261297 691 261355 697
rect 261496 700 271092 728
rect 251910 660 251916 672
rect 233252 632 251916 660
rect 251910 620 251916 632
rect 251968 620 251974 672
rect 252002 620 252008 672
rect 252060 660 252066 672
rect 252557 663 252615 669
rect 252557 660 252569 663
rect 252060 632 252569 660
rect 252060 620 252066 632
rect 252557 629 252569 632
rect 252603 629 252615 663
rect 252557 623 252615 629
rect 252830 620 252836 672
rect 252888 660 252894 672
rect 259270 660 259276 672
rect 252888 632 259276 660
rect 252888 620 252894 632
rect 259270 620 259276 632
rect 259328 620 259334 672
rect 259365 663 259423 669
rect 259365 629 259377 663
rect 259411 660 259423 663
rect 261496 660 261524 700
rect 259411 632 261524 660
rect 259411 629 259423 632
rect 259365 623 259423 629
rect 261570 620 261576 672
rect 261628 660 261634 672
rect 266998 660 267004 672
rect 261628 632 267004 660
rect 261628 620 261634 632
rect 266998 620 267004 632
rect 267056 620 267062 672
rect 267093 663 267151 669
rect 267093 629 267105 663
rect 267139 660 267151 663
rect 267182 660 267188 672
rect 267139 632 267188 660
rect 267139 629 267151 632
rect 267093 623 267151 629
rect 267182 620 267188 632
rect 267240 620 267246 672
rect 267277 663 267335 669
rect 267277 629 267289 663
rect 267323 660 267335 663
rect 270954 660 270960 672
rect 267323 632 270960 660
rect 267323 629 267335 632
rect 267277 623 267335 629
rect 270954 620 270960 632
rect 271012 620 271018 672
rect 271064 660 271092 700
rect 271138 688 271144 740
rect 271196 728 271202 740
rect 273257 731 273315 737
rect 273257 728 273269 731
rect 271196 700 273269 728
rect 271196 688 271202 700
rect 273257 697 273269 700
rect 273303 697 273315 731
rect 273257 691 273315 697
rect 273346 688 273352 740
rect 273404 728 273410 740
rect 279329 731 279387 737
rect 279329 728 279341 731
rect 273404 700 279341 728
rect 273404 688 273410 700
rect 279329 697 279341 700
rect 279375 697 279387 731
rect 279329 691 279387 697
rect 279789 731 279847 737
rect 279789 697 279801 731
rect 279835 728 279847 731
rect 281445 731 281503 737
rect 281445 728 281457 731
rect 279835 700 281457 728
rect 279835 697 279847 700
rect 279789 691 279847 697
rect 281445 697 281457 700
rect 281491 697 281503 731
rect 281445 691 281503 697
rect 281721 731 281779 737
rect 281721 697 281733 731
rect 281767 728 281779 731
rect 285493 731 285551 737
rect 285493 728 285505 731
rect 281767 700 285505 728
rect 281767 697 281779 700
rect 281721 691 281779 697
rect 285493 697 285505 700
rect 285539 697 285551 731
rect 285493 691 285551 697
rect 285769 731 285827 737
rect 285769 697 285781 731
rect 285815 728 285827 731
rect 290274 728 290280 740
rect 285815 700 290280 728
rect 285815 697 285827 700
rect 285769 691 285827 697
rect 290274 688 290280 700
rect 290332 688 290338 740
rect 290366 688 290372 740
rect 290424 728 290430 740
rect 295150 728 295156 740
rect 290424 700 295156 728
rect 290424 688 290430 700
rect 295150 688 295156 700
rect 295208 688 295214 740
rect 295245 731 295303 737
rect 295245 697 295257 731
rect 295291 728 295303 731
rect 319548 728 319576 836
rect 319625 833 319637 867
rect 319671 864 319683 867
rect 372724 864 372752 904
rect 319671 836 372752 864
rect 372801 867 372859 873
rect 319671 833 319683 836
rect 319625 827 319683 833
rect 372801 833 372813 867
rect 372847 864 372859 867
rect 372908 864 372936 904
rect 373902 892 373908 904
rect 373960 892 373966 944
rect 380158 892 380164 944
rect 380216 932 380222 944
rect 389358 932 389364 944
rect 380216 904 389364 932
rect 380216 892 380222 904
rect 389358 892 389364 904
rect 389416 892 389422 944
rect 511994 892 512000 944
rect 512052 932 512058 944
rect 516781 935 516839 941
rect 516781 932 516793 935
rect 512052 904 516793 932
rect 512052 892 512058 904
rect 516781 901 516793 904
rect 516827 901 516839 935
rect 516781 895 516839 901
rect 528189 935 528247 941
rect 528189 901 528201 935
rect 528235 932 528247 935
rect 538950 932 538956 944
rect 528235 904 538956 932
rect 528235 901 528247 904
rect 528189 895 528247 901
rect 538950 892 538956 904
rect 539008 892 539014 944
rect 559469 935 559527 941
rect 559469 901 559481 935
rect 559515 932 559527 935
rect 569402 932 569408 944
rect 559515 904 569408 932
rect 559515 901 559527 904
rect 559469 895 559527 901
rect 569402 892 569408 904
rect 569460 892 569466 944
rect 372847 836 372936 864
rect 372847 833 372859 836
rect 372801 827 372859 833
rect 373074 824 373080 876
rect 373132 864 373138 876
rect 378413 867 378471 873
rect 378413 864 378425 867
rect 373132 836 378425 864
rect 373132 824 373138 836
rect 378413 833 378425 836
rect 378459 833 378471 867
rect 378413 827 378471 833
rect 386509 867 386567 873
rect 386509 833 386521 867
rect 386555 864 386567 867
rect 404265 867 404323 873
rect 404265 864 404277 867
rect 386555 836 404277 864
rect 386555 833 386567 836
rect 386509 827 386567 833
rect 404265 833 404277 836
rect 404311 833 404323 867
rect 404265 827 404323 833
rect 425057 867 425115 873
rect 425057 833 425069 867
rect 425103 864 425115 867
rect 430853 867 430911 873
rect 430853 864 430865 867
rect 425103 836 430865 864
rect 425103 833 425115 836
rect 425057 827 425115 833
rect 430853 833 430865 836
rect 430899 833 430911 867
rect 430853 827 430911 833
rect 481085 867 481143 873
rect 481085 833 481097 867
rect 481131 864 481143 867
rect 508869 867 508927 873
rect 508869 864 508881 867
rect 481131 836 508881 864
rect 481131 833 481143 836
rect 481085 827 481143 833
rect 508869 833 508881 836
rect 508915 833 508927 867
rect 508869 827 508927 833
rect 538217 867 538275 873
rect 538217 833 538229 867
rect 538263 864 538275 867
rect 543093 867 543151 873
rect 543093 864 543105 867
rect 538263 836 543105 864
rect 538263 833 538275 836
rect 538217 827 538275 833
rect 543093 833 543105 836
rect 543139 833 543151 867
rect 543093 827 543151 833
rect 319714 756 319720 808
rect 319772 796 319778 808
rect 356425 799 356483 805
rect 356425 796 356437 799
rect 319772 768 356437 796
rect 319772 756 319778 768
rect 356425 765 356437 768
rect 356471 765 356483 799
rect 356425 759 356483 765
rect 356514 756 356520 808
rect 356572 796 356578 808
rect 372433 799 372491 805
rect 372433 796 372445 799
rect 356572 768 372445 796
rect 356572 756 356578 768
rect 372433 765 372445 768
rect 372479 765 372491 799
rect 372433 759 372491 765
rect 372522 756 372528 808
rect 372580 796 372586 808
rect 386325 799 386383 805
rect 386325 796 386337 799
rect 372580 768 386337 796
rect 372580 756 372586 768
rect 386325 765 386337 768
rect 386371 765 386383 799
rect 386325 759 386383 765
rect 386417 799 386475 805
rect 386417 765 386429 799
rect 386463 796 386475 799
rect 395985 799 396043 805
rect 395985 796 395997 799
rect 386463 768 395997 796
rect 386463 765 386475 768
rect 386417 759 386475 765
rect 395985 765 395997 768
rect 396031 765 396043 799
rect 395985 759 396043 765
rect 406102 756 406108 808
rect 406160 796 406166 808
rect 407022 796 407028 808
rect 406160 768 407028 796
rect 406160 756 406166 768
rect 407022 756 407028 768
rect 407080 756 407086 808
rect 411254 756 411260 808
rect 411312 796 411318 808
rect 425698 796 425704 808
rect 411312 768 425704 796
rect 411312 756 411318 768
rect 425698 756 425704 768
rect 425756 756 425762 808
rect 430761 799 430819 805
rect 430761 765 430773 799
rect 430807 796 430819 799
rect 436097 799 436155 805
rect 436097 796 436109 799
rect 430807 768 436109 796
rect 430807 765 430819 768
rect 430761 759 430819 765
rect 436097 765 436109 768
rect 436143 765 436155 799
rect 436097 759 436155 765
rect 463697 799 463755 805
rect 463697 765 463709 799
rect 463743 796 463755 799
rect 473173 799 473231 805
rect 473173 796 473185 799
rect 463743 768 473185 796
rect 463743 765 463755 768
rect 463697 759 463755 765
rect 473173 765 473185 768
rect 473219 765 473231 799
rect 473173 759 473231 765
rect 473357 799 473415 805
rect 473357 765 473369 799
rect 473403 796 473415 799
rect 473403 768 473676 796
rect 473403 765 473415 768
rect 473357 759 473415 765
rect 412177 731 412235 737
rect 412177 728 412189 731
rect 295291 700 319484 728
rect 319548 700 412189 728
rect 295291 697 295303 700
rect 295245 691 295303 697
rect 279973 663 280031 669
rect 279973 660 279985 663
rect 271064 632 279985 660
rect 279973 629 279985 632
rect 280019 629 280031 663
rect 279973 623 280031 629
rect 280062 620 280068 672
rect 280120 660 280126 672
rect 281534 660 281540 672
rect 280120 632 281540 660
rect 280120 620 280126 632
rect 281534 620 281540 632
rect 281592 620 281598 672
rect 281629 663 281687 669
rect 281629 629 281641 663
rect 281675 660 281687 663
rect 286042 660 286048 672
rect 281675 632 286048 660
rect 281675 629 281687 632
rect 281629 623 281687 629
rect 286042 620 286048 632
rect 286100 620 286106 672
rect 286137 663 286195 669
rect 286137 629 286149 663
rect 286183 660 286195 663
rect 289633 663 289691 669
rect 289633 660 289645 663
rect 286183 632 289645 660
rect 286183 629 286195 632
rect 286137 623 286195 629
rect 289633 629 289645 632
rect 289679 629 289691 663
rect 289633 623 289691 629
rect 289722 620 289728 672
rect 289780 660 289786 672
rect 290185 663 290243 669
rect 290185 660 290197 663
rect 289780 632 290197 660
rect 289780 620 289786 632
rect 290185 629 290197 632
rect 290231 629 290243 663
rect 290185 623 290243 629
rect 290645 663 290703 669
rect 290645 629 290657 663
rect 290691 660 290703 663
rect 296901 663 296959 669
rect 296901 660 296913 663
rect 290691 632 296913 660
rect 290691 629 290703 632
rect 290645 623 290703 629
rect 296901 629 296913 632
rect 296947 629 296959 663
rect 296901 623 296959 629
rect 296990 620 296996 672
rect 297048 660 297054 672
rect 300670 660 300676 672
rect 297048 632 300676 660
rect 297048 620 297054 632
rect 300670 620 300676 632
rect 300728 620 300734 672
rect 300762 620 300768 672
rect 300820 660 300826 672
rect 319349 663 319407 669
rect 319349 660 319361 663
rect 300820 632 319361 660
rect 300820 620 300826 632
rect 319349 629 319361 632
rect 319395 629 319407 663
rect 319456 660 319484 700
rect 412177 697 412189 700
rect 412223 697 412235 731
rect 412177 691 412235 697
rect 434990 688 434996 740
rect 435048 728 435054 740
rect 442810 728 442816 740
rect 435048 700 442816 728
rect 435048 688 435054 700
rect 442810 688 442816 700
rect 442868 688 442874 740
rect 335354 660 335360 672
rect 319456 632 335360 660
rect 319349 623 319407 629
rect 335354 620 335360 632
rect 335412 620 335418 672
rect 335538 620 335544 672
rect 335596 660 335602 672
rect 473357 663 473415 669
rect 473357 660 473369 663
rect 335596 632 473369 660
rect 335596 620 335602 632
rect 473357 629 473369 632
rect 473403 629 473415 663
rect 473648 660 473676 768
rect 476758 756 476764 808
rect 476816 796 476822 808
rect 486142 796 486148 808
rect 476816 768 486148 796
rect 476816 756 476822 768
rect 486142 756 486148 768
rect 486200 756 486206 808
rect 514757 799 514815 805
rect 514757 765 514769 799
rect 514803 796 514815 799
rect 518710 796 518716 808
rect 514803 768 518716 796
rect 514803 765 514815 768
rect 514757 759 514815 765
rect 518710 756 518716 768
rect 518768 756 518774 808
rect 476390 688 476396 740
rect 476448 728 476454 740
rect 490190 728 490196 740
rect 476448 700 490196 728
rect 476448 688 476454 700
rect 490190 688 490196 700
rect 490248 688 490254 740
rect 547230 660 547236 672
rect 473648 632 547236 660
rect 473357 623 473415 629
rect 547230 620 547236 632
rect 547288 620 547294 672
rect 183833 595 183891 601
rect 176580 564 183784 592
rect 176381 555 176439 561
rect 175875 496 176056 524
rect 175875 493 175887 496
rect 175829 487 175887 493
rect 176194 484 176200 536
rect 176252 524 176258 536
rect 176473 527 176531 533
rect 176252 496 176297 524
rect 176252 484 176258 496
rect 176473 493 176485 527
rect 176519 524 176531 527
rect 183649 527 183707 533
rect 183649 524 183661 527
rect 176519 496 183661 524
rect 176519 493 176531 496
rect 176473 487 176531 493
rect 183649 493 183661 496
rect 183695 493 183707 527
rect 183756 524 183784 564
rect 183833 561 183845 595
rect 183879 561 183891 595
rect 335449 595 335507 601
rect 335449 592 335461 595
rect 183833 555 183891 561
rect 183940 564 335461 592
rect 183940 524 183968 564
rect 335449 561 335461 564
rect 335495 561 335507 595
rect 335449 555 335507 561
rect 335725 595 335783 601
rect 335725 561 335737 595
rect 335771 592 335783 595
rect 347317 595 347375 601
rect 347317 592 347329 595
rect 335771 564 347329 592
rect 335771 561 335783 564
rect 335725 555 335783 561
rect 347317 561 347329 564
rect 347363 561 347375 595
rect 347317 555 347375 561
rect 347501 595 347559 601
rect 347501 561 347513 595
rect 347547 592 347559 595
rect 473449 595 473507 601
rect 473449 592 473461 595
rect 347547 564 473461 592
rect 347547 561 347559 564
rect 347501 555 347559 561
rect 473449 561 473461 564
rect 473495 561 473507 595
rect 473449 555 473507 561
rect 473541 595 473599 601
rect 473541 561 473553 595
rect 473587 592 473599 595
rect 480714 592 480720 604
rect 473587 564 480720 592
rect 473587 561 473599 564
rect 473541 555 473599 561
rect 480714 552 480720 564
rect 480772 552 480778 604
rect 509878 552 509884 604
rect 509936 592 509942 604
rect 516870 592 516876 604
rect 509936 564 516876 592
rect 509936 552 509942 564
rect 516870 552 516876 564
rect 516928 552 516934 604
rect 183756 496 183968 524
rect 183649 487 183707 493
rect 184014 484 184020 536
rect 184072 524 184078 536
rect 217502 524 217508 536
rect 184072 496 217508 524
rect 184072 484 184078 496
rect 217502 484 217508 496
rect 217560 484 217566 536
rect 217597 527 217655 533
rect 217597 493 217609 527
rect 217643 524 217655 527
rect 217686 524 217692 536
rect 217643 496 217692 524
rect 217643 493 217655 496
rect 217597 487 217655 493
rect 217686 484 217692 496
rect 217744 484 217750 536
rect 217778 484 217784 536
rect 217836 524 217842 536
rect 217873 527 217931 533
rect 217873 524 217885 527
rect 217836 496 217885 524
rect 217836 484 217842 496
rect 217873 493 217885 496
rect 217919 493 217931 527
rect 217873 487 217931 493
rect 217962 484 217968 536
rect 218020 524 218026 536
rect 241517 527 241575 533
rect 241517 524 241529 527
rect 218020 496 241529 524
rect 218020 484 218026 496
rect 241517 493 241529 496
rect 241563 493 241575 527
rect 241517 487 241575 493
rect 241790 484 241796 536
rect 241848 524 241854 536
rect 246574 524 246580 536
rect 241848 496 246580 524
rect 241848 484 241854 496
rect 246574 484 246580 496
rect 246632 484 246638 536
rect 247034 484 247040 536
rect 247092 524 247098 536
rect 247494 524 247500 536
rect 247092 496 247500 524
rect 247092 484 247098 496
rect 247494 484 247500 496
rect 247552 484 247558 536
rect 247589 527 247647 533
rect 247589 493 247601 527
rect 247635 524 247647 527
rect 251637 527 251695 533
rect 247635 496 251588 524
rect 247635 493 247647 496
rect 247589 487 247647 493
rect 111797 459 111855 465
rect 111797 456 111809 459
rect 97276 428 111809 456
rect 97169 419 97227 425
rect 111797 425 111809 428
rect 111843 425 111855 459
rect 111797 419 111855 425
rect 112257 459 112315 465
rect 112257 425 112269 459
rect 112303 456 112315 459
rect 135349 459 135407 465
rect 135349 456 135361 459
rect 112303 428 135361 456
rect 112303 425 112315 428
rect 112257 419 112315 425
rect 135349 425 135361 428
rect 135395 425 135407 459
rect 135349 419 135407 425
rect 135438 416 135444 468
rect 135496 456 135502 468
rect 142246 456 142252 468
rect 135496 428 142252 456
rect 135496 416 135502 428
rect 142246 416 142252 428
rect 142304 416 142310 468
rect 142338 416 142344 468
rect 142396 456 142402 468
rect 144730 456 144736 468
rect 142396 428 144736 456
rect 142396 416 142402 428
rect 144730 416 144736 428
rect 144788 416 144794 468
rect 144825 459 144883 465
rect 144825 425 144837 459
rect 144871 456 144883 459
rect 183465 459 183523 465
rect 183465 456 183477 459
rect 144871 428 183477 456
rect 144871 425 144883 428
rect 144825 419 144883 425
rect 183465 425 183477 428
rect 183511 425 183523 459
rect 193401 459 193459 465
rect 193401 456 193413 459
rect 183465 419 183523 425
rect 183664 428 193413 456
rect 74000 360 74304 388
rect 74353 391 74411 397
rect 73893 351 73951 357
rect 74353 357 74365 391
rect 74399 388 74411 391
rect 76561 391 76619 397
rect 76561 388 76573 391
rect 74399 360 76573 388
rect 74399 357 74411 360
rect 74353 351 74411 357
rect 76561 357 76573 360
rect 76607 357 76619 391
rect 76561 351 76619 357
rect 76653 391 76711 397
rect 76653 357 76665 391
rect 76699 388 76711 391
rect 89530 388 89536 400
rect 76699 360 89536 388
rect 76699 357 76711 360
rect 76653 351 76711 357
rect 89530 348 89536 360
rect 89588 348 89594 400
rect 89625 391 89683 397
rect 89625 357 89637 391
rect 89671 388 89683 391
rect 90726 388 90732 400
rect 89671 360 90732 388
rect 89671 357 89683 360
rect 89625 351 89683 357
rect 90726 348 90732 360
rect 90784 348 90790 400
rect 91094 348 91100 400
rect 91152 388 91158 400
rect 92661 391 92719 397
rect 92661 388 92673 391
rect 91152 360 92673 388
rect 91152 348 91158 360
rect 92661 357 92673 360
rect 92707 357 92719 391
rect 92661 351 92719 357
rect 92845 391 92903 397
rect 92845 357 92857 391
rect 92891 388 92903 391
rect 94222 388 94228 400
rect 92891 360 94228 388
rect 92891 357 92903 360
rect 92845 351 92903 357
rect 94222 348 94228 360
rect 94280 348 94286 400
rect 94317 391 94375 397
rect 94317 357 94329 391
rect 94363 388 94375 391
rect 95789 391 95847 397
rect 95789 388 95801 391
rect 94363 360 95801 388
rect 94363 357 94375 360
rect 94317 351 94375 357
rect 95789 357 95801 360
rect 95835 357 95847 391
rect 95789 351 95847 357
rect 95878 348 95884 400
rect 95936 388 95942 400
rect 111886 388 111892 400
rect 95936 360 111892 388
rect 95936 348 95942 360
rect 111886 348 111892 360
rect 111944 348 111950 400
rect 112070 348 112076 400
rect 112128 388 112134 400
rect 153194 388 153200 400
rect 112128 360 153200 388
rect 112128 348 112134 360
rect 153194 348 153200 360
rect 153252 348 153258 400
rect 153289 391 153347 397
rect 153289 357 153301 391
rect 153335 388 153347 391
rect 153746 388 153752 400
rect 153335 360 153752 388
rect 153335 357 153347 360
rect 153289 351 153347 357
rect 153746 348 153752 360
rect 153804 348 153810 400
rect 153841 391 153899 397
rect 153841 357 153853 391
rect 153887 388 153899 391
rect 154577 391 154635 397
rect 154577 388 154589 391
rect 153887 360 154589 388
rect 153887 357 153899 360
rect 153841 351 153899 357
rect 154577 357 154589 360
rect 154623 357 154635 391
rect 154577 351 154635 357
rect 154666 348 154672 400
rect 154724 388 154730 400
rect 157153 391 157211 397
rect 157153 388 157165 391
rect 154724 360 157165 388
rect 154724 348 154730 360
rect 157153 357 157165 360
rect 157199 357 157211 391
rect 157153 351 157211 357
rect 157242 348 157248 400
rect 157300 388 157306 400
rect 175921 391 175979 397
rect 175921 388 175933 391
rect 157300 360 175933 388
rect 157300 348 157306 360
rect 175921 357 175933 360
rect 175967 357 175979 391
rect 176286 388 176292 400
rect 176247 360 176292 388
rect 175921 351 175979 357
rect 176286 348 176292 360
rect 176344 348 176350 400
rect 183664 397 183692 428
rect 193401 425 193413 428
rect 193447 425 193459 459
rect 193401 419 193459 425
rect 193490 416 193496 468
rect 193548 456 193554 468
rect 198366 456 198372 468
rect 193548 428 198372 456
rect 193548 416 193554 428
rect 198366 416 198372 428
rect 198424 416 198430 468
rect 198458 416 198464 468
rect 198516 456 198522 468
rect 198516 428 198561 456
rect 198516 416 198522 428
rect 198734 416 198740 468
rect 198792 456 198798 468
rect 198921 459 198979 465
rect 198921 456 198933 459
rect 198792 428 198933 456
rect 198792 416 198798 428
rect 198921 425 198933 428
rect 198967 425 198979 459
rect 198921 419 198979 425
rect 199381 459 199439 465
rect 199381 425 199393 459
rect 199427 456 199439 459
rect 203061 459 203119 465
rect 203061 456 203073 459
rect 199427 428 203073 456
rect 199427 425 199439 428
rect 199381 419 199439 425
rect 203061 425 203073 428
rect 203107 425 203119 459
rect 203061 419 203119 425
rect 203150 416 203156 468
rect 203208 456 203214 468
rect 211982 456 211988 468
rect 203208 428 211988 456
rect 203208 416 203214 428
rect 211982 416 211988 428
rect 212040 416 212046 468
rect 212445 459 212503 465
rect 212445 425 212457 459
rect 212491 456 212503 459
rect 241609 459 241667 465
rect 241609 456 241621 459
rect 212491 428 241621 456
rect 212491 425 212503 428
rect 212445 419 212503 425
rect 241609 425 241621 428
rect 241655 425 241667 459
rect 241609 419 241667 425
rect 241698 416 241704 468
rect 241756 456 241762 468
rect 247218 456 247224 468
rect 241756 428 247224 456
rect 241756 416 241762 428
rect 247218 416 247224 428
rect 247276 416 247282 468
rect 250993 459 251051 465
rect 250993 425 251005 459
rect 251039 456 251051 459
rect 251361 459 251419 465
rect 251361 456 251373 459
rect 251039 428 251373 456
rect 251039 425 251051 428
rect 250993 419 251051 425
rect 251361 425 251373 428
rect 251407 425 251419 459
rect 251560 456 251588 496
rect 251637 493 251649 527
rect 251683 524 251695 527
rect 259641 527 259699 533
rect 259641 524 259653 527
rect 251683 496 259653 524
rect 251683 493 251695 496
rect 251637 487 251695 493
rect 259641 493 259653 496
rect 259687 493 259699 527
rect 260837 527 260895 533
rect 260837 524 260849 527
rect 259641 487 259699 493
rect 259748 496 260849 524
rect 251560 428 251680 456
rect 251361 419 251419 425
rect 176381 391 176439 397
rect 176381 357 176393 391
rect 176427 388 176439 391
rect 183557 391 183615 397
rect 183557 388 183569 391
rect 176427 360 183569 388
rect 176427 357 176439 360
rect 176381 351 176439 357
rect 183557 357 183569 360
rect 183603 357 183615 391
rect 183557 351 183615 357
rect 183649 391 183707 397
rect 183649 357 183661 391
rect 183695 357 183707 391
rect 193309 391 193367 397
rect 193309 388 193321 391
rect 183649 351 183707 357
rect 183756 360 193321 388
rect 35299 292 38792 320
rect 39025 323 39083 329
rect 35299 289 35311 292
rect 35253 283 35311 289
rect 39025 289 39037 323
rect 39071 320 39083 323
rect 39761 323 39819 329
rect 39761 320 39773 323
rect 39071 292 39773 320
rect 39071 289 39083 292
rect 39025 283 39083 289
rect 39761 289 39773 292
rect 39807 289 39819 323
rect 39761 283 39819 289
rect 39853 323 39911 329
rect 39853 289 39865 323
rect 39899 320 39911 323
rect 49142 320 49148 332
rect 39899 292 49148 320
rect 39899 289 39911 292
rect 39853 283 39911 289
rect 49142 280 49148 292
rect 49200 280 49206 332
rect 49237 323 49295 329
rect 49237 289 49249 323
rect 49283 320 49295 323
rect 58986 320 58992 332
rect 49283 292 58992 320
rect 49283 289 49295 292
rect 49237 283 49295 289
rect 58986 280 58992 292
rect 59044 280 59050 332
rect 183756 329 183784 360
rect 193309 357 193321 360
rect 193355 357 193367 391
rect 193309 351 193367 357
rect 193582 348 193588 400
rect 193640 388 193646 400
rect 196529 391 196587 397
rect 196529 388 196541 391
rect 193640 360 196541 388
rect 193640 348 193646 360
rect 196529 357 196541 360
rect 196575 357 196587 391
rect 196529 351 196587 357
rect 196618 348 196624 400
rect 196676 388 196682 400
rect 196897 391 196955 397
rect 196897 388 196909 391
rect 196676 360 196909 388
rect 196676 348 196682 360
rect 196897 357 196909 360
rect 196943 357 196955 391
rect 196897 351 196955 357
rect 196986 348 196992 400
rect 197044 388 197050 400
rect 198182 388 198188 400
rect 197044 360 198188 388
rect 197044 348 197050 360
rect 198182 348 198188 360
rect 198240 348 198246 400
rect 198274 348 198280 400
rect 198332 388 198338 400
rect 198645 391 198703 397
rect 198332 360 198377 388
rect 198332 348 198338 360
rect 198645 357 198657 391
rect 198691 388 198703 391
rect 199289 391 199347 397
rect 199289 388 199301 391
rect 198691 360 199301 388
rect 198691 357 198703 360
rect 198645 351 198703 357
rect 199289 357 199301 360
rect 199335 357 199347 391
rect 199289 351 199347 357
rect 199473 391 199531 397
rect 199473 357 199485 391
rect 199519 388 199531 391
rect 251545 391 251603 397
rect 251545 388 251557 391
rect 199519 360 251557 388
rect 199519 357 199531 360
rect 199473 351 199531 357
rect 251545 357 251557 360
rect 251591 357 251603 391
rect 251652 388 251680 428
rect 251726 416 251732 468
rect 251784 456 251790 468
rect 252830 456 252836 468
rect 251784 428 252836 456
rect 251784 416 251790 428
rect 252830 416 252836 428
rect 252888 416 252894 468
rect 253106 416 253112 468
rect 253164 456 253170 468
rect 259178 456 259184 468
rect 253164 428 259184 456
rect 253164 416 253170 428
rect 259178 416 259184 428
rect 259236 416 259242 468
rect 259748 388 259776 496
rect 260837 493 260849 496
rect 260883 493 260895 527
rect 260837 487 260895 493
rect 261754 484 261760 536
rect 261812 524 261818 536
rect 265434 524 265440 536
rect 261812 496 265440 524
rect 261812 484 261818 496
rect 265434 484 265440 496
rect 265492 484 265498 536
rect 265529 527 265587 533
rect 265529 493 265541 527
rect 265575 524 265587 527
rect 268841 527 268899 533
rect 268841 524 268853 527
rect 265575 496 268853 524
rect 265575 493 265587 496
rect 265529 487 265587 493
rect 268841 493 268853 496
rect 268887 493 268899 527
rect 268841 487 268899 493
rect 270405 527 270463 533
rect 270405 493 270417 527
rect 270451 524 270463 527
rect 270497 527 270555 533
rect 270497 524 270509 527
rect 270451 496 270509 524
rect 270451 493 270463 496
rect 270405 487 270463 493
rect 270497 493 270509 496
rect 270543 493 270555 527
rect 270497 487 270555 493
rect 270770 484 270776 536
rect 270828 524 270834 536
rect 270828 496 270873 524
rect 270828 484 270834 496
rect 271874 484 271880 536
rect 271932 524 271938 536
rect 279326 524 279332 536
rect 271932 496 279332 524
rect 271932 484 271938 496
rect 279326 484 279332 496
rect 279384 484 279390 536
rect 279789 527 279847 533
rect 279789 493 279801 527
rect 279835 493 279847 527
rect 279789 487 279847 493
rect 279896 496 290044 524
rect 260006 416 260012 468
rect 260064 456 260070 468
rect 260558 456 260564 468
rect 260064 428 260564 456
rect 260064 416 260070 428
rect 260558 416 260564 428
rect 260616 416 260622 468
rect 260653 459 260711 465
rect 260653 425 260665 459
rect 260699 456 260711 459
rect 260929 459 260987 465
rect 260929 456 260941 459
rect 260699 428 260941 456
rect 260699 425 260711 428
rect 260653 419 260711 425
rect 260929 425 260941 428
rect 260975 425 260987 459
rect 260929 419 260987 425
rect 261202 416 261208 468
rect 261260 456 261266 468
rect 262858 456 262864 468
rect 261260 428 262864 456
rect 261260 416 261266 428
rect 262858 416 262864 428
rect 262916 416 262922 468
rect 262950 416 262956 468
rect 263008 456 263014 468
rect 264882 456 264888 468
rect 263008 428 264888 456
rect 263008 416 263014 428
rect 264882 416 264888 428
rect 264940 416 264946 468
rect 265069 459 265127 465
rect 265069 425 265081 459
rect 265115 456 265127 459
rect 268933 459 268991 465
rect 268933 456 268945 459
rect 265115 428 268945 456
rect 265115 425 265127 428
rect 265069 419 265127 425
rect 268933 425 268945 428
rect 268979 425 268991 459
rect 268933 419 268991 425
rect 269022 416 269028 468
rect 269080 456 269086 468
rect 269482 456 269488 468
rect 269080 428 269488 456
rect 269080 416 269086 428
rect 269482 416 269488 428
rect 269540 416 269546 468
rect 270313 459 270371 465
rect 270313 425 270325 459
rect 270359 456 270371 459
rect 270589 459 270647 465
rect 270589 456 270601 459
rect 270359 428 270601 456
rect 270359 425 270371 428
rect 270313 419 270371 425
rect 270589 425 270601 428
rect 270635 425 270647 459
rect 270589 419 270647 425
rect 270678 416 270684 468
rect 270736 456 270742 468
rect 279804 456 279832 487
rect 270736 428 279832 456
rect 270736 416 270742 428
rect 251652 360 259776 388
rect 259825 391 259883 397
rect 251545 351 251603 357
rect 259825 357 259837 391
rect 259871 388 259883 391
rect 270497 391 270555 397
rect 270497 388 270509 391
rect 259871 360 270509 388
rect 259871 357 259883 360
rect 259825 351 259883 357
rect 270497 357 270509 360
rect 270543 357 270555 391
rect 270497 351 270555 357
rect 270770 348 270776 400
rect 270828 388 270834 400
rect 279896 388 279924 496
rect 279973 459 280031 465
rect 279973 425 279985 459
rect 280019 456 280031 459
rect 280249 459 280307 465
rect 280249 456 280261 459
rect 280019 428 280261 456
rect 280019 425 280031 428
rect 279973 419 280031 425
rect 280249 425 280261 428
rect 280295 425 280307 459
rect 280249 419 280307 425
rect 280338 416 280344 468
rect 280396 456 280402 468
rect 281534 456 281540 468
rect 280396 428 281540 456
rect 280396 416 280402 428
rect 281534 416 281540 428
rect 281592 416 281598 468
rect 281629 459 281687 465
rect 281629 425 281641 459
rect 281675 456 281687 459
rect 285493 459 285551 465
rect 285493 456 285505 459
rect 281675 428 285505 456
rect 281675 425 281687 428
rect 281629 419 281687 425
rect 285493 425 285505 428
rect 285539 425 285551 459
rect 285493 419 285551 425
rect 285582 416 285588 468
rect 285640 456 285646 468
rect 285674 456 285680 468
rect 285640 428 285680 456
rect 285640 416 285646 428
rect 285674 416 285680 428
rect 285732 416 285738 468
rect 285769 459 285827 465
rect 285769 425 285781 459
rect 285815 456 285827 459
rect 289909 459 289967 465
rect 289909 456 289921 459
rect 285815 428 289921 456
rect 285815 425 285827 428
rect 285769 419 285827 425
rect 289909 425 289921 428
rect 289955 425 289967 459
rect 289909 419 289967 425
rect 270828 360 279924 388
rect 280065 391 280123 397
rect 270828 348 270834 360
rect 280065 357 280077 391
rect 280111 388 280123 391
rect 289817 391 289875 397
rect 289817 388 289829 391
rect 280111 360 289829 388
rect 280111 357 280123 360
rect 280065 351 280123 357
rect 289817 357 289829 360
rect 289863 357 289875 391
rect 290016 388 290044 496
rect 290090 484 290096 536
rect 290148 524 290154 536
rect 293862 524 293868 536
rect 290148 496 293868 524
rect 290148 484 290154 496
rect 293862 484 293868 496
rect 293920 484 293926 536
rect 293957 527 294015 533
rect 293957 493 293969 527
rect 294003 524 294015 527
rect 296717 527 296775 533
rect 296717 524 296729 527
rect 294003 496 296729 524
rect 294003 493 294015 496
rect 293957 487 294015 493
rect 296717 493 296729 496
rect 296763 493 296775 527
rect 297453 527 297511 533
rect 297453 524 297465 527
rect 296717 487 296775 493
rect 296824 496 297465 524
rect 290182 416 290188 468
rect 290240 456 290246 468
rect 296824 456 296852 496
rect 297453 493 297465 496
rect 297499 493 297511 527
rect 297453 487 297511 493
rect 297545 527 297603 533
rect 297545 493 297557 527
rect 297591 524 297603 527
rect 318797 527 318855 533
rect 318797 524 318809 527
rect 297591 496 318809 524
rect 297591 493 297603 496
rect 297545 487 297603 493
rect 318797 493 318809 496
rect 318843 493 318855 527
rect 318797 487 318855 493
rect 321833 527 321891 533
rect 321833 493 321845 527
rect 321879 524 321891 527
rect 322937 527 322995 533
rect 322937 524 322949 527
rect 321879 496 322949 524
rect 321879 493 321891 496
rect 321833 487 321891 493
rect 322937 493 322949 496
rect 322983 493 322995 527
rect 322937 487 322995 493
rect 323397 527 323455 533
rect 323397 493 323409 527
rect 323443 524 323455 527
rect 327902 524 327908 536
rect 323443 496 327908 524
rect 323443 493 323455 496
rect 323397 487 323455 493
rect 327902 484 327908 496
rect 327960 484 327966 536
rect 327997 527 328055 533
rect 327997 493 328009 527
rect 328043 524 328055 527
rect 335541 527 335599 533
rect 335541 524 335553 527
rect 328043 496 335553 524
rect 328043 493 328055 496
rect 327997 487 328055 493
rect 335541 493 335553 496
rect 335587 493 335599 527
rect 336001 527 336059 533
rect 336001 524 336013 527
rect 335541 487 335599 493
rect 335648 496 336013 524
rect 290240 428 296852 456
rect 296993 459 297051 465
rect 290240 416 290246 428
rect 296993 425 297005 459
rect 297039 456 297051 459
rect 309229 459 309287 465
rect 309229 456 309241 459
rect 297039 428 309241 456
rect 297039 425 297051 428
rect 296993 419 297051 425
rect 309229 425 309241 428
rect 309275 425 309287 459
rect 309229 419 309287 425
rect 318613 459 318671 465
rect 318613 425 318625 459
rect 318659 456 318671 459
rect 318886 456 318892 468
rect 318659 428 318892 456
rect 318659 425 318671 428
rect 318613 419 318671 425
rect 318886 416 318892 428
rect 318944 416 318950 468
rect 318978 416 318984 468
rect 319036 456 319042 468
rect 323026 456 323032 468
rect 319036 428 323032 456
rect 319036 416 319042 428
rect 323026 416 323032 428
rect 323084 416 323090 468
rect 323213 459 323271 465
rect 323213 425 323225 459
rect 323259 456 323271 459
rect 335648 456 335676 496
rect 336001 493 336013 496
rect 336047 493 336059 527
rect 336001 487 336059 493
rect 336093 527 336151 533
rect 336093 493 336105 527
rect 336139 524 336151 527
rect 337473 527 337531 533
rect 337473 524 337485 527
rect 336139 496 337485 524
rect 336139 493 336151 496
rect 336093 487 336151 493
rect 337473 493 337485 496
rect 337519 493 337531 527
rect 337473 487 337531 493
rect 337565 527 337623 533
rect 337565 493 337577 527
rect 337611 524 337623 527
rect 338761 527 338819 533
rect 338761 524 338773 527
rect 337611 496 338773 524
rect 337611 493 337623 496
rect 337565 487 337623 493
rect 338761 493 338773 496
rect 338807 493 338819 527
rect 338761 487 338819 493
rect 338853 527 338911 533
rect 338853 493 338865 527
rect 338899 524 338911 527
rect 348329 527 348387 533
rect 348329 524 348341 527
rect 338899 496 348341 524
rect 338899 493 338911 496
rect 338853 487 338911 493
rect 348329 493 348341 496
rect 348375 493 348387 527
rect 348329 487 348387 493
rect 348513 527 348571 533
rect 348513 493 348525 527
rect 348559 524 348571 527
rect 352653 527 352711 533
rect 352653 524 352665 527
rect 348559 496 352665 524
rect 348559 493 348571 496
rect 348513 487 348571 493
rect 352653 493 352665 496
rect 352699 493 352711 527
rect 352653 487 352711 493
rect 352837 527 352895 533
rect 352837 493 352849 527
rect 352883 524 352895 527
rect 356517 527 356575 533
rect 356517 524 356529 527
rect 352883 496 356529 524
rect 352883 493 352895 496
rect 352837 487 352895 493
rect 356517 493 356529 496
rect 356563 493 356575 527
rect 356517 487 356575 493
rect 356609 527 356667 533
rect 356609 493 356621 527
rect 356655 524 356667 527
rect 376662 524 376668 536
rect 356655 496 376668 524
rect 356655 493 356667 496
rect 356609 487 356667 493
rect 376662 484 376668 496
rect 376720 484 376726 536
rect 381538 484 381544 536
rect 381596 524 381602 536
rect 386417 527 386475 533
rect 386417 524 386429 527
rect 381596 496 386429 524
rect 381596 484 381602 496
rect 386417 493 386429 496
rect 386463 493 386475 527
rect 386417 487 386475 493
rect 386509 527 386567 533
rect 386509 493 386521 527
rect 386555 524 386567 527
rect 393406 524 393412 536
rect 386555 496 393412 524
rect 386555 493 386567 496
rect 386509 487 386567 493
rect 393406 484 393412 496
rect 393464 484 393470 536
rect 395985 527 396043 533
rect 395985 493 395997 527
rect 396031 524 396043 527
rect 425057 527 425115 533
rect 425057 524 425069 527
rect 396031 496 425069 524
rect 396031 493 396043 496
rect 395985 487 396043 493
rect 425057 493 425069 496
rect 425103 493 425115 527
rect 425057 487 425115 493
rect 430853 527 430911 533
rect 430853 493 430865 527
rect 430899 524 430911 527
rect 463697 527 463755 533
rect 463697 524 463709 527
rect 430899 496 463709 524
rect 430899 493 430911 496
rect 430853 487 430911 493
rect 463697 493 463709 496
rect 463743 493 463755 527
rect 463697 487 463755 493
rect 473173 527 473231 533
rect 473173 493 473185 527
rect 473219 524 473231 527
rect 473357 527 473415 533
rect 473357 524 473369 527
rect 473219 496 473369 524
rect 473219 493 473231 496
rect 473173 487 473231 493
rect 473357 493 473369 496
rect 473403 493 473415 527
rect 473357 487 473415 493
rect 473633 527 473691 533
rect 473633 493 473645 527
rect 473679 524 473691 527
rect 481085 527 481143 533
rect 481085 524 481097 527
rect 473679 496 481097 524
rect 473679 493 473691 496
rect 473633 487 473691 493
rect 481085 493 481097 496
rect 481131 493 481143 527
rect 481085 487 481143 493
rect 508869 527 508927 533
rect 508869 493 508881 527
rect 508915 524 508927 527
rect 514757 527 514815 533
rect 514757 524 514769 527
rect 508915 496 514769 524
rect 508915 493 508927 496
rect 508869 487 508927 493
rect 514757 493 514769 496
rect 514803 493 514815 527
rect 514757 487 514815 493
rect 323259 428 335676 456
rect 335725 459 335783 465
rect 323259 425 323271 428
rect 323213 419 323271 425
rect 335725 425 335737 459
rect 335771 456 335783 459
rect 337838 456 337844 468
rect 335771 428 337844 456
rect 335771 425 335783 428
rect 335725 419 335783 425
rect 337838 416 337844 428
rect 337896 416 337902 468
rect 337933 459 337991 465
rect 337933 425 337945 459
rect 337979 456 337991 459
rect 372617 459 372675 465
rect 372617 456 372629 459
rect 337979 428 372629 456
rect 337979 425 337991 428
rect 337933 419 337991 425
rect 372617 425 372629 428
rect 372663 425 372675 459
rect 459557 459 459615 465
rect 459557 456 459569 459
rect 372617 419 372675 425
rect 372816 428 459569 456
rect 372816 397 372844 428
rect 459557 425 459569 428
rect 459603 425 459615 459
rect 459557 419 459615 425
rect 459741 459 459799 465
rect 459741 425 459753 459
rect 459787 456 459799 459
rect 473449 459 473507 465
rect 473449 456 473461 459
rect 459787 428 473461 456
rect 459787 425 459799 428
rect 459741 419 459799 425
rect 473449 425 473461 428
rect 473495 425 473507 459
rect 473449 419 473507 425
rect 473541 459 473599 465
rect 473541 425 473553 459
rect 473587 456 473599 459
rect 489822 456 489828 468
rect 473587 428 489828 456
rect 473587 425 473599 428
rect 473541 419 473599 425
rect 489822 416 489828 428
rect 489880 416 489886 468
rect 297545 391 297603 397
rect 297545 388 297557 391
rect 290016 360 297557 388
rect 289817 351 289875 357
rect 297545 357 297557 360
rect 297591 357 297603 391
rect 297545 351 297603 357
rect 297637 391 297695 397
rect 297637 357 297649 391
rect 297683 388 297695 391
rect 300673 391 300731 397
rect 300673 388 300685 391
rect 297683 360 300685 388
rect 297683 357 297695 360
rect 297637 351 297695 357
rect 300673 357 300685 360
rect 300719 357 300731 391
rect 300673 351 300731 357
rect 300765 391 300823 397
rect 300765 357 300777 391
rect 300811 388 300823 391
rect 322937 391 322995 397
rect 322937 388 322949 391
rect 300811 360 322949 388
rect 300811 357 300823 360
rect 300765 351 300823 357
rect 322937 357 322949 360
rect 322983 357 322995 391
rect 322937 351 322995 357
rect 323397 391 323455 397
rect 323397 357 323409 391
rect 323443 388 323455 391
rect 348237 391 348295 397
rect 348237 388 348249 391
rect 323443 360 348249 388
rect 323443 357 323455 360
rect 323397 351 323455 357
rect 348237 357 348249 360
rect 348283 357 348295 391
rect 348237 351 348295 357
rect 348329 391 348387 397
rect 348329 357 348341 391
rect 348375 388 348387 391
rect 356609 391 356667 397
rect 356609 388 356621 391
rect 348375 360 356621 388
rect 348375 357 348387 360
rect 348329 351 348387 357
rect 356609 357 356621 360
rect 356655 357 356667 391
rect 356609 351 356667 357
rect 356701 391 356759 397
rect 356701 357 356713 391
rect 356747 388 356759 391
rect 367097 391 367155 397
rect 367097 388 367109 391
rect 356747 360 367109 388
rect 356747 357 356759 360
rect 356701 351 356759 357
rect 367097 357 367109 360
rect 367143 357 367155 391
rect 372801 391 372859 397
rect 367097 351 367155 357
rect 368492 360 372476 388
rect 59081 323 59139 329
rect 59081 289 59093 323
rect 59127 320 59139 323
rect 60829 323 60887 329
rect 60829 320 60841 323
rect 59127 292 60841 320
rect 59127 289 59139 292
rect 59081 283 59139 289
rect 60829 289 60841 292
rect 60875 289 60887 323
rect 72973 323 73031 329
rect 72973 320 72985 323
rect 60829 283 60887 289
rect 60936 292 72985 320
rect 1394 212 1400 264
rect 1452 252 1458 264
rect 5629 255 5687 261
rect 5629 252 5641 255
rect 1452 224 5641 252
rect 1452 212 1458 224
rect 5629 221 5641 224
rect 5675 221 5687 255
rect 5629 215 5687 221
rect 5997 255 6055 261
rect 5997 221 6009 255
rect 6043 252 6055 255
rect 10410 252 10416 264
rect 6043 224 10416 252
rect 6043 221 6055 224
rect 5997 215 6055 221
rect 10410 212 10416 224
rect 10468 212 10474 264
rect 10505 255 10563 261
rect 10505 221 10517 255
rect 10551 252 10563 255
rect 25314 252 25320 264
rect 10551 224 25320 252
rect 10551 221 10563 224
rect 10505 215 10563 221
rect 25314 212 25320 224
rect 25372 212 25378 264
rect 38378 252 38384 264
rect 26252 224 38384 252
rect 3050 144 3056 196
rect 3108 184 3114 196
rect 5353 187 5411 193
rect 5353 184 5365 187
rect 3108 156 5365 184
rect 3108 144 3114 156
rect 5353 153 5365 156
rect 5399 153 5411 187
rect 5353 147 5411 153
rect 5537 187 5595 193
rect 5537 153 5549 187
rect 5583 184 5595 187
rect 26252 184 26280 224
rect 38378 212 38384 224
rect 38436 212 38442 264
rect 38657 255 38715 261
rect 38657 221 38669 255
rect 38703 252 38715 255
rect 53190 252 53196 264
rect 38703 224 53196 252
rect 38703 221 38715 224
rect 38657 215 38715 221
rect 53190 212 53196 224
rect 53248 212 53254 264
rect 53285 255 53343 261
rect 53285 221 53297 255
rect 53331 252 53343 255
rect 55582 252 55588 264
rect 53331 224 55588 252
rect 53331 221 53343 224
rect 53285 215 53343 221
rect 55582 212 55588 224
rect 55640 212 55646 264
rect 55674 212 55680 264
rect 55732 252 55738 264
rect 58161 255 58219 261
rect 58161 252 58173 255
rect 55732 224 58173 252
rect 55732 212 55738 224
rect 58161 221 58173 224
rect 58207 221 58219 255
rect 58161 215 58219 221
rect 58253 255 58311 261
rect 58253 221 58265 255
rect 58299 252 58311 255
rect 60936 252 60964 292
rect 72973 289 72985 292
rect 73019 289 73031 323
rect 72973 283 73031 289
rect 73065 323 73123 329
rect 73065 289 73077 323
rect 73111 320 73123 323
rect 107013 323 107071 329
rect 73111 292 106964 320
rect 73111 289 73123 292
rect 73065 283 73123 289
rect 58299 224 60964 252
rect 58299 221 58311 224
rect 58253 215 58311 221
rect 61010 212 61016 264
rect 61068 252 61074 264
rect 63497 255 63555 261
rect 63497 252 63509 255
rect 61068 224 63509 252
rect 61068 212 61074 224
rect 63497 221 63509 224
rect 63543 221 63555 255
rect 63497 215 63555 221
rect 63589 255 63647 261
rect 63589 221 63601 255
rect 63635 252 63647 255
rect 66898 252 66904 264
rect 63635 224 66904 252
rect 63635 221 63647 224
rect 63589 215 63647 221
rect 66898 212 66904 224
rect 66956 212 66962 264
rect 66990 212 66996 264
rect 67048 252 67054 264
rect 67269 255 67327 261
rect 67269 252 67281 255
rect 67048 224 67281 252
rect 67048 212 67054 224
rect 67269 221 67281 224
rect 67315 221 67327 255
rect 67269 215 67327 221
rect 67358 212 67364 264
rect 67416 252 67422 264
rect 73433 255 73491 261
rect 73433 252 73445 255
rect 67416 224 73445 252
rect 67416 212 67422 224
rect 73433 221 73445 224
rect 73479 221 73491 255
rect 73433 215 73491 221
rect 73522 212 73528 264
rect 73580 252 73586 264
rect 73709 255 73767 261
rect 73580 224 73625 252
rect 73580 212 73586 224
rect 73709 221 73721 255
rect 73755 252 73767 255
rect 106829 255 106887 261
rect 106829 252 106841 255
rect 73755 224 106841 252
rect 73755 221 73767 224
rect 73709 215 73767 221
rect 106829 221 106841 224
rect 106875 221 106887 255
rect 106936 252 106964 292
rect 107013 289 107025 323
rect 107059 320 107071 323
rect 111981 323 112039 329
rect 111981 320 111993 323
rect 107059 292 111993 320
rect 107059 289 107071 292
rect 107013 283 107071 289
rect 111981 289 111993 292
rect 112027 289 112039 323
rect 183741 323 183799 329
rect 111981 283 112039 289
rect 112180 292 183692 320
rect 112180 252 112208 292
rect 106936 224 112208 252
rect 112257 255 112315 261
rect 106829 215 106887 221
rect 112257 221 112269 255
rect 112303 252 112315 255
rect 151265 255 151323 261
rect 151265 252 151277 255
rect 112303 224 151277 252
rect 112303 221 112315 224
rect 112257 215 112315 221
rect 151265 221 151277 224
rect 151311 221 151323 255
rect 151265 215 151323 221
rect 151354 212 151360 264
rect 151412 252 151418 264
rect 151722 252 151728 264
rect 151412 224 151728 252
rect 151412 212 151418 224
rect 151722 212 151728 224
rect 151780 212 151786 264
rect 151817 255 151875 261
rect 151817 221 151829 255
rect 151863 252 151875 255
rect 183557 255 183615 261
rect 183557 252 183569 255
rect 151863 224 183569 252
rect 151863 221 151875 224
rect 151817 215 151875 221
rect 183557 221 183569 224
rect 183603 221 183615 255
rect 183664 252 183692 292
rect 183741 289 183753 323
rect 183787 289 183799 323
rect 183741 283 183799 289
rect 183833 323 183891 329
rect 183833 289 183845 323
rect 183879 320 183891 323
rect 184014 320 184020 332
rect 183879 292 184020 320
rect 183879 289 183891 292
rect 183833 283 183891 289
rect 184014 280 184020 292
rect 184072 280 184078 332
rect 285769 323 285827 329
rect 285769 320 285781 323
rect 184124 292 285781 320
rect 184124 252 184152 292
rect 285769 289 285781 292
rect 285815 289 285827 323
rect 285769 283 285827 289
rect 285861 323 285919 329
rect 285861 289 285873 323
rect 285907 320 285919 323
rect 288894 320 288900 332
rect 285907 292 288900 320
rect 285907 289 285919 292
rect 285861 283 285919 289
rect 288894 280 288900 292
rect 288952 280 288958 332
rect 289173 323 289231 329
rect 289173 289 289185 323
rect 289219 320 289231 323
rect 351917 323 351975 329
rect 351917 320 351929 323
rect 289219 292 351929 320
rect 289219 289 289231 292
rect 289173 283 289231 289
rect 351917 289 351929 292
rect 351963 289 351975 323
rect 351917 283 351975 289
rect 355965 323 356023 329
rect 355965 289 355977 323
rect 356011 320 356023 323
rect 368492 320 368520 360
rect 356011 292 368520 320
rect 368569 323 368627 329
rect 356011 289 356023 292
rect 355965 283 356023 289
rect 368569 289 368581 323
rect 368615 320 368627 323
rect 372341 323 372399 329
rect 372341 320 372353 323
rect 368615 292 372353 320
rect 368615 289 368627 292
rect 368569 283 368627 289
rect 372341 289 372353 292
rect 372387 289 372399 323
rect 372448 320 372476 360
rect 372801 357 372813 391
rect 372847 357 372859 391
rect 372801 351 372859 357
rect 373169 391 373227 397
rect 373169 357 373181 391
rect 373215 388 373227 391
rect 376662 388 376668 400
rect 373215 360 376668 388
rect 373215 357 373227 360
rect 373169 351 373227 357
rect 376662 348 376668 360
rect 376720 348 376726 400
rect 377030 348 377036 400
rect 377088 388 377094 400
rect 473357 391 473415 397
rect 473357 388 473369 391
rect 377088 360 473369 388
rect 377088 348 377094 360
rect 473357 357 473369 360
rect 473403 357 473415 391
rect 473357 351 473415 357
rect 473633 391 473691 397
rect 473633 357 473645 391
rect 473679 388 473691 391
rect 507765 391 507823 397
rect 507765 388 507777 391
rect 473679 360 507777 388
rect 473679 357 473691 360
rect 473633 351 473691 357
rect 507765 357 507777 360
rect 507811 357 507823 391
rect 507765 351 507823 357
rect 507857 391 507915 397
rect 507857 357 507869 391
rect 507903 388 507915 391
rect 528186 388 528192 400
rect 507903 360 528192 388
rect 507903 357 507915 360
rect 507857 351 507915 357
rect 528186 348 528192 360
rect 528244 348 528250 400
rect 473449 323 473507 329
rect 473449 320 473461 323
rect 372448 292 473461 320
rect 372341 283 372399 289
rect 473449 289 473461 292
rect 473495 289 473507 323
rect 473449 283 473507 289
rect 473725 323 473783 329
rect 473725 289 473737 323
rect 473771 320 473783 323
rect 499666 320 499672 332
rect 473771 292 499672 320
rect 473771 289 473783 292
rect 473725 283 473783 289
rect 499666 280 499672 292
rect 499724 280 499730 332
rect 183664 224 184152 252
rect 184201 255 184259 261
rect 183557 215 183615 221
rect 184201 221 184213 255
rect 184247 252 184259 255
rect 372525 255 372583 261
rect 372525 252 372537 255
rect 184247 224 372537 252
rect 184247 221 184259 224
rect 184201 215 184259 221
rect 372525 221 372537 224
rect 372571 221 372583 255
rect 372525 215 372583 221
rect 372985 255 373043 261
rect 372985 221 372997 255
rect 373031 252 373043 255
rect 509234 252 509240 264
rect 373031 224 509240 252
rect 373031 221 373043 224
rect 372985 215 373043 221
rect 509234 212 509240 224
rect 509292 212 509298 264
rect 5583 156 26280 184
rect 28169 187 28227 193
rect 5583 153 5595 156
rect 5537 147 5595 153
rect 28169 153 28181 187
rect 28215 184 28227 187
rect 38013 187 38071 193
rect 38013 184 38025 187
rect 28215 156 38025 184
rect 28215 153 28227 156
rect 28169 147 28227 153
rect 38013 153 38025 156
rect 38059 153 38071 187
rect 38013 147 38071 153
rect 38105 187 38163 193
rect 38105 153 38117 187
rect 38151 184 38163 187
rect 39669 187 39727 193
rect 39669 184 39681 187
rect 38151 156 39681 184
rect 38151 153 38163 156
rect 38105 147 38163 153
rect 39669 153 39681 156
rect 39715 153 39727 187
rect 39669 147 39727 153
rect 39761 187 39819 193
rect 39761 153 39773 187
rect 39807 184 39819 187
rect 49789 187 49847 193
rect 49789 184 49801 187
rect 39807 156 49801 184
rect 39807 153 39819 156
rect 39761 147 39819 153
rect 49789 153 49801 156
rect 49835 153 49847 187
rect 49789 147 49847 153
rect 49878 144 49884 196
rect 49936 184 49942 196
rect 58618 184 58624 196
rect 49936 156 58624 184
rect 49936 144 49942 156
rect 58618 144 58624 156
rect 58676 144 58682 196
rect 58986 144 58992 196
rect 59044 184 59050 196
rect 60737 187 60795 193
rect 60737 184 60749 187
rect 59044 156 60749 184
rect 59044 144 59050 156
rect 60737 153 60749 156
rect 60783 153 60795 187
rect 60737 147 60795 153
rect 60829 187 60887 193
rect 60829 153 60841 187
rect 60875 184 60887 187
rect 69290 184 69296 196
rect 60875 156 69296 184
rect 60875 153 60887 156
rect 60829 147 60887 153
rect 69290 144 69296 156
rect 69348 144 69354 196
rect 69385 187 69443 193
rect 69385 153 69397 187
rect 69431 184 69443 187
rect 72513 187 72571 193
rect 72513 184 72525 187
rect 69431 156 72525 184
rect 69431 153 69443 156
rect 69385 147 69443 153
rect 72513 153 72525 156
rect 72559 153 72571 187
rect 72513 147 72571 153
rect 72605 187 72663 193
rect 72605 153 72617 187
rect 72651 184 72663 187
rect 76469 187 76527 193
rect 76469 184 76481 187
rect 72651 156 76481 184
rect 72651 153 72663 156
rect 72605 147 72663 153
rect 76469 153 76481 156
rect 76515 153 76527 187
rect 76469 147 76527 153
rect 76561 187 76619 193
rect 76561 153 76573 187
rect 76607 184 76619 187
rect 83369 187 83427 193
rect 83369 184 83381 187
rect 76607 156 83381 184
rect 76607 153 76619 156
rect 76561 147 76619 153
rect 83369 153 83381 156
rect 83415 153 83427 187
rect 83369 147 83427 153
rect 83458 144 83464 196
rect 83516 184 83522 196
rect 84381 187 84439 193
rect 84381 184 84393 187
rect 83516 156 84393 184
rect 83516 144 83522 156
rect 84381 153 84393 156
rect 84427 153 84439 187
rect 84381 147 84439 153
rect 84470 144 84476 196
rect 84528 184 84534 196
rect 84565 187 84623 193
rect 84565 184 84577 187
rect 84528 156 84577 184
rect 84528 144 84534 156
rect 84565 153 84577 156
rect 84611 153 84623 187
rect 84565 147 84623 153
rect 84654 144 84660 196
rect 84712 184 84718 196
rect 87690 184 87696 196
rect 84712 156 87696 184
rect 84712 144 84718 156
rect 87690 144 87696 156
rect 87748 144 87754 196
rect 87785 187 87843 193
rect 87785 153 87797 187
rect 87831 184 87843 187
rect 91465 187 91523 193
rect 91465 184 91477 187
rect 87831 156 91477 184
rect 87831 153 87843 156
rect 87785 147 87843 153
rect 91465 153 91477 156
rect 91511 153 91523 187
rect 91465 147 91523 153
rect 91557 187 91615 193
rect 91557 153 91569 187
rect 91603 184 91615 187
rect 111797 187 111855 193
rect 111797 184 111809 187
rect 91603 156 111809 184
rect 91603 153 91615 156
rect 91557 147 91615 153
rect 111797 153 111809 156
rect 111843 153 111855 187
rect 111797 147 111855 153
rect 111889 187 111947 193
rect 111889 153 111901 187
rect 111935 184 111947 187
rect 112162 184 112168 196
rect 111935 156 112168 184
rect 111935 153 111947 156
rect 111889 147 111947 153
rect 112162 144 112168 156
rect 112220 144 112226 196
rect 112349 187 112407 193
rect 112349 153 112361 187
rect 112395 184 112407 187
rect 183462 184 183468 196
rect 112395 156 183468 184
rect 112395 153 112407 156
rect 112349 147 112407 153
rect 183462 144 183468 156
rect 183520 144 183526 196
rect 183741 187 183799 193
rect 183741 153 183753 187
rect 183787 184 183799 187
rect 183922 184 183928 196
rect 183787 156 183928 184
rect 183787 153 183799 156
rect 183741 147 183799 153
rect 183922 144 183928 156
rect 183980 144 183986 196
rect 184293 187 184351 193
rect 184293 153 184305 187
rect 184339 184 184351 187
rect 335357 187 335415 193
rect 335357 184 335369 187
rect 184339 156 335369 184
rect 184339 153 184351 156
rect 184293 147 184351 153
rect 335357 153 335369 156
rect 335403 153 335415 187
rect 335357 147 335415 153
rect 335633 187 335691 193
rect 335633 153 335645 187
rect 335679 184 335691 187
rect 347501 187 347559 193
rect 347501 184 347513 187
rect 335679 156 347513 184
rect 335679 153 335691 156
rect 335633 147 335691 153
rect 347501 153 347513 156
rect 347547 153 347559 187
rect 347501 147 347559 153
rect 347685 187 347743 193
rect 347685 153 347697 187
rect 347731 184 347743 187
rect 372341 187 372399 193
rect 372341 184 372353 187
rect 347731 156 372353 184
rect 347731 153 347743 156
rect 347685 147 347743 153
rect 372341 153 372353 156
rect 372387 153 372399 187
rect 372341 147 372399 153
rect 373261 187 373319 193
rect 373261 153 373273 187
rect 373307 184 373319 187
rect 376757 187 376815 193
rect 376757 184 376769 187
rect 373307 156 376769 184
rect 373307 153 373319 156
rect 373261 147 373319 153
rect 376757 153 376769 156
rect 376803 153 376815 187
rect 376757 147 376815 153
rect 376941 187 376999 193
rect 376941 153 376953 187
rect 376987 184 376999 187
rect 473449 187 473507 193
rect 473449 184 473461 187
rect 376987 156 473461 184
rect 376987 153 376999 156
rect 376941 147 376999 153
rect 473449 153 473461 156
rect 473495 153 473507 187
rect 473449 147 473507 153
rect 473633 187 473691 193
rect 473633 153 473645 187
rect 473679 184 473691 187
rect 569218 184 569224 196
rect 473679 156 569224 184
rect 473679 153 473691 156
rect 473633 147 473691 153
rect 569218 144 569224 156
rect 569276 144 569282 196
rect 5445 119 5503 125
rect 5445 116 5457 119
rect 5276 88 5457 116
rect 1765 51 1823 57
rect 1765 17 1777 51
rect 1811 48 1823 51
rect 5276 48 5304 88
rect 5445 85 5457 88
rect 5491 85 5503 119
rect 5445 79 5503 85
rect 5629 119 5687 125
rect 5629 85 5641 119
rect 5675 116 5687 119
rect 5997 119 6055 125
rect 5675 88 5948 116
rect 5675 85 5687 88
rect 5629 79 5687 85
rect 1811 20 5304 48
rect 5920 48 5948 88
rect 5997 85 6009 119
rect 6043 116 6055 119
rect 9769 119 9827 125
rect 9769 116 9781 119
rect 6043 88 9781 116
rect 6043 85 6055 88
rect 5997 79 6055 85
rect 9769 85 9781 88
rect 9815 85 9827 119
rect 9769 79 9827 85
rect 9858 76 9864 128
rect 9916 116 9922 128
rect 10505 119 10563 125
rect 10505 116 10517 119
rect 9916 88 10517 116
rect 9916 76 9922 88
rect 10505 85 10517 88
rect 10551 85 10563 119
rect 10505 79 10563 85
rect 10597 119 10655 125
rect 10597 85 10609 119
rect 10643 116 10655 119
rect 44358 116 44364 128
rect 10643 88 44364 116
rect 10643 85 10655 88
rect 10597 79 10655 85
rect 44358 76 44364 88
rect 44416 76 44422 128
rect 46290 76 46296 128
rect 46348 116 46354 128
rect 55309 119 55367 125
rect 55309 116 55321 119
rect 46348 88 55321 116
rect 46348 76 46354 88
rect 55309 85 55321 88
rect 55355 85 55367 119
rect 55309 79 55367 85
rect 55398 76 55404 128
rect 55456 116 55462 128
rect 92109 119 92167 125
rect 92109 116 92121 119
rect 55456 88 92121 116
rect 55456 76 55462 88
rect 92109 85 92121 88
rect 92155 85 92167 119
rect 92109 79 92167 85
rect 92477 119 92535 125
rect 92477 85 92489 119
rect 92523 116 92535 119
rect 183557 119 183615 125
rect 183557 116 183569 119
rect 92523 88 183569 116
rect 92523 85 92535 88
rect 92477 79 92535 85
rect 183557 85 183569 88
rect 183603 85 183615 119
rect 184017 119 184075 125
rect 183557 79 183615 85
rect 183664 88 183876 116
rect 13078 48 13084 60
rect 5920 20 13084 48
rect 1811 17 1823 20
rect 1765 11 1823 17
rect 13078 8 13084 20
rect 13136 8 13142 60
rect 13173 51 13231 57
rect 13173 17 13185 51
rect 13219 48 13231 51
rect 14461 51 14519 57
rect 14461 48 14473 51
rect 13219 20 14473 48
rect 13219 17 13231 20
rect 13173 11 13231 17
rect 14461 17 14473 20
rect 14507 17 14519 51
rect 14461 11 14519 17
rect 17402 8 17408 60
rect 17460 48 17466 60
rect 183664 48 183692 88
rect 17460 20 183692 48
rect 183848 48 183876 88
rect 184017 85 184029 119
rect 184063 116 184075 119
rect 335541 119 335599 125
rect 335541 116 335553 119
rect 184063 88 335553 116
rect 184063 85 184075 88
rect 184017 79 184075 85
rect 335541 85 335553 88
rect 335587 85 335599 119
rect 335541 79 335599 85
rect 335725 119 335783 125
rect 335725 85 335737 119
rect 335771 116 335783 119
rect 347409 119 347467 125
rect 347409 116 347421 119
rect 335771 88 347421 116
rect 335771 85 335783 88
rect 335725 79 335783 85
rect 347409 85 347421 88
rect 347455 85 347467 119
rect 347409 79 347467 85
rect 347593 119 347651 125
rect 347593 85 347605 119
rect 347639 116 347651 119
rect 372433 119 372491 125
rect 372433 116 372445 119
rect 347639 88 372445 116
rect 347639 85 347651 88
rect 347593 79 347651 85
rect 372433 85 372445 88
rect 372479 85 372491 119
rect 372433 79 372491 85
rect 372709 119 372767 125
rect 372709 85 372721 119
rect 372755 116 372767 119
rect 430761 119 430819 125
rect 430761 116 430773 119
rect 372755 88 430773 116
rect 372755 85 372767 88
rect 372709 79 372767 85
rect 430761 85 430773 88
rect 430807 85 430819 119
rect 430761 79 430819 85
rect 436097 119 436155 125
rect 436097 85 436109 119
rect 436143 116 436155 119
rect 568850 116 568856 128
rect 436143 88 568856 116
rect 436143 85 436155 88
rect 436097 79 436155 85
rect 568850 76 568856 88
rect 568908 76 568914 128
rect 335449 51 335507 57
rect 335449 48 335461 51
rect 183848 20 335461 48
rect 17460 8 17466 20
rect 335449 17 335461 20
rect 335495 17 335507 51
rect 335449 11 335507 17
rect 335633 51 335691 57
rect 335633 17 335645 51
rect 335679 48 335691 51
rect 347317 51 347375 57
rect 347317 48 347329 51
rect 335679 20 347329 48
rect 335679 17 335691 20
rect 335633 11 335691 17
rect 347317 17 347329 20
rect 347363 17 347375 51
rect 347317 11 347375 17
rect 347685 51 347743 57
rect 347685 17 347697 51
rect 347731 48 347743 51
rect 473354 48 473360 60
rect 347731 20 473360 48
rect 347731 17 347743 20
rect 347685 11 347743 17
rect 473354 8 473360 20
rect 473412 8 473418 60
rect 473722 8 473728 60
rect 473780 48 473786 60
rect 568301 51 568359 57
rect 568301 48 568313 51
rect 473780 20 568313 48
rect 473780 8 473786 20
rect 568301 17 568313 20
rect 568347 17 568359 51
rect 568301 11 568359 17
<< via1 >>
rect 129648 700680 129700 700732
rect 170312 700680 170364 700732
rect 105452 700612 105504 700664
rect 106188 700612 106240 700664
rect 110328 700612 110380 700664
rect 235172 700612 235224 700664
rect 89628 700544 89680 700596
rect 300124 700544 300176 700596
rect 40500 700476 40552 700528
rect 41328 700476 41380 700528
rect 70308 700476 70360 700528
rect 364984 700476 365036 700528
rect 50988 700408 51040 700460
rect 429844 700408 429896 700460
rect 31668 700340 31720 700392
rect 494796 700340 494848 700392
rect 10968 700272 11020 700324
rect 559656 700272 559708 700324
rect 30380 684428 30432 684480
rect 31668 684428 31720 684480
rect 50068 684428 50120 684480
rect 50988 684428 51040 684480
rect 128636 684428 128688 684480
rect 129648 684428 129700 684480
rect 109040 684020 109092 684072
rect 110328 684020 110380 684072
rect 106188 683816 106240 683868
rect 148324 683816 148376 683868
rect 41328 683748 41380 683800
rect 168012 683748 168064 683800
rect 285956 683204 286008 683256
rect 295248 683204 295300 683256
rect 364524 683204 364576 683256
rect 375380 683204 375432 683256
rect 384212 683204 384264 683256
rect 391204 683204 391256 683256
rect 403900 683204 403952 683256
rect 408408 683204 408460 683256
rect 462872 683204 462924 683256
rect 471980 683204 472032 683256
rect 482468 683204 482520 683256
rect 494060 683204 494112 683256
rect 187608 683136 187660 683188
rect 569868 683136 569920 683188
rect 305920 680960 305972 681012
rect 327632 680960 327684 681012
rect 379428 680552 379480 680604
rect 381636 680552 381688 680604
rect 557448 680552 557500 680604
rect 563244 680552 563296 680604
rect 226708 680348 226760 680400
rect 246212 680348 246264 680400
rect 207020 680323 207072 680332
rect 207020 680289 207029 680323
rect 207029 680289 207063 680323
rect 207063 680289 207072 680323
rect 207020 680280 207072 680289
rect 1952 679804 2004 679856
rect 3424 679736 3476 679788
rect 2504 679600 2556 679652
rect 265900 680348 265952 680400
rect 380072 680391 380124 680400
rect 380072 680357 380081 680391
rect 380081 680357 380115 680391
rect 380115 680357 380124 680391
rect 380072 680348 380124 680357
rect 391204 680348 391256 680400
rect 394700 680391 394752 680400
rect 394700 680357 394709 680391
rect 394709 680357 394743 680391
rect 394743 680357 394752 680391
rect 394700 680348 394752 680357
rect 403164 680391 403216 680400
rect 403164 680357 403173 680391
rect 403173 680357 403207 680391
rect 403207 680357 403216 680391
rect 403164 680348 403216 680357
rect 295248 680280 295300 680332
rect 296720 680280 296772 680332
rect 327632 680280 327684 680332
rect 364800 680323 364852 680332
rect 364800 680289 364809 680323
rect 364809 680289 364843 680323
rect 364843 680289 364852 680323
rect 364800 680280 364852 680289
rect 370228 680323 370280 680332
rect 370228 680289 370237 680323
rect 370237 680289 370271 680323
rect 370271 680289 370280 680323
rect 370228 680280 370280 680289
rect 375380 680280 375432 680332
rect 408408 680280 408460 680332
rect 463792 680416 463844 680468
rect 466644 680416 466696 680468
rect 559380 680416 559432 680468
rect 412732 680391 412784 680400
rect 412732 680357 412741 680391
rect 412741 680357 412775 680391
rect 412775 680357 412784 680391
rect 412732 680348 412784 680357
rect 418620 680391 418672 680400
rect 418620 680357 418629 680391
rect 418629 680357 418663 680391
rect 418663 680357 418672 680391
rect 418620 680348 418672 680357
rect 423588 680348 423640 680400
rect 428188 680391 428240 680400
rect 428188 680357 428197 680391
rect 428197 680357 428231 680391
rect 428231 680357 428240 680391
rect 428188 680348 428240 680357
rect 437756 680391 437808 680400
rect 437756 680357 437765 680391
rect 437765 680357 437799 680391
rect 437799 680357 437808 680391
rect 437756 680348 437808 680357
rect 443552 680391 443604 680400
rect 443552 680357 443561 680391
rect 443561 680357 443595 680391
rect 443595 680357 443604 680391
rect 443552 680348 443604 680357
rect 451372 680391 451424 680400
rect 451372 680357 451381 680391
rect 451381 680357 451415 680391
rect 451415 680357 451424 680391
rect 451372 680348 451424 680357
rect 457168 680391 457220 680400
rect 457168 680357 457177 680391
rect 457177 680357 457211 680391
rect 457211 680357 457220 680391
rect 457168 680348 457220 680357
rect 466552 680391 466604 680400
rect 466552 680357 466561 680391
rect 466561 680357 466595 680391
rect 466595 680357 466604 680391
rect 466552 680348 466604 680357
rect 471980 680348 472032 680400
rect 494060 680391 494112 680400
rect 494060 680357 494069 680391
rect 494069 680357 494103 680391
rect 494103 680357 494112 680391
rect 494060 680348 494112 680357
rect 495440 680391 495492 680400
rect 495440 680357 495449 680391
rect 495449 680357 495483 680391
rect 495483 680357 495492 680391
rect 502248 680391 502300 680400
rect 495440 680348 495492 680357
rect 502248 680357 502257 680391
rect 502257 680357 502291 680391
rect 502291 680357 502300 680391
rect 502248 680348 502300 680357
rect 505928 680391 505980 680400
rect 505928 680357 505937 680391
rect 505937 680357 505971 680391
rect 505971 680357 505980 680391
rect 505928 680348 505980 680357
rect 515404 680391 515456 680400
rect 515404 680357 515413 680391
rect 515413 680357 515447 680391
rect 515447 680357 515456 680391
rect 515404 680348 515456 680357
rect 522120 680391 522172 680400
rect 522120 680357 522129 680391
rect 522129 680357 522163 680391
rect 522163 680357 522172 680391
rect 522120 680348 522172 680357
rect 524420 680391 524472 680400
rect 524420 680357 524429 680391
rect 524429 680357 524463 680391
rect 524463 680357 524472 680391
rect 534356 680391 534408 680400
rect 524420 680348 524472 680357
rect 534356 680357 534365 680391
rect 534365 680357 534399 680391
rect 534399 680357 534408 680391
rect 534356 680348 534408 680357
rect 541808 680348 541860 680400
rect 544016 680391 544068 680400
rect 544016 680357 544025 680391
rect 544025 680357 544059 680391
rect 544059 680357 544068 680391
rect 544016 680348 544068 680357
rect 481180 680323 481232 680332
rect 481180 680289 481189 680323
rect 481189 680289 481223 680323
rect 481223 680289 481232 680323
rect 481180 680280 481232 680289
rect 485780 680323 485832 680332
rect 485780 680289 485789 680323
rect 485789 680289 485823 680323
rect 485823 680289 485832 680323
rect 485780 680280 485832 680289
rect 554780 680280 554832 680332
rect 554872 680323 554924 680332
rect 554872 680289 554881 680323
rect 554881 680289 554915 680323
rect 554915 680289 554924 680323
rect 554872 680280 554924 680289
rect 558552 680280 558604 680332
rect 559196 680323 559248 680332
rect 559196 680289 559205 680323
rect 559205 680289 559239 680323
rect 559239 680289 559248 680323
rect 559196 680280 559248 680289
rect 560760 680323 560812 680332
rect 560760 680289 560769 680323
rect 560769 680289 560803 680323
rect 560803 680289 560812 680323
rect 560760 680280 560812 680289
rect 561588 680323 561640 680332
rect 561588 680289 561597 680323
rect 561597 680289 561631 680323
rect 561631 680289 561640 680323
rect 561588 680280 561640 680289
rect 561772 680323 561824 680332
rect 561772 680289 561781 680323
rect 561781 680289 561815 680323
rect 561815 680289 561824 680323
rect 561772 680280 561824 680289
rect 561864 680323 561916 680332
rect 561864 680289 561873 680323
rect 561873 680289 561907 680323
rect 561907 680289 561916 680323
rect 562508 680323 562560 680332
rect 561864 680280 561916 680289
rect 562508 680289 562517 680323
rect 562517 680289 562551 680323
rect 562551 680289 562560 680323
rect 562508 680280 562560 680289
rect 566372 680280 566424 680332
rect 568396 679600 568448 679652
rect 3700 679124 3752 679176
rect 572720 679124 572772 679176
rect 2228 679056 2280 679108
rect 569224 679056 569276 679108
rect 1860 678988 1912 679040
rect 571432 678988 571484 679040
rect 204 677492 256 677544
rect 1400 677492 1452 677544
rect 571432 677492 571484 677544
rect 578148 677492 578200 677544
rect 1952 676132 2004 676184
rect 1952 675996 2004 676048
rect 578148 674772 578200 674824
rect 580172 674772 580224 674824
rect 569960 659243 570012 659252
rect 569960 659209 569969 659243
rect 569969 659209 570003 659243
rect 570003 659209 570012 659243
rect 569960 659200 570012 659209
rect 569960 654168 570012 654220
rect 577504 654168 577556 654220
rect 569960 654075 570012 654084
rect 569960 654041 569969 654075
rect 569969 654041 570003 654075
rect 570003 654041 570012 654075
rect 569960 654032 570012 654041
rect 1860 648592 1912 648644
rect 1952 648592 2004 648644
rect 1952 648091 2004 648100
rect 1952 648057 1961 648091
rect 1961 648057 1995 648091
rect 1995 648057 2004 648091
rect 1952 648048 2004 648057
rect 1952 642608 2004 642660
rect 1952 641792 2004 641844
rect 1952 641588 2004 641640
rect 1952 639319 2004 639328
rect 1952 639285 1961 639319
rect 1961 639285 1995 639319
rect 1995 639285 2004 639319
rect 1952 639276 2004 639285
rect 1860 633471 1912 633480
rect 1860 633437 1869 633471
rect 1869 633437 1903 633471
rect 1903 633437 1912 633471
rect 1860 633428 1912 633437
rect 569960 630164 570012 630216
rect 572720 630164 572772 630216
rect 577504 627852 577556 627904
rect 579712 627852 579764 627904
rect 1584 618264 1636 618316
rect 1676 618264 1728 618316
rect 1860 618264 1912 618316
rect 1952 618264 2004 618316
rect 569960 609628 570012 609680
rect 570328 609628 570380 609680
rect 569960 609220 570012 609272
rect 570052 609220 570104 609272
rect 1952 608676 2004 608728
rect 1860 608540 1912 608592
rect 1952 602352 2004 602404
rect 1952 602123 2004 602132
rect 1952 602089 1961 602123
rect 1961 602089 1995 602123
rect 1995 602089 2004 602123
rect 1952 602080 2004 602089
rect 1952 601944 2004 601996
rect 1952 601060 2004 601112
rect 1584 600924 1636 600976
rect 1952 600924 2004 600976
rect 1952 600516 2004 600568
rect 1952 599879 2004 599888
rect 1952 599845 1961 599879
rect 1961 599845 1995 599879
rect 1995 599845 2004 599879
rect 1952 599836 2004 599845
rect 1952 599700 2004 599752
rect 1952 596980 2004 597032
rect 1676 591948 1728 592000
rect 1860 591948 1912 592000
rect 1952 580456 2004 580508
rect 1952 580227 2004 580236
rect 1952 580193 1961 580227
rect 1961 580193 1995 580227
rect 1995 580193 2004 580227
rect 1952 580184 2004 580193
rect 1584 577260 1636 577312
rect 1952 577260 2004 577312
rect 574744 574744 574796 574796
rect 580264 574744 580316 574796
rect 569960 571344 570012 571396
rect 572720 571344 572772 571396
rect 1952 569304 2004 569356
rect 1768 569100 1820 569152
rect 1860 566627 1912 566636
rect 1860 566593 1869 566627
rect 1869 566593 1903 566627
rect 1903 566593 1912 566627
rect 1860 566584 1912 566593
rect 1952 565496 2004 565548
rect 1952 564408 2004 564460
rect 1308 564068 1360 564120
rect 1952 564068 2004 564120
rect 1860 563728 1912 563780
rect 1952 563388 2004 563440
rect 1952 563116 2004 563168
rect 569960 563048 570012 563100
rect 574744 563048 574796 563100
rect 1952 561076 2004 561128
rect 1584 556180 1636 556232
rect 1952 556180 2004 556232
rect 569960 552075 570012 552084
rect 569960 552041 569969 552075
rect 569969 552041 570003 552075
rect 570003 552041 570012 552075
rect 569960 552032 570012 552041
rect 569960 551828 570012 551880
rect 572720 551828 572772 551880
rect 569960 551055 570012 551064
rect 569960 551021 569969 551055
rect 569969 551021 570003 551055
rect 570003 551021 570012 551055
rect 569960 551012 570012 551021
rect 1860 547680 1912 547732
rect 1860 534012 1912 534064
rect 1860 533808 1912 533860
rect 573364 532720 573416 532772
rect 580172 532720 580224 532772
rect 569960 531088 570012 531140
rect 569960 530995 570012 531004
rect 569960 530961 569969 530995
rect 569969 530961 570003 530995
rect 570003 530961 570012 530995
rect 569960 530952 570012 530961
rect 1952 529227 2004 529236
rect 1952 529193 1961 529227
rect 1961 529193 1995 529227
rect 1995 529193 2004 529227
rect 1952 529184 2004 529193
rect 569960 528887 570012 528896
rect 569960 528853 569969 528887
rect 569969 528853 570003 528887
rect 570003 528853 570012 528887
rect 569960 528844 570012 528853
rect 569960 528708 570012 528760
rect 1952 527688 2004 527740
rect 1952 527144 2004 527196
rect 1676 527119 1728 527128
rect 1676 527085 1685 527119
rect 1685 527085 1719 527119
rect 1719 527085 1728 527119
rect 1676 527076 1728 527085
rect 1768 526940 1820 526992
rect 1952 526464 2004 526516
rect 1584 526328 1636 526380
rect 1952 526328 2004 526380
rect 1952 526124 2004 526176
rect 569960 522631 570012 522640
rect 569960 522597 569969 522631
rect 569969 522597 570003 522631
rect 570003 522597 570012 522631
rect 569960 522588 570012 522597
rect 1952 522452 2004 522504
rect 569960 522452 570012 522504
rect 1952 522316 2004 522368
rect 569960 522316 570012 522368
rect 573364 522316 573416 522368
rect 569960 521024 570012 521076
rect 569960 518483 570012 518492
rect 569960 518449 569969 518483
rect 569969 518449 570003 518483
rect 570003 518449 570012 518483
rect 569960 518440 570012 518449
rect 1952 510663 2004 510672
rect 1952 510629 1961 510663
rect 1961 510629 1995 510663
rect 1995 510629 2004 510663
rect 1952 510620 2004 510629
rect 1952 510051 2004 510060
rect 1952 510017 1961 510051
rect 1961 510017 1995 510051
rect 1995 510017 2004 510051
rect 1952 510008 2004 510017
rect 1768 509872 1820 509924
rect 1952 509872 2004 509924
rect 1676 509532 1728 509584
rect 1952 507288 2004 507340
rect 1952 507152 2004 507204
rect 1952 506064 2004 506116
rect 1584 505180 1636 505232
rect 1952 505180 2004 505232
rect 569960 505155 570012 505164
rect 569960 505121 569969 505155
rect 569969 505121 570003 505155
rect 570003 505121 570012 505155
rect 569960 505112 570012 505121
rect 1952 504772 2004 504824
rect 1860 504475 1912 504484
rect 1860 504441 1869 504475
rect 1869 504441 1903 504475
rect 1903 504441 1912 504475
rect 1860 504432 1912 504441
rect 569960 504160 570012 504212
rect 1768 504135 1820 504144
rect 1768 504101 1777 504135
rect 1777 504101 1811 504135
rect 1811 504101 1820 504135
rect 1768 504092 1820 504101
rect 569960 503140 570012 503192
rect 569960 503047 570012 503056
rect 569960 503013 569969 503047
rect 569969 503013 570003 503047
rect 570003 503013 570012 503047
rect 569960 503004 570012 503013
rect 1676 502299 1728 502308
rect 1676 502265 1685 502299
rect 1685 502265 1719 502299
rect 1719 502265 1728 502299
rect 1676 502256 1728 502265
rect 1952 502188 2004 502240
rect 1952 501780 2004 501832
rect 1768 497539 1820 497548
rect 1768 497505 1777 497539
rect 1777 497505 1811 497539
rect 1811 497505 1820 497539
rect 1768 497496 1820 497505
rect 1952 497539 2004 497548
rect 1952 497505 1961 497539
rect 1961 497505 1995 497539
rect 1995 497505 2004 497539
rect 1952 497496 2004 497505
rect 1860 493348 1912 493400
rect 569960 487092 570012 487144
rect 579804 487092 579856 487144
rect 569960 486956 570012 487008
rect 570144 486956 570196 487008
rect 1768 483692 1820 483744
rect 1952 479544 2004 479596
rect 1952 479340 2004 479392
rect 1952 474691 2004 474700
rect 1952 474657 1961 474691
rect 1961 474657 1995 474691
rect 1995 474657 2004 474691
rect 1952 474648 2004 474657
rect 1860 474079 1912 474088
rect 1860 474045 1869 474079
rect 1869 474045 1903 474079
rect 1903 474045 1912 474079
rect 1860 474036 1912 474045
rect 1676 472744 1728 472796
rect 1952 472744 2004 472796
rect 1768 472107 1820 472116
rect 1768 472073 1777 472107
rect 1777 472073 1811 472107
rect 1811 472073 1820 472107
rect 1768 472064 1820 472073
rect 1032 469752 1084 469804
rect 1952 469752 2004 469804
rect 569960 468571 570012 468580
rect 569960 468537 569969 468571
rect 569969 468537 570003 468571
rect 570003 468537 570012 468571
rect 569960 468528 570012 468537
rect 1952 468256 2004 468308
rect 569960 468256 570012 468308
rect 1952 468052 2004 468104
rect 1952 467576 2004 467628
rect 569960 467576 570012 467628
rect 570052 467075 570104 467084
rect 570052 467041 570061 467075
rect 570061 467041 570095 467075
rect 570095 467041 570104 467075
rect 570052 467032 570104 467041
rect 570052 466828 570104 466880
rect 570052 465332 570104 465384
rect 569960 465196 570012 465248
rect 570144 465196 570196 465248
rect 570144 465060 570196 465112
rect 1952 464924 2004 464976
rect 569868 464244 569920 464296
rect 570052 464108 570104 464160
rect 569960 463972 570012 464024
rect 569960 463836 570012 463888
rect 569960 463700 570012 463752
rect 569960 463564 570012 463616
rect 570052 462748 570104 462800
rect 1952 462383 2004 462392
rect 1952 462349 1961 462383
rect 1961 462349 1995 462383
rect 1995 462349 2004 462383
rect 1952 462340 2004 462349
rect 569960 461703 570012 461712
rect 569960 461669 569969 461703
rect 569969 461669 570003 461703
rect 570003 461669 570012 461703
rect 569960 461660 570012 461669
rect 569960 461431 570012 461440
rect 569960 461397 569969 461431
rect 569969 461397 570003 461431
rect 570003 461397 570012 461431
rect 569960 461388 570012 461397
rect 1400 459824 1452 459876
rect 1860 459824 1912 459876
rect 1952 454631 2004 454640
rect 1952 454597 1961 454631
rect 1961 454597 1995 454631
rect 1995 454597 2004 454631
rect 1952 454588 2004 454597
rect 1768 450848 1820 450900
rect 1952 450848 2004 450900
rect 1952 450712 2004 450764
rect 1952 450032 2004 450084
rect 1952 449896 2004 449948
rect 569960 449352 570012 449404
rect 1860 449191 1912 449200
rect 1860 449157 1869 449191
rect 1869 449157 1903 449191
rect 1903 449157 1912 449191
rect 1860 449148 1912 449157
rect 569960 449148 570012 449200
rect 1860 449012 1912 449064
rect 1952 448740 2004 448792
rect 1676 448715 1728 448724
rect 1676 448681 1685 448715
rect 1685 448681 1719 448715
rect 1719 448681 1728 448715
rect 1676 448672 1728 448681
rect 1400 448604 1452 448656
rect 1952 448604 2004 448656
rect 1952 448468 2004 448520
rect 1952 447924 2004 447976
rect 1952 447788 2004 447840
rect 1860 442280 1912 442332
rect 569960 441600 570012 441652
rect 1952 441396 2004 441448
rect 1860 440963 1912 440972
rect 1860 440929 1869 440963
rect 1869 440929 1903 440963
rect 1903 440929 1912 440963
rect 1860 440920 1912 440929
rect 1952 439195 2004 439204
rect 1952 439161 1961 439195
rect 1961 439161 1995 439195
rect 1995 439161 2004 439195
rect 1952 439152 2004 439161
rect 574744 438880 574796 438932
rect 580172 438880 580224 438932
rect 570052 436815 570104 436824
rect 570052 436781 570061 436815
rect 570061 436781 570095 436815
rect 570095 436781 570104 436815
rect 570052 436772 570104 436781
rect 1952 434231 2004 434240
rect 1952 434197 1961 434231
rect 1961 434197 1995 434231
rect 1995 434197 2004 434231
rect 1952 434188 2004 434197
rect 569960 432531 570012 432540
rect 569960 432497 569969 432531
rect 569969 432497 570003 432531
rect 570003 432497 570012 432531
rect 569960 432488 570012 432497
rect 1676 432216 1728 432268
rect 1952 432216 2004 432268
rect 1952 425731 2004 425740
rect 1952 425697 1961 425731
rect 1961 425697 1995 425731
rect 1995 425697 2004 425731
rect 1952 425688 2004 425697
rect 1400 425552 1452 425604
rect 1768 425552 1820 425604
rect 1400 419840 1452 419892
rect 1676 419840 1728 419892
rect 569960 418276 570012 418328
rect 569960 418183 570012 418192
rect 569960 418149 569969 418183
rect 569969 418149 570003 418183
rect 570003 418149 570012 418183
rect 569960 418140 570012 418149
rect 1860 414944 1912 414996
rect 1952 414987 2004 414996
rect 1952 414953 1961 414987
rect 1961 414953 1995 414987
rect 1995 414953 2004 414987
rect 1952 414944 2004 414953
rect 1860 414740 1912 414792
rect 1400 414604 1452 414656
rect 1676 414604 1728 414656
rect 570604 411952 570656 412004
rect 572720 411952 572772 412004
rect 1952 407303 2004 407312
rect 1952 407269 1961 407303
rect 1961 407269 1995 407303
rect 1995 407269 2004 407303
rect 1952 407260 2004 407269
rect 569960 407056 570012 407108
rect 570052 407056 570104 407108
rect 1952 405671 2004 405680
rect 1952 405637 1961 405671
rect 1961 405637 1995 405671
rect 1995 405637 2004 405671
rect 1952 405628 2004 405637
rect 1860 405603 1912 405612
rect 1860 405569 1869 405603
rect 1869 405569 1903 405603
rect 1903 405569 1912 405603
rect 1860 405560 1912 405569
rect 1400 405424 1452 405476
rect 1768 405424 1820 405476
rect 569960 402271 570012 402280
rect 569960 402237 569969 402271
rect 569969 402237 570003 402271
rect 570003 402237 570012 402271
rect 569960 402228 570012 402237
rect 569960 401616 570012 401668
rect 570604 401616 570656 401668
rect 570052 399508 570104 399560
rect 1400 398420 1452 398472
rect 1768 398420 1820 398472
rect 569960 396788 570012 396840
rect 569960 394952 570012 395004
rect 570052 394612 570104 394664
rect 570236 394612 570288 394664
rect 1860 393975 1912 393984
rect 1860 393941 1869 393975
rect 1869 393941 1903 393975
rect 1903 393941 1912 393975
rect 1860 393932 1912 393941
rect 569960 393796 570012 393848
rect 569960 393703 570012 393712
rect 569960 393669 569969 393703
rect 569969 393669 570003 393703
rect 570003 393669 570012 393703
rect 569960 393660 570012 393669
rect 1952 393499 2004 393508
rect 1952 393465 1961 393499
rect 1961 393465 1995 393499
rect 1995 393465 2004 393499
rect 1952 393456 2004 393465
rect 569960 393116 570012 393168
rect 569960 392912 570012 392964
rect 569960 392708 570012 392760
rect 569960 392572 570012 392624
rect 570328 392572 570380 392624
rect 569960 392300 570012 392352
rect 574836 391960 574888 392012
rect 580172 391960 580224 392012
rect 569960 389988 570012 390040
rect 569960 389895 570012 389904
rect 569960 389861 569969 389895
rect 569969 389861 570003 389895
rect 570003 389861 570012 389895
rect 569960 389852 570012 389861
rect 569960 389036 570012 389088
rect 569960 388492 570012 388544
rect 569960 388356 570012 388408
rect 570236 388356 570288 388408
rect 1952 387336 2004 387388
rect 1952 387200 2004 387252
rect 1400 387107 1452 387116
rect 1400 387073 1409 387107
rect 1409 387073 1443 387107
rect 1443 387073 1452 387107
rect 1400 387064 1452 387073
rect 1768 387064 1820 387116
rect 1952 387107 2004 387116
rect 1952 387073 1961 387107
rect 1961 387073 1995 387107
rect 1995 387073 2004 387107
rect 1952 387064 2004 387073
rect 1400 386928 1452 386980
rect 1768 386928 1820 386980
rect 1952 386928 2004 386980
rect 569960 382823 570012 382832
rect 569960 382789 569969 382823
rect 569969 382789 570003 382823
rect 570003 382789 570012 382823
rect 569960 382780 570012 382789
rect 569960 382644 570012 382696
rect 569960 381828 570012 381880
rect 1952 381148 2004 381200
rect 1768 380672 1820 380724
rect 1952 380672 2004 380724
rect 1400 380536 1452 380588
rect 1768 380536 1820 380588
rect 1952 379108 2004 379160
rect 1952 378972 2004 379024
rect 1952 376728 2004 376780
rect 569960 376703 570012 376712
rect 569960 376669 569969 376703
rect 569969 376669 570003 376703
rect 570003 376669 570012 376703
rect 569960 376660 570012 376669
rect 570144 376660 570196 376712
rect 569960 376524 570012 376576
rect 1952 370651 2004 370660
rect 1952 370617 1961 370651
rect 1961 370617 1995 370651
rect 1995 370617 2004 370651
rect 1952 370608 2004 370617
rect 1676 370515 1728 370524
rect 1676 370481 1685 370515
rect 1685 370481 1719 370515
rect 1719 370481 1728 370515
rect 1676 370472 1728 370481
rect 1952 370336 2004 370388
rect 1952 370200 2004 370252
rect 569960 369724 570012 369776
rect 569960 369427 570012 369436
rect 569960 369393 569969 369427
rect 569969 369393 570003 369427
rect 570003 369393 570012 369427
rect 569960 369384 570012 369393
rect 1952 369248 2004 369300
rect 569960 368339 570012 368348
rect 569960 368305 569969 368339
rect 569969 368305 570003 368339
rect 570003 368305 570012 368339
rect 569960 368296 570012 368305
rect 569960 368024 570012 368076
rect 570144 368024 570196 368076
rect 1676 367795 1728 367804
rect 1676 367761 1685 367795
rect 1685 367761 1719 367795
rect 1719 367761 1728 367795
rect 1676 367752 1728 367761
rect 569960 367752 570012 367804
rect 570052 362312 570104 362364
rect 570236 362312 570288 362364
rect 569960 360000 570012 360052
rect 570328 360000 570380 360052
rect 569960 359864 570012 359916
rect 569960 359524 570012 359576
rect 569960 359116 570012 359168
rect 569960 358844 570012 358896
rect 569960 358708 570012 358760
rect 570236 358708 570288 358760
rect 569960 358572 570012 358624
rect 1400 358368 1452 358420
rect 1768 358368 1820 358420
rect 1860 358232 1912 358284
rect 569960 358232 570012 358284
rect 1860 358139 1912 358148
rect 1860 358105 1869 358139
rect 1869 358105 1903 358139
rect 1903 358105 1912 358139
rect 1860 358096 1912 358105
rect 1768 358028 1820 358080
rect 570052 358096 570104 358148
rect 570144 358096 570196 358148
rect 570236 358028 570288 358080
rect 570052 357892 570104 357944
rect 570144 357892 570196 357944
rect 569960 357824 570012 357876
rect 569960 353991 570012 354000
rect 569960 353957 569969 353991
rect 569969 353957 570003 353991
rect 570003 353957 570012 353991
rect 569960 353948 570012 353957
rect 569960 353744 570012 353796
rect 569960 353651 570012 353660
rect 569960 353617 569969 353651
rect 569969 353617 570003 353651
rect 570003 353617 570012 353651
rect 569960 353608 570012 353617
rect 570328 353268 570380 353320
rect 1952 353200 2004 353252
rect 569868 353200 569920 353252
rect 1768 353064 1820 353116
rect 1952 353064 2004 353116
rect 1400 352928 1452 352980
rect 1768 352928 1820 352980
rect 1952 352928 2004 352980
rect 570052 352588 570104 352640
rect 569960 352316 570012 352368
rect 569960 348959 570012 348968
rect 569960 348925 569969 348959
rect 569969 348925 570003 348959
rect 570003 348925 570012 348959
rect 569960 348916 570012 348925
rect 569960 347964 570012 348016
rect 569960 347692 570012 347744
rect 1952 345720 2004 345772
rect 1860 345652 1912 345704
rect 574928 345040 574980 345092
rect 580172 345040 580224 345092
rect 569960 344879 570012 344888
rect 569960 344845 569969 344879
rect 569969 344845 570003 344879
rect 570003 344845 570012 344879
rect 569960 344836 570012 344845
rect 569960 342227 570012 342236
rect 569960 342193 569969 342227
rect 569969 342193 570003 342227
rect 570003 342193 570012 342227
rect 569960 342184 570012 342193
rect 1952 340824 2004 340876
rect 1952 340688 2004 340740
rect 1952 340255 2004 340264
rect 1952 340221 1961 340255
rect 1961 340221 1995 340255
rect 1995 340221 2004 340255
rect 1952 340212 2004 340221
rect 1400 340144 1452 340196
rect 1768 340144 1820 340196
rect 1952 338079 2004 338088
rect 1952 338045 1961 338079
rect 1961 338045 1995 338079
rect 1995 338045 2004 338079
rect 1952 338036 2004 338045
rect 1952 334160 2004 334212
rect 1952 334024 2004 334076
rect 1308 333684 1360 333736
rect 1952 333684 2004 333736
rect 1952 333412 2004 333464
rect 1952 331780 2004 331832
rect 1400 331508 1452 331560
rect 1768 331508 1820 331560
rect 569960 331279 570012 331288
rect 569960 331245 569969 331279
rect 569969 331245 570003 331279
rect 570003 331245 570012 331279
rect 569960 331236 570012 331245
rect 569960 331075 570012 331084
rect 569960 331041 569969 331075
rect 569969 331041 570003 331075
rect 570003 331041 570012 331075
rect 569960 331032 570012 331041
rect 569960 330488 570012 330540
rect 1952 329740 2004 329792
rect 569960 329672 570012 329724
rect 569960 329536 570012 329588
rect 569960 329400 570012 329452
rect 569960 329264 570012 329316
rect 1952 329171 2004 329180
rect 1952 329137 1961 329171
rect 1961 329137 1995 329171
rect 1995 329137 2004 329171
rect 1952 329128 2004 329137
rect 569960 327768 570012 327820
rect 569960 327632 570012 327684
rect 572720 327632 572772 327684
rect 569960 327156 570012 327208
rect 569960 327020 570012 327072
rect 569960 325660 570012 325712
rect 570144 325524 570196 325576
rect 570052 325023 570104 325032
rect 570052 324989 570061 325023
rect 570061 324989 570095 325023
rect 570095 324989 570104 325023
rect 570052 324980 570104 324989
rect 569960 320968 570012 321020
rect 570144 320968 570196 321020
rect 569960 320875 570012 320884
rect 569960 320841 569969 320875
rect 569969 320841 570003 320875
rect 570003 320841 570012 320875
rect 569960 320832 570012 320841
rect 570052 320696 570104 320748
rect 1952 319175 2004 319184
rect 1952 319141 1961 319175
rect 1961 319141 1995 319175
rect 1995 319141 2004 319175
rect 1952 319132 2004 319141
rect 1952 318928 2004 318980
rect 569960 317951 570012 317960
rect 569960 317917 569969 317951
rect 569969 317917 570003 317951
rect 570003 317917 570012 317951
rect 569960 317908 570012 317917
rect 570052 315800 570104 315852
rect 570328 315800 570380 315852
rect 569960 315639 570012 315648
rect 569960 315605 569969 315639
rect 569969 315605 570003 315639
rect 570003 315605 570012 315639
rect 569960 315596 570012 315605
rect 570236 315596 570288 315648
rect 570052 315528 570104 315580
rect 570236 315503 570288 315512
rect 570236 315469 570245 315503
rect 570245 315469 570279 315503
rect 570279 315469 570288 315503
rect 570236 315460 570288 315469
rect 1952 315120 2004 315172
rect 1952 315027 2004 315036
rect 1952 314993 1961 315027
rect 1961 314993 1995 315027
rect 1995 314993 2004 315027
rect 1952 314984 2004 314993
rect 1952 312536 2004 312588
rect 1952 312400 2004 312452
rect 1952 312264 2004 312316
rect 1952 312128 2004 312180
rect 1952 311992 2004 312044
rect 1952 311788 2004 311840
rect 1952 311652 2004 311704
rect 1952 311516 2004 311568
rect 1952 309859 2004 309868
rect 1952 309825 1961 309859
rect 1961 309825 1995 309859
rect 1995 309825 2004 309859
rect 1952 309816 2004 309825
rect 1952 309612 2004 309664
rect 569960 309068 570012 309120
rect 569960 306960 570012 307012
rect 1952 306663 2004 306672
rect 1952 306629 1961 306663
rect 1961 306629 1995 306663
rect 1995 306629 2004 306663
rect 1952 306620 2004 306629
rect 569960 306187 570012 306196
rect 569960 306153 569969 306187
rect 569969 306153 570003 306187
rect 570003 306153 570012 306187
rect 569960 306144 570012 306153
rect 1952 305600 2004 305652
rect 1952 305464 2004 305516
rect 1952 305328 2004 305380
rect 1952 304512 2004 304564
rect 1952 304376 2004 304428
rect 570052 304240 570104 304292
rect 1952 304104 2004 304156
rect 1952 303968 2004 304020
rect 570236 303832 570288 303884
rect 1952 303356 2004 303408
rect 1952 303220 2004 303272
rect 569960 302744 570012 302796
rect 3332 301792 3384 301844
rect 3700 301792 3752 301844
rect 1952 301452 2004 301504
rect 569960 301112 570012 301164
rect 569960 300883 570012 300892
rect 569960 300849 569969 300883
rect 569969 300849 570003 300883
rect 570003 300849 570012 300883
rect 569960 300840 570012 300849
rect 570420 300364 570472 300416
rect 570328 300228 570380 300280
rect 570144 300092 570196 300144
rect 569960 300067 570012 300076
rect 569960 300033 569969 300067
rect 569969 300033 570003 300067
rect 570003 300033 570012 300067
rect 569960 300024 570012 300033
rect 569960 298571 570012 298580
rect 569960 298537 569969 298571
rect 569969 298537 570003 298571
rect 570003 298537 570012 298571
rect 569960 298528 570012 298537
rect 569960 298392 570012 298444
rect 575020 298120 575072 298172
rect 580172 298120 580224 298172
rect 1308 296216 1360 296268
rect 570052 296148 570104 296200
rect 1952 296080 2004 296132
rect 569960 296080 570012 296132
rect 570236 296012 570288 296064
rect 1400 295944 1452 295996
rect 1952 295808 2004 295860
rect 570328 295128 570380 295180
rect 480 294584 532 294636
rect 1952 293360 2004 293412
rect 1952 293088 2004 293140
rect 570236 292748 570288 292800
rect 570420 292544 570472 292596
rect 569960 292408 570012 292460
rect 569960 289620 570012 289672
rect 570328 288260 570380 288312
rect 20 286968 72 287020
rect 570236 285472 570288 285524
rect 569960 285336 570012 285388
rect 569960 285175 570012 285184
rect 569960 285141 569969 285175
rect 569969 285141 570003 285175
rect 570003 285141 570012 285175
rect 569960 285132 570012 285141
rect 569960 284928 570012 284980
rect 569960 284792 570012 284844
rect 1952 284724 2004 284776
rect 1952 284588 2004 284640
rect 569960 284588 570012 284640
rect 570512 284588 570564 284640
rect 1952 284316 2004 284368
rect 1400 283951 1452 283960
rect 1400 283917 1409 283951
rect 1409 283917 1443 283951
rect 1443 283917 1452 283951
rect 1400 283908 1452 283917
rect 1952 283908 2004 283960
rect 569960 283840 570012 283892
rect 569960 283747 570012 283756
rect 569960 283713 569969 283747
rect 569969 283713 570003 283747
rect 570003 283713 570012 283747
rect 569960 283704 570012 283713
rect 1952 283364 2004 283416
rect 569960 283500 570012 283552
rect 570052 283432 570104 283484
rect 569960 283364 570012 283416
rect 570052 283296 570104 283348
rect 1952 283228 2004 283280
rect 569960 277924 570012 277976
rect 570328 277924 570380 277976
rect 569960 277516 570012 277568
rect 570144 277516 570196 277568
rect 569960 277244 570012 277296
rect 569960 274456 570012 274508
rect 1952 273912 2004 273964
rect 569960 274184 570012 274236
rect 570052 273708 570104 273760
rect 569960 273071 570012 273080
rect 569960 273037 569969 273071
rect 569969 273037 570003 273071
rect 570003 273037 570012 273071
rect 569960 273028 570012 273037
rect 569960 272892 570012 272944
rect 569960 272756 570012 272808
rect 572720 272756 572772 272808
rect 569960 272552 570012 272604
rect 570420 272552 570472 272604
rect 569868 272348 569920 272400
rect 569960 271575 570012 271584
rect 569960 271541 569969 271575
rect 569969 271541 570003 271575
rect 570003 271541 570012 271575
rect 569960 271532 570012 271541
rect 569960 270988 570012 271040
rect 569960 270852 570012 270904
rect 570144 270852 570196 270904
rect 569960 270580 570012 270632
rect 570328 270580 570380 270632
rect 569960 270444 570012 270496
rect 569960 270308 570012 270360
rect 1952 270172 2004 270224
rect 569960 270172 570012 270224
rect 570236 270172 570288 270224
rect 569960 270036 570012 270088
rect 569960 269900 570012 269952
rect 1952 269764 2004 269816
rect 569960 269764 570012 269816
rect 1952 269399 2004 269408
rect 1952 269365 1961 269399
rect 1961 269365 1995 269399
rect 1995 269365 2004 269399
rect 1952 269356 2004 269365
rect 569960 267291 570012 267300
rect 569960 267257 569969 267291
rect 569969 267257 570003 267291
rect 570003 267257 570012 267291
rect 569960 267248 570012 267257
rect 1952 266568 2004 266620
rect 1952 266432 2004 266484
rect 569960 266364 570012 266416
rect 296 266296 348 266348
rect 1952 266296 2004 266348
rect 569960 265888 570012 265940
rect 1952 264707 2004 264716
rect 1952 264673 1961 264707
rect 1961 264673 1995 264707
rect 1995 264673 2004 264707
rect 1952 264664 2004 264673
rect 388 264256 440 264308
rect 1952 264256 2004 264308
rect 1952 264120 2004 264172
rect 1308 263984 1360 264036
rect 1952 263984 2004 264036
rect 569960 263984 570012 264036
rect 1400 261536 1452 261588
rect 1124 261511 1176 261520
rect 1124 261477 1133 261511
rect 1133 261477 1167 261511
rect 1167 261477 1176 261511
rect 1124 261468 1176 261477
rect 1860 261468 1912 261520
rect 1124 260720 1176 260772
rect 1768 260720 1820 260772
rect 569960 259879 570012 259888
rect 569960 259845 569969 259879
rect 569969 259845 570003 259879
rect 570003 259845 570012 259879
rect 569960 259836 570012 259845
rect 569960 259564 570012 259616
rect 1400 258204 1452 258256
rect 1768 258204 1820 258256
rect 756 257388 808 257440
rect 1400 257388 1452 257440
rect 572 257252 624 257304
rect 1952 257252 2004 257304
rect 569960 256504 570012 256556
rect 570236 256504 570288 256556
rect 570052 254736 570104 254788
rect 572 251855 624 251864
rect 572 251821 581 251855
rect 581 251821 615 251855
rect 615 251821 624 251855
rect 572 251812 624 251821
rect 848 251855 900 251864
rect 848 251821 857 251855
rect 857 251821 891 251855
rect 891 251821 900 251855
rect 848 251812 900 251821
rect 1860 251812 1912 251864
rect 569960 251744 570012 251796
rect 570144 251744 570196 251796
rect 574744 251200 574796 251252
rect 580172 251200 580224 251252
rect 569960 250928 570012 250980
rect 569960 250792 570012 250844
rect 570328 250792 570380 250844
rect 569960 250588 570012 250640
rect 569960 250452 570012 250504
rect 1952 250248 2004 250300
rect 1952 250155 2004 250164
rect 1952 250121 1961 250155
rect 1961 250121 1995 250155
rect 1995 250121 2004 250155
rect 1952 250112 2004 250121
rect 1308 248956 1360 249008
rect 1952 248956 2004 249008
rect 569960 247256 570012 247308
rect 570052 246687 570104 246696
rect 570052 246653 570061 246687
rect 570061 246653 570095 246687
rect 570095 246653 570104 246687
rect 570052 246644 570104 246653
rect 570052 246508 570104 246560
rect 569960 243652 570012 243704
rect 569960 243516 570012 243568
rect 1952 243083 2004 243092
rect 1952 243049 1961 243083
rect 1961 243049 1995 243083
rect 1995 243049 2004 243083
rect 1952 243040 2004 243049
rect 1952 242947 2004 242956
rect 1952 242913 1961 242947
rect 1961 242913 1995 242947
rect 1995 242913 2004 242947
rect 1952 242904 2004 242913
rect 1952 242539 2004 242548
rect 1952 242505 1961 242539
rect 1961 242505 1995 242539
rect 1995 242505 2004 242539
rect 1952 242496 2004 242505
rect 1860 242224 1912 242276
rect 1952 242224 2004 242276
rect 1768 242199 1820 242208
rect 1768 242165 1777 242199
rect 1777 242165 1811 242199
rect 1811 242165 1820 242199
rect 1768 242156 1820 242165
rect 1768 242020 1820 242072
rect 480 241612 532 241664
rect 1952 241612 2004 241664
rect 570144 239436 570196 239488
rect 1952 238416 2004 238468
rect 1952 238280 2004 238332
rect 1768 238144 1820 238196
rect 1952 238144 2004 238196
rect 1860 237940 1912 237992
rect 569960 236036 570012 236088
rect 480 235424 532 235476
rect 1768 235424 1820 235476
rect 569960 233656 570012 233708
rect 569960 233520 570012 233572
rect 570144 233520 570196 233572
rect 569960 230231 570012 230240
rect 569960 230197 569969 230231
rect 569969 230197 570003 230231
rect 570003 230197 570012 230231
rect 569960 230188 570012 230197
rect 569960 229984 570012 230036
rect 570144 229984 570196 230036
rect 570420 229848 570472 229900
rect 569960 229780 570012 229832
rect 570328 229780 570380 229832
rect 570144 229712 570196 229764
rect 570052 229644 570104 229696
rect 569960 229236 570012 229288
rect 1768 228395 1820 228404
rect 1768 228361 1777 228395
rect 1777 228361 1811 228395
rect 1811 228361 1820 228395
rect 1768 228352 1820 228361
rect 570052 227035 570104 227044
rect 570052 227001 570061 227035
rect 570061 227001 570095 227035
rect 570095 227001 570104 227035
rect 570052 226992 570104 227001
rect 570236 226856 570288 226908
rect 569960 225972 570012 226024
rect 570236 225972 570288 226024
rect 569960 225768 570012 225820
rect 1952 221688 2004 221740
rect 756 221620 808 221672
rect 1400 221620 1452 221672
rect 1308 221527 1360 221536
rect 1308 221493 1317 221527
rect 1317 221493 1351 221527
rect 1351 221493 1360 221527
rect 1308 221484 1360 221493
rect 1400 221484 1452 221536
rect 388 221348 440 221400
rect 1400 221280 1452 221332
rect 1952 221008 2004 221060
rect 1952 219920 2004 219972
rect 1952 218288 2004 218340
rect 1952 217676 2004 217728
rect 1400 217404 1452 217456
rect 112 216792 164 216844
rect 569960 215636 570012 215688
rect 569960 215364 570012 215416
rect 569960 214616 570012 214668
rect 570144 214591 570196 214600
rect 570144 214557 570153 214591
rect 570153 214557 570187 214591
rect 570187 214557 570196 214591
rect 570144 214548 570196 214557
rect 1400 214276 1452 214328
rect 1952 214276 2004 214328
rect 572 214140 624 214192
rect 1952 214140 2004 214192
rect 569960 214004 570012 214056
rect 570236 214004 570288 214056
rect 1952 212848 2004 212900
rect 848 209924 900 209976
rect 570144 208360 570196 208412
rect 570420 208360 570472 208412
rect 1216 207723 1268 207732
rect 1216 207689 1225 207723
rect 1225 207689 1259 207723
rect 1259 207689 1268 207723
rect 1216 207680 1268 207689
rect 572 205028 624 205080
rect 1216 205028 1268 205080
rect 1400 204892 1452 204944
rect 569960 205028 570012 205080
rect 570236 205028 570288 205080
rect 1952 204824 2004 204876
rect 1400 204756 1452 204808
rect 569960 204756 570012 204808
rect 1952 204688 2004 204740
rect 570052 204416 570104 204468
rect 574836 204280 574888 204332
rect 580172 204280 580224 204332
rect 569960 203668 570012 203720
rect 569960 203532 570012 203584
rect 569960 203396 570012 203448
rect 570236 203396 570288 203448
rect 569960 203124 570012 203176
rect 569960 202988 570012 203040
rect 569960 202623 570012 202632
rect 569960 202589 569969 202623
rect 569969 202589 570003 202623
rect 570003 202589 570012 202623
rect 569960 202580 570012 202589
rect 1952 201832 2004 201884
rect 572 200200 624 200252
rect 1400 200200 1452 200252
rect 296 199495 348 199504
rect 296 199461 305 199495
rect 305 199461 339 199495
rect 339 199461 348 199495
rect 296 199452 348 199461
rect 848 199495 900 199504
rect 848 199461 857 199495
rect 857 199461 891 199495
rect 891 199461 900 199495
rect 848 199452 900 199461
rect 1400 198228 1452 198280
rect 1952 198160 2004 198212
rect 1400 198067 1452 198076
rect 1400 198033 1409 198067
rect 1409 198033 1443 198067
rect 1443 198033 1452 198067
rect 1400 198024 1452 198033
rect 1952 197752 2004 197804
rect 940 197659 992 197668
rect 940 197625 949 197659
rect 949 197625 983 197659
rect 983 197625 992 197659
rect 940 197616 992 197625
rect 1952 197659 2004 197668
rect 1952 197625 1961 197659
rect 1961 197625 1995 197659
rect 1995 197625 2004 197659
rect 1952 197616 2004 197625
rect 940 197480 992 197532
rect 1952 196367 2004 196376
rect 1952 196333 1961 196367
rect 1961 196333 1995 196367
rect 1995 196333 2004 196367
rect 1952 196324 2004 196333
rect 1952 196188 2004 196240
rect 1952 196052 2004 196104
rect 1952 195916 2004 195968
rect 1952 195780 2004 195832
rect 1492 195644 1544 195696
rect 1308 195508 1360 195560
rect 1492 195508 1544 195560
rect 664 195100 716 195152
rect 1952 195032 2004 195084
rect 1216 194896 1268 194948
rect 1952 194896 2004 194948
rect 1952 194692 2004 194744
rect 664 193987 716 193996
rect 664 193953 673 193987
rect 673 193953 707 193987
rect 707 193953 716 193987
rect 664 193944 716 193953
rect 1952 193944 2004 193996
rect 569960 193876 570012 193928
rect 569960 192720 570012 192772
rect 569960 192491 570012 192500
rect 569960 192457 569969 192491
rect 569969 192457 570003 192491
rect 570003 192457 570012 192491
rect 569960 192448 570012 192457
rect 569960 192176 570012 192228
rect 569960 192040 570012 192092
rect 570052 191972 570104 192024
rect 569960 191904 570012 191956
rect 569960 191700 570012 191752
rect 570052 191700 570104 191752
rect 569960 191564 570012 191616
rect 570328 191564 570380 191616
rect 570144 191496 570196 191548
rect 569960 191428 570012 191480
rect 1952 189728 2004 189780
rect 1952 189592 2004 189644
rect 1952 189184 2004 189236
rect 1952 188912 2004 188964
rect 1952 188640 2004 188692
rect 569960 188572 570012 188624
rect 570236 188572 570288 188624
rect 1952 188504 2004 188556
rect 569960 188368 570012 188420
rect 1952 186464 2004 186516
rect 1216 182860 1268 182912
rect 296 182835 348 182844
rect 296 182801 305 182835
rect 305 182801 339 182835
rect 339 182801 348 182835
rect 296 182792 348 182801
rect 569960 180412 570012 180464
rect 569960 179800 570012 179852
rect 1860 179639 1912 179648
rect 1860 179605 1869 179639
rect 1869 179605 1903 179639
rect 1903 179605 1912 179639
rect 1860 179596 1912 179605
rect 1860 179052 1912 179104
rect 1768 178415 1820 178424
rect 1768 178381 1777 178415
rect 1777 178381 1811 178415
rect 1811 178381 1820 178415
rect 1768 178372 1820 178381
rect 569960 177692 570012 177744
rect 570328 177692 570380 177744
rect 1952 177667 2004 177676
rect 1952 177633 1961 177667
rect 1961 177633 1995 177667
rect 1995 177633 2004 177667
rect 1952 177624 2004 177633
rect 570144 177284 570196 177336
rect 1860 176944 1912 176996
rect 569960 176808 570012 176860
rect 1952 176740 2004 176792
rect 1952 176604 2004 176656
rect 1952 176468 2004 176520
rect 1952 176332 2004 176384
rect 1768 176239 1820 176248
rect 1768 176205 1777 176239
rect 1777 176205 1811 176239
rect 1811 176205 1820 176239
rect 1768 176196 1820 176205
rect 1952 176239 2004 176248
rect 1952 176205 1961 176239
rect 1961 176205 1995 176239
rect 1995 176205 2004 176239
rect 1952 176196 2004 176205
rect 388 176060 440 176112
rect 1952 175924 2004 175976
rect 1216 175584 1268 175636
rect 569960 175176 570012 175228
rect 569960 174947 570012 174956
rect 569960 174913 569969 174947
rect 569969 174913 570003 174947
rect 570003 174913 570012 174947
rect 569960 174904 570012 174913
rect 204 174607 256 174616
rect 204 174573 213 174607
rect 213 174573 247 174607
rect 247 174573 256 174607
rect 204 174564 256 174573
rect 204 174428 256 174480
rect 1492 174428 1544 174480
rect 569960 173612 570012 173664
rect 570144 173612 570196 173664
rect 1492 173136 1544 173188
rect 1860 173136 1912 173188
rect 1860 173000 1912 173052
rect 1216 171912 1268 171964
rect 1400 171912 1452 171964
rect 570052 171912 570104 171964
rect 112 170960 164 171012
rect 480 170323 532 170332
rect 480 170289 489 170323
rect 489 170289 523 170323
rect 523 170289 532 170323
rect 480 170280 532 170289
rect 569960 169328 570012 169380
rect 569960 169124 570012 169176
rect 1952 169099 2004 169108
rect 1952 169065 1961 169099
rect 1961 169065 1995 169099
rect 1995 169065 2004 169099
rect 1952 169056 2004 169065
rect 569960 168988 570012 169040
rect 570144 168988 570196 169040
rect 1952 167968 2004 168020
rect 1952 167764 2004 167816
rect 388 167628 440 167680
rect 1952 167628 2004 167680
rect 1952 167356 2004 167408
rect 1032 167220 1084 167272
rect 1952 167220 2004 167272
rect 1952 166880 2004 166932
rect 1032 166744 1084 166796
rect 1952 166744 2004 166796
rect 1952 166404 2004 166456
rect 480 166132 532 166184
rect 388 165860 440 165912
rect 1952 166268 2004 166320
rect 1400 165996 1452 166048
rect 1952 165996 2004 166048
rect 1952 165860 2004 165912
rect 1952 165452 2004 165504
rect 480 163888 532 163940
rect 1492 163888 1544 163940
rect 1032 163752 1084 163804
rect 1492 163752 1544 163804
rect 569960 163727 570012 163736
rect 569960 163693 569969 163727
rect 569969 163693 570003 163727
rect 570003 163693 570012 163727
rect 569960 163684 570012 163693
rect 569960 163523 570012 163532
rect 569960 163489 569969 163523
rect 569969 163489 570003 163523
rect 570003 163489 570012 163523
rect 569960 163480 570012 163489
rect 756 163276 808 163328
rect 570420 162231 570472 162240
rect 570420 162197 570429 162231
rect 570429 162197 570463 162231
rect 570463 162197 570472 162231
rect 570420 162188 570472 162197
rect 570052 161984 570104 162036
rect 756 161576 808 161628
rect 1308 161576 1360 161628
rect 1492 160080 1544 160132
rect 1492 159944 1544 159996
rect 1952 159944 2004 159996
rect 1952 159808 2004 159860
rect 1492 159672 1544 159724
rect 1952 159672 2004 159724
rect 1032 159536 1084 159588
rect 1492 159332 1544 159384
rect 1952 159264 2004 159316
rect 1952 159128 2004 159180
rect 756 159060 808 159112
rect 569960 157879 570012 157888
rect 569960 157845 569969 157879
rect 569969 157845 570003 157879
rect 570003 157845 570012 157879
rect 569960 157836 570012 157845
rect 570144 157632 570196 157684
rect 569960 157496 570012 157548
rect 570144 157496 570196 157548
rect 569960 157360 570012 157412
rect 574928 157360 574980 157412
rect 580172 157360 580224 157412
rect 1584 156340 1636 156392
rect 1400 156204 1452 156256
rect 1584 156204 1636 156256
rect 569960 155864 570012 155916
rect 570236 155728 570288 155780
rect 570052 155592 570104 155644
rect 480 155388 532 155440
rect 1308 155388 1360 155440
rect 569960 155184 570012 155236
rect 569868 155116 569920 155168
rect 570052 155048 570104 155100
rect 569960 154980 570012 155032
rect 569960 154844 570012 154896
rect 1400 154776 1452 154828
rect 1952 154028 2004 154080
rect 570052 153892 570104 153944
rect 388 153867 440 153876
rect 388 153833 397 153867
rect 397 153833 431 153867
rect 431 153833 440 153867
rect 388 153824 440 153833
rect 569960 153824 570012 153876
rect 570236 153824 570288 153876
rect 1860 153756 1912 153808
rect 570236 153459 570288 153468
rect 570236 153425 570245 153459
rect 570245 153425 570279 153459
rect 570279 153425 570288 153459
rect 570236 153416 570288 153425
rect 112 151988 164 152040
rect 388 151988 440 152040
rect 570052 149540 570104 149592
rect 570052 149404 570104 149456
rect 570328 149404 570380 149456
rect 569960 149311 570012 149320
rect 569960 149277 569969 149311
rect 569969 149277 570003 149311
rect 570003 149277 570012 149311
rect 569960 149268 570012 149277
rect 570236 149064 570288 149116
rect 570420 149064 570472 149116
rect 480 148724 532 148776
rect 1400 148588 1452 148640
rect 569960 148452 570012 148504
rect 570052 148316 570104 148368
rect 569960 147908 570012 147960
rect 569960 147772 570012 147824
rect 570144 147772 570196 147824
rect 569960 147636 570012 147688
rect 112 147092 164 147144
rect 388 147092 440 147144
rect 1584 147092 1636 147144
rect 1952 147092 2004 147144
rect 388 146999 440 147008
rect 388 146965 397 146999
rect 397 146965 431 146999
rect 431 146965 440 146999
rect 388 146956 440 146965
rect 756 146999 808 147008
rect 756 146965 765 146999
rect 765 146965 799 146999
rect 799 146965 808 146999
rect 756 146956 808 146965
rect 1952 146999 2004 147008
rect 1952 146965 1961 146999
rect 1961 146965 1995 146999
rect 1995 146965 2004 146999
rect 1952 146956 2004 146965
rect 569960 146956 570012 147008
rect 1584 146344 1636 146396
rect 572 146208 624 146260
rect 1216 145936 1268 145988
rect 1860 145911 1912 145920
rect 1860 145877 1869 145911
rect 1869 145877 1903 145911
rect 1903 145877 1912 145911
rect 1860 145868 1912 145877
rect 1952 145800 2004 145852
rect 1860 145664 1912 145716
rect 296 145639 348 145648
rect 296 145605 305 145639
rect 305 145605 339 145639
rect 339 145605 348 145639
rect 296 145596 348 145605
rect 1952 145596 2004 145648
rect 569960 144236 570012 144288
rect 570328 144236 570380 144288
rect 2780 143624 2832 143676
rect 3148 143624 3200 143676
rect 1860 143123 1912 143132
rect 1860 143089 1869 143123
rect 1869 143089 1903 143123
rect 1903 143089 1912 143123
rect 1860 143080 1912 143089
rect 1032 142944 1084 142996
rect 1584 142944 1636 142996
rect 1032 142808 1084 142860
rect 664 141856 716 141908
rect 848 141856 900 141908
rect 572 141720 624 141772
rect 848 141720 900 141772
rect 572 141627 624 141636
rect 572 141593 581 141627
rect 581 141593 615 141627
rect 615 141593 624 141627
rect 572 141584 624 141593
rect 1492 141491 1544 141500
rect 1492 141457 1501 141491
rect 1501 141457 1535 141491
rect 1535 141457 1544 141491
rect 1492 141448 1544 141457
rect 1952 141312 2004 141364
rect 1860 141244 1912 141296
rect 1952 141176 2004 141228
rect 1860 141108 1912 141160
rect 1952 139952 2004 140004
rect 1952 139068 2004 139120
rect 1952 138864 2004 138916
rect 1492 138796 1544 138848
rect 756 138728 808 138780
rect 1308 138660 1360 138712
rect 1492 138592 1544 138644
rect 1952 138592 2004 138644
rect 204 138524 256 138576
rect 664 138524 716 138576
rect 1952 138252 2004 138304
rect 1952 137912 2004 137964
rect 569960 134920 570012 134972
rect 569960 134716 570012 134768
rect 940 134648 992 134700
rect 1400 134648 1452 134700
rect 1860 134580 1912 134632
rect 1032 134512 1084 134564
rect 1676 134555 1728 134564
rect 1676 134521 1685 134555
rect 1685 134521 1719 134555
rect 1719 134521 1728 134555
rect 1676 134512 1728 134521
rect 570052 134512 570104 134564
rect 1952 134444 2004 134496
rect 940 134376 992 134428
rect 569960 134308 570012 134360
rect 570236 134308 570288 134360
rect 569960 134172 570012 134224
rect 1768 133467 1820 133476
rect 1768 133433 1777 133467
rect 1777 133433 1811 133467
rect 1811 133433 1820 133467
rect 1768 133424 1820 133433
rect 1032 133288 1084 133340
rect 569960 133084 570012 133136
rect 1952 132064 2004 132116
rect 1952 130840 2004 130892
rect 1952 130568 2004 130620
rect 1952 129412 2004 129464
rect 1952 129140 2004 129192
rect 848 128868 900 128920
rect 1860 128324 1912 128376
rect 1768 126624 1820 126676
rect 1860 126352 1912 126404
rect 388 126284 440 126336
rect 848 126284 900 126336
rect 1584 126216 1636 126268
rect 388 126080 440 126132
rect 1952 126080 2004 126132
rect 1676 126012 1728 126064
rect 1860 124967 1912 124976
rect 1860 124933 1869 124967
rect 1869 124933 1903 124967
rect 1903 124933 1912 124967
rect 1860 124924 1912 124933
rect 1952 124967 2004 124976
rect 1952 124933 1961 124967
rect 1961 124933 1995 124967
rect 1995 124933 2004 124967
rect 1952 124924 2004 124933
rect 1676 124899 1728 124908
rect 1676 124865 1685 124899
rect 1685 124865 1719 124899
rect 1719 124865 1728 124899
rect 1676 124856 1728 124865
rect 1400 124720 1452 124772
rect 1768 124763 1820 124772
rect 1768 124729 1777 124763
rect 1777 124729 1811 124763
rect 1811 124729 1820 124763
rect 1768 124720 1820 124729
rect 756 124584 808 124636
rect 1400 124584 1452 124636
rect 572720 124040 572772 124092
rect 574836 124040 574888 124092
rect 756 121184 808 121236
rect 940 121184 992 121236
rect 940 121048 992 121100
rect 1216 121048 1268 121100
rect 1952 118031 2004 118040
rect 1952 117997 1961 118031
rect 1961 117997 1995 118031
rect 1995 117997 2004 118031
rect 1952 117988 2004 117997
rect 1952 117784 2004 117836
rect 1216 117512 1268 117564
rect 1952 117512 2004 117564
rect 1952 117376 2004 117428
rect 1308 116424 1360 116476
rect 1216 115064 1268 115116
rect 1952 110984 2004 111036
rect 574744 110440 574796 110492
rect 580172 110440 580224 110492
rect 1216 110032 1268 110084
rect 1952 110032 2004 110084
rect 1952 109692 2004 109744
rect 1952 109420 2004 109472
rect 1952 109284 2004 109336
rect 1952 109148 2004 109200
rect 1952 108876 2004 108928
rect 1952 108740 2004 108792
rect 1952 108604 2004 108656
rect 1952 108468 2004 108520
rect 1952 108332 2004 108384
rect 1216 108060 1268 108112
rect 1952 108060 2004 108112
rect 1952 107652 2004 107704
rect 1308 107312 1360 107364
rect 1952 107312 2004 107364
rect 1952 107176 2004 107228
rect 1952 107083 2004 107092
rect 1952 107049 1961 107083
rect 1961 107049 1995 107083
rect 1995 107049 2004 107083
rect 1952 107040 2004 107049
rect 1216 102552 1268 102604
rect 1952 98404 2004 98456
rect 1308 98311 1360 98320
rect 1308 98277 1317 98311
rect 1317 98277 1351 98311
rect 1351 98277 1360 98311
rect 1308 98268 1360 98277
rect 1952 98268 2004 98320
rect 388 98132 440 98184
rect 1308 98132 1360 98184
rect 1952 98175 2004 98184
rect 1952 98141 1961 98175
rect 1961 98141 1995 98175
rect 1995 98141 2004 98175
rect 1952 98132 2004 98141
rect 572720 96500 572772 96552
rect 574928 96500 574980 96552
rect 480 96228 532 96280
rect 1860 94775 1912 94784
rect 1860 94741 1869 94775
rect 1869 94741 1903 94775
rect 1903 94741 1912 94775
rect 1860 94732 1912 94741
rect 1952 94664 2004 94716
rect 1952 93984 2004 94036
rect 1952 93576 2004 93628
rect 1860 93440 1912 93492
rect 1952 93372 2004 93424
rect 1860 93279 1912 93288
rect 1860 93245 1869 93279
rect 1869 93245 1903 93279
rect 1903 93245 1912 93279
rect 1860 93236 1912 93245
rect 1952 93236 2004 93288
rect 572 93100 624 93152
rect 1952 92148 2004 92200
rect 1952 92012 2004 92064
rect 1952 91876 2004 91928
rect 1952 91740 2004 91792
rect 1952 91604 2004 91656
rect 1952 91468 2004 91520
rect 1952 91332 2004 91384
rect 1952 91196 2004 91248
rect 1952 86411 2004 86420
rect 1952 86377 1961 86411
rect 1961 86377 1995 86411
rect 1995 86377 2004 86411
rect 1952 86368 2004 86377
rect 1860 86300 1912 86352
rect 1952 86164 2004 86216
rect 1860 86096 1912 86148
rect 1952 84736 2004 84788
rect 1952 84600 2004 84652
rect 1952 83784 2004 83836
rect 1952 83580 2004 83632
rect 1308 83444 1360 83496
rect 1860 83444 1912 83496
rect 1952 82084 2004 82136
rect 572 80928 624 80980
rect 1952 80724 2004 80776
rect 569960 77256 570012 77308
rect 569960 76712 570012 76764
rect 569960 76576 570012 76628
rect 569960 76440 570012 76492
rect 570144 76440 570196 76492
rect 569960 76347 570012 76356
rect 569960 76313 569969 76347
rect 569969 76313 570003 76347
rect 570003 76313 570012 76347
rect 569960 76304 570012 76313
rect 569960 76168 570012 76220
rect 569960 74808 570012 74860
rect 569960 74672 570012 74724
rect 570236 74672 570288 74724
rect 569960 73720 570012 73772
rect 569960 73584 570012 73636
rect 569960 73380 570012 73432
rect 569960 73244 570012 73296
rect 570236 73244 570288 73296
rect 569960 73108 570012 73160
rect 569960 72972 570012 73024
rect 572 72564 624 72616
rect 1860 72564 1912 72616
rect 1860 72471 1912 72480
rect 1860 72437 1869 72471
rect 1869 72437 1903 72471
rect 1903 72437 1912 72471
rect 1860 72428 1912 72437
rect 569960 72428 570012 72480
rect 1308 72156 1360 72208
rect 1952 72156 2004 72208
rect 1952 71952 2004 72004
rect 1216 71000 1268 71052
rect 1952 71000 2004 71052
rect 1308 69300 1360 69352
rect 569960 68348 570012 68400
rect 570236 68348 570288 68400
rect 569960 68008 570012 68060
rect 569960 67872 570012 67924
rect 570144 67872 570196 67924
rect 1952 67464 2004 67516
rect 1308 67328 1360 67380
rect 1952 67328 2004 67380
rect 1952 67192 2004 67244
rect 204 66920 256 66972
rect 1952 66716 2004 66768
rect 1952 66580 2004 66632
rect 1952 66487 2004 66496
rect 1952 66453 1961 66487
rect 1961 66453 1995 66487
rect 1995 66453 2004 66487
rect 1952 66444 2004 66453
rect 570144 66104 570196 66156
rect 570052 65968 570104 66020
rect 1676 65875 1728 65884
rect 1676 65841 1685 65875
rect 1685 65841 1719 65875
rect 1719 65841 1728 65875
rect 1676 65832 1728 65841
rect 1216 65424 1268 65476
rect 2044 65424 2096 65476
rect 1308 65220 1360 65272
rect 569960 64948 570012 65000
rect 1676 64787 1728 64796
rect 1676 64753 1685 64787
rect 1685 64753 1719 64787
rect 1719 64753 1728 64787
rect 1676 64744 1728 64753
rect 1952 64744 2004 64796
rect 1952 64608 2004 64660
rect 574744 63520 574796 63572
rect 580172 63520 580224 63572
rect 1216 63316 1268 63368
rect 1952 63316 2004 63368
rect 1952 63112 2004 63164
rect 1952 62976 2004 63028
rect 1952 62840 2004 62892
rect 1952 62228 2004 62280
rect 569960 61684 570012 61736
rect 569960 61548 570012 61600
rect 570144 61548 570196 61600
rect 570052 61276 570104 61328
rect 569960 60732 570012 60784
rect 569960 59916 570012 59968
rect 569960 58828 570012 58880
rect 569960 58692 570012 58744
rect 1308 57876 1360 57928
rect 1952 57060 2004 57112
rect 569960 56967 570012 56976
rect 569960 56933 569969 56967
rect 569969 56933 570003 56967
rect 570003 56933 570012 56967
rect 569960 56924 570012 56933
rect 1952 56856 2004 56908
rect 1952 56720 2004 56772
rect 569960 56652 570012 56704
rect 1952 56584 2004 56636
rect 569960 56516 570012 56568
rect 1952 55836 2004 55888
rect 1952 55156 2004 55208
rect 569960 53728 570012 53780
rect 1952 52708 2004 52760
rect 1952 52572 2004 52624
rect 1032 50371 1084 50380
rect 1032 50337 1041 50371
rect 1041 50337 1075 50371
rect 1075 50337 1084 50371
rect 1032 50328 1084 50337
rect 112 47472 164 47524
rect 569960 45500 570012 45552
rect 570328 45500 570380 45552
rect 569960 43256 570012 43308
rect 1952 43052 2004 43104
rect 1952 42780 2004 42832
rect 569960 42347 570012 42356
rect 569960 42313 569969 42347
rect 569969 42313 570003 42347
rect 570003 42313 570012 42347
rect 569960 42304 570012 42313
rect 569960 42168 570012 42220
rect 569960 41760 570012 41812
rect 569960 41624 570012 41676
rect 569960 41080 570012 41132
rect 569960 40987 570012 40996
rect 569960 40953 569969 40987
rect 569969 40953 570003 40987
rect 570003 40953 570012 40987
rect 569960 40944 570012 40953
rect 569960 40672 570012 40724
rect 569960 40400 570012 40452
rect 569960 40264 570012 40316
rect 569960 40128 570012 40180
rect 569960 39992 570012 40044
rect 569960 39856 570012 39908
rect 569960 39695 570012 39704
rect 569960 39661 569969 39695
rect 569969 39661 570003 39695
rect 570003 39661 570012 39695
rect 569960 39652 570012 39661
rect 1952 39448 2004 39500
rect 569960 39380 570012 39432
rect 1492 39312 1544 39364
rect 1952 39312 2004 39364
rect 1952 39176 2004 39228
rect 570236 39040 570288 39092
rect 1308 38496 1360 38548
rect 1860 38496 1912 38548
rect 1032 37043 1084 37052
rect 1032 37009 1041 37043
rect 1041 37009 1075 37043
rect 1075 37009 1084 37043
rect 1032 37000 1084 37009
rect 1952 35640 2004 35692
rect 1952 35504 2004 35556
rect 1952 35368 2004 35420
rect 388 35232 440 35284
rect 1952 35232 2004 35284
rect 20 35003 72 35012
rect 20 34969 29 35003
rect 29 34969 63 35003
rect 63 34969 72 35003
rect 20 34960 72 34969
rect 570328 34756 570380 34808
rect 664 33575 716 33584
rect 664 33541 673 33575
rect 673 33541 707 33575
rect 707 33541 716 33575
rect 664 33532 716 33541
rect 570144 31016 570196 31068
rect 112 29860 164 29912
rect 1860 29724 1912 29776
rect 1768 29656 1820 29708
rect 1768 29520 1820 29572
rect 1492 29495 1544 29504
rect 1492 29461 1501 29495
rect 1501 29461 1535 29495
rect 1535 29461 1544 29495
rect 1492 29452 1544 29461
rect 1952 28296 2004 28348
rect 1492 27956 1544 28008
rect 1952 27956 2004 28008
rect 1952 27208 2004 27260
rect 1216 27072 1268 27124
rect 1952 27072 2004 27124
rect 1216 26936 1268 26988
rect 1952 26936 2004 26988
rect 1492 26800 1544 26852
rect 1952 26800 2004 26852
rect 569960 26460 570012 26512
rect 569960 25712 570012 25764
rect 569960 25508 570012 25560
rect 569960 25100 570012 25152
rect 570236 25100 570288 25152
rect 569960 24284 570012 24336
rect 570328 24284 570380 24336
rect 112 24259 164 24268
rect 112 24225 121 24259
rect 121 24225 155 24259
rect 155 24225 164 24259
rect 112 24216 164 24225
rect 569960 24148 570012 24200
rect 1492 24012 1544 24064
rect 1492 23740 1544 23792
rect 569960 23740 570012 23792
rect 569960 23536 570012 23588
rect 570236 23536 570288 23588
rect 569960 23196 570012 23248
rect 1952 22176 2004 22228
rect 1952 22040 2004 22092
rect 1308 21564 1360 21616
rect 112 20136 164 20188
rect 1400 20136 1452 20188
rect 1032 20000 1084 20052
rect 1400 19932 1452 19984
rect 756 19796 808 19848
rect 1308 18844 1360 18896
rect 1400 18708 1452 18760
rect 1400 18572 1452 18624
rect 1952 18436 2004 18488
rect 1032 18368 1084 18420
rect 480 18232 532 18284
rect 1860 17892 1912 17944
rect 569960 17620 570012 17672
rect 1124 16668 1176 16720
rect 1860 16532 1912 16584
rect 1860 16396 1912 16448
rect 1952 16260 2004 16312
rect 1860 16056 1912 16108
rect 1400 15920 1452 15972
rect 1492 15716 1544 15768
rect 1952 15716 2004 15768
rect 1124 15580 1176 15632
rect 1952 15580 2004 15632
rect 1952 15444 2004 15496
rect 1952 15308 2004 15360
rect 1492 15104 1544 15156
rect 1492 14968 1544 15020
rect 1768 14968 1820 15020
rect 1952 15104 2004 15156
rect 571616 15104 571668 15156
rect 580172 15104 580224 15156
rect 1124 14807 1176 14816
rect 1124 14773 1133 14807
rect 1133 14773 1167 14807
rect 1167 14773 1176 14807
rect 1124 14764 1176 14773
rect 1860 14764 1912 14816
rect 570328 14696 570380 14748
rect 1124 14628 1176 14680
rect 1952 13472 2004 13524
rect 1952 13336 2004 13388
rect 1124 12996 1176 13048
rect 1952 12996 2004 13048
rect 1124 12792 1176 12844
rect 1952 12792 2004 12844
rect 1492 12452 1544 12504
rect 1952 12452 2004 12504
rect 1124 12316 1176 12368
rect 1308 12180 1360 12232
rect 1308 12044 1360 12096
rect 848 11840 900 11892
rect 848 10480 900 10532
rect 572 10387 624 10396
rect 572 10353 581 10387
rect 581 10353 615 10387
rect 615 10353 624 10387
rect 572 10344 624 10353
rect 664 10344 716 10396
rect 1032 10387 1084 10396
rect 1032 10353 1041 10387
rect 1041 10353 1075 10387
rect 1075 10353 1084 10387
rect 1032 10344 1084 10353
rect 480 10140 532 10192
rect 940 10208 992 10260
rect 1032 10072 1084 10124
rect 1308 9392 1360 9444
rect 1584 8712 1636 8764
rect 480 8687 532 8696
rect 480 8653 489 8687
rect 489 8653 523 8687
rect 523 8653 532 8687
rect 480 8644 532 8653
rect 569960 8576 570012 8628
rect 570328 8576 570380 8628
rect 569960 8143 570012 8152
rect 569960 8109 569969 8143
rect 569969 8109 570003 8143
rect 570003 8109 570012 8143
rect 569960 8100 570012 8109
rect 569960 7828 570012 7880
rect 848 7488 900 7540
rect 756 4700 808 4752
rect 1952 4700 2004 4752
rect 756 3723 808 3732
rect 756 3689 765 3723
rect 765 3689 799 3723
rect 799 3689 808 3723
rect 756 3680 808 3689
rect 1860 3723 1912 3732
rect 1860 3689 1869 3723
rect 1869 3689 1903 3723
rect 1903 3689 1912 3723
rect 1860 3680 1912 3689
rect 1216 3315 1268 3324
rect 1216 3281 1225 3315
rect 1225 3281 1259 3315
rect 1259 3281 1268 3315
rect 1216 3272 1268 3281
rect 124312 3111 124364 3120
rect 124312 3077 124321 3111
rect 124321 3077 124355 3111
rect 124355 3077 124364 3111
rect 177948 3111 178000 3120
rect 124312 3068 124364 3077
rect 177948 3077 177957 3111
rect 177957 3077 177991 3111
rect 177991 3077 178000 3111
rect 177948 3068 178000 3077
rect 268384 3111 268436 3120
rect 268384 3077 268393 3111
rect 268393 3077 268427 3111
rect 268427 3077 268436 3111
rect 268384 3068 268436 3077
rect 1492 1776 1544 1828
rect 1676 1708 1728 1760
rect 1492 1640 1544 1692
rect 20 1572 72 1624
rect 3792 1708 3844 1760
rect 7656 1708 7708 1760
rect 2964 1640 3016 1692
rect 4068 1640 4120 1692
rect 5448 1683 5500 1692
rect 5448 1649 5457 1683
rect 5457 1649 5491 1683
rect 5491 1649 5500 1683
rect 5448 1640 5500 1649
rect 22100 1708 22152 1760
rect 22192 1708 22244 1760
rect 26424 1708 26476 1760
rect 18328 1640 18380 1692
rect 19340 1640 19392 1692
rect 26608 1640 26660 1692
rect 37740 1640 37792 1692
rect 39028 1640 39080 1692
rect 42708 1640 42760 1692
rect 10416 1572 10468 1624
rect 42524 1572 42576 1624
rect 45560 1640 45612 1692
rect 48688 1751 48740 1760
rect 48688 1717 48697 1751
rect 48697 1717 48731 1751
rect 48731 1717 48740 1751
rect 48688 1708 48740 1717
rect 48872 1708 48924 1760
rect 50620 1708 50672 1760
rect 50804 1751 50856 1760
rect 50804 1717 50813 1751
rect 50813 1717 50847 1751
rect 50847 1717 50856 1751
rect 50804 1708 50856 1717
rect 56416 1708 56468 1760
rect 56692 1708 56744 1760
rect 111984 1708 112036 1760
rect 56784 1683 56836 1692
rect 56784 1649 56793 1683
rect 56793 1649 56827 1683
rect 56827 1649 56836 1683
rect 56784 1640 56836 1649
rect 57888 1640 57940 1692
rect 71780 1640 71832 1692
rect 128268 1751 128320 1760
rect 128268 1717 128277 1751
rect 128277 1717 128311 1751
rect 128311 1717 128320 1751
rect 128268 1708 128320 1717
rect 124588 1640 124640 1692
rect 111340 1572 111392 1624
rect 112168 1572 112220 1624
rect 115204 1572 115256 1624
rect 125784 1572 125836 1624
rect 134524 1640 134576 1692
rect 135168 1640 135220 1692
rect 137192 1640 137244 1692
rect 138296 1640 138348 1692
rect 138388 1640 138440 1692
rect 138756 1640 138808 1692
rect 138940 1708 138992 1760
rect 145564 1708 145616 1760
rect 145840 1708 145892 1760
rect 146208 1708 146260 1760
rect 147036 1708 147088 1760
rect 148324 1708 148376 1760
rect 148600 1708 148652 1760
rect 149244 1708 149296 1760
rect 149336 1708 149388 1760
rect 149980 1708 150032 1760
rect 128820 1572 128872 1624
rect 150164 1640 150216 1692
rect 156788 1708 156840 1760
rect 144736 1572 144788 1624
rect 148968 1572 149020 1624
rect 150624 1640 150676 1692
rect 161572 1708 161624 1760
rect 169484 1708 169536 1760
rect 170956 1708 171008 1760
rect 171048 1708 171100 1760
rect 174268 1708 174320 1760
rect 175280 1708 175332 1760
rect 177856 1708 177908 1760
rect 1584 1436 1636 1488
rect 3516 1436 3568 1488
rect 6828 1436 6880 1488
rect 17960 1504 18012 1556
rect 18052 1504 18104 1556
rect 28356 1504 28408 1556
rect 36176 1504 36228 1556
rect 39580 1504 39632 1556
rect 41144 1504 41196 1556
rect 45468 1504 45520 1556
rect 56600 1504 56652 1556
rect 58072 1504 58124 1556
rect 59268 1504 59320 1556
rect 59360 1504 59412 1556
rect 66904 1504 66956 1556
rect 940 1368 992 1420
rect 5264 1368 5316 1420
rect 5908 1368 5960 1420
rect 6460 1368 6512 1420
rect 10692 1368 10744 1420
rect 4988 1300 5040 1352
rect 5356 1300 5408 1352
rect 3148 1232 3200 1284
rect 8852 1232 8904 1284
rect 10600 1300 10652 1352
rect 29092 1368 29144 1420
rect 14464 1300 14516 1352
rect 14556 1300 14608 1352
rect 18052 1300 18104 1352
rect 48964 1436 49016 1488
rect 57980 1436 58032 1488
rect 60740 1436 60792 1488
rect 78588 1436 78640 1488
rect 101680 1504 101732 1556
rect 102232 1504 102284 1556
rect 103336 1504 103388 1556
rect 103704 1504 103756 1556
rect 47032 1300 47084 1352
rect 62304 1368 62356 1420
rect 68836 1368 68888 1420
rect 68928 1368 68980 1420
rect 71872 1368 71924 1420
rect 74448 1368 74500 1420
rect 74540 1368 74592 1420
rect 27896 1232 27948 1284
rect 24308 1164 24360 1216
rect 4988 1096 5040 1148
rect 5080 1028 5132 1080
rect 33876 1096 33928 1148
rect 55036 1300 55088 1352
rect 58256 1300 58308 1352
rect 59176 1300 59228 1352
rect 78864 1368 78916 1420
rect 81348 1368 81400 1420
rect 81808 1368 81860 1420
rect 76656 1300 76708 1352
rect 47952 1232 48004 1284
rect 48688 1232 48740 1284
rect 39396 1164 39448 1216
rect 56692 1164 56744 1216
rect 57980 1164 58032 1216
rect 63684 1232 63736 1284
rect 78772 1232 78824 1284
rect 82360 1232 82412 1284
rect 85672 1368 85724 1420
rect 85856 1368 85908 1420
rect 86316 1300 86368 1352
rect 86868 1300 86920 1352
rect 63592 1164 63644 1216
rect 66904 1164 66956 1216
rect 78864 1096 78916 1148
rect 84936 1164 84988 1216
rect 91928 1232 91980 1284
rect 92572 1232 92624 1284
rect 92664 1232 92716 1284
rect 106924 1436 106976 1488
rect 111248 1436 111300 1488
rect 109868 1368 109920 1420
rect 111432 1368 111484 1420
rect 115204 1368 115256 1420
rect 119436 1368 119488 1420
rect 119804 1368 119856 1420
rect 120356 1368 120408 1420
rect 121000 1368 121052 1420
rect 122012 1368 122064 1420
rect 122748 1436 122800 1488
rect 125968 1436 126020 1488
rect 127992 1436 128044 1488
rect 128452 1436 128504 1488
rect 142528 1504 142580 1556
rect 142896 1504 142948 1556
rect 152004 1504 152056 1556
rect 157064 1572 157116 1624
rect 157156 1547 157208 1556
rect 157156 1513 157165 1547
rect 157165 1513 157199 1547
rect 157199 1513 157208 1547
rect 157156 1504 157208 1513
rect 157340 1547 157392 1556
rect 157340 1513 157349 1547
rect 157349 1513 157383 1547
rect 157383 1513 157392 1547
rect 157340 1504 157392 1513
rect 158904 1640 158956 1692
rect 158812 1572 158864 1624
rect 159364 1572 159416 1624
rect 169116 1640 169168 1692
rect 169576 1640 169628 1692
rect 157984 1504 158036 1556
rect 160284 1504 160336 1556
rect 160928 1504 160980 1556
rect 183744 1708 183796 1760
rect 190368 1708 190420 1760
rect 191012 1708 191064 1760
rect 191196 1751 191248 1760
rect 191196 1717 191205 1751
rect 191205 1717 191239 1751
rect 191239 1717 191248 1751
rect 191196 1708 191248 1717
rect 191748 1708 191800 1760
rect 179052 1640 179104 1692
rect 179144 1640 179196 1692
rect 179328 1640 179380 1692
rect 179512 1640 179564 1692
rect 178684 1572 178736 1624
rect 178776 1615 178828 1624
rect 178776 1581 178785 1615
rect 178785 1581 178819 1615
rect 178819 1581 178828 1615
rect 178776 1572 178828 1581
rect 183928 1572 183980 1624
rect 169852 1504 169904 1556
rect 102232 1343 102284 1352
rect 102232 1309 102241 1343
rect 102241 1309 102275 1343
rect 102275 1309 102284 1343
rect 102232 1300 102284 1309
rect 100300 1232 100352 1284
rect 101956 1232 102008 1284
rect 102784 1232 102836 1284
rect 103336 1232 103388 1284
rect 106648 1232 106700 1284
rect 106832 1232 106884 1284
rect 110420 1232 110472 1284
rect 110604 1232 110656 1284
rect 111156 1232 111208 1284
rect 111892 1232 111944 1284
rect 116492 1232 116544 1284
rect 116676 1275 116728 1284
rect 116676 1241 116685 1275
rect 116685 1241 116719 1275
rect 116719 1241 116728 1275
rect 116676 1232 116728 1241
rect 116768 1232 116820 1284
rect 121368 1232 121420 1284
rect 126152 1232 126204 1284
rect 128636 1300 128688 1352
rect 128912 1343 128964 1352
rect 128544 1232 128596 1284
rect 128912 1309 128921 1343
rect 128921 1309 128955 1343
rect 128955 1309 128964 1343
rect 128912 1300 128964 1309
rect 129280 1300 129332 1352
rect 145564 1479 145616 1488
rect 145564 1445 145573 1479
rect 145573 1445 145607 1479
rect 145607 1445 145616 1479
rect 145564 1436 145616 1445
rect 134800 1368 134852 1420
rect 135812 1368 135864 1420
rect 138756 1368 138808 1420
rect 139124 1368 139176 1420
rect 139216 1368 139268 1420
rect 140320 1368 140372 1420
rect 140412 1368 140464 1420
rect 141148 1368 141200 1420
rect 144184 1368 144236 1420
rect 145104 1368 145156 1420
rect 145196 1368 145248 1420
rect 149244 1436 149296 1488
rect 149428 1436 149480 1488
rect 152556 1436 152608 1488
rect 148876 1368 148928 1420
rect 162860 1368 162912 1420
rect 169392 1436 169444 1488
rect 171508 1436 171560 1488
rect 184204 1572 184256 1624
rect 166816 1368 166868 1420
rect 167276 1368 167328 1420
rect 167368 1368 167420 1420
rect 169208 1368 169260 1420
rect 173624 1368 173676 1420
rect 177856 1436 177908 1488
rect 189908 1504 189960 1556
rect 190000 1504 190052 1556
rect 190092 1504 190144 1556
rect 190552 1504 190604 1556
rect 214196 1572 214248 1624
rect 214472 1572 214524 1624
rect 214932 1572 214984 1624
rect 216588 1572 216640 1624
rect 216772 1640 216824 1692
rect 220176 1640 220228 1692
rect 197820 1504 197872 1556
rect 198556 1504 198608 1556
rect 199108 1504 199160 1556
rect 182640 1436 182692 1488
rect 190368 1479 190420 1488
rect 190368 1445 190377 1479
rect 190377 1445 190411 1479
rect 190411 1445 190420 1479
rect 190368 1436 190420 1445
rect 191012 1436 191064 1488
rect 191288 1436 191340 1488
rect 191656 1479 191708 1488
rect 191656 1445 191665 1479
rect 191665 1445 191699 1479
rect 191699 1445 191708 1479
rect 191656 1436 191708 1445
rect 191840 1436 191892 1488
rect 192116 1436 192168 1488
rect 196532 1436 196584 1488
rect 196992 1436 197044 1488
rect 200212 1436 200264 1488
rect 204628 1504 204680 1556
rect 204536 1436 204588 1488
rect 233516 1708 233568 1760
rect 236552 1708 236604 1760
rect 240140 1708 240192 1760
rect 241520 1708 241572 1760
rect 250168 1708 250220 1760
rect 253664 1708 253716 1760
rect 257068 1708 257120 1760
rect 258448 1640 258500 1692
rect 260748 1640 260800 1692
rect 261300 1640 261352 1692
rect 261760 1640 261812 1692
rect 262312 1751 262364 1760
rect 262312 1717 262321 1751
rect 262321 1717 262355 1751
rect 262355 1717 262364 1751
rect 262312 1708 262364 1717
rect 280068 1708 280120 1760
rect 280252 1708 280304 1760
rect 290280 1708 290332 1760
rect 337844 1708 337896 1760
rect 352932 1708 352984 1760
rect 366364 1708 366416 1760
rect 569040 1776 569092 1828
rect 569224 1776 569276 1828
rect 375932 1708 375984 1760
rect 404452 1708 404504 1760
rect 474924 1708 474976 1760
rect 481272 1708 481324 1760
rect 489000 1708 489052 1760
rect 501788 1708 501840 1760
rect 512368 1708 512420 1760
rect 529388 1708 529440 1760
rect 559104 1708 559156 1760
rect 567292 1708 567344 1760
rect 568304 1751 568356 1760
rect 568304 1717 568313 1751
rect 568313 1717 568347 1751
rect 568347 1717 568356 1751
rect 568304 1708 568356 1717
rect 296812 1640 296864 1692
rect 299940 1640 299992 1692
rect 314752 1640 314804 1692
rect 319720 1640 319772 1692
rect 348700 1640 348752 1692
rect 358176 1640 358228 1692
rect 413836 1640 413888 1692
rect 415676 1640 415728 1692
rect 418804 1640 418856 1692
rect 432328 1640 432380 1692
rect 443644 1640 443696 1692
rect 453304 1640 453356 1692
rect 462872 1640 462924 1692
rect 509056 1640 509108 1692
rect 558000 1640 558052 1692
rect 569776 1640 569828 1692
rect 232044 1572 232096 1624
rect 232504 1572 232556 1624
rect 234068 1572 234120 1624
rect 237932 1572 237984 1624
rect 238116 1572 238168 1624
rect 238668 1572 238720 1624
rect 238760 1572 238812 1624
rect 262312 1572 262364 1624
rect 272156 1572 272208 1624
rect 273904 1572 273956 1624
rect 273996 1572 274048 1624
rect 280252 1572 280304 1624
rect 280528 1572 280580 1624
rect 290372 1572 290424 1624
rect 290924 1572 290976 1624
rect 293684 1572 293736 1624
rect 204812 1436 204864 1488
rect 211344 1436 211396 1488
rect 177488 1368 177540 1420
rect 179788 1368 179840 1420
rect 179880 1411 179932 1420
rect 179880 1377 179889 1411
rect 179889 1377 179923 1411
rect 179923 1377 179932 1411
rect 179880 1368 179932 1377
rect 217692 1368 217744 1420
rect 218060 1368 218112 1420
rect 218428 1368 218480 1420
rect 150256 1300 150308 1352
rect 134616 1232 134668 1284
rect 134800 1232 134852 1284
rect 140780 1232 140832 1284
rect 142804 1232 142856 1284
rect 151912 1300 151964 1352
rect 152096 1232 152148 1284
rect 152648 1232 152700 1284
rect 87880 1207 87932 1216
rect 87880 1173 87889 1207
rect 87889 1173 87923 1207
rect 87923 1173 87932 1207
rect 87880 1164 87932 1173
rect 88156 1164 88208 1216
rect 88524 1164 88576 1216
rect 88616 1164 88668 1216
rect 92204 1164 92256 1216
rect 93124 1164 93176 1216
rect 104624 1164 104676 1216
rect 106556 1164 106608 1216
rect 110512 1164 110564 1216
rect 111984 1207 112036 1216
rect 111984 1173 111993 1207
rect 111993 1173 112027 1207
rect 112027 1173 112036 1207
rect 111984 1164 112036 1173
rect 119344 1164 119396 1216
rect 139492 1164 139544 1216
rect 144828 1164 144880 1216
rect 144920 1164 144972 1216
rect 83188 1096 83240 1148
rect 83372 1096 83424 1148
rect 83556 1096 83608 1148
rect 5540 1028 5592 1080
rect 62304 1028 62356 1080
rect 62396 1028 62448 1080
rect 66628 1028 66680 1080
rect 66720 1028 66772 1080
rect 68836 1028 68888 1080
rect 3240 960 3292 1012
rect 83004 1028 83056 1080
rect 92020 1028 92072 1080
rect 103980 1096 104032 1148
rect 104808 1096 104860 1148
rect 105820 1096 105872 1148
rect 115940 1096 115992 1148
rect 122840 1096 122892 1148
rect 123208 1096 123260 1148
rect 134800 1096 134852 1148
rect 140228 1096 140280 1148
rect 142344 1096 142396 1148
rect 147588 1096 147640 1148
rect 92756 1028 92808 1080
rect 92848 1028 92900 1080
rect 121184 1028 121236 1080
rect 116216 960 116268 1012
rect 120080 960 120132 1012
rect 122472 960 122524 1012
rect 123944 960 123996 1012
rect 147496 1028 147548 1080
rect 149796 1164 149848 1216
rect 152464 1164 152516 1216
rect 149980 1096 150032 1148
rect 156420 1232 156472 1284
rect 157432 1232 157484 1284
rect 158168 1232 158220 1284
rect 158628 1232 158680 1284
rect 158812 1232 158864 1284
rect 159456 1232 159508 1284
rect 162308 1232 162360 1284
rect 163688 1232 163740 1284
rect 169944 1232 169996 1284
rect 176016 1232 176068 1284
rect 177672 1275 177724 1284
rect 177672 1241 177681 1275
rect 177681 1241 177715 1275
rect 177715 1241 177724 1275
rect 177672 1232 177724 1241
rect 178040 1232 178092 1284
rect 178132 1232 178184 1284
rect 190184 1300 190236 1352
rect 190828 1300 190880 1352
rect 191472 1300 191524 1352
rect 195244 1300 195296 1352
rect 197268 1300 197320 1352
rect 198464 1300 198516 1352
rect 199200 1343 199252 1352
rect 199200 1309 199209 1343
rect 199209 1309 199243 1343
rect 199243 1309 199252 1343
rect 199200 1300 199252 1309
rect 202972 1300 203024 1352
rect 211160 1300 211212 1352
rect 214380 1300 214432 1352
rect 214748 1300 214800 1352
rect 218796 1368 218848 1420
rect 232596 1436 232648 1488
rect 233148 1436 233200 1488
rect 238944 1436 238996 1488
rect 241336 1436 241388 1488
rect 249892 1436 249944 1488
rect 250720 1436 250772 1488
rect 285772 1504 285824 1556
rect 289728 1504 289780 1556
rect 298560 1504 298612 1556
rect 394884 1572 394936 1624
rect 395436 1572 395488 1624
rect 398656 1572 398708 1624
rect 399576 1572 399628 1624
rect 403716 1572 403768 1624
rect 432972 1572 433024 1624
rect 443460 1572 443512 1624
rect 453212 1572 453264 1624
rect 515588 1572 515640 1624
rect 528836 1572 528888 1624
rect 549260 1572 549312 1624
rect 568304 1572 568356 1624
rect 568672 1572 568724 1624
rect 305552 1504 305604 1556
rect 305644 1504 305696 1556
rect 318892 1504 318944 1556
rect 423404 1504 423456 1556
rect 425060 1504 425112 1556
rect 568488 1504 568540 1556
rect 568764 1504 568816 1556
rect 259092 1368 259144 1420
rect 259184 1368 259236 1420
rect 263048 1436 263100 1488
rect 265164 1436 265216 1488
rect 265440 1479 265492 1488
rect 265440 1445 265449 1479
rect 265449 1445 265483 1479
rect 265483 1445 265492 1479
rect 265440 1436 265492 1445
rect 265624 1436 265676 1488
rect 268660 1436 268712 1488
rect 268844 1479 268896 1488
rect 268844 1445 268853 1479
rect 268853 1445 268887 1479
rect 268887 1445 268896 1479
rect 268844 1436 268896 1445
rect 269488 1436 269540 1488
rect 271328 1436 271380 1488
rect 272248 1436 272300 1488
rect 272340 1436 272392 1488
rect 273812 1436 273864 1488
rect 279516 1479 279568 1488
rect 279516 1445 279525 1479
rect 279525 1445 279559 1479
rect 279559 1445 279568 1479
rect 279516 1436 279568 1445
rect 280252 1436 280304 1488
rect 281724 1436 281776 1488
rect 282092 1436 282144 1488
rect 282184 1436 282236 1488
rect 289360 1436 289412 1488
rect 290372 1436 290424 1488
rect 293960 1436 294012 1488
rect 294788 1436 294840 1488
rect 295340 1436 295392 1488
rect 296812 1436 296864 1488
rect 299940 1436 299992 1488
rect 309232 1436 309284 1488
rect 309968 1436 310020 1488
rect 318432 1479 318484 1488
rect 318432 1445 318441 1479
rect 318441 1445 318475 1479
rect 318475 1445 318484 1479
rect 318432 1436 318484 1445
rect 320272 1436 320324 1488
rect 329748 1436 329800 1488
rect 356336 1436 356388 1488
rect 385316 1436 385368 1488
rect 451924 1436 451976 1488
rect 309324 1368 309376 1420
rect 309784 1368 309836 1420
rect 356796 1368 356848 1420
rect 565820 1368 565872 1420
rect 225512 1300 225564 1352
rect 153844 1164 153896 1216
rect 154212 1096 154264 1148
rect 157524 1096 157576 1148
rect 158444 1096 158496 1148
rect 160560 1096 160612 1148
rect 161112 1164 161164 1216
rect 161296 1164 161348 1216
rect 178960 1164 179012 1216
rect 179236 1164 179288 1216
rect 183928 1164 183980 1216
rect 189448 1164 189500 1216
rect 190552 1164 190604 1216
rect 190920 1164 190972 1216
rect 224776 1164 224828 1216
rect 232412 1232 232464 1284
rect 233056 1232 233108 1284
rect 233148 1232 233200 1284
rect 238116 1232 238168 1284
rect 239128 1275 239180 1284
rect 239128 1241 239137 1275
rect 239137 1241 239171 1275
rect 239171 1241 239180 1275
rect 239312 1275 239364 1284
rect 239128 1232 239180 1241
rect 239312 1241 239321 1275
rect 239321 1241 239355 1275
rect 239355 1241 239364 1275
rect 239312 1232 239364 1241
rect 239772 1232 239824 1284
rect 239864 1232 239916 1284
rect 241244 1232 241296 1284
rect 241336 1232 241388 1284
rect 253112 1232 253164 1284
rect 253296 1232 253348 1284
rect 254032 1232 254084 1284
rect 254124 1232 254176 1284
rect 256516 1232 256568 1284
rect 256608 1232 256660 1284
rect 260380 1232 260432 1284
rect 260472 1232 260524 1284
rect 271328 1232 271380 1284
rect 272156 1232 272208 1284
rect 272340 1275 272392 1284
rect 272340 1241 272349 1275
rect 272349 1241 272383 1275
rect 272383 1241 272392 1275
rect 272340 1232 272392 1241
rect 273812 1275 273864 1284
rect 273812 1241 273821 1275
rect 273821 1241 273855 1275
rect 273855 1241 273864 1275
rect 273812 1232 273864 1241
rect 273904 1232 273956 1284
rect 279516 1232 279568 1284
rect 296720 1232 296772 1284
rect 238024 1164 238076 1216
rect 238392 1164 238444 1216
rect 238576 1164 238628 1216
rect 238944 1164 238996 1216
rect 251364 1164 251416 1216
rect 260564 1164 260616 1216
rect 270592 1164 270644 1216
rect 270776 1164 270828 1216
rect 279884 1164 279936 1216
rect 281908 1164 281960 1216
rect 290188 1164 290240 1216
rect 290556 1164 290608 1216
rect 291016 1164 291068 1216
rect 300676 1164 300728 1216
rect 318432 1164 318484 1216
rect 327540 1232 327592 1284
rect 329656 1232 329708 1284
rect 357992 1232 358044 1284
rect 365260 1232 365312 1284
rect 338304 1164 338356 1216
rect 354036 1164 354088 1216
rect 356980 1164 357032 1216
rect 424968 1232 425020 1284
rect 480168 1232 480220 1284
rect 492496 1232 492548 1284
rect 492680 1232 492732 1284
rect 512000 1232 512052 1284
rect 535368 1232 535420 1284
rect 549168 1232 549220 1284
rect 568304 1300 568356 1352
rect 564440 1232 564492 1284
rect 493968 1164 494020 1216
rect 494244 1164 494296 1216
rect 569500 1164 569552 1216
rect 161020 1096 161072 1148
rect 166908 1096 166960 1148
rect 169024 1096 169076 1148
rect 217968 1096 218020 1148
rect 223764 1096 223816 1148
rect 223856 1139 223908 1148
rect 223856 1105 223865 1139
rect 223865 1105 223899 1139
rect 223899 1105 223908 1139
rect 223856 1096 223908 1105
rect 224040 1096 224092 1148
rect 225052 1096 225104 1148
rect 225236 1096 225288 1148
rect 225512 1139 225564 1148
rect 225512 1105 225521 1139
rect 225521 1105 225555 1139
rect 225555 1105 225564 1139
rect 225512 1096 225564 1105
rect 148876 1028 148928 1080
rect 239220 1071 239272 1080
rect 239220 1037 239229 1071
rect 239229 1037 239263 1071
rect 239263 1037 239272 1071
rect 239220 1028 239272 1037
rect 245568 1028 245620 1080
rect 247132 1028 247184 1080
rect 247500 1028 247552 1080
rect 248236 1028 248288 1080
rect 125600 960 125652 1012
rect 3332 892 3384 944
rect 56784 892 56836 944
rect 58072 892 58124 944
rect 61200 892 61252 944
rect 62948 892 63000 944
rect 64880 892 64932 944
rect 68928 892 68980 944
rect 70676 892 70728 944
rect 1124 824 1176 876
rect 4988 824 5040 876
rect 28264 824 28316 876
rect 42156 824 42208 876
rect 46664 824 46716 876
rect 3056 756 3108 808
rect 19432 799 19484 808
rect 19432 765 19441 799
rect 19441 765 19475 799
rect 19475 765 19484 799
rect 19432 756 19484 765
rect 29736 756 29788 808
rect 38200 756 38252 808
rect 42064 756 42116 808
rect 43352 756 43404 808
rect 63776 824 63828 876
rect 63868 824 63920 876
rect 76472 892 76524 944
rect 97264 892 97316 944
rect 76840 824 76892 876
rect 82544 824 82596 876
rect 82728 824 82780 876
rect 48044 756 48096 808
rect 55220 756 55272 808
rect 79048 756 79100 808
rect 83832 824 83884 876
rect 84752 824 84804 876
rect 87880 824 87932 876
rect 93492 824 93544 876
rect 94044 824 94096 876
rect 97080 824 97132 876
rect 101680 892 101732 944
rect 116584 892 116636 944
rect 117136 892 117188 944
rect 122564 892 122616 944
rect 123484 892 123536 944
rect 123576 892 123628 944
rect 131672 960 131724 1012
rect 129096 935 129148 944
rect 129096 901 129105 935
rect 129105 901 129139 935
rect 129139 901 129148 935
rect 129096 892 129148 901
rect 129464 892 129516 944
rect 140504 935 140556 944
rect 140504 901 140513 935
rect 140513 901 140547 935
rect 140547 901 140556 935
rect 140504 892 140556 901
rect 142436 892 142488 944
rect 146116 960 146168 1012
rect 149520 892 149572 944
rect 152372 892 152424 944
rect 154120 892 154172 944
rect 154396 892 154448 944
rect 155132 892 155184 944
rect 83648 756 83700 808
rect 848 688 900 740
rect 13268 688 13320 740
rect 15200 688 15252 740
rect 17960 688 18012 740
rect 92664 756 92716 808
rect 92848 756 92900 808
rect 93032 756 93084 808
rect 101404 756 101456 808
rect 103428 824 103480 876
rect 106464 824 106516 876
rect 108856 824 108908 876
rect 101956 756 102008 808
rect 106924 756 106976 808
rect 107016 756 107068 808
rect 83832 688 83884 740
rect 100760 688 100812 740
rect 102416 688 102468 740
rect 102692 688 102744 740
rect 107844 688 107896 740
rect 108028 756 108080 808
rect 109408 824 109460 876
rect 109960 824 110012 876
rect 110052 824 110104 876
rect 111524 688 111576 740
rect 111616 688 111668 740
rect 112352 756 112404 808
rect 112812 756 112864 808
rect 113548 756 113600 808
rect 113732 756 113784 808
rect 120540 756 120592 808
rect 120724 799 120776 808
rect 120724 765 120733 799
rect 120733 765 120767 799
rect 120767 765 120776 799
rect 120724 756 120776 765
rect 122472 756 122524 808
rect 122564 756 122616 808
rect 152096 756 152148 808
rect 153476 756 153528 808
rect 112076 688 112128 740
rect 152188 688 152240 740
rect 1308 620 1360 672
rect 112 552 164 604
rect 4896 552 4948 604
rect 7380 620 7432 672
rect 10508 552 10560 604
rect 13452 552 13504 604
rect 22192 552 22244 604
rect 26700 620 26752 672
rect 46756 620 46808 672
rect 46940 620 46992 672
rect 59360 620 59412 672
rect 60004 620 60056 672
rect 75644 620 75696 672
rect 52828 552 52880 604
rect 3608 484 3660 536
rect 1032 416 1084 468
rect 4988 484 5040 536
rect 73252 484 73304 536
rect 93400 595 93452 604
rect 93400 561 93409 595
rect 93409 561 93443 595
rect 93443 561 93452 595
rect 93400 552 93452 561
rect 93860 552 93912 604
rect 103060 552 103112 604
rect 122196 620 122248 672
rect 150256 663 150308 672
rect 150256 629 150265 663
rect 150265 629 150299 663
rect 150299 629 150308 663
rect 150256 620 150308 629
rect 153568 688 153620 740
rect 156604 731 156656 740
rect 156604 697 156613 731
rect 156613 697 156647 731
rect 156647 697 156656 731
rect 156604 688 156656 697
rect 156788 731 156840 740
rect 156788 697 156797 731
rect 156797 697 156831 731
rect 156831 697 156840 731
rect 156788 688 156840 697
rect 241980 960 242032 1012
rect 296904 960 296956 1012
rect 306932 960 306984 1012
rect 318616 960 318668 1012
rect 319444 960 319496 1012
rect 319536 960 319588 1012
rect 327724 960 327776 1012
rect 327816 960 327868 1012
rect 329564 960 329616 1012
rect 162584 892 162636 944
rect 160836 756 160888 808
rect 160744 688 160796 740
rect 169484 756 169536 808
rect 163228 688 163280 740
rect 163872 688 163924 740
rect 163964 688 164016 740
rect 26884 280 26936 332
rect 35164 280 35216 332
rect 92572 416 92624 468
rect 92756 416 92808 468
rect 157340 620 157392 672
rect 157616 663 157668 672
rect 157616 629 157625 663
rect 157625 629 157659 663
rect 157659 629 157668 663
rect 157616 620 157668 629
rect 157800 620 157852 672
rect 159456 620 159508 672
rect 160928 620 160980 672
rect 163136 620 163188 672
rect 166172 620 166224 672
rect 166632 620 166684 672
rect 175648 756 175700 808
rect 177580 824 177632 876
rect 177764 824 177816 876
rect 179604 824 179656 876
rect 179696 824 179748 876
rect 180616 824 180668 876
rect 180708 824 180760 876
rect 317696 892 317748 944
rect 328736 892 328788 944
rect 328828 892 328880 944
rect 331680 960 331732 1012
rect 331772 960 331824 1012
rect 335728 960 335780 1012
rect 335820 960 335872 1012
rect 329748 892 329800 944
rect 343088 892 343140 944
rect 352196 1028 352248 1080
rect 372804 1028 372856 1080
rect 413652 1028 413704 1080
rect 453304 1028 453356 1080
rect 480168 1028 480220 1080
rect 501328 1028 501380 1080
rect 512644 1028 512696 1080
rect 535368 1028 535420 1080
rect 349528 892 349580 944
rect 356244 892 356296 944
rect 568212 960 568264 1012
rect 169668 688 169720 740
rect 175924 688 175976 740
rect 176016 688 176068 740
rect 183744 756 183796 808
rect 208216 756 208268 808
rect 213828 756 213880 808
rect 219348 756 219400 808
rect 219440 756 219492 808
rect 232964 756 233016 808
rect 178316 688 178368 740
rect 180156 688 180208 740
rect 180248 688 180300 740
rect 184020 688 184072 740
rect 221372 688 221424 740
rect 176108 620 176160 672
rect 175924 595 175976 604
rect 175924 561 175933 595
rect 175933 561 175967 595
rect 175967 561 175976 595
rect 175924 552 175976 561
rect 175740 484 175792 536
rect 176660 620 176712 672
rect 177120 620 177172 672
rect 177948 620 178000 672
rect 183560 620 183612 672
rect 204352 620 204404 672
rect 207756 620 207808 672
rect 207848 620 207900 672
rect 214104 620 214156 672
rect 215024 620 215076 672
rect 217600 620 217652 672
rect 219440 620 219492 672
rect 219624 620 219676 672
rect 221096 620 221148 672
rect 224224 620 224276 672
rect 224408 663 224460 672
rect 224408 629 224417 663
rect 224417 629 224451 663
rect 224451 629 224460 663
rect 224408 620 224460 629
rect 224592 620 224644 672
rect 225328 620 225380 672
rect 231492 620 231544 672
rect 238484 756 238536 808
rect 239220 756 239272 808
rect 286232 824 286284 876
rect 287520 824 287572 876
rect 289636 824 289688 876
rect 293776 824 293828 876
rect 306748 824 306800 876
rect 309968 824 310020 876
rect 310060 824 310112 876
rect 231676 620 231728 672
rect 233148 620 233200 672
rect 251916 620 251968 672
rect 252008 620 252060 672
rect 252836 620 252888 672
rect 259276 620 259328 672
rect 261576 620 261628 672
rect 267004 620 267056 672
rect 267188 620 267240 672
rect 270960 620 271012 672
rect 271144 688 271196 740
rect 273352 688 273404 740
rect 290280 688 290332 740
rect 290372 688 290424 740
rect 295156 688 295208 740
rect 373908 892 373960 944
rect 380164 892 380216 944
rect 389364 892 389416 944
rect 512000 892 512052 944
rect 538956 892 539008 944
rect 569408 892 569460 944
rect 373080 824 373132 876
rect 319720 756 319772 808
rect 356520 756 356572 808
rect 372528 756 372580 808
rect 406108 756 406160 808
rect 407028 756 407080 808
rect 411260 756 411312 808
rect 425704 756 425756 808
rect 280068 620 280120 672
rect 281540 620 281592 672
rect 286048 620 286100 672
rect 289728 620 289780 672
rect 296996 620 297048 672
rect 300676 620 300728 672
rect 300768 620 300820 672
rect 434996 688 435048 740
rect 442816 688 442868 740
rect 335360 620 335412 672
rect 335544 620 335596 672
rect 476764 756 476816 808
rect 486148 756 486200 808
rect 518716 756 518768 808
rect 476396 688 476448 740
rect 490196 688 490248 740
rect 547236 620 547288 672
rect 176200 527 176252 536
rect 176200 493 176209 527
rect 176209 493 176243 527
rect 176243 493 176252 527
rect 176200 484 176252 493
rect 480720 552 480772 604
rect 509884 552 509936 604
rect 516876 552 516928 604
rect 184020 484 184072 536
rect 217508 484 217560 536
rect 217692 484 217744 536
rect 217784 484 217836 536
rect 217968 484 218020 536
rect 241796 484 241848 536
rect 246580 484 246632 536
rect 247040 484 247092 536
rect 247500 484 247552 536
rect 135444 416 135496 468
rect 142252 416 142304 468
rect 142344 416 142396 468
rect 144736 416 144788 468
rect 89536 348 89588 400
rect 90732 348 90784 400
rect 91100 348 91152 400
rect 94228 348 94280 400
rect 95884 348 95936 400
rect 111892 348 111944 400
rect 112076 348 112128 400
rect 153200 348 153252 400
rect 153752 348 153804 400
rect 154672 348 154724 400
rect 157248 348 157300 400
rect 176292 391 176344 400
rect 176292 357 176301 391
rect 176301 357 176335 391
rect 176335 357 176344 391
rect 176292 348 176344 357
rect 193496 416 193548 468
rect 198372 416 198424 468
rect 198464 459 198516 468
rect 198464 425 198473 459
rect 198473 425 198507 459
rect 198507 425 198516 459
rect 198464 416 198516 425
rect 198740 416 198792 468
rect 203156 416 203208 468
rect 211988 416 212040 468
rect 241704 416 241756 468
rect 247224 416 247276 468
rect 49148 280 49200 332
rect 58992 280 59044 332
rect 193588 348 193640 400
rect 196624 348 196676 400
rect 196992 348 197044 400
rect 198188 348 198240 400
rect 198280 391 198332 400
rect 198280 357 198289 391
rect 198289 357 198323 391
rect 198323 357 198332 391
rect 198280 348 198332 357
rect 251732 416 251784 468
rect 252836 416 252888 468
rect 253112 416 253164 468
rect 259184 416 259236 468
rect 261760 484 261812 536
rect 265440 484 265492 536
rect 270776 527 270828 536
rect 270776 493 270785 527
rect 270785 493 270819 527
rect 270819 493 270828 527
rect 270776 484 270828 493
rect 271880 484 271932 536
rect 279332 484 279384 536
rect 260012 416 260064 468
rect 260564 416 260616 468
rect 261208 416 261260 468
rect 262864 416 262916 468
rect 262956 416 263008 468
rect 264888 416 264940 468
rect 269028 416 269080 468
rect 269488 416 269540 468
rect 270684 416 270736 468
rect 270776 348 270828 400
rect 280344 416 280396 468
rect 281540 416 281592 468
rect 285588 416 285640 468
rect 285680 416 285732 468
rect 290096 484 290148 536
rect 293868 484 293920 536
rect 290188 416 290240 468
rect 327908 484 327960 536
rect 318892 416 318944 468
rect 318984 416 319036 468
rect 323032 416 323084 468
rect 376668 484 376720 536
rect 381544 484 381596 536
rect 393412 484 393464 536
rect 337844 416 337896 468
rect 489828 416 489880 468
rect 1400 212 1452 264
rect 10416 212 10468 264
rect 25320 212 25372 264
rect 3056 144 3108 196
rect 38384 212 38436 264
rect 53196 212 53248 264
rect 55588 212 55640 264
rect 55680 212 55732 264
rect 61016 212 61068 264
rect 66904 212 66956 264
rect 66996 212 67048 264
rect 67364 212 67416 264
rect 73528 255 73580 264
rect 73528 221 73537 255
rect 73537 221 73571 255
rect 73571 221 73580 255
rect 73528 212 73580 221
rect 151360 212 151412 264
rect 151728 212 151780 264
rect 184020 280 184072 332
rect 288900 280 288952 332
rect 376668 348 376720 400
rect 377036 348 377088 400
rect 528192 348 528244 400
rect 499672 280 499724 332
rect 509240 212 509292 264
rect 49884 144 49936 196
rect 58624 144 58676 196
rect 58992 144 59044 196
rect 69296 144 69348 196
rect 83464 144 83516 196
rect 84476 144 84528 196
rect 84660 144 84712 196
rect 87696 144 87748 196
rect 112168 144 112220 196
rect 183468 144 183520 196
rect 183928 144 183980 196
rect 569224 144 569276 196
rect 9864 76 9916 128
rect 44364 76 44416 128
rect 46296 76 46348 128
rect 55404 76 55456 128
rect 13084 8 13136 60
rect 17408 8 17460 60
rect 568856 76 568908 128
rect 473360 8 473412 60
rect 473728 8 473780 60
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 40512 700534 40540 703520
rect 105464 700670 105492 703520
rect 170324 700738 170352 703520
rect 129648 700732 129700 700738
rect 129648 700674 129700 700680
rect 170312 700732 170364 700738
rect 170312 700674 170364 700680
rect 105452 700664 105504 700670
rect 105452 700606 105504 700612
rect 106188 700664 106240 700670
rect 106188 700606 106240 700612
rect 110328 700664 110380 700670
rect 110328 700606 110380 700612
rect 89628 700596 89680 700602
rect 89628 700538 89680 700544
rect 40500 700528 40552 700534
rect 40500 700470 40552 700476
rect 41328 700528 41380 700534
rect 41328 700470 41380 700476
rect 70308 700528 70360 700534
rect 70308 700470 70360 700476
rect 31668 700392 31720 700398
rect 31668 700334 31720 700340
rect 10968 700324 11020 700330
rect 10968 700266 11020 700272
rect 1398 682272 1454 682281
rect 1398 682207 1454 682216
rect 1412 677550 1440 682207
rect 10980 680898 11008 700266
rect 31680 684486 31708 700334
rect 30380 684480 30432 684486
rect 30380 684422 30432 684428
rect 31668 684480 31720 684486
rect 31668 684422 31720 684428
rect 10810 680870 11008 680898
rect 30392 680884 30420 684422
rect 41340 683806 41368 700470
rect 50988 700460 51040 700466
rect 50988 700402 51040 700408
rect 51000 684486 51028 700402
rect 50068 684480 50120 684486
rect 50068 684422 50120 684428
rect 50988 684480 51040 684486
rect 50988 684422 51040 684428
rect 41328 683800 41380 683806
rect 41328 683742 41380 683748
rect 50080 680884 50108 684422
rect 70320 680762 70348 700470
rect 89640 680898 89668 700538
rect 106200 683874 106228 700606
rect 110340 684078 110368 700606
rect 129660 684486 129688 700674
rect 235184 700670 235212 703520
rect 235172 700664 235224 700670
rect 235172 700606 235224 700612
rect 300136 700602 300164 703520
rect 300124 700596 300176 700602
rect 300124 700538 300176 700544
rect 364996 700534 365024 703520
rect 364984 700528 365036 700534
rect 364984 700470 365036 700476
rect 429856 700466 429884 703520
rect 429844 700460 429896 700466
rect 429844 700402 429896 700408
rect 494808 700398 494836 703520
rect 494796 700392 494848 700398
rect 494796 700334 494848 700340
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 128636 684480 128688 684486
rect 128636 684422 128688 684428
rect 129648 684480 129700 684486
rect 129648 684422 129700 684428
rect 109040 684072 109092 684078
rect 109040 684014 109092 684020
rect 110328 684072 110380 684078
rect 110328 684014 110380 684020
rect 106188 683868 106240 683874
rect 106188 683810 106240 683816
rect 89378 680870 89668 680898
rect 109052 680884 109080 684014
rect 128648 680884 128676 684422
rect 148324 683868 148376 683874
rect 148324 683810 148376 683816
rect 148336 680884 148364 683810
rect 168012 683800 168064 683806
rect 168012 683742 168064 683748
rect 168024 680884 168052 683742
rect 285956 683256 286008 683262
rect 285956 683198 286008 683204
rect 295248 683256 295300 683262
rect 295248 683198 295300 683204
rect 364524 683256 364576 683262
rect 364524 683198 364576 683204
rect 375380 683256 375432 683262
rect 375380 683198 375432 683204
rect 384212 683256 384264 683262
rect 384212 683198 384264 683204
rect 391204 683256 391256 683262
rect 391204 683198 391256 683204
rect 403900 683256 403952 683262
rect 403900 683198 403952 683204
rect 408408 683256 408460 683262
rect 408408 683198 408460 683204
rect 462872 683256 462924 683262
rect 462872 683198 462924 683204
rect 471980 683256 472032 683262
rect 471980 683198 472032 683204
rect 482468 683256 482520 683262
rect 482468 683198 482520 683204
rect 494060 683256 494112 683262
rect 494060 683198 494112 683204
rect 187608 683188 187660 683194
rect 187608 683130 187660 683136
rect 187620 680884 187648 683130
rect 285968 680884 285996 683198
rect 69690 680734 70348 680762
rect 226708 680400 226760 680406
rect 207032 680338 207322 680354
rect 246212 680400 246264 680406
rect 226760 680348 227010 680354
rect 226708 680342 227010 680348
rect 265900 680400 265952 680406
rect 246264 680348 246606 680354
rect 246212 680342 246606 680348
rect 265952 680348 266294 680354
rect 265900 680342 266294 680348
rect 207020 680332 207322 680338
rect 207072 680326 207322 680332
rect 226720 680326 227010 680342
rect 246224 680326 246606 680342
rect 265912 680326 266294 680342
rect 295260 680338 295288 683198
rect 305920 681012 305972 681018
rect 305920 680954 305972 680960
rect 327632 681012 327684 681018
rect 327632 680954 327684 680960
rect 305932 680898 305960 680954
rect 305578 680870 305960 680898
rect 325606 680504 325662 680513
rect 325266 680462 325606 680490
rect 325606 680439 325662 680448
rect 296718 680368 296774 680377
rect 295248 680332 295300 680338
rect 207020 680274 207072 680280
rect 327644 680338 327672 680954
rect 364536 680884 364564 683198
rect 345018 680640 345074 680649
rect 344954 680598 345018 680626
rect 345018 680575 345074 680584
rect 364798 680368 364854 680377
rect 296718 680303 296720 680312
rect 295248 680274 295300 680280
rect 296772 680303 296774 680312
rect 327632 680332 327684 680338
rect 296720 680274 296772 680280
rect 364798 680303 364800 680312
rect 327632 680274 327684 680280
rect 364852 680303 364854 680312
rect 370226 680368 370282 680377
rect 375392 680338 375420 683198
rect 384224 680884 384252 683198
rect 379426 680640 379482 680649
rect 379426 680575 379428 680584
rect 379480 680575 379482 680584
rect 381636 680604 381688 680610
rect 379428 680546 379480 680552
rect 381636 680546 381688 680552
rect 380072 680400 380124 680406
rect 380070 680368 380072 680377
rect 381648 680377 381676 680546
rect 391216 680406 391244 683198
rect 403912 680884 403940 683198
rect 391204 680400 391256 680406
rect 380124 680368 380126 680377
rect 370226 680303 370228 680312
rect 364800 680274 364852 680280
rect 370280 680303 370282 680312
rect 375380 680332 375432 680338
rect 370228 680274 370280 680280
rect 380070 680303 380126 680312
rect 381634 680368 381690 680377
rect 394700 680400 394752 680406
rect 391204 680342 391256 680348
rect 394698 680368 394700 680377
rect 403164 680400 403216 680406
rect 394752 680368 394754 680377
rect 381634 680303 381690 680312
rect 394698 680303 394754 680312
rect 403162 680368 403164 680377
rect 403216 680368 403218 680377
rect 408420 680338 408448 683198
rect 439502 680912 439558 680921
rect 462884 680884 462912 683198
rect 439502 680847 439558 680856
rect 412732 680400 412784 680406
rect 412730 680368 412732 680377
rect 418620 680400 418672 680406
rect 412784 680368 412786 680377
rect 403162 680303 403218 680312
rect 408408 680332 408460 680338
rect 375380 680274 375432 680280
rect 412730 680303 412786 680312
rect 418618 680368 418620 680377
rect 423588 680400 423640 680406
rect 418672 680368 418674 680377
rect 423522 680348 423588 680354
rect 428188 680400 428240 680406
rect 423522 680342 423640 680348
rect 428186 680368 428188 680377
rect 437756 680400 437808 680406
rect 428240 680368 428242 680377
rect 423522 680326 423628 680342
rect 418618 680303 418674 680312
rect 428186 680303 428242 680312
rect 437754 680368 437756 680377
rect 439516 680377 439544 680847
rect 466642 680504 466698 680513
rect 463792 680468 463844 680474
rect 466642 680439 466644 680448
rect 463792 680410 463844 680416
rect 466696 680439 466698 680448
rect 466644 680410 466696 680416
rect 443552 680400 443604 680406
rect 437808 680368 437810 680377
rect 437754 680303 437810 680312
rect 439502 680368 439558 680377
rect 443210 680348 443552 680354
rect 451372 680400 451424 680406
rect 443210 680342 443604 680348
rect 451370 680368 451372 680377
rect 457168 680400 457220 680406
rect 451424 680368 451426 680377
rect 443210 680326 443592 680342
rect 439502 680303 439558 680312
rect 451370 680303 451426 680312
rect 457166 680368 457168 680377
rect 457220 680368 457222 680377
rect 457166 680303 457222 680312
rect 463698 680368 463754 680377
rect 463804 680354 463832 680410
rect 471992 680406 472020 683198
rect 482480 680884 482508 683198
rect 494072 680406 494100 683198
rect 569868 683188 569920 683194
rect 569868 683130 569920 683136
rect 564714 681048 564770 681057
rect 564714 680983 564770 680992
rect 543830 680640 543886 680649
rect 543830 680575 543886 680584
rect 557446 680640 557502 680649
rect 557446 680575 557448 680584
rect 466552 680400 466604 680406
rect 463754 680326 463832 680354
rect 466550 680368 466552 680377
rect 471980 680400 472032 680406
rect 466604 680368 466606 680377
rect 463698 680303 463754 680312
rect 494060 680400 494112 680406
rect 471980 680342 472032 680348
rect 481178 680368 481234 680377
rect 466550 680303 466606 680312
rect 481178 680303 481180 680312
rect 408408 680274 408460 680280
rect 481232 680303 481234 680312
rect 485778 680368 485834 680377
rect 495440 680400 495492 680406
rect 494060 680342 494112 680348
rect 495438 680368 495440 680377
rect 502248 680400 502300 680406
rect 495492 680368 495494 680377
rect 485778 680303 485780 680312
rect 481180 680274 481232 680280
rect 485832 680303 485834 680312
rect 502182 680348 502248 680354
rect 505928 680400 505980 680406
rect 502182 680342 502300 680348
rect 505926 680368 505928 680377
rect 515404 680400 515456 680406
rect 505980 680368 505982 680377
rect 502182 680326 502288 680342
rect 495438 680303 495494 680312
rect 505926 680303 505982 680312
rect 515402 680368 515404 680377
rect 522120 680400 522172 680406
rect 515456 680368 515458 680377
rect 521870 680348 522120 680354
rect 524420 680400 524472 680406
rect 521870 680342 522172 680348
rect 524418 680368 524420 680377
rect 534356 680400 534408 680406
rect 524472 680368 524474 680377
rect 521870 680326 522160 680342
rect 515402 680303 515458 680312
rect 524418 680303 524474 680312
rect 534354 680368 534356 680377
rect 541808 680400 541860 680406
rect 534408 680368 534410 680377
rect 541466 680348 541808 680354
rect 543844 680377 543872 680575
rect 557500 680575 557502 680584
rect 559378 680640 559434 680649
rect 559378 680575 559434 680584
rect 563244 680604 563296 680610
rect 557448 680546 557500 680552
rect 554778 680504 554834 680513
rect 554778 680439 554834 680448
rect 559194 680504 559250 680513
rect 559392 680474 559420 680575
rect 563244 680546 563296 680552
rect 563256 680513 563284 680546
rect 564728 680513 564756 680983
rect 561586 680504 561642 680513
rect 559194 680439 559250 680448
rect 559380 680468 559432 680474
rect 544016 680400 544068 680406
rect 541466 680342 541860 680348
rect 543830 680368 543886 680377
rect 541466 680326 541848 680342
rect 534354 680303 534410 680312
rect 543830 680303 543886 680312
rect 544014 680368 544016 680377
rect 544068 680368 544070 680377
rect 554792 680338 554820 680439
rect 554870 680368 554926 680377
rect 544014 680303 544070 680312
rect 554780 680332 554832 680338
rect 485780 680274 485832 680280
rect 554870 680303 554872 680312
rect 554780 680274 554832 680280
rect 554924 680303 554926 680312
rect 558550 680368 558606 680377
rect 559208 680338 559236 680439
rect 561586 680439 561642 680448
rect 561770 680504 561826 680513
rect 561770 680439 561826 680448
rect 563242 680504 563298 680513
rect 563242 680439 563298 680448
rect 564714 680504 564770 680513
rect 564714 680439 564770 680448
rect 559380 680410 559432 680416
rect 560758 680368 560814 680377
rect 558550 680303 558552 680312
rect 554872 680274 554924 680280
rect 558604 680303 558606 680312
rect 559196 680332 559248 680338
rect 558552 680274 558604 680280
rect 561218 680368 561274 680377
rect 561154 680326 561218 680354
rect 560758 680303 560760 680312
rect 559196 680274 559248 680280
rect 560812 680303 560814 680312
rect 561600 680338 561628 680439
rect 561784 680338 561812 680439
rect 561862 680368 561918 680377
rect 561218 680303 561274 680312
rect 561588 680332 561640 680338
rect 560760 680274 560812 680280
rect 561588 680274 561640 680280
rect 561772 680332 561824 680338
rect 561862 680303 561864 680312
rect 561772 680274 561824 680280
rect 561916 680303 561918 680312
rect 562506 680368 562562 680377
rect 562506 680303 562508 680312
rect 561864 680274 561916 680280
rect 562560 680303 562562 680312
rect 566370 680368 566426 680377
rect 566370 680303 566372 680312
rect 562508 680274 562560 680280
rect 566424 680303 566426 680312
rect 566372 680274 566424 680280
rect 1952 679856 2004 679862
rect 1952 679798 2004 679804
rect 1860 679040 1912 679046
rect 1860 678982 1912 678988
rect 204 677544 256 677550
rect 204 677486 256 677492
rect 1400 677544 1452 677550
rect 1400 677486 1452 677492
rect 18 624608 74 624617
rect 18 624543 74 624552
rect 32 287026 60 624543
rect 110 352200 166 352209
rect 110 352135 166 352144
rect 20 287020 72 287026
rect 20 286962 72 286968
rect 124 216850 152 352135
rect 112 216844 164 216850
rect 112 216786 164 216792
rect 18 215792 74 215801
rect 18 215727 74 215736
rect 32 36145 60 215727
rect 216 174622 244 677486
rect 1872 672466 1900 678982
rect 1964 676190 1992 679798
rect 3424 679788 3476 679794
rect 3424 679730 3476 679736
rect 2504 679652 2556 679658
rect 2504 679594 2556 679600
rect 2228 679108 2280 679114
rect 2228 679050 2280 679056
rect 1952 676184 2004 676190
rect 1952 676126 2004 676132
rect 1952 676048 2004 676054
rect 1952 675990 2004 675996
rect 1964 674370 1992 675990
rect 1964 674342 2176 674370
rect 1872 672438 2084 672466
rect 1122 669488 1178 669497
rect 1122 669423 1178 669432
rect 1032 469804 1084 469810
rect 1032 469746 1084 469752
rect 754 442368 810 442377
rect 754 442303 810 442312
rect 570 374368 626 374377
rect 570 374303 626 374312
rect 480 294636 532 294642
rect 480 294578 532 294584
rect 296 266348 348 266354
rect 296 266290 348 266296
rect 308 221218 336 266290
rect 388 264308 440 264314
rect 388 264250 440 264256
rect 400 221406 428 264250
rect 492 241670 520 294578
rect 584 257310 612 374303
rect 662 329080 718 329089
rect 662 329015 718 329024
rect 572 257304 624 257310
rect 572 257246 624 257252
rect 572 251864 624 251870
rect 572 251806 624 251812
rect 480 241664 532 241670
rect 480 241606 532 241612
rect 480 235476 532 235482
rect 480 235418 532 235424
rect 388 221400 440 221406
rect 388 221342 440 221348
rect 308 221190 428 221218
rect 296 199504 348 199510
rect 296 199446 348 199452
rect 308 182850 336 199446
rect 296 182844 348 182850
rect 296 182786 348 182792
rect 400 176118 428 221190
rect 388 176112 440 176118
rect 388 176054 440 176060
rect 204 174616 256 174622
rect 492 174570 520 235418
rect 584 214198 612 251806
rect 572 214192 624 214198
rect 572 214134 624 214140
rect 570 208176 626 208185
rect 570 208111 626 208120
rect 584 205086 612 208111
rect 572 205080 624 205086
rect 572 205022 624 205028
rect 572 200252 624 200258
rect 572 200194 624 200200
rect 204 174558 256 174564
rect 400 174542 520 174570
rect 204 174480 256 174486
rect 204 174422 256 174428
rect 112 171012 164 171018
rect 112 170954 164 170960
rect 124 152046 152 170954
rect 112 152040 164 152046
rect 112 151982 164 151988
rect 112 147144 164 147150
rect 112 147086 164 147092
rect 124 47530 152 147086
rect 216 138582 244 174422
rect 400 167686 428 174542
rect 480 170332 532 170338
rect 480 170274 532 170280
rect 388 167680 440 167686
rect 388 167622 440 167628
rect 492 166190 520 170274
rect 480 166184 532 166190
rect 480 166126 532 166132
rect 388 165912 440 165918
rect 388 165854 440 165860
rect 400 153882 428 165854
rect 480 163940 532 163946
rect 480 163882 532 163888
rect 492 155446 520 163882
rect 480 155440 532 155446
rect 480 155382 532 155388
rect 388 153876 440 153882
rect 388 153818 440 153824
rect 388 152040 440 152046
rect 388 151982 440 151988
rect 400 147150 428 151982
rect 480 148776 532 148782
rect 480 148718 532 148724
rect 388 147144 440 147150
rect 388 147086 440 147092
rect 388 147008 440 147014
rect 388 146950 440 146956
rect 296 145648 348 145654
rect 296 145590 348 145596
rect 204 138576 256 138582
rect 204 138518 256 138524
rect 204 66972 256 66978
rect 204 66914 256 66920
rect 112 47524 164 47530
rect 112 47466 164 47472
rect 18 36136 74 36145
rect 18 36071 74 36080
rect 20 35012 72 35018
rect 20 34954 72 34960
rect 32 1630 60 34954
rect 112 29912 164 29918
rect 112 29854 164 29860
rect 124 24274 152 29854
rect 112 24268 164 24274
rect 112 24210 164 24216
rect 112 20188 164 20194
rect 112 20130 164 20136
rect 20 1624 72 1630
rect 20 1566 72 1572
rect 124 610 152 20130
rect 216 649 244 66914
rect 202 640 258 649
rect 112 604 164 610
rect 202 575 258 584
rect 112 546 164 552
rect 308 377 336 145590
rect 400 126342 428 146950
rect 388 126336 440 126342
rect 388 126278 440 126284
rect 388 126132 440 126138
rect 388 126074 440 126080
rect 400 98190 428 126074
rect 492 103465 520 148718
rect 584 146266 612 200194
rect 676 195158 704 329015
rect 768 257446 796 442303
rect 938 397352 994 397361
rect 938 397287 994 397296
rect 756 257440 808 257446
rect 756 257382 808 257388
rect 848 251864 900 251870
rect 848 251806 900 251812
rect 756 221672 808 221678
rect 756 221614 808 221620
rect 664 195152 716 195158
rect 664 195094 716 195100
rect 664 193996 716 194002
rect 664 193938 716 193944
rect 572 146260 624 146266
rect 572 146202 624 146208
rect 676 146146 704 193938
rect 768 163334 796 221614
rect 860 209982 888 251806
rect 848 209976 900 209982
rect 848 209918 900 209924
rect 848 199504 900 199510
rect 848 199446 900 199452
rect 756 163328 808 163334
rect 756 163270 808 163276
rect 756 161628 808 161634
rect 756 161570 808 161576
rect 768 159118 796 161570
rect 756 159112 808 159118
rect 756 159054 808 159060
rect 756 147008 808 147014
rect 756 146950 808 146956
rect 584 146118 704 146146
rect 584 141778 612 146118
rect 664 141908 716 141914
rect 664 141850 716 141856
rect 572 141772 624 141778
rect 572 141714 624 141720
rect 572 141636 624 141642
rect 572 141578 624 141584
rect 478 103456 534 103465
rect 478 103391 534 103400
rect 388 98184 440 98190
rect 388 98126 440 98132
rect 480 96280 532 96286
rect 480 96222 532 96228
rect 388 35284 440 35290
rect 388 35226 440 35232
rect 400 513 428 35226
rect 492 18290 520 96222
rect 584 93158 612 141578
rect 676 138666 704 141850
rect 768 138786 796 146950
rect 860 141914 888 199446
rect 952 197674 980 397287
rect 940 197668 992 197674
rect 940 197610 992 197616
rect 940 197532 992 197538
rect 940 197474 992 197480
rect 848 141908 900 141914
rect 848 141850 900 141856
rect 848 141772 900 141778
rect 848 141714 900 141720
rect 756 138780 808 138786
rect 756 138722 808 138728
rect 676 138638 796 138666
rect 664 138576 716 138582
rect 664 138518 716 138524
rect 572 93152 624 93158
rect 572 93094 624 93100
rect 572 80980 624 80986
rect 572 80922 624 80928
rect 584 78985 612 80922
rect 570 78976 626 78985
rect 570 78911 626 78920
rect 572 72616 624 72622
rect 572 72558 624 72564
rect 480 18284 532 18290
rect 480 18226 532 18232
rect 478 18048 534 18057
rect 478 17983 534 17992
rect 492 10282 520 17983
rect 584 10402 612 72558
rect 676 33590 704 138518
rect 768 124642 796 138638
rect 860 128926 888 141714
rect 952 134706 980 197474
rect 1044 167278 1072 469746
rect 1136 261526 1164 669423
rect 2056 658186 2084 672438
rect 1964 658158 2084 658186
rect 1964 648650 1992 658158
rect 1860 648644 1912 648650
rect 1860 648586 1912 648592
rect 1952 648644 2004 648650
rect 1952 648586 2004 648592
rect 1872 647986 1900 648586
rect 1952 648100 2004 648106
rect 2148 648088 2176 674342
rect 2004 648060 2176 648088
rect 1952 648042 2004 648048
rect 1872 647958 1992 647986
rect 1214 646776 1270 646785
rect 1214 646711 1270 646720
rect 1124 261520 1176 261526
rect 1124 261462 1176 261468
rect 1124 260772 1176 260778
rect 1124 260714 1176 260720
rect 1032 167272 1084 167278
rect 1032 167214 1084 167220
rect 1032 166796 1084 166802
rect 1032 166738 1084 166744
rect 1044 163810 1072 166738
rect 1032 163804 1084 163810
rect 1032 163746 1084 163752
rect 1032 159588 1084 159594
rect 1032 159530 1084 159536
rect 1044 143002 1072 159530
rect 1032 142996 1084 143002
rect 1032 142938 1084 142944
rect 1032 142860 1084 142866
rect 1032 142802 1084 142808
rect 940 134700 992 134706
rect 940 134642 992 134648
rect 1044 134570 1072 142802
rect 1032 134564 1084 134570
rect 1032 134506 1084 134512
rect 940 134428 992 134434
rect 940 134370 992 134376
rect 848 128920 900 128926
rect 848 128862 900 128868
rect 848 126336 900 126342
rect 848 126278 900 126284
rect 756 124636 808 124642
rect 756 124578 808 124584
rect 756 121236 808 121242
rect 756 121178 808 121184
rect 664 33584 716 33590
rect 664 33526 716 33532
rect 662 32328 718 32337
rect 662 32263 718 32272
rect 676 10402 704 32263
rect 768 19961 796 121178
rect 754 19952 810 19961
rect 754 19887 810 19896
rect 756 19848 808 19854
rect 756 19790 808 19796
rect 572 10396 624 10402
rect 572 10338 624 10344
rect 664 10396 716 10402
rect 664 10338 716 10344
rect 492 10254 704 10282
rect 480 10192 532 10198
rect 480 10134 532 10140
rect 492 8702 520 10134
rect 480 8696 532 8702
rect 480 8638 532 8644
rect 570 7848 626 7857
rect 570 7783 626 7792
rect 386 504 442 513
rect 584 480 612 7783
rect 676 785 704 10254
rect 768 4758 796 19790
rect 860 11898 888 126278
rect 952 121242 980 134370
rect 1032 133340 1084 133346
rect 1032 133282 1084 133288
rect 940 121236 992 121242
rect 940 121178 992 121184
rect 940 121100 992 121106
rect 940 121042 992 121048
rect 848 11892 900 11898
rect 848 11834 900 11840
rect 848 10532 900 10538
rect 848 10474 900 10480
rect 860 10146 888 10474
rect 952 10266 980 121042
rect 1044 50386 1072 133282
rect 1032 50380 1084 50386
rect 1032 50322 1084 50328
rect 1032 37052 1084 37058
rect 1032 36994 1084 37000
rect 1044 20058 1072 36994
rect 1032 20052 1084 20058
rect 1032 19994 1084 20000
rect 1032 18420 1084 18426
rect 1032 18362 1084 18368
rect 1044 10402 1072 18362
rect 1136 16726 1164 260714
rect 1228 207738 1256 646711
rect 1964 642666 1992 647958
rect 2240 646898 2268 679050
rect 2516 677090 2544 679594
rect 2332 677062 2544 677090
rect 2332 652746 2360 677062
rect 3436 655194 3464 679730
rect 568224 679658 568436 679674
rect 568224 679652 568448 679658
rect 568224 679646 568396 679652
rect 3700 679176 3752 679182
rect 3700 679118 3752 679124
rect 3712 676274 3740 679118
rect 3712 676246 3832 676274
rect 3804 666618 3832 676246
rect 568224 673418 568252 679646
rect 568396 679594 568448 679600
rect 569224 679108 569276 679114
rect 569224 679050 569276 679056
rect 568224 673390 568344 673418
rect 3620 666590 3832 666618
rect 3620 659682 3648 666590
rect 568316 663898 568344 673390
rect 568316 663870 568528 663898
rect 3620 659654 3832 659682
rect 3344 655166 3464 655194
rect 3344 653426 3372 655166
rect 3344 653398 3556 653426
rect 2332 652718 2544 652746
rect 2056 646870 2268 646898
rect 1952 642660 2004 642666
rect 1952 642602 2004 642608
rect 2056 641866 2084 646870
rect 1964 641850 2084 641866
rect 1952 641844 2084 641850
rect 2004 641838 2084 641844
rect 1952 641786 2004 641792
rect 2516 641730 2544 652718
rect 3528 648666 3556 653398
rect 3804 648666 3832 659654
rect 568500 659002 568528 663870
rect 569236 659138 569264 679050
rect 569880 674812 569908 683130
rect 572720 679176 572772 679182
rect 572720 679118 572772 679124
rect 571432 679040 571484 679046
rect 571432 678982 571484 678988
rect 571444 677550 571472 678982
rect 571432 677544 571484 677550
rect 571432 677486 571484 677492
rect 569788 674784 569908 674812
rect 569788 663762 569816 674784
rect 572732 667457 572760 679118
rect 578148 677544 578200 677550
rect 578148 677486 578200 677492
rect 578160 674830 578188 677486
rect 578148 674824 578200 674830
rect 578148 674766 578200 674772
rect 580172 674824 580224 674830
rect 580172 674766 580224 674772
rect 580184 674665 580212 674766
rect 580170 674656 580226 674665
rect 580170 674591 580226 674600
rect 572718 667448 572774 667457
rect 572718 667383 572774 667392
rect 569788 663734 569908 663762
rect 569880 659274 569908 663734
rect 569880 659258 570000 659274
rect 569880 659252 570012 659258
rect 569880 659246 569960 659252
rect 569960 659194 570012 659200
rect 569236 659110 570000 659138
rect 3528 648638 3648 648666
rect 1872 641702 2544 641730
rect 1872 641050 1900 641702
rect 1952 641640 2004 641646
rect 1952 641582 2004 641588
rect 1964 641186 1992 641582
rect 1964 641158 2360 641186
rect 1872 641022 2176 641050
rect 1952 639328 2004 639334
rect 1952 639270 2004 639276
rect 1860 633480 1912 633486
rect 1860 633422 1912 633428
rect 1582 623792 1638 623801
rect 1582 623727 1638 623736
rect 1596 618322 1624 623727
rect 1872 618322 1900 633422
rect 1964 632482 1992 639270
rect 2148 632618 2176 641022
rect 2332 632890 2360 641158
rect 3620 639146 3648 648638
rect 3436 639118 3648 639146
rect 3712 648638 3832 648666
rect 568316 658974 568528 659002
rect 3436 639010 3464 639118
rect 3344 638982 3464 639010
rect 3344 635474 3372 638982
rect 3068 635446 3372 635474
rect 2332 632862 2636 632890
rect 2148 632590 2360 632618
rect 1964 632454 2176 632482
rect 2148 618882 2176 632454
rect 2148 618854 2268 618882
rect 2240 618610 2268 618854
rect 2148 618582 2268 618610
rect 1584 618316 1636 618322
rect 1584 618258 1636 618264
rect 1676 618316 1728 618322
rect 1676 618258 1728 618264
rect 1860 618316 1912 618322
rect 1860 618258 1912 618264
rect 1952 618316 2004 618322
rect 1952 618258 2004 618264
rect 1582 601080 1638 601089
rect 1582 601015 1638 601024
rect 1596 600982 1624 601015
rect 1584 600976 1636 600982
rect 1584 600918 1636 600924
rect 1688 592006 1716 618258
rect 1964 608734 1992 618258
rect 1952 608728 2004 608734
rect 1952 608670 2004 608676
rect 1860 608592 1912 608598
rect 1860 608534 1912 608540
rect 1872 596306 1900 608534
rect 2148 602562 2176 618582
rect 1964 602534 2176 602562
rect 1964 602410 1992 602534
rect 1952 602404 2004 602410
rect 1952 602346 2004 602352
rect 2332 602154 2360 632590
rect 2608 618338 2636 632862
rect 3068 622826 3096 635446
rect 3712 634658 3740 648638
rect 568316 640370 568344 658974
rect 569972 654226 570000 659110
rect 569960 654220 570012 654226
rect 569960 654162 570012 654168
rect 577504 654220 577556 654226
rect 577504 654162 577556 654168
rect 569960 654084 570012 654090
rect 569960 654026 570012 654032
rect 569972 653970 570000 654026
rect 569696 653942 570000 653970
rect 569696 647170 569724 653942
rect 569604 647142 569724 647170
rect 568316 640342 568436 640370
rect 3620 634630 3740 634658
rect 3620 623778 3648 634630
rect 3528 623750 3648 623778
rect 3068 622798 3372 622826
rect 1964 602138 2360 602154
rect 1952 602132 2360 602138
rect 2004 602126 2360 602132
rect 2424 618310 2636 618338
rect 1952 602074 2004 602080
rect 2424 602018 2452 618310
rect 1964 602002 2452 602018
rect 1952 601996 2452 602002
rect 2004 601990 2452 601996
rect 1952 601938 2004 601944
rect 3344 601882 3372 622798
rect 3528 613578 3556 623750
rect 568408 621058 568436 640342
rect 569604 630442 569632 647142
rect 572718 640248 572774 640257
rect 572718 640183 572774 640192
rect 569604 630414 570092 630442
rect 569960 630216 570012 630222
rect 568224 621030 568436 621058
rect 568868 630164 569960 630170
rect 568868 630158 570012 630164
rect 568868 630142 570000 630158
rect 3528 613550 3740 613578
rect 3712 612762 3740 613550
rect 568224 613442 568252 621030
rect 568868 620922 568896 630142
rect 570064 625274 570092 630414
rect 572732 630222 572760 640183
rect 572720 630216 572772 630222
rect 572720 630158 572772 630164
rect 577516 627910 577544 654162
rect 577504 627904 577556 627910
rect 577504 627846 577556 627852
rect 579712 627904 579764 627910
rect 579712 627846 579764 627852
rect 579724 627745 579752 627846
rect 579710 627736 579766 627745
rect 579710 627671 579766 627680
rect 568776 620894 568896 620922
rect 569788 625246 570092 625274
rect 568224 613414 568344 613442
rect 3712 612734 3832 612762
rect 3804 602426 3832 612734
rect 568316 604330 568344 613414
rect 568776 610994 568804 620894
rect 569788 613034 569816 625246
rect 569788 613006 570092 613034
rect 568776 610966 568896 610994
rect 568868 610722 568896 610966
rect 568776 610694 568896 610722
rect 568316 604302 568620 604330
rect 1964 601854 3372 601882
rect 3620 602398 3832 602426
rect 1964 601118 1992 601854
rect 1952 601112 2004 601118
rect 1952 601054 2004 601060
rect 1952 600976 2004 600982
rect 2004 600936 2176 600964
rect 1952 600918 2004 600924
rect 2148 600794 2176 600936
rect 2148 600766 2544 600794
rect 2516 600658 2544 600766
rect 2976 600766 3372 600794
rect 2976 600658 3004 600766
rect 2516 600630 3004 600658
rect 1952 600568 2004 600574
rect 2004 600516 2360 600522
rect 1952 600510 2360 600516
rect 1964 600494 2360 600510
rect 2332 599978 2360 600494
rect 2332 599950 2728 599978
rect 1952 599888 2004 599894
rect 2004 599848 2636 599876
rect 1952 599830 2004 599836
rect 1952 599752 2004 599758
rect 1952 599694 2004 599700
rect 1964 599162 1992 599694
rect 1964 599134 2452 599162
rect 2424 597258 2452 599134
rect 2608 598890 2636 599848
rect 2240 597230 2452 597258
rect 2516 598862 2636 598890
rect 1952 597032 2004 597038
rect 1952 596974 2004 596980
rect 1964 596578 1992 596974
rect 2240 596578 2268 597230
rect 1964 596550 2176 596578
rect 2240 596550 2452 596578
rect 2148 596306 2176 596550
rect 1872 596278 1992 596306
rect 2148 596278 2360 596306
rect 1676 592000 1728 592006
rect 1676 591942 1728 591948
rect 1860 592000 1912 592006
rect 1860 591942 1912 591948
rect 1872 580258 1900 591942
rect 1964 580514 1992 596278
rect 2332 591954 2360 596278
rect 2424 591988 2452 596550
rect 2516 593450 2544 598862
rect 2700 598074 2728 599950
rect 2700 598046 2820 598074
rect 2516 593422 2728 593450
rect 2424 591960 2544 591988
rect 2148 591926 2360 591954
rect 1952 580508 2004 580514
rect 1952 580450 2004 580456
rect 2148 580258 2176 591926
rect 1780 580230 1900 580258
rect 1964 580242 2176 580258
rect 1952 580236 2176 580242
rect 1582 578368 1638 578377
rect 1582 578303 1638 578312
rect 1596 577318 1624 578303
rect 1584 577312 1636 577318
rect 1584 577254 1636 577260
rect 1780 569242 1808 580230
rect 2004 580230 2176 580236
rect 1952 580178 2004 580184
rect 2516 578354 2544 591960
rect 1688 569214 1808 569242
rect 1872 578326 2544 578354
rect 1872 569242 1900 578326
rect 1952 577312 2004 577318
rect 2004 577272 2636 577300
rect 1952 577254 2004 577260
rect 1964 569362 2268 569378
rect 1952 569356 2268 569362
rect 2004 569350 2268 569356
rect 1952 569298 2004 569304
rect 2240 569242 2268 569350
rect 2608 569242 2636 577272
rect 1872 569214 2176 569242
rect 2240 569214 2636 569242
rect 1306 567352 1362 567361
rect 1306 567287 1362 567296
rect 1320 564126 1348 567287
rect 1308 564120 1360 564126
rect 1308 564062 1360 564068
rect 1584 556232 1636 556238
rect 1582 556200 1584 556209
rect 1636 556200 1638 556209
rect 1582 556135 1638 556144
rect 1582 533080 1638 533089
rect 1582 533015 1638 533024
rect 1596 526386 1624 533015
rect 1688 527134 1716 569214
rect 1768 569152 1820 569158
rect 1768 569094 1820 569100
rect 1780 563530 1808 569094
rect 2148 567202 2176 569214
rect 2148 567174 2268 567202
rect 1860 566636 1912 566642
rect 1860 566578 1912 566584
rect 1872 563786 1900 566578
rect 2240 565570 2268 567174
rect 1964 565554 2268 565570
rect 1952 565548 2268 565554
rect 2004 565542 2268 565548
rect 1952 565490 2004 565496
rect 2700 565434 2728 593422
rect 2792 579714 2820 598046
rect 3344 594810 3372 600766
rect 3252 594782 3372 594810
rect 3252 592906 3280 594782
rect 3252 592878 3464 592906
rect 2792 579686 2912 579714
rect 2884 579578 2912 579686
rect 2884 579550 3188 579578
rect 3160 576722 3188 579550
rect 3068 576694 3188 576722
rect 3068 576586 3096 576694
rect 2976 576558 3096 576586
rect 2976 572370 3004 576558
rect 3436 572370 3464 592878
rect 3620 591988 3648 602398
rect 568592 595082 568620 604302
rect 568316 595054 568620 595082
rect 568316 594946 568344 595054
rect 568224 594918 568344 594946
rect 3620 591960 3740 591988
rect 3712 591818 3740 591960
rect 3712 591790 3832 591818
rect 2884 572342 3004 572370
rect 3252 572342 3464 572370
rect 2884 570466 2912 572342
rect 3252 570738 3280 572342
rect 3068 570710 3280 570738
rect 2884 570438 3004 570466
rect 2976 570058 3004 570438
rect 3068 570194 3096 570710
rect 3068 570166 3188 570194
rect 3160 570058 3188 570166
rect 2976 570030 3740 570058
rect 3160 565978 3188 570030
rect 3160 565950 3372 565978
rect 1964 565406 2728 565434
rect 1964 564466 1992 565406
rect 1952 564460 2004 564466
rect 1952 564402 2004 564408
rect 1952 564120 2004 564126
rect 2004 564068 2728 564074
rect 1952 564062 2728 564068
rect 1964 564046 2728 564062
rect 1860 563780 1912 563786
rect 1860 563722 1912 563728
rect 1780 563502 2544 563530
rect 1952 563440 2004 563446
rect 1952 563382 2004 563388
rect 1964 563258 1992 563382
rect 1964 563230 2452 563258
rect 1952 563168 2004 563174
rect 2004 563116 2268 563122
rect 1952 563110 2268 563116
rect 1964 563094 2268 563110
rect 1952 561128 2004 561134
rect 2004 561076 2176 561082
rect 1952 561070 2176 561076
rect 1964 561054 2176 561070
rect 1952 556232 2004 556238
rect 1952 556174 2004 556180
rect 1860 547732 1912 547738
rect 1860 547674 1912 547680
rect 1872 534070 1900 547674
rect 1860 534064 1912 534070
rect 1860 534006 1912 534012
rect 1860 533860 1912 533866
rect 1860 533802 1912 533808
rect 1676 527128 1728 527134
rect 1676 527070 1728 527076
rect 1768 526992 1820 526998
rect 1768 526934 1820 526940
rect 1584 526380 1636 526386
rect 1584 526322 1636 526328
rect 1490 510640 1546 510649
rect 1490 510575 1546 510584
rect 1398 465080 1454 465089
rect 1398 465015 1454 465024
rect 1412 459882 1440 465015
rect 1400 459876 1452 459882
rect 1400 459818 1452 459824
rect 1398 452432 1454 452441
rect 1398 452367 1454 452376
rect 1412 448662 1440 452367
rect 1400 448656 1452 448662
rect 1400 448598 1452 448604
rect 1400 425604 1452 425610
rect 1400 425546 1452 425552
rect 1412 419898 1440 425546
rect 1400 419892 1452 419898
rect 1400 419834 1452 419840
rect 1398 419792 1454 419801
rect 1398 419727 1454 419736
rect 1412 414662 1440 419727
rect 1400 414656 1452 414662
rect 1400 414598 1452 414604
rect 1400 405476 1452 405482
rect 1400 405418 1452 405424
rect 1412 398478 1440 405418
rect 1400 398472 1452 398478
rect 1400 398414 1452 398420
rect 1398 395040 1454 395049
rect 1398 394975 1454 394984
rect 1412 387122 1440 394975
rect 1400 387116 1452 387122
rect 1400 387058 1452 387064
rect 1400 386980 1452 386986
rect 1400 386922 1452 386928
rect 1412 380594 1440 386922
rect 1400 380588 1452 380594
rect 1400 380530 1452 380536
rect 1400 358420 1452 358426
rect 1400 358362 1452 358368
rect 1412 352986 1440 358362
rect 1400 352980 1452 352986
rect 1400 352922 1452 352928
rect 1400 340196 1452 340202
rect 1400 340138 1452 340144
rect 1306 337512 1362 337521
rect 1306 337447 1362 337456
rect 1320 333742 1348 337447
rect 1308 333736 1360 333742
rect 1308 333678 1360 333684
rect 1412 331566 1440 340138
rect 1400 331560 1452 331566
rect 1400 331502 1452 331508
rect 1398 306368 1454 306377
rect 1398 306303 1454 306312
rect 1308 296268 1360 296274
rect 1308 296210 1360 296216
rect 1320 264042 1348 296210
rect 1412 296002 1440 306303
rect 1400 295996 1452 296002
rect 1400 295938 1452 295944
rect 1398 294400 1454 294409
rect 1398 294335 1454 294344
rect 1412 283966 1440 294335
rect 1400 283960 1452 283966
rect 1400 283902 1452 283908
rect 1398 283792 1454 283801
rect 1398 283727 1454 283736
rect 1308 264036 1360 264042
rect 1308 263978 1360 263984
rect 1412 261594 1440 283727
rect 1400 261588 1452 261594
rect 1400 261530 1452 261536
rect 1398 261080 1454 261089
rect 1398 261015 1454 261024
rect 1412 258262 1440 261015
rect 1400 258256 1452 258262
rect 1400 258198 1452 258204
rect 1400 257440 1452 257446
rect 1400 257382 1452 257388
rect 1412 251818 1440 257382
rect 1320 251790 1440 251818
rect 1320 249014 1348 251790
rect 1398 251288 1454 251297
rect 1398 251223 1454 251232
rect 1308 249008 1360 249014
rect 1308 248950 1360 248956
rect 1306 238368 1362 238377
rect 1306 238303 1362 238312
rect 1320 221542 1348 238303
rect 1412 221678 1440 251223
rect 1400 221672 1452 221678
rect 1400 221614 1452 221620
rect 1308 221536 1360 221542
rect 1400 221536 1452 221542
rect 1308 221478 1360 221484
rect 1398 221504 1400 221513
rect 1452 221504 1454 221513
rect 1398 221439 1454 221448
rect 1400 221332 1452 221338
rect 1400 221274 1452 221280
rect 1412 217462 1440 221274
rect 1400 217456 1452 217462
rect 1400 217398 1452 217404
rect 1306 214568 1362 214577
rect 1306 214503 1362 214512
rect 1216 207732 1268 207738
rect 1216 207674 1268 207680
rect 1216 205080 1268 205086
rect 1216 205022 1268 205028
rect 1228 194954 1256 205022
rect 1320 195566 1348 214503
rect 1400 214328 1452 214334
rect 1400 214270 1452 214276
rect 1412 204950 1440 214270
rect 1400 204944 1452 204950
rect 1400 204886 1452 204892
rect 1400 204808 1452 204814
rect 1400 204750 1452 204756
rect 1412 200258 1440 204750
rect 1400 200252 1452 200258
rect 1400 200194 1452 200200
rect 1400 198280 1452 198286
rect 1398 198248 1400 198257
rect 1452 198248 1454 198257
rect 1398 198183 1454 198192
rect 1400 198076 1452 198082
rect 1400 198018 1452 198024
rect 1308 195560 1360 195566
rect 1308 195502 1360 195508
rect 1216 194948 1268 194954
rect 1216 194890 1268 194896
rect 1306 193080 1362 193089
rect 1306 193015 1362 193024
rect 1216 182912 1268 182918
rect 1216 182854 1268 182860
rect 1228 175642 1256 182854
rect 1216 175636 1268 175642
rect 1216 175578 1268 175584
rect 1216 171964 1268 171970
rect 1216 171906 1268 171912
rect 1228 146962 1256 171906
rect 1320 161634 1348 193015
rect 1412 171970 1440 198018
rect 1504 195702 1532 510575
rect 1582 509960 1638 509969
rect 1780 509930 1808 526934
rect 1582 509895 1638 509904
rect 1768 509924 1820 509930
rect 1596 505238 1624 509895
rect 1768 509866 1820 509872
rect 1872 509810 1900 533802
rect 1964 529242 1992 556174
rect 1952 529236 2004 529242
rect 1952 529178 2004 529184
rect 2148 527762 2176 561054
rect 2240 556050 2268 563094
rect 2240 556022 2360 556050
rect 2332 541090 2360 556022
rect 1964 527746 2176 527762
rect 1952 527740 2176 527746
rect 2004 527734 2176 527740
rect 2240 541062 2360 541090
rect 1952 527682 2004 527688
rect 2240 527218 2268 541062
rect 2424 536738 2452 563230
rect 2516 550746 2544 563502
rect 2700 554826 2728 564046
rect 2700 554798 3096 554826
rect 2516 550718 3004 550746
rect 2976 550474 3004 550718
rect 3068 550610 3096 554798
rect 3068 550582 3280 550610
rect 1964 527202 2268 527218
rect 1952 527196 2268 527202
rect 2004 527190 2268 527196
rect 2332 536710 2452 536738
rect 2792 550446 3004 550474
rect 1952 527138 2004 527144
rect 2332 526538 2360 536710
rect 1964 526522 2360 526538
rect 1952 526516 2360 526522
rect 2004 526510 2360 526516
rect 1952 526458 2004 526464
rect 1964 526386 2728 526402
rect 1952 526380 2728 526386
rect 2004 526374 2728 526380
rect 1952 526322 2004 526328
rect 1952 526176 2004 526182
rect 2004 526124 2544 526130
rect 1952 526118 2544 526124
rect 1964 526102 2544 526118
rect 1952 522504 2004 522510
rect 2004 522452 2268 522458
rect 1952 522446 2268 522452
rect 1964 522430 2268 522446
rect 1952 522368 2004 522374
rect 2004 522316 2176 522322
rect 1952 522310 2176 522316
rect 1964 522294 2176 522310
rect 1952 510672 2004 510678
rect 2004 510620 2084 510626
rect 1952 510614 2084 510620
rect 1964 510598 2084 510614
rect 2056 510082 2084 510598
rect 1964 510066 2084 510082
rect 1952 510060 2084 510066
rect 2004 510054 2084 510060
rect 1952 510002 2004 510008
rect 1952 509924 2004 509930
rect 2148 509912 2176 522294
rect 2004 509884 2176 509912
rect 1952 509866 2004 509872
rect 1780 509782 1900 509810
rect 1676 509584 1728 509590
rect 1676 509526 1728 509532
rect 1584 505232 1636 505238
rect 1584 505174 1636 505180
rect 1688 502314 1716 509526
rect 1780 504150 1808 509782
rect 2240 507362 2268 522430
rect 2516 514842 2544 526102
rect 2700 516202 2728 526374
rect 1964 507346 2268 507362
rect 1952 507340 2268 507346
rect 2004 507334 2268 507340
rect 2332 514814 2544 514842
rect 2608 516174 2728 516202
rect 1952 507282 2004 507288
rect 2332 507226 2360 514814
rect 1964 507210 2360 507226
rect 1952 507204 2360 507210
rect 2004 507198 2360 507204
rect 1952 507146 2004 507152
rect 2608 506546 2636 516174
rect 1964 506518 2636 506546
rect 1964 506122 1992 506518
rect 1952 506116 2004 506122
rect 1952 506058 2004 506064
rect 2792 505458 2820 550446
rect 3252 545714 3280 550582
rect 3068 545686 3280 545714
rect 3068 510762 3096 545686
rect 3068 510734 3280 510762
rect 1872 505430 2820 505458
rect 1872 504914 1900 505430
rect 1952 505232 2004 505238
rect 2004 505180 3004 505186
rect 1952 505174 3004 505180
rect 1964 505158 3004 505174
rect 1872 504886 2820 504914
rect 1952 504824 2004 504830
rect 2004 504784 2084 504812
rect 1952 504766 2004 504772
rect 1860 504484 1912 504490
rect 1860 504426 1912 504432
rect 1768 504144 1820 504150
rect 1768 504086 1820 504092
rect 1676 502308 1728 502314
rect 1676 502250 1728 502256
rect 1872 497842 1900 504426
rect 1952 502240 2004 502246
rect 1952 502182 2004 502188
rect 1964 501922 1992 502182
rect 2056 502058 2084 504784
rect 2056 502030 2728 502058
rect 1964 501894 2544 501922
rect 1952 501832 2004 501838
rect 2004 501780 2360 501786
rect 1952 501774 2360 501780
rect 1964 501758 2360 501774
rect 1872 497814 2176 497842
rect 1768 497548 1820 497554
rect 1768 497490 1820 497496
rect 1952 497548 2004 497554
rect 1952 497490 2004 497496
rect 1582 487792 1638 487801
rect 1582 487727 1638 487736
rect 1492 195696 1544 195702
rect 1492 195638 1544 195644
rect 1492 195560 1544 195566
rect 1492 195502 1544 195508
rect 1504 174486 1532 195502
rect 1492 174480 1544 174486
rect 1492 174422 1544 174428
rect 1492 173188 1544 173194
rect 1492 173130 1544 173136
rect 1504 173097 1532 173130
rect 1490 173088 1546 173097
rect 1490 173023 1546 173032
rect 1400 171964 1452 171970
rect 1400 171906 1452 171912
rect 1490 170368 1546 170377
rect 1490 170303 1546 170312
rect 1398 167648 1454 167657
rect 1398 167583 1454 167592
rect 1412 166054 1440 167583
rect 1400 166048 1452 166054
rect 1400 165990 1452 165996
rect 1398 165064 1454 165073
rect 1398 164999 1454 165008
rect 1308 161628 1360 161634
rect 1308 161570 1360 161576
rect 1412 156262 1440 164999
rect 1504 163946 1532 170303
rect 1492 163940 1544 163946
rect 1492 163882 1544 163888
rect 1492 163804 1544 163810
rect 1492 163746 1544 163752
rect 1504 160138 1532 163746
rect 1492 160132 1544 160138
rect 1492 160074 1544 160080
rect 1492 159996 1544 160002
rect 1492 159938 1544 159944
rect 1504 159730 1532 159938
rect 1492 159724 1544 159730
rect 1492 159666 1544 159672
rect 1492 159384 1544 159390
rect 1492 159326 1544 159332
rect 1400 156256 1452 156262
rect 1400 156198 1452 156204
rect 1308 155440 1360 155446
rect 1308 155382 1360 155388
rect 1320 147098 1348 155382
rect 1400 154828 1452 154834
rect 1400 154770 1452 154776
rect 1412 148646 1440 154770
rect 1400 148640 1452 148646
rect 1400 148582 1452 148588
rect 1320 147070 1440 147098
rect 1228 146934 1348 146962
rect 1216 145988 1268 145994
rect 1216 145930 1268 145936
rect 1228 121106 1256 145930
rect 1320 138718 1348 146934
rect 1308 138712 1360 138718
rect 1308 138654 1360 138660
rect 1412 134858 1440 147070
rect 1504 142882 1532 159326
rect 1596 156398 1624 487727
rect 1780 483750 1808 497490
rect 1860 493400 1912 493406
rect 1860 493342 1912 493348
rect 1768 483744 1820 483750
rect 1768 483686 1820 483692
rect 1872 483562 1900 493342
rect 1780 483534 1900 483562
rect 1676 472796 1728 472802
rect 1676 472738 1728 472744
rect 1688 467786 1716 472738
rect 1780 472122 1808 483534
rect 1964 479602 1992 497490
rect 2148 489138 2176 497814
rect 2056 489110 2176 489138
rect 2056 487642 2084 489110
rect 2332 489002 2360 501758
rect 2148 488974 2360 489002
rect 2148 487778 2176 488974
rect 2516 488866 2544 501894
rect 2700 489002 2728 502030
rect 2792 489274 2820 504886
rect 2976 495394 3004 505158
rect 2976 495366 3096 495394
rect 2792 489246 3004 489274
rect 2976 489002 3004 489246
rect 3068 489138 3096 495366
rect 3252 489274 3280 510734
rect 3160 489246 3280 489274
rect 3160 489138 3188 489246
rect 3068 489110 3280 489138
rect 2700 488974 3004 489002
rect 2976 488866 3004 488974
rect 2332 488838 3004 488866
rect 2148 487750 2268 487778
rect 2056 487614 2176 487642
rect 1952 479596 2004 479602
rect 1952 479538 2004 479544
rect 1952 479392 2004 479398
rect 1952 479334 2004 479340
rect 1964 474706 1992 479334
rect 1952 474700 2004 474706
rect 1952 474642 2004 474648
rect 2148 474586 2176 487614
rect 1872 474558 2176 474586
rect 1872 474094 1900 474558
rect 1860 474088 1912 474094
rect 1860 474030 1912 474036
rect 1952 472796 2004 472802
rect 2240 472784 2268 487750
rect 2004 472756 2268 472784
rect 1952 472738 2004 472744
rect 2332 472410 2360 488838
rect 2516 487778 2544 488838
rect 2976 488594 3004 488838
rect 2884 488566 3004 488594
rect 2516 487750 2636 487778
rect 2608 478122 2636 487750
rect 2884 482882 2912 488566
rect 3160 487914 3188 489110
rect 2976 487886 3188 487914
rect 2976 487098 3004 487886
rect 2976 487070 3096 487098
rect 3068 483018 3096 487070
rect 3068 482990 3188 483018
rect 2700 482854 2912 482882
rect 2700 478258 2728 482854
rect 3160 482474 3188 482990
rect 3068 482446 3188 482474
rect 2700 478230 3004 478258
rect 2608 478094 2728 478122
rect 1872 472382 2360 472410
rect 1768 472116 1820 472122
rect 1768 472058 1820 472064
rect 1872 468194 1900 472382
rect 2700 472274 2728 478094
rect 2976 473362 3004 478230
rect 1964 472246 2728 472274
rect 2792 473334 3004 473362
rect 1964 469810 1992 472246
rect 2792 472138 2820 473334
rect 2424 472110 2820 472138
rect 2424 469962 2452 472110
rect 2056 469934 2452 469962
rect 1952 469804 2004 469810
rect 1952 469746 2004 469752
rect 2056 468330 2084 469934
rect 1964 468314 2084 468330
rect 1952 468308 2084 468314
rect 2004 468302 2084 468308
rect 2148 468302 2820 468330
rect 1952 468250 2004 468256
rect 2148 468194 2176 468302
rect 1872 468166 2176 468194
rect 1952 468104 2004 468110
rect 2004 468052 2452 468058
rect 1952 468046 2452 468052
rect 1964 468030 2452 468046
rect 1688 467758 2268 467786
rect 1952 467628 2004 467634
rect 2004 467588 2176 467616
rect 1952 467570 2004 467576
rect 1952 464976 2004 464982
rect 2004 464936 2084 464964
rect 1952 464918 2004 464924
rect 1952 462392 2004 462398
rect 1952 462334 2004 462340
rect 1860 459876 1912 459882
rect 1860 459818 1912 459824
rect 1768 450900 1820 450906
rect 1768 450842 1820 450848
rect 1676 448724 1728 448730
rect 1676 448666 1728 448672
rect 1688 442082 1716 448666
rect 1780 442218 1808 450842
rect 1872 449206 1900 459818
rect 1964 454646 1992 462334
rect 1952 454640 2004 454646
rect 1952 454582 2004 454588
rect 2056 450922 2084 464936
rect 1964 450906 2084 450922
rect 1952 450900 2084 450906
rect 2004 450894 2084 450900
rect 1952 450842 2004 450848
rect 2148 450786 2176 467588
rect 1964 450770 2176 450786
rect 1952 450764 2176 450770
rect 2004 450758 2176 450764
rect 1952 450706 2004 450712
rect 2240 450106 2268 467758
rect 2424 467106 2452 468030
rect 1964 450090 2268 450106
rect 1952 450084 2268 450090
rect 2004 450078 2268 450084
rect 2332 467078 2452 467106
rect 1952 450026 2004 450032
rect 2332 449970 2360 467078
rect 2792 460034 2820 468302
rect 3068 463026 3096 482446
rect 3252 474178 3280 489110
rect 2516 460006 2820 460034
rect 2976 462998 3096 463026
rect 3160 474150 3280 474178
rect 2516 454050 2544 460006
rect 1964 449954 2360 449970
rect 1952 449948 2360 449954
rect 2004 449942 2360 449948
rect 2424 454022 2544 454050
rect 1952 449890 2004 449896
rect 2424 449834 2452 454022
rect 2976 451330 3004 462998
rect 3160 455274 3188 474150
rect 3344 474076 3372 565950
rect 3712 554826 3740 570030
rect 3620 554798 3740 554826
rect 3620 545850 3648 554798
rect 3804 549250 3832 591790
rect 568224 588962 568252 594918
rect 568776 594810 568804 610694
rect 569960 609680 570012 609686
rect 568592 594782 568804 594810
rect 569420 609628 569960 609634
rect 569420 609622 570012 609628
rect 569420 609606 570000 609622
rect 568592 592770 568620 594782
rect 569420 592770 569448 609606
rect 570064 609278 570092 613006
rect 570326 612504 570382 612513
rect 570326 612439 570382 612448
rect 570340 609686 570368 612439
rect 570328 609680 570380 609686
rect 570328 609622 570380 609628
rect 569960 609272 570012 609278
rect 569788 609220 569960 609226
rect 569788 609214 570012 609220
rect 570052 609272 570104 609278
rect 570052 609214 570104 609220
rect 569788 609198 570000 609214
rect 569788 604466 569816 609198
rect 569788 604438 569908 604466
rect 568592 592742 568804 592770
rect 569420 592742 569540 592770
rect 568776 589098 568804 592742
rect 568684 589070 568804 589098
rect 568224 588934 568436 588962
rect 568408 584474 568436 588934
rect 568316 584446 568436 584474
rect 568316 579578 568344 584446
rect 568224 579550 568344 579578
rect 568224 576722 568252 579550
rect 568224 576694 568344 576722
rect 568316 554146 568344 576694
rect 568684 568426 568712 589070
rect 569512 574682 569540 592742
rect 569880 588010 569908 604438
rect 569696 587982 569908 588010
rect 569696 574954 569724 587982
rect 572718 585848 572774 585857
rect 572718 585783 572774 585792
rect 569696 574926 570092 574954
rect 569236 574654 569540 574682
rect 568684 568398 568804 568426
rect 568316 554118 568528 554146
rect 568500 553330 568528 554118
rect 3436 545822 3648 545850
rect 3712 549222 3832 549250
rect 568408 553302 568528 553330
rect 568408 549250 568436 553302
rect 568408 549222 568528 549250
rect 3436 536738 3464 545822
rect 3436 536710 3648 536738
rect 3620 526504 3648 536710
rect 3712 534018 3740 549222
rect 568500 540818 568528 549222
rect 568776 543538 568804 568398
rect 568592 543510 568804 543538
rect 568592 540954 568620 543510
rect 569236 543266 569264 574654
rect 569960 571396 570012 571402
rect 569052 543238 569264 543266
rect 569328 571356 569960 571384
rect 569052 540954 569080 543238
rect 568592 540926 568712 540954
rect 569052 540926 569264 540954
rect 568316 540790 568528 540818
rect 568316 535922 568344 540790
rect 568316 535894 568436 535922
rect 3712 533990 3832 534018
rect 3436 526476 3648 526504
rect 3436 521642 3464 526476
rect 3436 521614 3648 521642
rect 3620 512122 3648 521614
rect 3436 512094 3648 512122
rect 3436 497570 3464 512094
rect 3436 497542 3740 497570
rect 3712 487098 3740 497542
rect 3620 487070 3740 487098
rect 3620 483018 3648 487070
rect 3528 482990 3648 483018
rect 3528 478938 3556 482990
rect 3436 478910 3556 478938
rect 3436 474858 3464 478910
rect 3436 474830 3740 474858
rect 3344 474048 3464 474076
rect 3436 473906 3464 474048
rect 3344 473878 3464 473906
rect 3160 455246 3280 455274
rect 2976 451302 3188 451330
rect 3160 451194 3188 451302
rect 3252 451194 3280 455246
rect 2976 451166 3280 451194
rect 2976 450752 3004 451166
rect 1964 449806 2452 449834
rect 2700 450724 3004 450752
rect 1860 449200 1912 449206
rect 1860 449142 1912 449148
rect 1860 449064 1912 449070
rect 1860 449006 1912 449012
rect 1872 442338 1900 449006
rect 1964 448798 1992 449806
rect 1952 448792 2004 448798
rect 1952 448734 2004 448740
rect 1952 448656 2004 448662
rect 2004 448616 2360 448644
rect 1952 448598 2004 448604
rect 1952 448520 2004 448526
rect 2004 448480 2176 448508
rect 1952 448462 2004 448468
rect 1952 447976 2004 447982
rect 2004 447936 2084 447964
rect 1952 447918 2004 447924
rect 1952 447840 2004 447846
rect 1952 447782 2004 447788
rect 1964 442354 1992 447782
rect 2056 444666 2084 447936
rect 2148 444802 2176 448480
rect 2332 444938 2360 448616
rect 2332 444910 2636 444938
rect 2148 444774 2544 444802
rect 2056 444638 2452 444666
rect 1860 442332 1912 442338
rect 1964 442326 2176 442354
rect 1860 442274 1912 442280
rect 1780 442190 1900 442218
rect 1688 442054 1808 442082
rect 1676 432268 1728 432274
rect 1676 432210 1728 432216
rect 1688 425490 1716 432210
rect 1780 425610 1808 442054
rect 1872 441266 1900 442190
rect 2148 441538 2176 442326
rect 2148 441510 2360 441538
rect 1952 441448 2004 441454
rect 2004 441396 2176 441402
rect 1952 441390 2176 441396
rect 1964 441374 2176 441390
rect 1872 441238 2084 441266
rect 1860 440972 1912 440978
rect 1860 440914 1912 440920
rect 1768 425604 1820 425610
rect 1768 425546 1820 425552
rect 1688 425462 1808 425490
rect 1676 419892 1728 419898
rect 1676 419834 1728 419840
rect 1688 414746 1716 419834
rect 1780 414882 1808 425462
rect 1872 415002 1900 440914
rect 1952 439204 2004 439210
rect 1952 439146 2004 439152
rect 1964 434246 1992 439146
rect 1952 434240 2004 434246
rect 1952 434182 2004 434188
rect 2056 432290 2084 441238
rect 1964 432274 2084 432290
rect 1952 432268 2084 432274
rect 2004 432262 2084 432268
rect 1952 432210 2004 432216
rect 1952 425740 2004 425746
rect 1952 425682 2004 425688
rect 1964 415002 1992 425682
rect 1860 414996 1912 415002
rect 1860 414938 1912 414944
rect 1952 414996 2004 415002
rect 1952 414938 2004 414944
rect 1780 414854 2084 414882
rect 1860 414792 1912 414798
rect 1688 414718 1808 414746
rect 1860 414734 1912 414740
rect 1676 414656 1728 414662
rect 1676 414598 1728 414604
rect 1688 370530 1716 414598
rect 1780 405482 1808 414718
rect 1872 405618 1900 414734
rect 1952 407312 2004 407318
rect 1952 407254 2004 407260
rect 1964 405686 1992 407254
rect 1952 405680 2004 405686
rect 1952 405622 2004 405628
rect 1860 405612 1912 405618
rect 1860 405554 1912 405560
rect 1768 405476 1820 405482
rect 1768 405418 1820 405424
rect 2056 402506 2084 414854
rect 1780 402478 2084 402506
rect 1780 398562 1808 402478
rect 1780 398534 2084 398562
rect 1768 398472 1820 398478
rect 1768 398414 1820 398420
rect 1780 387122 1808 398414
rect 1860 393984 1912 393990
rect 1860 393926 1912 393932
rect 1768 387116 1820 387122
rect 1768 387058 1820 387064
rect 1768 386980 1820 386986
rect 1768 386922 1820 386928
rect 1780 380730 1808 386922
rect 1768 380724 1820 380730
rect 1768 380666 1820 380672
rect 1768 380588 1820 380594
rect 1768 380530 1820 380536
rect 1676 370524 1728 370530
rect 1676 370466 1728 370472
rect 1676 367804 1728 367810
rect 1676 367746 1728 367752
rect 1584 156392 1636 156398
rect 1584 156334 1636 156340
rect 1584 156256 1636 156262
rect 1584 156198 1636 156204
rect 1596 148753 1624 156198
rect 1582 148744 1638 148753
rect 1582 148679 1638 148688
rect 1584 147144 1636 147150
rect 1584 147086 1636 147092
rect 1596 146985 1624 147086
rect 1582 146976 1638 146985
rect 1582 146911 1638 146920
rect 1584 146396 1636 146402
rect 1584 146338 1636 146344
rect 1596 143002 1624 146338
rect 1584 142996 1636 143002
rect 1584 142938 1636 142944
rect 1504 142854 1624 142882
rect 1492 141500 1544 141506
rect 1492 141442 1544 141448
rect 1504 138854 1532 141442
rect 1492 138848 1544 138854
rect 1492 138790 1544 138796
rect 1490 138680 1546 138689
rect 1490 138615 1492 138624
rect 1544 138615 1546 138624
rect 1492 138586 1544 138592
rect 1320 134830 1440 134858
rect 1320 122097 1348 134830
rect 1400 134700 1452 134706
rect 1400 134642 1452 134648
rect 1412 124778 1440 134642
rect 1596 134450 1624 142854
rect 1688 134570 1716 367746
rect 1780 358426 1808 380530
rect 1768 358420 1820 358426
rect 1768 358362 1820 358368
rect 1872 358290 1900 393926
rect 1952 393508 2004 393514
rect 1952 393450 2004 393456
rect 1964 387394 1992 393450
rect 1952 387388 2004 387394
rect 1952 387330 2004 387336
rect 2056 387274 2084 398534
rect 1964 387258 2084 387274
rect 1952 387252 2084 387258
rect 2004 387246 2084 387252
rect 1952 387194 2004 387200
rect 2148 387138 2176 441374
rect 2332 418146 2360 441510
rect 1964 387122 2176 387138
rect 1952 387116 2176 387122
rect 2004 387110 2176 387116
rect 2240 418118 2360 418146
rect 1952 387058 2004 387064
rect 2240 387002 2268 418118
rect 2424 409170 2452 444638
rect 2516 441538 2544 444774
rect 2608 441674 2636 444910
rect 2700 443986 2728 450724
rect 3160 450650 3188 451166
rect 3068 450622 3188 450650
rect 2700 443958 2912 443986
rect 2608 441646 2728 441674
rect 2516 441510 2636 441538
rect 2608 419506 2636 441510
rect 2700 439362 2728 441646
rect 2700 439334 2820 439362
rect 2792 424402 2820 439334
rect 2884 424674 2912 443958
rect 3068 439226 3096 450622
rect 3344 448066 3372 473878
rect 3712 463570 3740 474830
rect 3436 463542 3740 463570
rect 3436 459490 3464 463542
rect 3436 459462 3740 459490
rect 3712 454050 3740 459462
rect 3436 454022 3740 454050
rect 3436 448338 3464 454022
rect 3804 453914 3832 533990
rect 568408 524498 568436 535894
rect 568684 528578 568712 540926
rect 568316 524470 568436 524498
rect 568592 528550 568712 528578
rect 568316 485738 568344 524470
rect 568592 514842 568620 528550
rect 568592 514814 568712 514842
rect 568684 507770 568712 514814
rect 569236 514706 569264 540926
rect 568960 514678 569264 514706
rect 568684 507742 568804 507770
rect 568776 503690 568804 507742
rect 568592 503662 568804 503690
rect 568592 494170 568620 503662
rect 568960 498930 568988 514678
rect 569328 514570 569356 571356
rect 569960 571338 570012 571344
rect 570064 569514 570092 574926
rect 572732 571402 572760 585783
rect 580262 580816 580318 580825
rect 580262 580751 580318 580760
rect 580276 574802 580304 580751
rect 574744 574796 574796 574802
rect 574744 574738 574796 574744
rect 580264 574796 580316 574802
rect 580264 574738 580316 574744
rect 572720 571396 572772 571402
rect 572720 571338 572772 571344
rect 569880 569486 570092 569514
rect 569880 567882 569908 569486
rect 569788 567854 569908 567882
rect 569788 551970 569816 567854
rect 574756 563106 574784 574738
rect 569960 563100 570012 563106
rect 569960 563042 570012 563048
rect 574744 563100 574796 563106
rect 574744 563042 574796 563048
rect 569972 562986 570000 563042
rect 569880 562958 570000 562986
rect 569880 552106 569908 562958
rect 572718 558648 572774 558657
rect 572718 558583 572774 558592
rect 569880 552090 570000 552106
rect 569880 552084 570012 552090
rect 569880 552078 569960 552084
rect 569960 552026 570012 552032
rect 569788 551942 570092 551970
rect 569960 551880 570012 551886
rect 569880 551840 569960 551868
rect 569880 551698 569908 551840
rect 569960 551822 570012 551828
rect 569236 514542 569356 514570
rect 569420 551670 569908 551698
rect 568960 498902 569080 498930
rect 568592 494142 568804 494170
rect 568776 485738 568804 494142
rect 568316 485710 568528 485738
rect 568500 481522 568528 485710
rect 3620 453886 3832 453914
rect 568316 481494 568528 481522
rect 568684 485710 568804 485738
rect 3620 449834 3648 453886
rect 3620 449806 3832 449834
rect 3436 448310 3740 448338
rect 3344 448038 3556 448066
rect 3528 447658 3556 448038
rect 3436 447630 3556 447658
rect 3436 439498 3464 447630
rect 3712 444938 3740 448310
rect 3528 444910 3740 444938
rect 3528 439634 3556 444910
rect 3528 439606 3740 439634
rect 3436 439470 3556 439498
rect 3068 439198 3464 439226
rect 2884 424646 3096 424674
rect 2792 424374 2912 424402
rect 2332 409142 2452 409170
rect 2516 419478 2636 419506
rect 2332 398018 2360 409142
rect 2516 399514 2544 419478
rect 2884 416650 2912 424374
rect 3068 422634 3096 424646
rect 3436 422634 3464 439198
rect 2976 422606 3464 422634
rect 2976 416650 3004 422606
rect 3068 416786 3096 422606
rect 3528 422362 3556 439470
rect 3436 422334 3556 422362
rect 3436 422090 3464 422334
rect 3712 422090 3740 439606
rect 3344 422062 3464 422090
rect 3528 422062 3740 422090
rect 3068 416758 3280 416786
rect 2884 416622 3096 416650
rect 2976 416378 3004 416622
rect 2608 416350 3004 416378
rect 2608 399650 2636 416350
rect 3068 413522 3096 416622
rect 3252 415290 3280 416758
rect 3160 415262 3280 415290
rect 3160 413658 3188 415262
rect 3344 413930 3372 422062
rect 3528 421954 3556 422062
rect 3436 421926 3556 421954
rect 3436 414202 3464 421926
rect 3436 414174 3740 414202
rect 3344 413902 3556 413930
rect 3160 413630 3464 413658
rect 2976 413494 3096 413522
rect 2608 399622 2728 399650
rect 2700 399514 2728 399622
rect 2516 399486 2636 399514
rect 2700 399486 2912 399514
rect 2608 399378 2636 399486
rect 2608 399350 2728 399378
rect 2332 397990 2452 398018
rect 1964 386986 2268 387002
rect 1952 386980 2268 386986
rect 2004 386974 2268 386980
rect 1952 386922 2004 386928
rect 2424 386866 2452 397990
rect 2700 394754 2728 399350
rect 2056 386838 2452 386866
rect 2516 394726 2728 394754
rect 2056 382378 2084 386838
rect 2516 386594 2544 394726
rect 2884 394618 2912 399486
rect 2148 386566 2544 386594
rect 2608 394590 2912 394618
rect 2976 394618 3004 413494
rect 3436 404410 3464 413630
rect 3068 404382 3464 404410
rect 3068 394754 3096 404382
rect 3528 402778 3556 413902
rect 3344 402750 3556 402778
rect 3344 400330 3372 402750
rect 3344 400302 3556 400330
rect 3528 399922 3556 400302
rect 3344 399894 3556 399922
rect 3344 395978 3372 399894
rect 3344 395950 3556 395978
rect 3068 394726 3372 394754
rect 2976 394590 3188 394618
rect 2148 382514 2176 386566
rect 2608 386458 2636 394590
rect 3160 394346 3188 394590
rect 3068 394318 3188 394346
rect 3068 394074 3096 394318
rect 2976 394046 3096 394074
rect 2976 391218 3004 394046
rect 3344 393972 3372 394726
rect 3160 393944 3372 393972
rect 2976 391190 3096 391218
rect 2332 386430 2636 386458
rect 2332 382650 2360 386430
rect 3068 386322 3096 391190
rect 2884 386294 3096 386322
rect 3160 386322 3188 393944
rect 3528 386968 3556 395950
rect 3528 386940 3648 386968
rect 3160 386294 3280 386322
rect 2884 386186 2912 386294
rect 2700 386158 2912 386186
rect 2700 382922 2728 386158
rect 3252 385778 3280 386294
rect 3068 385750 3280 385778
rect 3068 385506 3096 385750
rect 3068 385478 3280 385506
rect 3252 385098 3280 385478
rect 3252 385070 3464 385098
rect 2700 382894 3004 382922
rect 2332 382622 2912 382650
rect 2148 382486 2820 382514
rect 2056 382350 2636 382378
rect 1952 381200 2004 381206
rect 2004 381148 2544 381154
rect 1952 381142 2544 381148
rect 1964 381126 2544 381142
rect 1952 380724 2004 380730
rect 2004 380684 2360 380712
rect 1952 380666 2004 380672
rect 2332 379250 2360 380684
rect 2332 379222 2452 379250
rect 1952 379160 2004 379166
rect 2004 379108 2176 379114
rect 1952 379102 2176 379108
rect 1964 379086 2176 379102
rect 1952 379024 2004 379030
rect 2004 378972 2084 378978
rect 1952 378966 2084 378972
rect 1964 378950 2084 378966
rect 1952 376780 2004 376786
rect 1952 376722 2004 376728
rect 1964 370666 1992 376722
rect 1952 370660 2004 370666
rect 1952 370602 2004 370608
rect 2056 370546 2084 378950
rect 1964 370518 2084 370546
rect 1964 370394 1992 370518
rect 2148 370410 2176 379086
rect 2424 375306 2452 379222
rect 1952 370388 2004 370394
rect 1952 370330 2004 370336
rect 2056 370382 2176 370410
rect 2332 375278 2452 375306
rect 2056 370274 2084 370382
rect 2332 370376 2360 375278
rect 2332 370348 2452 370376
rect 1964 370258 2084 370274
rect 1952 370252 2084 370258
rect 2004 370246 2084 370252
rect 1952 370194 2004 370200
rect 2424 370002 2452 370348
rect 1964 369974 2452 370002
rect 1964 369306 1992 369974
rect 2516 369594 2544 381126
rect 2056 369566 2544 369594
rect 1952 369300 2004 369306
rect 1952 369242 2004 369248
rect 2056 362114 2084 369566
rect 2608 368234 2636 382350
rect 2792 370512 2820 382486
rect 1964 362086 2084 362114
rect 2240 368206 2636 368234
rect 2700 370484 2820 370512
rect 1860 358284 1912 358290
rect 1860 358226 1912 358232
rect 1860 358148 1912 358154
rect 1860 358090 1912 358096
rect 1768 358080 1820 358086
rect 1768 358022 1820 358028
rect 1780 353122 1808 358022
rect 1768 353116 1820 353122
rect 1768 353058 1820 353064
rect 1768 352980 1820 352986
rect 1768 352922 1820 352928
rect 1780 340202 1808 352922
rect 1872 351234 1900 358090
rect 1964 353258 1992 362086
rect 1952 353252 2004 353258
rect 1952 353194 2004 353200
rect 1952 353116 2004 353122
rect 2004 353076 2084 353104
rect 1952 353058 2004 353064
rect 2056 353002 2084 353076
rect 1952 352980 2004 352986
rect 2056 352974 2176 353002
rect 1952 352922 2004 352928
rect 1964 351370 1992 352922
rect 1964 351342 2084 351370
rect 1872 351206 1992 351234
rect 1964 345778 1992 351206
rect 1952 345772 2004 345778
rect 1952 345714 2004 345720
rect 1860 345704 1912 345710
rect 1860 345646 1912 345652
rect 1768 340196 1820 340202
rect 1768 340138 1820 340144
rect 1872 336410 1900 345646
rect 2056 340898 2084 351342
rect 1964 340882 2084 340898
rect 1952 340876 2084 340882
rect 2004 340870 2084 340876
rect 1952 340818 2004 340824
rect 2148 340762 2176 352974
rect 2240 347018 2268 368206
rect 2700 364970 2728 370484
rect 2516 364942 2728 364970
rect 2516 364426 2544 364942
rect 2884 364834 2912 382622
rect 2792 364806 2912 364834
rect 2792 364426 2820 364806
rect 2516 364398 2912 364426
rect 2792 363882 2820 364398
rect 2332 363854 2820 363882
rect 2332 363066 2360 363854
rect 2884 363338 2912 364398
rect 2976 363474 3004 382894
rect 3436 382650 3464 385070
rect 3344 382622 3464 382650
rect 3344 378026 3372 382622
rect 3068 377998 3372 378026
rect 3068 364970 3096 377998
rect 3620 376258 3648 386940
rect 3252 376230 3648 376258
rect 3252 375714 3280 376230
rect 3252 375686 3372 375714
rect 3344 365514 3372 375686
rect 3344 365486 3556 365514
rect 3068 364942 3464 364970
rect 2976 363446 3096 363474
rect 2792 363310 2912 363338
rect 2332 363038 2452 363066
rect 2240 346990 2360 347018
rect 1964 340746 2176 340762
rect 1952 340740 2176 340746
rect 2004 340734 2176 340740
rect 1952 340682 2004 340688
rect 2332 340626 2360 346990
rect 2424 346066 2452 363038
rect 2792 346610 2820 363310
rect 3068 352322 3096 363446
rect 3436 363338 3464 364942
rect 2884 352294 3096 352322
rect 3252 363310 3464 363338
rect 2884 350010 2912 352294
rect 3252 352186 3280 363310
rect 3528 361298 3556 365486
rect 3068 352158 3280 352186
rect 3344 361270 3556 361298
rect 2884 349982 3004 350010
rect 2516 346582 2820 346610
rect 2516 346066 2544 346582
rect 2424 346038 2728 346066
rect 2516 344978 2544 346038
rect 2700 345522 2728 346038
rect 2700 345494 2912 345522
rect 2516 344950 2728 344978
rect 2148 340598 2360 340626
rect 1952 340264 2004 340270
rect 1952 340206 2004 340212
rect 1964 338094 1992 340206
rect 1952 338088 2004 338094
rect 1952 338030 2004 338036
rect 2148 336546 2176 340598
rect 2700 339674 2728 344950
rect 1780 336382 1900 336410
rect 1964 336518 2176 336546
rect 2240 339646 2728 339674
rect 1780 333418 1808 336382
rect 1964 334218 1992 336518
rect 2240 336410 2268 339646
rect 2056 336382 2268 336410
rect 1952 334212 2004 334218
rect 1952 334154 2004 334160
rect 1952 334076 2004 334082
rect 2056 334064 2084 336382
rect 2884 334064 2912 345494
rect 2976 344978 3004 349982
rect 3068 345386 3096 352158
rect 3344 346202 3372 361270
rect 3712 354498 3740 414174
rect 3528 354470 3740 354498
rect 3528 347426 3556 354470
rect 3528 347398 3740 347426
rect 3344 346174 3648 346202
rect 3068 345358 3464 345386
rect 3436 345250 3464 345358
rect 3620 345250 3648 346174
rect 3344 345222 3648 345250
rect 2976 344950 3096 344978
rect 2004 334036 2084 334064
rect 2148 334036 2912 334064
rect 3068 334064 3096 344950
rect 3344 344570 3372 345222
rect 3436 345114 3464 345222
rect 3436 345086 3648 345114
rect 3252 344542 3372 344570
rect 3252 344298 3280 344542
rect 3252 344270 3372 344298
rect 3146 339688 3202 339697
rect 3344 339674 3372 344270
rect 3202 339646 3372 339674
rect 3146 339623 3202 339632
rect 3620 334064 3648 345086
rect 3068 334036 3188 334064
rect 1952 334018 2004 334024
rect 2148 333826 2176 334036
rect 1872 333798 2176 333826
rect 1872 333554 1900 333798
rect 1952 333736 2004 333742
rect 2004 333684 2912 333690
rect 1952 333678 2912 333684
rect 1964 333662 2912 333678
rect 2884 333656 2912 333662
rect 2884 333628 3004 333656
rect 1872 333526 2912 333554
rect 1952 333464 2004 333470
rect 1780 333390 1900 333418
rect 1952 333406 2004 333412
rect 1768 331560 1820 331566
rect 1768 331502 1820 331508
rect 1780 260778 1808 331502
rect 1872 261526 1900 333390
rect 1964 332058 1992 333406
rect 1964 332030 2820 332058
rect 1952 331832 2004 331838
rect 2004 331780 2636 331786
rect 1952 331774 2636 331780
rect 1964 331758 2636 331774
rect 1952 329792 2004 329798
rect 2004 329740 2268 329746
rect 1952 329734 2268 329740
rect 1964 329718 2268 329734
rect 1952 329180 2004 329186
rect 1952 329122 2004 329128
rect 1964 319190 1992 329122
rect 2240 325394 2268 329718
rect 2056 325366 2268 325394
rect 1952 319184 2004 319190
rect 1952 319126 2004 319132
rect 1952 318980 2004 318986
rect 2056 318968 2084 325366
rect 2608 324986 2636 331758
rect 2004 318940 2084 318968
rect 2148 324958 2636 324986
rect 1952 318922 2004 318928
rect 2148 318866 2176 324958
rect 2792 324850 2820 332030
rect 2516 324822 2820 324850
rect 2516 321042 2544 324822
rect 2884 324714 2912 333526
rect 2608 324686 2912 324714
rect 2608 321178 2636 324686
rect 2608 321150 2820 321178
rect 2516 321014 2636 321042
rect 1964 318838 2176 318866
rect 1964 315178 1992 318838
rect 2608 317914 2636 321014
rect 2792 318050 2820 321150
rect 2976 318458 3004 333628
rect 3160 327434 3188 334036
rect 3528 334036 3648 334064
rect 3160 327406 3280 327434
rect 3252 327162 3280 327406
rect 3068 327134 3280 327162
rect 3068 321178 3096 327134
rect 3528 322130 3556 334036
rect 3436 322102 3556 322130
rect 3068 321150 3280 321178
rect 3146 321056 3202 321065
rect 3146 320991 3202 321000
rect 2976 318430 3096 318458
rect 3068 318050 3096 318430
rect 2792 318022 2912 318050
rect 2056 317886 2636 317914
rect 1952 315172 2004 315178
rect 1952 315114 2004 315120
rect 1952 315036 2004 315042
rect 1952 314978 2004 314984
rect 1964 312594 1992 314978
rect 1952 312588 2004 312594
rect 1952 312530 2004 312536
rect 1952 312452 2004 312458
rect 2056 312440 2084 317886
rect 2884 317778 2912 318022
rect 2608 317750 2912 317778
rect 2976 318022 3096 318050
rect 2608 317642 2636 317750
rect 2004 312412 2084 312440
rect 2424 317614 2636 317642
rect 1952 312394 2004 312400
rect 2424 312338 2452 317614
rect 2976 317234 3004 318022
rect 2792 317206 3004 317234
rect 2792 314106 2820 317206
rect 1964 312322 2452 312338
rect 1952 312316 2452 312322
rect 2004 312310 2452 312316
rect 2608 314078 2820 314106
rect 1952 312258 2004 312264
rect 2608 312202 2636 314078
rect 3160 313834 3188 320991
rect 1964 312186 2636 312202
rect 1952 312180 2636 312186
rect 2004 312174 2636 312180
rect 2976 313806 3188 313834
rect 1952 312122 2004 312128
rect 2976 312066 3004 313806
rect 1964 312050 2452 312066
rect 1952 312044 2452 312050
rect 2004 312038 2452 312044
rect 1952 311986 2004 311992
rect 1952 311840 2004 311846
rect 2004 311788 2360 311794
rect 1952 311782 2360 311788
rect 1964 311766 2360 311782
rect 1952 311704 2004 311710
rect 2004 311652 2268 311658
rect 1952 311646 2268 311652
rect 1964 311630 2268 311646
rect 1952 311568 2004 311574
rect 2004 311516 2176 311522
rect 1952 311510 2176 311516
rect 1964 311494 2176 311510
rect 1952 309868 2004 309874
rect 1952 309810 2004 309816
rect 1964 309754 1992 309810
rect 1964 309726 2084 309754
rect 1952 309664 2004 309670
rect 1952 309606 2004 309612
rect 1964 306678 1992 309606
rect 1952 306672 2004 306678
rect 1952 306614 2004 306620
rect 1952 305652 2004 305658
rect 2056 305640 2084 309726
rect 2004 305612 2084 305640
rect 1952 305594 2004 305600
rect 1952 305516 2004 305522
rect 2148 305504 2176 311494
rect 2004 305476 2176 305504
rect 1952 305458 2004 305464
rect 2240 305402 2268 311630
rect 1964 305386 2268 305402
rect 1952 305380 2268 305386
rect 2004 305374 2268 305380
rect 1952 305322 2004 305328
rect 2332 304586 2360 311766
rect 1964 304570 2360 304586
rect 1952 304564 2360 304570
rect 2004 304558 2360 304564
rect 1952 304506 2004 304512
rect 2424 304450 2452 312038
rect 2608 312038 3004 312066
rect 2608 310434 2636 312038
rect 3252 310570 3280 321150
rect 3436 320498 3464 322102
rect 3344 320470 3464 320498
rect 3344 314786 3372 320470
rect 3712 320362 3740 347398
rect 3436 320334 3740 320362
rect 3436 320090 3464 320334
rect 3436 320062 3740 320090
rect 3712 315058 3740 320062
rect 3436 315030 3740 315058
rect 3436 314786 3464 315030
rect 3344 314758 3556 314786
rect 3252 310542 3372 310570
rect 3344 310434 3372 310542
rect 2608 310406 2820 310434
rect 1964 304434 2452 304450
rect 1952 304428 2452 304434
rect 2004 304422 2452 304428
rect 1952 304370 2004 304376
rect 1964 304286 2360 304314
rect 1964 304162 1992 304286
rect 1952 304156 2004 304162
rect 1952 304098 2004 304104
rect 1952 304020 2004 304026
rect 1952 303962 2004 303968
rect 1964 303906 1992 303962
rect 1964 303878 2268 303906
rect 1952 303408 2004 303414
rect 2240 303362 2268 303878
rect 2004 303356 2268 303362
rect 1952 303350 2268 303356
rect 1964 303334 2268 303350
rect 1952 303272 2004 303278
rect 1952 303214 2004 303220
rect 1964 302138 1992 303214
rect 1964 302110 2176 302138
rect 1952 301504 2004 301510
rect 1952 301446 2004 301452
rect 1964 296138 1992 301446
rect 1952 296132 2004 296138
rect 1952 296074 2004 296080
rect 2148 295882 2176 302110
rect 1964 295866 2176 295882
rect 1952 295860 2176 295866
rect 2004 295854 2176 295860
rect 1952 295802 2004 295808
rect 2332 295746 2360 304286
rect 1964 295718 2360 295746
rect 1964 293418 1992 295718
rect 2792 295474 2820 310406
rect 2976 310406 3372 310434
rect 2976 305130 3004 310406
rect 3436 305810 3464 314758
rect 3252 305782 3464 305810
rect 2976 305102 3188 305130
rect 3160 298738 3188 305102
rect 3252 301832 3280 305782
rect 3332 301844 3384 301850
rect 3252 301804 3332 301832
rect 3332 301786 3384 301792
rect 3528 301730 3556 314758
rect 3804 302682 3832 449806
rect 568316 418418 568344 481494
rect 568684 466426 568712 485710
rect 569052 480978 569080 498902
rect 569236 490634 569264 514542
rect 569144 490606 569264 490634
rect 569144 485738 569172 490606
rect 569144 485710 569264 485738
rect 569236 485602 569264 485710
rect 569236 485574 569356 485602
rect 569052 480950 569172 480978
rect 569144 474722 569172 480950
rect 568592 466398 568712 466426
rect 569052 474694 569172 474722
rect 568592 455410 568620 466398
rect 569052 464930 569080 474694
rect 569328 465032 569356 485574
rect 569420 465236 569448 551670
rect 570064 551426 570092 551942
rect 572732 551886 572760 558583
rect 572720 551880 572772 551886
rect 572720 551822 572772 551828
rect 569788 551398 570092 551426
rect 569788 531026 569816 551398
rect 569960 551064 570012 551070
rect 569880 551012 569960 551018
rect 569880 551006 570012 551012
rect 569880 550990 570000 551006
rect 569880 533338 569908 550990
rect 580170 533896 580226 533905
rect 580170 533831 580226 533840
rect 569880 533310 570000 533338
rect 569972 531146 570000 533310
rect 580184 532778 580212 533831
rect 573364 532772 573416 532778
rect 573364 532714 573416 532720
rect 580172 532772 580224 532778
rect 580172 532714 580224 532720
rect 569960 531140 570012 531146
rect 569960 531082 570012 531088
rect 569788 531010 570000 531026
rect 569788 531004 570012 531010
rect 569788 530998 569960 531004
rect 569960 530946 570012 530952
rect 570326 530904 570382 530913
rect 570064 530862 570326 530890
rect 570064 530040 570092 530862
rect 570326 530839 570382 530848
rect 569604 530012 570092 530040
rect 569604 524498 569632 530012
rect 569960 528896 570012 528902
rect 569788 528844 569960 528850
rect 569788 528838 570012 528844
rect 569788 528822 570000 528838
rect 569604 524470 569724 524498
rect 569696 523682 569724 524470
rect 569512 523654 569724 523682
rect 569512 466868 569540 523654
rect 569788 522730 569816 528822
rect 569960 528760 570012 528766
rect 569880 528708 569960 528714
rect 569880 528702 570012 528708
rect 569880 528686 570000 528702
rect 569880 527082 569908 528686
rect 569880 527054 570000 527082
rect 569696 522702 569816 522730
rect 569696 522458 569724 522702
rect 569972 522646 570000 527054
rect 569960 522640 570012 522646
rect 569960 522582 570012 522588
rect 569960 522504 570012 522510
rect 569696 522452 569960 522458
rect 569696 522446 570012 522452
rect 569696 522430 570000 522446
rect 573376 522374 573404 532714
rect 569960 522368 570012 522374
rect 569604 522316 569960 522322
rect 569604 522310 570012 522316
rect 573364 522368 573416 522374
rect 573364 522310 573416 522316
rect 569604 522294 570000 522310
rect 569604 468058 569632 522294
rect 569960 521076 570012 521082
rect 569960 521018 570012 521024
rect 569972 520962 570000 521018
rect 569788 520934 570000 520962
rect 569788 504234 569816 520934
rect 569960 518492 570012 518498
rect 569960 518434 570012 518440
rect 569972 517426 570000 518434
rect 569880 517398 570000 517426
rect 569880 507770 569908 517398
rect 569880 507742 570000 507770
rect 569972 505170 570000 507742
rect 569960 505164 570012 505170
rect 569960 505106 570012 505112
rect 569788 504218 570000 504234
rect 569788 504212 570012 504218
rect 569788 504206 569960 504212
rect 569960 504154 570012 504160
rect 570326 503704 570382 503713
rect 569696 503662 570326 503690
rect 569696 468330 569724 503662
rect 570326 503639 570382 503648
rect 569960 503192 570012 503198
rect 569788 503140 569960 503146
rect 569788 503134 570012 503140
rect 569788 503118 570000 503134
rect 569788 491042 569816 503118
rect 569960 503056 570012 503062
rect 569880 503004 569960 503010
rect 569880 502998 570012 503004
rect 569880 502982 570000 502998
rect 569880 491314 569908 502982
rect 569880 491286 570184 491314
rect 569788 491014 570000 491042
rect 569972 487150 570000 491014
rect 569960 487144 570012 487150
rect 569960 487086 570012 487092
rect 570156 487014 570184 491286
rect 579804 487144 579856 487150
rect 579804 487086 579856 487092
rect 569960 487008 570012 487014
rect 569788 486956 569960 486962
rect 569788 486950 570012 486956
rect 570144 487008 570196 487014
rect 570144 486950 570196 486956
rect 569788 486934 570000 486950
rect 569788 468602 569816 486934
rect 579816 486849 579844 487086
rect 579802 486840 579858 486849
rect 579802 486775 579858 486784
rect 570326 476504 570382 476513
rect 570064 476462 570326 476490
rect 569788 468586 570000 468602
rect 569788 468580 570012 468586
rect 569788 468574 569960 468580
rect 569960 468522 570012 468528
rect 569696 468314 570000 468330
rect 569696 468308 570012 468314
rect 569696 468302 569960 468308
rect 569960 468250 570012 468256
rect 569604 468030 570000 468058
rect 569972 467634 570000 468030
rect 569960 467628 570012 467634
rect 569960 467570 570012 467576
rect 570064 467090 570092 476462
rect 570326 476439 570382 476448
rect 570052 467084 570104 467090
rect 570052 467026 570104 467032
rect 569972 466942 570184 466970
rect 569972 466868 570000 466942
rect 569512 466840 570000 466868
rect 570052 466880 570104 466886
rect 570052 466822 570104 466828
rect 570064 465390 570092 466822
rect 570052 465384 570104 465390
rect 570052 465326 570104 465332
rect 570156 465254 570184 466942
rect 569960 465248 570012 465254
rect 569420 465208 569960 465236
rect 569960 465190 570012 465196
rect 570144 465248 570196 465254
rect 570144 465190 570196 465196
rect 570144 465112 570196 465118
rect 570144 465054 570196 465060
rect 569328 465004 570092 465032
rect 569052 464902 570000 464930
rect 569868 464296 569920 464302
rect 569868 464238 569920 464244
rect 569880 463978 569908 464238
rect 569972 464030 570000 464902
rect 570064 464166 570092 465004
rect 570052 464160 570104 464166
rect 570052 464102 570104 464108
rect 568776 463950 569908 463978
rect 569960 464024 570012 464030
rect 569960 463966 570012 463972
rect 568592 455382 568712 455410
rect 568684 452010 568712 455382
rect 568592 451982 568712 452010
rect 568592 449018 568620 451982
rect 568776 451058 568804 463950
rect 569960 463888 570012 463894
rect 568960 463836 569960 463842
rect 568960 463830 570012 463836
rect 568960 463814 570000 463830
rect 568960 455410 568988 463814
rect 569960 463752 570012 463758
rect 569328 463700 569960 463706
rect 569328 463694 570012 463700
rect 569328 463678 570000 463694
rect 568960 455382 569264 455410
rect 568684 451030 568804 451058
rect 568684 449698 568712 451030
rect 568684 449670 569172 449698
rect 569144 449426 569172 449670
rect 569236 449426 569264 455382
rect 569052 449398 569264 449426
rect 568592 448990 568896 449018
rect 568868 443306 568896 448990
rect 568408 443278 568896 443306
rect 568408 434058 568436 443278
rect 569052 442762 569080 449398
rect 568592 442734 569080 442762
rect 568408 434030 568528 434058
rect 568500 419506 568528 434030
rect 568592 420730 568620 442734
rect 569144 442490 569172 449398
rect 569328 442490 569356 463678
rect 569960 463616 570012 463622
rect 569960 463558 570012 463564
rect 569972 463026 570000 463558
rect 570156 463026 570184 465054
rect 568684 442462 569356 442490
rect 569420 462998 570000 463026
rect 570064 462998 570184 463026
rect 568684 440858 568712 442462
rect 569144 442354 569172 442462
rect 569144 442326 569264 442354
rect 569236 442082 569264 442326
rect 569236 442054 569356 442082
rect 568684 440830 568896 440858
rect 568868 434058 568896 440830
rect 568868 434030 569172 434058
rect 569144 422226 569172 434030
rect 568868 422198 569172 422226
rect 568868 421954 568896 422198
rect 568868 421926 568988 421954
rect 568960 421682 568988 421926
rect 568868 421654 568988 421682
rect 568868 421138 568896 421654
rect 568776 421110 568896 421138
rect 568776 420866 568804 421110
rect 568776 420838 568896 420866
rect 568868 420730 568896 420838
rect 568592 420702 569172 420730
rect 568868 420594 568896 420702
rect 568868 420566 568988 420594
rect 568500 419478 568896 419506
rect 568316 418390 568436 418418
rect 568408 418180 568436 418390
rect 568316 418152 568436 418180
rect 568316 411346 568344 418152
rect 568224 411318 568344 411346
rect 568224 399548 568252 411318
rect 568868 406858 568896 419478
rect 568592 406830 568896 406858
rect 568592 406586 568620 406830
rect 568408 406558 568620 406586
rect 568408 405634 568436 406558
rect 568960 405906 568988 420566
rect 569144 413386 569172 420702
rect 568684 405878 568988 405906
rect 569052 413358 569172 413386
rect 568408 405606 568528 405634
rect 568500 400738 568528 405606
rect 568684 400874 568712 405878
rect 569052 405498 569080 413358
rect 569052 405470 569264 405498
rect 568684 400846 568896 400874
rect 568500 400710 568804 400738
rect 568224 399520 568436 399548
rect 568408 394074 568436 399520
rect 568316 394046 568436 394074
rect 568316 390402 568344 394046
rect 568776 393938 568804 400710
rect 568224 390374 568344 390402
rect 568408 393910 568804 393938
rect 568224 374490 568252 390374
rect 568408 389076 568436 393910
rect 568868 393836 568896 400846
rect 568684 393808 568896 393836
rect 568684 392850 568712 393808
rect 569236 393122 569264 405470
rect 569328 393666 569356 442054
rect 569420 393836 569448 462998
rect 570064 462890 570092 462998
rect 569512 462862 570092 462890
rect 569512 394890 569540 462862
rect 570052 462800 570104 462806
rect 570052 462742 570104 462748
rect 569960 461712 570012 461718
rect 569696 461672 569960 461700
rect 569696 457586 569724 461672
rect 569960 461654 570012 461660
rect 570064 461530 570092 462742
rect 569604 457558 569724 457586
rect 569880 461502 570092 461530
rect 569604 399378 569632 457558
rect 569880 457450 569908 461502
rect 569960 461440 570012 461446
rect 569960 461382 570012 461388
rect 569696 457422 569908 457450
rect 569696 399514 569724 457422
rect 569972 449410 570000 461382
rect 569960 449404 570012 449410
rect 569960 449346 570012 449352
rect 570326 449304 570382 449313
rect 569788 449262 570326 449290
rect 569788 439498 569816 449262
rect 570326 449239 570382 449248
rect 569960 449200 570012 449206
rect 569960 449142 570012 449148
rect 569972 447930 570000 449142
rect 569880 447902 570000 447930
rect 569880 441674 569908 447902
rect 569880 441658 570000 441674
rect 569880 441652 570012 441658
rect 569880 441646 569960 441652
rect 569960 441594 570012 441600
rect 580170 439920 580226 439929
rect 580170 439855 580226 439864
rect 569788 439470 569908 439498
rect 569880 432562 569908 439470
rect 580184 438938 580212 439855
rect 574744 438932 574796 438938
rect 574744 438874 574796 438880
rect 580172 438932 580224 438938
rect 580172 438874 580224 438880
rect 570052 436824 570104 436830
rect 570052 436766 570104 436772
rect 569880 432546 570000 432562
rect 569880 432540 570012 432546
rect 569880 432534 569960 432540
rect 569960 432482 570012 432488
rect 570064 428754 570092 436766
rect 569880 428726 570092 428754
rect 569880 428482 569908 428726
rect 569788 428454 569908 428482
rect 569788 418418 569816 428454
rect 572718 422648 572774 422657
rect 572718 422583 572774 422592
rect 569788 418390 570000 418418
rect 569972 418334 570000 418390
rect 569960 418328 570012 418334
rect 569960 418270 570012 418276
rect 569960 418192 570012 418198
rect 569960 418134 570012 418140
rect 569972 407114 570000 418134
rect 572732 412010 572760 422583
rect 570604 412004 570656 412010
rect 570604 411946 570656 411952
rect 572720 412004 572772 412010
rect 572720 411946 572772 411952
rect 569960 407108 570012 407114
rect 569960 407050 570012 407056
rect 570052 407108 570104 407114
rect 570052 407050 570104 407056
rect 569960 402280 570012 402286
rect 569880 402228 569960 402234
rect 569880 402222 570012 402228
rect 569880 402206 570000 402222
rect 569696 399486 569816 399514
rect 569604 399350 569724 399378
rect 569696 394992 569724 399350
rect 569788 396386 569816 399486
rect 569880 396658 569908 402206
rect 569960 401668 570012 401674
rect 569960 401610 570012 401616
rect 569972 396846 570000 401610
rect 570064 399566 570092 407050
rect 570616 401674 570644 411946
rect 570604 401668 570656 401674
rect 570604 401610 570656 401616
rect 570052 399560 570104 399566
rect 570052 399502 570104 399508
rect 569960 396840 570012 396846
rect 569960 396782 570012 396788
rect 569880 396630 570092 396658
rect 570064 396488 570092 396630
rect 570064 396460 570184 396488
rect 569788 396358 570092 396386
rect 569960 395004 570012 395010
rect 569696 394964 569960 394992
rect 569960 394946 570012 394952
rect 569512 394862 570000 394890
rect 569972 393854 570000 394862
rect 570064 394670 570092 396358
rect 570052 394664 570104 394670
rect 570052 394606 570104 394612
rect 569960 393848 570012 393854
rect 569420 393808 569908 393836
rect 569880 393700 569908 393808
rect 569960 393790 570012 393796
rect 569960 393712 570012 393718
rect 569880 393672 569960 393700
rect 569328 393638 569816 393666
rect 569960 393654 570012 393660
rect 569788 393258 569816 393638
rect 569788 393230 570000 393258
rect 569972 393174 570000 393230
rect 569960 393168 570012 393174
rect 569236 393094 569908 393122
rect 569960 393110 570012 393116
rect 569880 392986 569908 393094
rect 569880 392970 570000 392986
rect 569880 392964 570012 392970
rect 569880 392958 569960 392964
rect 569960 392906 570012 392912
rect 568684 392822 570092 392850
rect 569960 392760 570012 392766
rect 568592 392720 569960 392748
rect 568592 389076 568620 392720
rect 569960 392702 570012 392708
rect 569960 392624 570012 392630
rect 569960 392566 570012 392572
rect 569972 392442 570000 392566
rect 569144 392414 570000 392442
rect 569144 389858 569172 392414
rect 569960 392352 570012 392358
rect 569420 392312 569960 392340
rect 569420 392306 569448 392312
rect 568776 389830 569172 389858
rect 569236 392278 569448 392306
rect 569960 392294 570012 392300
rect 568408 389048 568528 389076
rect 568592 389048 568712 389076
rect 568500 388770 568528 389048
rect 568500 388742 568620 388770
rect 568592 374626 568620 388742
rect 568684 376666 568712 389048
rect 568776 377210 568804 389830
rect 569236 389722 569264 392278
rect 570064 392170 570092 392822
rect 569052 389694 569264 389722
rect 569512 392142 570092 392170
rect 569052 381154 569080 389694
rect 569512 389586 569540 392142
rect 569960 390040 570012 390046
rect 568960 381126 569080 381154
rect 569236 389558 569540 389586
rect 569604 389988 569960 389994
rect 569604 389982 570012 389988
rect 569604 389966 570000 389982
rect 568960 380882 568988 381126
rect 568960 380854 569080 380882
rect 568776 377182 568988 377210
rect 568684 376638 568896 376666
rect 568316 374598 568620 374626
rect 568316 374490 568344 374598
rect 568224 374462 568804 374490
rect 568316 374082 568344 374462
rect 568224 374054 568344 374082
rect 568224 362930 568252 374054
rect 568776 373130 568804 374462
rect 568316 373102 568804 373130
rect 568316 371498 568344 373102
rect 568316 371470 568528 371498
rect 568500 364154 568528 371470
rect 568500 364126 568620 364154
rect 568592 363202 568620 364126
rect 568868 363882 568896 376638
rect 568960 364018 568988 377182
rect 569052 367554 569080 380854
rect 569236 378162 569264 389558
rect 569604 389314 569632 389966
rect 569960 389904 570012 389910
rect 569960 389846 570012 389852
rect 569144 378134 569264 378162
rect 569328 389286 569632 389314
rect 569144 367690 569172 378134
rect 569328 378026 569356 389286
rect 569972 389178 570000 389846
rect 569236 377998 569356 378026
rect 569420 389150 570000 389178
rect 569420 378026 569448 389150
rect 569960 389088 570012 389094
rect 569512 389036 569960 389042
rect 569512 389030 570012 389036
rect 569512 389014 570000 389030
rect 569512 378298 569540 389014
rect 569960 388544 570012 388550
rect 569604 388492 569960 388498
rect 569604 388486 570012 388492
rect 569604 388470 570000 388486
rect 569604 378434 569632 388470
rect 569960 388408 570012 388414
rect 569788 388356 569960 388362
rect 569788 388350 570012 388356
rect 569788 388334 570000 388350
rect 569788 382922 569816 388334
rect 569788 382894 570000 382922
rect 569972 382838 570000 382894
rect 569960 382832 570012 382838
rect 569960 382774 570012 382780
rect 569960 382696 570012 382702
rect 569788 382644 569960 382650
rect 569788 382638 570012 382644
rect 569788 382622 570000 382638
rect 569788 382242 569816 382622
rect 569788 382214 570000 382242
rect 569972 381886 570000 382214
rect 569960 381880 570012 381886
rect 569960 381822 570012 381828
rect 569604 378406 569908 378434
rect 569512 378270 569816 378298
rect 569420 377998 569540 378026
rect 569236 367962 569264 377998
rect 569512 377346 569540 377998
rect 569420 377318 569540 377346
rect 569420 368064 569448 377318
rect 569788 377210 569816 378270
rect 569512 377182 569816 377210
rect 569512 368336 569540 377182
rect 569880 377074 569908 378406
rect 569604 377046 569908 377074
rect 569604 369458 569632 377046
rect 570156 376718 570184 396460
rect 570326 394904 570382 394913
rect 570326 394839 570382 394848
rect 570236 394664 570288 394670
rect 570236 394606 570288 394612
rect 570248 388414 570276 394606
rect 570340 392630 570368 394839
rect 570328 392624 570380 392630
rect 570328 392566 570380 392572
rect 570236 388408 570288 388414
rect 570236 388350 570288 388356
rect 569960 376712 570012 376718
rect 569788 376672 569960 376700
rect 569788 376394 569816 376672
rect 569960 376654 570012 376660
rect 570144 376712 570196 376718
rect 570144 376654 570196 376660
rect 569960 376576 570012 376582
rect 569960 376518 570012 376524
rect 569696 376366 569816 376394
rect 569696 369594 569724 376366
rect 569972 369782 570000 376518
rect 569960 369776 570012 369782
rect 569960 369718 570012 369724
rect 569696 369566 570092 369594
rect 569604 369442 570000 369458
rect 569604 369436 570012 369442
rect 569604 369430 569960 369436
rect 569960 369378 570012 369384
rect 569960 368348 570012 368354
rect 569512 368308 569960 368336
rect 569960 368290 570012 368296
rect 569960 368076 570012 368082
rect 569420 368036 569960 368064
rect 569960 368018 570012 368024
rect 569236 367934 569448 367962
rect 569420 367792 569448 367934
rect 569960 367804 570012 367810
rect 569420 367764 569960 367792
rect 569960 367746 570012 367752
rect 569144 367662 570000 367690
rect 569052 367526 569632 367554
rect 568960 363990 569448 364018
rect 568868 363854 568988 363882
rect 568960 363610 568988 363854
rect 568960 363582 569356 363610
rect 568592 363174 568804 363202
rect 568776 362930 568804 363174
rect 568224 362902 569080 362930
rect 568776 362794 568804 362902
rect 568592 362766 568804 362794
rect 568592 358714 568620 362766
rect 569052 358884 569080 362902
rect 569328 362794 569356 363582
rect 569144 362766 569356 362794
rect 569144 359156 569172 362766
rect 569420 359564 569448 363990
rect 569604 359904 569632 367526
rect 569972 360058 570000 367662
rect 570064 362370 570092 369566
rect 570144 368076 570196 368082
rect 570144 368018 570196 368024
rect 570052 362364 570104 362370
rect 570052 362306 570104 362312
rect 570156 362250 570184 368018
rect 570326 367704 570382 367713
rect 570326 367639 570382 367648
rect 570236 362364 570288 362370
rect 570236 362306 570288 362312
rect 570064 362222 570184 362250
rect 569960 360052 570012 360058
rect 569960 359994 570012 360000
rect 569960 359916 570012 359922
rect 569604 359876 569960 359904
rect 569960 359858 570012 359864
rect 569960 359576 570012 359582
rect 569420 359536 569960 359564
rect 569960 359518 570012 359524
rect 569960 359168 570012 359174
rect 569144 359128 569960 359156
rect 569960 359110 570012 359116
rect 569960 358896 570012 358902
rect 569052 358856 569960 358884
rect 569960 358838 570012 358844
rect 569960 358760 570012 358766
rect 568224 358686 568620 358714
rect 568684 358720 569960 358748
rect 568224 339130 568252 358686
rect 568408 358550 568620 358578
rect 568408 358442 568436 358550
rect 568316 358414 568436 358442
rect 568592 358442 568620 358550
rect 568684 358442 568712 358720
rect 569960 358702 570012 358708
rect 569960 358624 570012 358630
rect 568592 358414 568712 358442
rect 569880 358584 569960 358612
rect 568316 339402 568344 358414
rect 569880 358272 569908 358584
rect 569960 358566 570012 358572
rect 568592 358244 569908 358272
rect 569960 358284 570012 358290
rect 568592 343754 568620 358244
rect 569960 358226 570012 358232
rect 569972 358136 570000 358226
rect 570064 358154 570092 362222
rect 570248 362114 570276 362306
rect 570156 362086 570276 362114
rect 570156 358154 570184 362086
rect 570340 360176 570368 367639
rect 570248 360148 570368 360176
rect 570248 358766 570276 360148
rect 570328 360052 570380 360058
rect 570328 359994 570380 360000
rect 570236 358760 570288 358766
rect 570236 358702 570288 358708
rect 568868 358108 570000 358136
rect 570052 358148 570104 358154
rect 568868 356946 568896 358108
rect 570052 358090 570104 358096
rect 570144 358148 570196 358154
rect 570144 358090 570196 358096
rect 570236 358080 570288 358086
rect 568684 356918 568896 356946
rect 569236 358028 570236 358034
rect 569236 358022 570288 358028
rect 569236 358006 570276 358022
rect 568684 344026 568712 356918
rect 569236 356674 569264 358006
rect 570052 357944 570104 357950
rect 570052 357886 570104 357892
rect 570144 357944 570196 357950
rect 570144 357886 570196 357892
rect 569960 357876 570012 357882
rect 569960 357818 570012 357824
rect 568960 356646 569264 356674
rect 568960 349602 568988 356646
rect 568868 349574 568988 349602
rect 569052 354334 569632 354362
rect 568868 344842 568896 349574
rect 569052 349466 569080 354334
rect 569604 353784 569632 354334
rect 569972 354006 570000 357818
rect 569960 354000 570012 354006
rect 569960 353942 570012 353948
rect 569960 353796 570012 353802
rect 569604 353756 569960 353784
rect 569960 353738 570012 353744
rect 569960 353660 570012 353666
rect 569960 353602 570012 353608
rect 569868 353252 569920 353258
rect 569868 353194 569920 353200
rect 568960 349438 569080 349466
rect 568960 344842 568988 349438
rect 569880 349194 569908 353194
rect 569972 352458 570000 353602
rect 570064 352646 570092 357886
rect 570052 352640 570104 352646
rect 570052 352582 570104 352588
rect 569972 352430 570092 352458
rect 569960 352368 570012 352374
rect 569960 352310 570012 352316
rect 568776 344814 568988 344842
rect 569236 349166 569908 349194
rect 568776 344162 568804 344814
rect 568868 344298 568896 344814
rect 568868 344270 569080 344298
rect 568776 344134 568896 344162
rect 568684 343998 568804 344026
rect 568592 343726 568712 343754
rect 568316 339374 568620 339402
rect 568224 339102 568528 339130
rect 568500 337498 568528 339102
rect 568316 337470 568528 337498
rect 568316 337362 568344 337470
rect 568592 337362 568620 339374
rect 568224 337334 568620 337362
rect 568224 315568 568252 337334
rect 568316 320226 568344 337334
rect 568684 332738 568712 343726
rect 568592 332710 568712 332738
rect 568592 332602 568620 332710
rect 568776 332602 568804 343998
rect 568500 332574 568620 332602
rect 568684 332574 568804 332602
rect 568500 327808 568528 332574
rect 568684 327978 568712 332574
rect 568868 328930 568896 344134
rect 569052 337634 569080 344270
rect 569236 339674 569264 349166
rect 569972 349058 570000 352310
rect 569420 349030 570000 349058
rect 569420 348378 569448 349030
rect 569960 348968 570012 348974
rect 569328 348350 569448 348378
rect 569604 348928 569960 348956
rect 569328 339810 569356 348350
rect 569604 348242 569632 348928
rect 569960 348910 570012 348916
rect 569420 348214 569632 348242
rect 569420 339946 569448 348214
rect 570064 348140 570092 352430
rect 569512 348112 570092 348140
rect 569512 340082 569540 348112
rect 569960 348016 570012 348022
rect 569604 347976 569960 348004
rect 569604 340218 569632 347976
rect 569960 347958 570012 347964
rect 570156 347868 570184 357886
rect 570340 353326 570368 359994
rect 570328 353320 570380 353326
rect 570328 353262 570380 353268
rect 569696 347840 570184 347868
rect 569696 340320 569724 347840
rect 569960 347744 570012 347750
rect 569880 347704 569960 347732
rect 569880 340490 569908 347704
rect 569960 347686 570012 347692
rect 569960 344888 570012 344894
rect 569960 344830 570012 344836
rect 569972 342242 570000 344830
rect 569960 342236 570012 342242
rect 569960 342178 570012 342184
rect 572718 341048 572774 341057
rect 572718 340983 572774 340992
rect 569880 340462 570000 340490
rect 569696 340292 569908 340320
rect 569604 340190 569816 340218
rect 569512 340054 569724 340082
rect 569420 339918 569632 339946
rect 569328 339782 569540 339810
rect 569236 339646 569448 339674
rect 569420 337634 569448 339646
rect 568960 337606 569080 337634
rect 569144 337606 569448 337634
rect 568960 329338 568988 337606
rect 568960 329310 569080 329338
rect 569052 329066 569080 329310
rect 569144 329202 569172 337606
rect 569512 337362 569540 339782
rect 569328 337334 569540 337362
rect 569328 329610 569356 337334
rect 569604 337226 569632 339918
rect 569420 337198 569632 337226
rect 569420 330018 569448 337198
rect 569696 337090 569724 340054
rect 569512 337062 569724 337090
rect 569512 330290 569540 337062
rect 569788 336002 569816 340190
rect 569604 335974 569816 336002
rect 569604 330426 569632 335974
rect 569880 335866 569908 340292
rect 569696 335838 569908 335866
rect 569696 330698 569724 335838
rect 569972 333282 570000 340462
rect 569788 333254 570000 333282
rect 569788 330970 569816 333254
rect 569960 331288 570012 331294
rect 569880 331236 569960 331242
rect 569880 331230 570012 331236
rect 569880 331214 570000 331230
rect 569880 331106 569908 331214
rect 569880 331090 570000 331106
rect 569880 331084 570012 331090
rect 569880 331078 569960 331084
rect 569960 331026 570012 331032
rect 569788 330942 570276 330970
rect 569696 330670 570000 330698
rect 569972 330546 570000 330670
rect 569960 330540 570012 330546
rect 569960 330482 570012 330488
rect 569604 330398 570184 330426
rect 569512 330262 570092 330290
rect 569420 329990 570000 330018
rect 569972 329730 570000 329990
rect 569960 329724 570012 329730
rect 569960 329666 570012 329672
rect 569328 329594 570000 329610
rect 569328 329588 570012 329594
rect 569328 329582 569960 329588
rect 569960 329530 570012 329536
rect 569420 329458 570000 329474
rect 569420 329452 570012 329458
rect 569420 329446 569960 329452
rect 569420 329202 569448 329446
rect 569960 329394 570012 329400
rect 569144 329174 569448 329202
rect 569512 329322 570000 329338
rect 569512 329316 570012 329322
rect 569512 329310 569960 329316
rect 569512 329066 569540 329310
rect 569960 329258 570012 329264
rect 569052 329038 569540 329066
rect 568868 328902 569080 328930
rect 568684 327950 568896 327978
rect 568408 327780 568528 327808
rect 568408 324442 568436 327780
rect 568408 324414 568620 324442
rect 568316 320198 568436 320226
rect 568408 315840 568436 320198
rect 568592 317948 568620 324414
rect 568868 324170 568896 327950
rect 569052 327808 569080 328902
rect 569960 327820 570012 327826
rect 569052 327780 569960 327808
rect 569960 327762 570012 327768
rect 569236 327678 569632 327706
rect 568868 324142 568988 324170
rect 568960 322946 568988 324142
rect 569236 322946 569264 327678
rect 569604 327672 569632 327678
rect 569960 327684 570012 327690
rect 569604 327644 569960 327672
rect 569960 327626 570012 327632
rect 569960 327208 570012 327214
rect 568684 322918 568988 322946
rect 569052 322918 569264 322946
rect 569512 327168 569960 327196
rect 568684 320090 568712 322918
rect 569052 321586 569080 322918
rect 569052 321558 569264 321586
rect 568684 320062 569172 320090
rect 568592 317920 568804 317948
rect 568408 315812 568712 315840
rect 568224 315540 568344 315568
rect 568316 315500 568344 315540
rect 568224 315472 568344 315500
rect 568224 315194 568252 315472
rect 568224 315166 568344 315194
rect 568316 314786 568344 315166
rect 568684 314786 568712 315812
rect 2240 295446 2820 295474
rect 2976 298710 3188 298738
rect 3344 301702 3556 301730
rect 3620 302654 3832 302682
rect 568224 314758 568712 314786
rect 568776 314786 568804 317920
rect 569144 315194 569172 320062
rect 569236 315500 569264 321558
rect 569512 320090 569540 327168
rect 569960 327150 570012 327156
rect 569960 327072 570012 327078
rect 569788 327032 569960 327060
rect 569788 320736 569816 327032
rect 569960 327014 570012 327020
rect 569960 325712 570012 325718
rect 569880 325672 569960 325700
rect 569880 320906 569908 325672
rect 569960 325654 570012 325660
rect 570064 325122 570092 330262
rect 570156 325582 570184 330398
rect 570144 325576 570196 325582
rect 570144 325518 570196 325524
rect 569972 325094 570092 325122
rect 569972 321026 570000 325094
rect 570052 325032 570104 325038
rect 570052 324974 570104 324980
rect 569960 321020 570012 321026
rect 569960 320962 570012 320968
rect 569880 320890 570000 320906
rect 569880 320884 570012 320890
rect 569880 320878 569960 320884
rect 569960 320826 570012 320832
rect 570064 320754 570092 324974
rect 570144 321020 570196 321026
rect 570144 320962 570196 320968
rect 570052 320748 570104 320754
rect 569788 320708 569908 320736
rect 569880 320498 569908 320708
rect 570052 320690 570104 320696
rect 570156 320634 570184 320962
rect 569788 320470 569908 320498
rect 570064 320606 570184 320634
rect 569512 320062 569632 320090
rect 569236 315472 569540 315500
rect 569144 315166 569264 315194
rect 568776 314758 568896 314786
rect 1952 293412 2004 293418
rect 1952 293354 2004 293360
rect 1952 293140 2004 293146
rect 1952 293082 2004 293088
rect 1964 284866 1992 293082
rect 2240 288130 2268 295446
rect 2976 288266 3004 298710
rect 3344 298058 3372 301702
rect 3344 298030 3464 298058
rect 3436 296698 3464 298030
rect 3160 296670 3464 296698
rect 3160 296120 3188 296670
rect 3620 296562 3648 302654
rect 3700 301844 3752 301850
rect 3752 301804 3832 301832
rect 3700 301786 3752 301792
rect 3344 296534 3648 296562
rect 3344 296120 3372 296534
rect 3068 296092 3372 296120
rect 3068 295202 3096 296092
rect 3160 296018 3188 296092
rect 3160 295990 3464 296018
rect 3436 295984 3464 295990
rect 3436 295956 3648 295984
rect 3068 295174 3188 295202
rect 2976 288238 3096 288266
rect 2240 288102 3004 288130
rect 1964 284838 2912 284866
rect 1952 284776 2004 284782
rect 2004 284736 2820 284764
rect 1952 284718 2004 284724
rect 1952 284640 2004 284646
rect 2004 284600 2544 284628
rect 1952 284582 2004 284588
rect 1952 284368 2004 284374
rect 2004 284316 2452 284322
rect 1952 284310 2452 284316
rect 1964 284294 2452 284310
rect 1952 283960 2004 283966
rect 2004 283920 2176 283948
rect 1952 283902 2004 283908
rect 1952 283416 2004 283422
rect 2004 283364 2084 283370
rect 1952 283358 2084 283364
rect 1964 283342 2084 283358
rect 1952 283280 2004 283286
rect 1952 283222 2004 283228
rect 1964 273970 1992 283222
rect 1952 273964 2004 273970
rect 1952 273906 2004 273912
rect 2056 270314 2084 283342
rect 2148 273306 2176 283920
rect 2424 276706 2452 284294
rect 2516 276842 2544 284600
rect 2516 276814 2728 276842
rect 2240 276678 2452 276706
rect 2240 274938 2268 276678
rect 2700 276570 2728 276814
rect 2608 276542 2728 276570
rect 2608 276434 2636 276542
rect 2516 276406 2636 276434
rect 2516 275754 2544 276406
rect 2792 276162 2820 284736
rect 2884 281602 2912 284838
rect 2976 281738 3004 288102
rect 3068 282554 3096 288238
rect 3160 283404 3188 295174
rect 3620 283404 3648 295956
rect 3804 283404 3832 301804
rect 568224 300370 568252 314758
rect 568316 309856 568344 314758
rect 568868 314654 568896 314758
rect 568868 314626 568988 314654
rect 568960 310570 568988 314626
rect 568408 310542 568988 310570
rect 568408 309856 568436 310542
rect 568316 309828 568528 309856
rect 568408 309754 568436 309828
rect 568316 309726 568436 309754
rect 568316 308394 568344 309726
rect 568500 309346 568528 309828
rect 568408 309318 568528 309346
rect 568592 309318 568988 309346
rect 568408 308530 568436 309318
rect 568592 309108 568620 309318
rect 568960 309108 568988 309318
rect 568500 309080 568620 309108
rect 568868 309080 568988 309108
rect 568500 308530 568528 309080
rect 568868 308666 568896 309080
rect 568868 308638 569080 308666
rect 568408 308502 568988 308530
rect 568500 308394 568528 308502
rect 568316 308366 568712 308394
rect 568500 300642 568528 308366
rect 568684 301050 568712 308366
rect 568960 302818 568988 308502
rect 569052 304994 569080 308638
rect 569236 304994 569264 315166
rect 569512 314650 569540 315472
rect 569604 315330 569632 320062
rect 569788 315636 569816 320470
rect 569960 317960 570012 317966
rect 569880 317908 569960 317914
rect 569880 317902 570012 317908
rect 569880 317886 570000 317902
rect 569880 315772 569908 317886
rect 570064 315858 570092 320606
rect 570052 315852 570104 315858
rect 570052 315794 570104 315800
rect 569880 315744 570000 315772
rect 569972 315738 570000 315744
rect 569972 315710 570184 315738
rect 569960 315648 570012 315654
rect 569788 315608 569960 315636
rect 569960 315590 570012 315596
rect 570052 315580 570104 315586
rect 570052 315522 570104 315528
rect 569604 315302 570000 315330
rect 569420 314622 569540 314650
rect 569420 309856 569448 314622
rect 569052 304966 569264 304994
rect 569328 309828 569448 309856
rect 568960 302790 569172 302818
rect 569144 301050 569172 302790
rect 568684 301022 569264 301050
rect 569144 300880 569172 301022
rect 569052 300852 569172 300880
rect 568500 300614 568712 300642
rect 568224 300342 568528 300370
rect 568500 300132 568528 300342
rect 568684 300234 568712 300614
rect 568592 300206 568712 300234
rect 568592 300132 568620 300206
rect 3160 283376 3464 283404
rect 3436 282962 3464 283376
rect 3528 283376 3832 283404
rect 568224 300104 568620 300132
rect 3528 282962 3556 283376
rect 3620 283098 3648 283376
rect 3620 283070 3740 283098
rect 3712 282962 3740 283070
rect 3436 282934 3832 282962
rect 3068 282526 3464 282554
rect 3436 282146 3464 282526
rect 3528 282282 3556 282934
rect 3528 282254 3648 282282
rect 3344 282118 3464 282146
rect 3344 282010 3372 282118
rect 3252 281982 3372 282010
rect 2976 281710 3188 281738
rect 2884 281574 3096 281602
rect 3068 281466 3096 281574
rect 2884 281438 3096 281466
rect 2884 276298 2912 281438
rect 3160 277930 3188 281710
rect 3252 277930 3280 281982
rect 2976 277902 3280 277930
rect 2976 276706 3004 277902
rect 3160 277522 3188 277902
rect 3160 277494 3464 277522
rect 2976 276678 3280 276706
rect 2884 276270 3004 276298
rect 2608 276134 2820 276162
rect 2608 275754 2636 276134
rect 2516 275726 2912 275754
rect 2608 275346 2636 275726
rect 2608 275318 2820 275346
rect 2240 274910 2728 274938
rect 2148 273278 2636 273306
rect 2056 270286 2360 270314
rect 1952 270224 2004 270230
rect 2004 270172 2268 270178
rect 1952 270166 2268 270172
rect 1964 270150 2268 270166
rect 1952 269816 2004 269822
rect 2004 269776 2176 269804
rect 1952 269758 2004 269764
rect 1952 269408 2004 269414
rect 1952 269350 2004 269356
rect 1964 266626 1992 269350
rect 2148 266642 2176 269776
rect 1952 266620 2004 266626
rect 1952 266562 2004 266568
rect 2056 266614 2176 266642
rect 2056 266506 2084 266614
rect 1964 266490 2084 266506
rect 1952 266484 2084 266490
rect 2004 266478 2084 266484
rect 1952 266426 2004 266432
rect 1952 266348 2004 266354
rect 2240 266336 2268 270150
rect 2004 266308 2268 266336
rect 1952 266290 2004 266296
rect 2332 264738 2360 270286
rect 1964 264722 2360 264738
rect 1952 264716 2360 264722
rect 2004 264710 2360 264716
rect 1952 264658 2004 264664
rect 2608 264466 2636 273278
rect 1964 264438 2636 264466
rect 1964 264314 1992 264438
rect 1952 264308 2004 264314
rect 1952 264250 2004 264256
rect 1964 264178 2176 264194
rect 1952 264172 2176 264178
rect 2004 264166 2176 264172
rect 1952 264114 2004 264120
rect 1952 264036 2004 264042
rect 1952 263978 2004 263984
rect 1860 261520 1912 261526
rect 1860 261462 1912 261468
rect 1768 260772 1820 260778
rect 1768 260714 1820 260720
rect 1768 258256 1820 258262
rect 1768 258198 1820 258204
rect 1780 242214 1808 258198
rect 1964 257530 1992 263978
rect 2148 261474 2176 264166
rect 2700 263922 2728 274910
rect 2424 263894 2728 263922
rect 2424 262154 2452 263894
rect 2792 263650 2820 275318
rect 2884 267186 2912 275726
rect 2976 269090 3004 276270
rect 3252 269226 3280 276678
rect 3436 276434 3464 277494
rect 3160 269198 3280 269226
rect 3344 276406 3464 276434
rect 3160 269090 3188 269198
rect 2976 269062 3280 269090
rect 3160 268682 3188 269062
rect 3068 268654 3188 268682
rect 3068 268274 3096 268654
rect 2976 268246 3096 268274
rect 2976 268002 3004 268246
rect 2976 267974 3096 268002
rect 3068 267186 3096 267974
rect 2884 267158 3188 267186
rect 2608 263622 2820 263650
rect 2608 262154 2636 263622
rect 3068 263378 3096 267158
rect 2792 263350 3096 263378
rect 2792 262290 2820 263350
rect 3160 262562 3188 267158
rect 3068 262534 3188 262562
rect 2792 262262 3004 262290
rect 2976 262154 3004 262262
rect 3068 262154 3096 262534
rect 2424 262126 2544 262154
rect 2608 262126 2820 262154
rect 2976 262126 3188 262154
rect 2516 262018 2544 262126
rect 2516 261990 2636 262018
rect 2056 261446 2176 261474
rect 2056 258210 2084 261446
rect 2608 258210 2636 261990
rect 2056 258182 2728 258210
rect 1964 257502 2452 257530
rect 1952 257304 2004 257310
rect 2004 257252 2084 257258
rect 1952 257246 2084 257252
rect 1964 257230 2084 257246
rect 2056 256986 2084 257230
rect 2056 256958 2268 256986
rect 2240 251954 2268 256958
rect 2056 251926 2268 251954
rect 1860 251864 1912 251870
rect 1860 251806 1912 251812
rect 1872 242282 1900 251806
rect 2056 250322 2084 251926
rect 1964 250306 2084 250322
rect 1952 250300 2084 250306
rect 2004 250294 2084 250300
rect 1952 250242 2004 250248
rect 1952 250164 2004 250170
rect 1952 250106 2004 250112
rect 1964 249098 1992 250106
rect 1964 249070 2084 249098
rect 1952 249008 2004 249014
rect 1952 248950 2004 248956
rect 1964 243098 1992 248950
rect 1952 243092 2004 243098
rect 1952 243034 2004 243040
rect 1952 242956 2004 242962
rect 1952 242898 2004 242904
rect 1964 242554 1992 242898
rect 1952 242548 2004 242554
rect 1952 242490 2004 242496
rect 2056 242298 2084 249070
rect 2424 247738 2452 257502
rect 1964 242282 2084 242298
rect 1860 242276 1912 242282
rect 1860 242218 1912 242224
rect 1952 242276 2084 242282
rect 2004 242270 2084 242276
rect 2148 247710 2452 247738
rect 1952 242218 2004 242224
rect 1768 242208 1820 242214
rect 2148 242162 2176 247710
rect 2608 242978 2636 258182
rect 1768 242150 1820 242156
rect 1872 242134 2176 242162
rect 2332 242950 2636 242978
rect 1768 242072 1820 242078
rect 1768 242014 1820 242020
rect 1780 238202 1808 242014
rect 1768 238196 1820 238202
rect 1768 238138 1820 238144
rect 1872 238082 1900 242134
rect 1952 241664 2004 241670
rect 2004 241624 2084 241652
rect 1952 241606 2004 241612
rect 1952 238468 2004 238474
rect 2056 238456 2084 241624
rect 2004 238428 2084 238456
rect 1952 238410 2004 238416
rect 1952 238332 2004 238338
rect 2004 238292 2268 238320
rect 1952 238274 2004 238280
rect 1952 238196 2004 238202
rect 1952 238138 2004 238144
rect 1780 238054 1900 238082
rect 1780 235482 1808 238054
rect 1860 237992 1912 237998
rect 1860 237934 1912 237940
rect 1768 235476 1820 235482
rect 1768 235418 1820 235424
rect 1768 228404 1820 228410
rect 1768 228346 1820 228352
rect 1780 178430 1808 228346
rect 1872 179654 1900 237934
rect 1964 221746 1992 238138
rect 2240 226114 2268 238292
rect 2148 226086 2268 226114
rect 1952 221740 2004 221746
rect 1952 221682 2004 221688
rect 2148 221082 2176 226086
rect 1964 221066 2176 221082
rect 1952 221060 2176 221066
rect 2004 221054 2176 221060
rect 1952 221002 2004 221008
rect 1952 219972 2004 219978
rect 2332 219960 2360 242950
rect 2700 234274 2728 258182
rect 2424 234246 2728 234274
rect 2424 233730 2452 234246
rect 2792 234002 2820 262126
rect 3068 256986 3096 262126
rect 2884 256958 3096 256986
rect 2884 234002 2912 256958
rect 3160 256850 3188 262126
rect 2700 233974 2912 234002
rect 2976 256822 3188 256850
rect 2700 233866 2728 233974
rect 2608 233838 2728 233866
rect 2792 233866 2820 233974
rect 2792 233838 2912 233866
rect 2608 233730 2636 233838
rect 2424 233702 2820 233730
rect 2608 232234 2636 233702
rect 2004 219932 2360 219960
rect 2516 232206 2636 232234
rect 1952 219914 2004 219920
rect 2516 218362 2544 232206
rect 1964 218346 2544 218362
rect 1952 218340 2544 218346
rect 2004 218334 2544 218340
rect 1952 218282 2004 218288
rect 1952 217728 2004 217734
rect 2004 217676 2360 217682
rect 1952 217670 2360 217676
rect 1964 217654 2360 217670
rect 2332 217444 2360 217654
rect 2332 217416 2452 217444
rect 2424 216594 2452 217416
rect 2792 217410 2820 233702
rect 1964 216566 2452 216594
rect 2608 217382 2820 217410
rect 1964 214334 1992 216566
rect 1952 214328 2004 214334
rect 1952 214270 2004 214276
rect 1952 214192 2004 214198
rect 2004 214140 2084 214146
rect 1952 214134 2084 214140
rect 1964 214118 2084 214134
rect 1952 212900 2004 212906
rect 1952 212842 2004 212848
rect 1964 204882 1992 212842
rect 1952 204876 2004 204882
rect 1952 204818 2004 204824
rect 2056 204762 2084 214118
rect 2608 207890 2636 217382
rect 1964 204746 2084 204762
rect 1952 204740 2084 204746
rect 2004 204734 2084 204740
rect 2148 207862 2636 207890
rect 1952 204682 2004 204688
rect 2148 203674 2176 207862
rect 2884 203946 2912 233838
rect 2976 232642 3004 256822
rect 3252 256714 3280 269062
rect 3068 256686 3280 256714
rect 3068 255218 3096 256686
rect 3344 256000 3372 276406
rect 3620 274394 3648 282254
rect 3160 255972 3372 256000
rect 3436 274366 3648 274394
rect 3160 255354 3188 255972
rect 3160 255326 3372 255354
rect 3344 255218 3372 255326
rect 3436 255218 3464 274366
rect 3712 274258 3740 282934
rect 3528 274230 3740 274258
rect 3528 263378 3556 274230
rect 3528 263350 3648 263378
rect 3620 262970 3648 263350
rect 3620 262942 3740 262970
rect 3712 262698 3740 262942
rect 3804 262698 3832 282934
rect 568224 274224 568252 300104
rect 568500 284050 568528 300104
rect 569052 300098 569080 300852
rect 568684 300070 569080 300098
rect 568684 300064 568712 300070
rect 568592 300036 568712 300064
rect 568592 284322 568620 300036
rect 569236 295168 569264 301022
rect 569144 295140 569264 295168
rect 569144 284628 569172 295140
rect 569328 295066 569356 309828
rect 569972 309210 570000 315302
rect 569788 309182 570000 309210
rect 569788 309074 569816 309182
rect 569512 309046 569816 309074
rect 569960 309120 570012 309126
rect 569960 309062 570012 309068
rect 569512 301186 569540 309046
rect 569972 307850 570000 309062
rect 569880 307822 570000 307850
rect 569880 307578 569908 307822
rect 569880 307550 570000 307578
rect 569972 307018 570000 307550
rect 569960 307012 570012 307018
rect 569960 306954 570012 306960
rect 569960 306196 570012 306202
rect 569604 306156 569960 306184
rect 569604 302784 569632 306156
rect 569960 306138 570012 306144
rect 570064 304298 570092 315522
rect 570052 304292 570104 304298
rect 570052 304234 570104 304240
rect 569960 302796 570012 302802
rect 569604 302756 569960 302784
rect 569960 302738 570012 302744
rect 569512 301170 570000 301186
rect 569512 301164 570012 301170
rect 569512 301158 569960 301164
rect 569960 301106 570012 301112
rect 569960 300892 570012 300898
rect 569960 300834 570012 300840
rect 569972 300082 570000 300834
rect 570156 300150 570184 315710
rect 570248 315654 570276 330942
rect 572732 327690 572760 340983
rect 572720 327684 572772 327690
rect 572720 327626 572772 327632
rect 570328 315852 570380 315858
rect 570328 315794 570380 315800
rect 570236 315648 570288 315654
rect 570236 315590 570288 315596
rect 570236 315512 570288 315518
rect 570236 315454 570288 315460
rect 570248 303890 570276 315454
rect 570236 303884 570288 303890
rect 570236 303826 570288 303832
rect 570340 302954 570368 315794
rect 572718 313848 572774 313857
rect 572718 313783 572774 313792
rect 570248 302926 570368 302954
rect 570144 300144 570196 300150
rect 570144 300086 570196 300092
rect 569960 300076 570012 300082
rect 569960 300018 570012 300024
rect 569960 298580 570012 298586
rect 569604 298540 569960 298568
rect 569604 296426 569632 298540
rect 569960 298522 570012 298528
rect 569960 298444 570012 298450
rect 569960 298386 570012 298392
rect 569236 295038 569356 295066
rect 569512 296398 569632 296426
rect 569236 291530 569264 295038
rect 569512 294250 569540 296398
rect 569972 296290 570000 298386
rect 569420 294222 569540 294250
rect 569604 296262 570000 296290
rect 569236 291502 569356 291530
rect 569328 284866 569356 291502
rect 569420 285002 569448 294222
rect 569604 293706 569632 296262
rect 570052 296200 570104 296206
rect 570052 296142 570104 296148
rect 569960 296132 570012 296138
rect 569960 296074 570012 296080
rect 569972 296018 570000 296074
rect 569512 293678 569632 293706
rect 569696 295990 570000 296018
rect 569512 285172 569540 293678
rect 569696 292890 569724 295990
rect 570064 293298 570092 296142
rect 570248 296070 570276 302926
rect 570420 300416 570472 300422
rect 570420 300358 570472 300364
rect 570328 300280 570380 300286
rect 570328 300222 570380 300228
rect 570236 296064 570288 296070
rect 570236 296006 570288 296012
rect 570340 295186 570368 300222
rect 570328 295180 570380 295186
rect 570328 295122 570380 295128
rect 569604 292862 569724 292890
rect 569788 293270 570092 293298
rect 569604 285274 569632 292862
rect 569788 287858 569816 293270
rect 570236 292800 570288 292806
rect 570236 292742 570288 292748
rect 569960 292460 570012 292466
rect 569960 292402 570012 292408
rect 569972 289678 570000 292402
rect 569960 289672 570012 289678
rect 569960 289614 570012 289620
rect 569788 287830 570000 287858
rect 569972 285394 570000 287830
rect 570248 285530 570276 292742
rect 570432 292602 570460 300358
rect 570420 292596 570472 292602
rect 570420 292538 570472 292544
rect 570328 288312 570380 288318
rect 570328 288254 570380 288260
rect 570236 285524 570288 285530
rect 570236 285466 570288 285472
rect 569960 285388 570012 285394
rect 569960 285330 570012 285336
rect 569604 285246 570092 285274
rect 569960 285184 570012 285190
rect 569512 285144 569960 285172
rect 569960 285126 570012 285132
rect 569420 284986 570000 285002
rect 569420 284980 570012 284986
rect 569420 284974 569960 284980
rect 569960 284922 570012 284928
rect 569328 284850 570000 284866
rect 569328 284844 570012 284850
rect 569328 284838 569960 284844
rect 569960 284786 570012 284792
rect 569960 284640 570012 284646
rect 569144 284600 569960 284628
rect 569960 284582 570012 284588
rect 568592 284294 570000 284322
rect 568500 284022 568712 284050
rect 568684 283642 568712 284022
rect 569972 283898 570000 284294
rect 569960 283892 570012 283898
rect 569960 283834 570012 283840
rect 569960 283756 570012 283762
rect 569960 283698 570012 283704
rect 569972 283642 570000 283698
rect 568500 283614 568712 283642
rect 569052 283614 570000 283642
rect 568500 276842 568528 283614
rect 569052 277386 569080 283614
rect 569960 283552 570012 283558
rect 569144 283500 569960 283506
rect 569144 283494 570012 283500
rect 569144 283478 570000 283494
rect 570064 283490 570092 285246
rect 570052 283484 570104 283490
rect 569144 277556 569172 283478
rect 570052 283426 570104 283432
rect 569960 283416 570012 283422
rect 569236 283376 569960 283404
rect 569236 277964 569264 283376
rect 570340 283370 570368 288254
rect 570418 286104 570474 286113
rect 570418 286039 570474 286048
rect 569960 283358 570012 283364
rect 570052 283348 570104 283354
rect 570052 283290 570104 283296
rect 570156 283342 570368 283370
rect 569960 277976 570012 277982
rect 569236 277936 569960 277964
rect 569960 277918 570012 277924
rect 569960 277568 570012 277574
rect 569144 277528 569960 277556
rect 569960 277510 570012 277516
rect 569052 277358 569264 277386
rect 569236 277284 569264 277358
rect 569960 277296 570012 277302
rect 569236 277256 569960 277284
rect 569960 277238 570012 277244
rect 568500 276814 570000 276842
rect 569972 274514 570000 276814
rect 569960 274508 570012 274514
rect 569960 274450 570012 274456
rect 569960 274236 570012 274242
rect 568224 274196 569960 274224
rect 569960 274178 570012 274184
rect 570064 274122 570092 283290
rect 570156 277658 570184 283342
rect 570328 277976 570380 277982
rect 570328 277918 570380 277924
rect 570156 277630 570276 277658
rect 570144 277568 570196 277574
rect 570144 277510 570196 277516
rect 569972 274094 570092 274122
rect 569972 273086 570000 274094
rect 570052 273760 570104 273766
rect 570052 273702 570104 273708
rect 569960 273080 570012 273086
rect 569960 273022 570012 273028
rect 569960 272944 570012 272950
rect 3528 262670 3832 262698
rect 568224 272892 569960 272898
rect 568224 272886 570012 272892
rect 568224 272870 570000 272886
rect 3528 257258 3556 262670
rect 3712 257394 3740 262670
rect 3712 257366 3832 257394
rect 3528 257230 3740 257258
rect 3068 255190 3648 255218
rect 3344 251410 3372 255190
rect 3068 251382 3372 251410
rect 3068 232778 3096 251382
rect 3436 245834 3464 255190
rect 3160 245806 3464 245834
rect 3160 239850 3188 245806
rect 3620 241346 3648 255190
rect 3344 241318 3648 241346
rect 3344 240122 3372 241318
rect 3712 240938 3740 257230
rect 3620 240910 3740 240938
rect 3620 240666 3648 240910
rect 3804 240802 3832 257366
rect 3712 240774 3832 240802
rect 3712 240666 3740 240774
rect 3620 240638 3832 240666
rect 3344 240094 3648 240122
rect 3160 239822 3556 239850
rect 3528 239714 3556 239822
rect 3620 239714 3648 240094
rect 3252 239686 3648 239714
rect 3252 234138 3280 239686
rect 3528 239442 3556 239686
rect 3712 239442 3740 240638
rect 3436 239414 3740 239442
rect 3436 234410 3464 239414
rect 3160 234110 3280 234138
rect 3344 234382 3464 234410
rect 3160 233730 3188 234110
rect 3344 234002 3372 234382
rect 3528 234002 3556 239414
rect 3252 233974 3556 234002
rect 3252 233730 3280 233974
rect 3344 233866 3372 233974
rect 3344 233838 3556 233866
rect 3160 233702 3464 233730
rect 3252 232778 3280 233702
rect 3068 232750 3372 232778
rect 2976 232614 3188 232642
rect 3160 225978 3188 232614
rect 1964 203646 2176 203674
rect 2240 203918 2912 203946
rect 2976 225950 3188 225978
rect 1964 201890 1992 203646
rect 1952 201884 2004 201890
rect 1952 201826 2004 201832
rect 2240 198234 2268 203918
rect 2976 203538 3004 225950
rect 3252 225706 3280 232750
rect 3160 225678 3280 225706
rect 3160 225434 3188 225678
rect 3344 225570 3372 232750
rect 3436 226386 3464 233702
rect 3528 226386 3556 233838
rect 3804 231690 3832 240638
rect 568224 236858 568252 272870
rect 569960 272808 570012 272814
rect 568500 272768 569960 272796
rect 568394 248432 568450 248441
rect 568316 248390 568394 248418
rect 568316 236994 568344 248390
rect 568394 248367 568450 248376
rect 568500 243794 568528 272768
rect 569960 272750 570012 272756
rect 569960 272604 570012 272610
rect 569960 272546 570012 272552
rect 569868 272400 569920 272406
rect 569868 272342 569920 272348
rect 569880 271810 569908 272342
rect 568684 271782 569908 271810
rect 568684 253858 568712 271782
rect 569972 271674 570000 272546
rect 568868 271646 570000 271674
rect 568868 271402 568896 271646
rect 569960 271584 570012 271590
rect 569960 271526 570012 271532
rect 568776 271374 568896 271402
rect 568776 262834 568804 271374
rect 569972 271266 570000 271526
rect 568868 271238 570000 271266
rect 568868 262970 568896 271238
rect 570064 271164 570092 273702
rect 568960 271136 570092 271164
rect 568960 263106 568988 271136
rect 569960 271040 570012 271046
rect 569052 270988 569960 270994
rect 569052 270982 570012 270988
rect 569052 270966 570000 270982
rect 569052 263242 569080 270966
rect 570156 270910 570184 277510
rect 569960 270904 570012 270910
rect 569144 270852 569960 270858
rect 569144 270846 570012 270852
rect 570144 270904 570196 270910
rect 570144 270846 570196 270852
rect 569144 270830 570000 270846
rect 569144 263378 569172 270830
rect 569960 270632 570012 270638
rect 569236 270580 569960 270586
rect 569236 270574 570012 270580
rect 569236 270558 570000 270574
rect 569236 263514 569264 270558
rect 569960 270496 570012 270502
rect 569328 270444 569960 270450
rect 569328 270438 570012 270444
rect 569328 270422 570000 270438
rect 569328 263650 569356 270422
rect 569960 270360 570012 270366
rect 569420 270308 569960 270314
rect 569420 270302 570012 270308
rect 569420 270286 570000 270302
rect 569420 264024 569448 270286
rect 570248 270230 570276 277630
rect 570340 270638 570368 277918
rect 570432 272610 570460 286039
rect 570512 284640 570564 284646
rect 570510 284608 570512 284617
rect 570564 284608 570566 284617
rect 570510 284543 570566 284552
rect 572732 272814 572760 313783
rect 572720 272808 572772 272814
rect 572720 272750 572772 272756
rect 570420 272604 570472 272610
rect 570420 272546 570472 272552
rect 570328 270632 570380 270638
rect 570328 270574 570380 270580
rect 569960 270224 570012 270230
rect 569512 270172 569960 270178
rect 569512 270166 570012 270172
rect 570236 270224 570288 270230
rect 570236 270166 570288 270172
rect 569512 270150 570000 270166
rect 569512 264194 569540 270150
rect 569960 270088 570012 270094
rect 569604 270036 569960 270042
rect 569604 270030 570012 270036
rect 569604 270014 570000 270030
rect 569604 266336 569632 270014
rect 569960 269952 570012 269958
rect 569696 269900 569960 269906
rect 569696 269894 570012 269900
rect 569696 269878 570000 269894
rect 569696 267050 569724 269878
rect 569960 269816 570012 269822
rect 569788 269764 569960 269770
rect 569788 269758 570012 269764
rect 569788 269742 570000 269758
rect 569788 267288 569816 269742
rect 569960 267300 570012 267306
rect 569788 267260 569960 267288
rect 569960 267242 570012 267248
rect 569696 267022 570000 267050
rect 569972 266422 570000 267022
rect 569960 266416 570012 266422
rect 569960 266358 570012 266364
rect 569604 266308 569816 266336
rect 569788 266234 569816 266308
rect 569788 266206 569908 266234
rect 569880 265928 569908 266206
rect 569960 265940 570012 265946
rect 569880 265900 569960 265928
rect 569960 265882 570012 265888
rect 569512 264166 570092 264194
rect 569960 264036 570012 264042
rect 569420 263996 569960 264024
rect 569960 263978 570012 263984
rect 569328 263622 569724 263650
rect 569236 263486 569540 263514
rect 569144 263350 569448 263378
rect 569052 263214 569356 263242
rect 568960 263078 569264 263106
rect 568868 262942 569172 262970
rect 568776 262806 568896 262834
rect 568592 253830 568712 253858
rect 568592 250186 568620 253830
rect 568868 250492 568896 262806
rect 569144 256034 569172 262942
rect 569236 260137 569264 263078
rect 569222 260128 569278 260137
rect 569222 260063 569278 260072
rect 568960 256006 569172 256034
rect 568960 250628 568988 256006
rect 569328 254674 569356 263214
rect 569052 254646 569356 254674
rect 569052 250730 569080 254646
rect 569420 254538 569448 263350
rect 569144 254510 569448 254538
rect 569144 250866 569172 254510
rect 569512 251682 569540 263486
rect 569696 252498 569724 263622
rect 570064 260012 570092 264166
rect 569788 259984 570092 260012
rect 569788 256442 569816 259984
rect 569960 259888 570012 259894
rect 569960 259830 570012 259836
rect 569972 259706 570000 259830
rect 569880 259678 570000 259706
rect 569880 256578 569908 259678
rect 569960 259616 570012 259622
rect 569960 259558 570012 259564
rect 569972 257258 570000 259558
rect 574756 259457 574784 438874
rect 580170 393000 580226 393009
rect 580170 392935 580226 392944
rect 580184 392018 580212 392935
rect 574836 392012 574888 392018
rect 574836 391954 574888 391960
rect 580172 392012 580224 392018
rect 580172 391954 580224 391960
rect 574742 259448 574798 259457
rect 574742 259383 574798 259392
rect 569972 257230 570092 257258
rect 569880 256562 570000 256578
rect 569880 256556 570012 256562
rect 569880 256550 569960 256556
rect 569960 256498 570012 256504
rect 569788 256414 570000 256442
rect 569972 254674 570000 256414
rect 570064 254794 570092 257230
rect 570236 256556 570288 256562
rect 570236 256498 570288 256504
rect 570052 254788 570104 254794
rect 570052 254730 570104 254736
rect 569972 254646 570092 254674
rect 569696 252470 570000 252498
rect 569972 251802 570000 252470
rect 569960 251796 570012 251802
rect 569960 251738 570012 251744
rect 569512 251654 570000 251682
rect 569972 250986 570000 251654
rect 569960 250980 570012 250986
rect 569960 250922 570012 250928
rect 569144 250850 570000 250866
rect 569144 250844 570012 250850
rect 569144 250838 569960 250844
rect 569960 250786 570012 250792
rect 569052 250702 569448 250730
rect 569420 250628 569448 250702
rect 569960 250640 570012 250646
rect 568960 250600 569356 250628
rect 569420 250600 569960 250628
rect 568868 250464 569264 250492
rect 568592 250158 569172 250186
rect 568408 243766 568528 243794
rect 568408 242978 568436 243766
rect 569144 243556 569172 250158
rect 569052 243528 569172 243556
rect 568408 242950 568712 242978
rect 568684 242842 568712 242950
rect 568684 242814 568988 242842
rect 568960 240666 568988 242814
rect 569052 240666 569080 243528
rect 569236 240802 569264 250464
rect 569328 240938 569356 250600
rect 569960 250582 570012 250588
rect 569960 250504 570012 250510
rect 569788 250452 569960 250458
rect 569788 250446 570012 250452
rect 569788 250430 570000 250446
rect 569788 248282 569816 250430
rect 569788 248254 570000 248282
rect 569972 247314 570000 248254
rect 569960 247308 570012 247314
rect 569960 247250 570012 247256
rect 570064 246702 570092 254646
rect 570144 251796 570196 251802
rect 570144 251738 570196 251744
rect 570052 246696 570104 246702
rect 570052 246638 570104 246644
rect 570052 246560 570104 246566
rect 570052 246502 570104 246508
rect 569960 243704 570012 243710
rect 569788 243664 569960 243692
rect 569788 242842 569816 243664
rect 569960 243646 570012 243652
rect 569960 243568 570012 243574
rect 569960 243510 570012 243516
rect 569696 242814 569816 242842
rect 569328 240910 569632 240938
rect 569236 240774 569540 240802
rect 568960 240638 569264 240666
rect 569052 240394 569080 240638
rect 569236 240530 569264 240638
rect 569236 240502 569448 240530
rect 569052 240366 569264 240394
rect 569236 237674 569264 240366
rect 568592 237646 569264 237674
rect 568592 236994 568620 237646
rect 568316 236966 568712 236994
rect 568224 236830 568528 236858
rect 568500 236586 568528 236830
rect 568408 236558 568528 236586
rect 568408 236178 568436 236558
rect 568408 236150 568528 236178
rect 568500 235362 568528 236150
rect 568316 235334 568528 235362
rect 568316 235226 568344 235334
rect 568592 235226 568620 236966
rect 568684 236450 568712 236966
rect 568684 236422 568804 236450
rect 3620 231662 3832 231690
rect 568224 235198 568620 235226
rect 3620 226522 3648 231662
rect 3620 226494 3832 226522
rect 3436 226358 3740 226386
rect 3528 226250 3556 226358
rect 3528 226222 3648 226250
rect 1964 198218 2268 198234
rect 1952 198212 2268 198218
rect 2004 198206 2268 198212
rect 2332 203510 3004 203538
rect 3068 225406 3188 225434
rect 3252 225542 3372 225570
rect 1952 198154 2004 198160
rect 2332 197826 2360 203510
rect 3068 203130 3096 225406
rect 3252 225298 3280 225542
rect 3160 225270 3280 225298
rect 3160 218770 3188 225270
rect 3620 219858 3648 226222
rect 3436 219830 3648 219858
rect 3436 219586 3464 219830
rect 3252 219558 3464 219586
rect 3252 219042 3280 219558
rect 3252 219014 3372 219042
rect 3344 218770 3372 219014
rect 3436 219014 3648 219042
rect 3436 218770 3464 219014
rect 3160 218742 3464 218770
rect 3344 218226 3372 218742
rect 3252 218198 3372 218226
rect 3252 210882 3280 218198
rect 3252 210854 3464 210882
rect 3436 203130 3464 210854
rect 1964 197810 2360 197826
rect 1952 197804 2360 197810
rect 2004 197798 2360 197804
rect 2976 203102 3096 203130
rect 3252 203102 3464 203130
rect 1952 197746 2004 197752
rect 2976 197690 3004 203102
rect 3252 202994 3280 203102
rect 3620 202994 3648 219014
rect 1964 197674 3004 197690
rect 1952 197668 3004 197674
rect 2004 197662 3004 197668
rect 3068 202966 3280 202994
rect 3436 202966 3648 202994
rect 1952 197610 2004 197616
rect 1952 196376 2004 196382
rect 2004 196324 2912 196330
rect 1952 196318 2912 196324
rect 1964 196302 2912 196318
rect 1952 196240 2004 196246
rect 2004 196200 2820 196228
rect 1952 196182 2004 196188
rect 1952 196104 2004 196110
rect 2004 196052 2728 196058
rect 1952 196046 2728 196052
rect 1964 196030 2728 196046
rect 1952 195968 2004 195974
rect 2004 195916 2636 195922
rect 1952 195910 2636 195916
rect 1964 195894 2636 195910
rect 1952 195832 2004 195838
rect 2004 195780 2176 195786
rect 1952 195774 2176 195780
rect 1964 195758 2176 195774
rect 2148 195242 2176 195758
rect 2148 195214 2544 195242
rect 1964 195090 2452 195106
rect 1952 195084 2452 195090
rect 2004 195078 2452 195084
rect 1952 195026 2004 195032
rect 1952 194948 2004 194954
rect 1952 194890 2004 194896
rect 1964 194834 1992 194890
rect 1964 194806 2360 194834
rect 1952 194744 2004 194750
rect 2004 194704 2176 194732
rect 1952 194686 2004 194692
rect 1952 193996 2004 194002
rect 2004 193956 2084 193984
rect 1952 193938 2004 193944
rect 2056 189938 2084 193956
rect 1964 189910 2084 189938
rect 1964 189786 1992 189910
rect 1952 189780 2004 189786
rect 1952 189722 2004 189728
rect 1952 189644 2004 189650
rect 2148 189632 2176 194704
rect 2004 189604 2176 189632
rect 1952 189586 2004 189592
rect 2332 189530 2360 194806
rect 2148 189502 2360 189530
rect 1952 189236 2004 189242
rect 2148 189224 2176 189502
rect 2424 189394 2452 195078
rect 2004 189196 2176 189224
rect 2332 189366 2452 189394
rect 1952 189178 2004 189184
rect 1952 188964 2004 188970
rect 2332 188952 2360 189366
rect 2516 189224 2544 195214
rect 2004 188924 2360 188952
rect 2424 189196 2544 189224
rect 1952 188906 2004 188912
rect 1952 188692 2004 188698
rect 2424 188680 2452 189196
rect 2608 188952 2636 195894
rect 2004 188652 2452 188680
rect 2516 188924 2636 188952
rect 1952 188634 2004 188640
rect 1952 188556 2004 188562
rect 2004 188516 2084 188544
rect 1952 188498 2004 188504
rect 1952 186516 2004 186522
rect 1952 186458 2004 186464
rect 1860 179648 1912 179654
rect 1860 179590 1912 179596
rect 1860 179104 1912 179110
rect 1860 179046 1912 179052
rect 1768 178424 1820 178430
rect 1768 178366 1820 178372
rect 1872 177002 1900 179046
rect 1964 177682 1992 186458
rect 1952 177676 2004 177682
rect 1952 177618 2004 177624
rect 1860 176996 1912 177002
rect 1860 176938 1912 176944
rect 2056 176882 2084 188516
rect 2516 186266 2544 188924
rect 2700 186266 2728 196030
rect 2240 186238 2544 186266
rect 2608 186238 2728 186266
rect 2240 177018 2268 186238
rect 2608 186130 2636 186238
rect 2332 186102 2636 186130
rect 2332 177290 2360 186102
rect 2792 185994 2820 196200
rect 2700 185966 2820 185994
rect 2700 177970 2728 185966
rect 2884 185586 2912 196302
rect 3068 193338 3096 202966
rect 3436 193338 3464 202966
rect 3712 195650 3740 226358
rect 2976 193310 3464 193338
rect 3620 195622 3740 195650
rect 2976 192114 3004 193310
rect 3068 192250 3096 193310
rect 3068 192222 3556 192250
rect 2976 192086 3188 192114
rect 2884 185558 3096 185586
rect 2870 185328 2926 185337
rect 2870 185263 2926 185272
rect 2700 177942 2820 177970
rect 2332 177262 2728 177290
rect 2240 176990 2636 177018
rect 1872 176854 2084 176882
rect 1768 176248 1820 176254
rect 1768 176190 1820 176196
rect 1676 134564 1728 134570
rect 1676 134506 1728 134512
rect 1596 134422 1716 134450
rect 1688 132410 1716 134422
rect 1780 133482 1808 176190
rect 1872 173194 1900 176854
rect 1952 176792 2004 176798
rect 2004 176740 2452 176746
rect 1952 176734 2452 176740
rect 1964 176718 2452 176734
rect 1952 176656 2004 176662
rect 2424 176610 2452 176718
rect 2004 176604 2360 176610
rect 1952 176598 2360 176604
rect 1964 176582 2360 176598
rect 2424 176582 2544 176610
rect 1952 176520 2004 176526
rect 2332 176508 2360 176582
rect 2004 176480 2268 176508
rect 2332 176480 2452 176508
rect 1952 176462 2004 176468
rect 1952 176384 2004 176390
rect 2240 176372 2268 176480
rect 2004 176344 2176 176372
rect 2240 176344 2360 176372
rect 1952 176326 2004 176332
rect 1952 176248 2004 176254
rect 2148 176236 2176 176344
rect 2004 176208 2084 176236
rect 2148 176208 2268 176236
rect 1952 176190 2004 176196
rect 2056 176100 2084 176208
rect 2056 176072 2176 176100
rect 1952 175976 2004 175982
rect 1952 175918 2004 175924
rect 1860 173188 1912 173194
rect 1860 173130 1912 173136
rect 1860 173052 1912 173058
rect 1860 172994 1912 173000
rect 1872 168994 1900 172994
rect 1964 169114 1992 175918
rect 1952 169108 2004 169114
rect 1952 169050 2004 169056
rect 1872 168966 2084 168994
rect 1952 168020 2004 168026
rect 2056 168008 2084 168966
rect 2004 167980 2084 168008
rect 1952 167962 2004 167968
rect 1952 167816 2004 167822
rect 2148 167804 2176 176072
rect 2004 167776 2176 167804
rect 1952 167758 2004 167764
rect 1952 167680 2004 167686
rect 2240 167668 2268 176208
rect 2004 167640 2268 167668
rect 1952 167622 2004 167628
rect 2332 167498 2360 176344
rect 1964 167470 2360 167498
rect 1964 167414 1992 167470
rect 1952 167408 2004 167414
rect 1952 167350 2004 167356
rect 1952 167272 2004 167278
rect 2424 167260 2452 176480
rect 2004 167232 2452 167260
rect 1952 167214 2004 167220
rect 2516 167090 2544 176582
rect 1872 167062 2544 167090
rect 1872 153814 1900 167062
rect 2608 166954 2636 176990
rect 1964 166938 2636 166954
rect 1952 166932 2636 166938
rect 2004 166926 2636 166932
rect 1952 166874 2004 166880
rect 2700 166818 2728 177262
rect 1964 166802 2728 166818
rect 1952 166796 2728 166802
rect 2004 166790 2728 166796
rect 1952 166738 2004 166744
rect 2792 166682 2820 177942
rect 1964 166654 2820 166682
rect 1964 166462 1992 166654
rect 1952 166456 2004 166462
rect 1952 166398 2004 166404
rect 1952 166320 2004 166326
rect 2004 166268 2360 166274
rect 1952 166262 2360 166268
rect 1964 166246 2360 166262
rect 1952 166048 2004 166054
rect 2332 166002 2360 166246
rect 2884 166002 2912 185263
rect 3068 185178 3096 185558
rect 2976 185150 3096 185178
rect 2976 172666 3004 185150
rect 3160 184226 3188 192086
rect 3528 191298 3556 192222
rect 3344 191270 3556 191298
rect 3344 191162 3372 191270
rect 3068 184198 3188 184226
rect 3252 191134 3372 191162
rect 3068 172802 3096 184198
rect 3252 183002 3280 191134
rect 3620 189122 3648 195622
rect 3804 195378 3832 226494
rect 568224 208978 568252 235198
rect 568316 234138 568344 235198
rect 568316 234110 568620 234138
rect 568592 231146 568620 234110
rect 568776 232098 568804 236422
rect 568776 232070 569080 232098
rect 568500 231118 568620 231146
rect 568500 223666 568528 231118
rect 569052 225706 569080 232070
rect 569420 231690 569448 240502
rect 568960 225678 569080 225706
rect 569236 231662 569448 231690
rect 568500 223638 568712 223666
rect 568224 208950 568344 208978
rect 568316 208400 568344 208950
rect 568684 208400 568712 223638
rect 568854 222320 568910 222329
rect 568960 222306 568988 225678
rect 569236 225570 569264 231662
rect 569512 231554 569540 240774
rect 569604 233594 569632 240910
rect 569696 233730 569724 242814
rect 569972 236094 570000 243510
rect 569960 236088 570012 236094
rect 569960 236030 570012 236036
rect 569696 233714 570000 233730
rect 569696 233708 570012 233714
rect 569696 233702 569960 233708
rect 569960 233650 570012 233656
rect 569604 233578 570000 233594
rect 569604 233572 570012 233578
rect 569604 233566 569960 233572
rect 569960 233514 570012 233520
rect 568910 222278 568988 222306
rect 569052 225542 569264 225570
rect 569328 231526 569540 231554
rect 568854 222255 568910 222264
rect 569052 220538 569080 225542
rect 568868 220510 569080 220538
rect 568868 209522 568896 220510
rect 569328 218770 569356 231526
rect 569960 230240 570012 230246
rect 569512 230188 569960 230194
rect 569512 230182 570012 230188
rect 569512 230166 570000 230182
rect 569512 223938 569540 230166
rect 569960 230036 570012 230042
rect 569960 229978 570012 229984
rect 569972 229922 570000 229978
rect 569696 229894 570000 229922
rect 569696 224346 569724 229894
rect 569960 229832 570012 229838
rect 569788 229780 569960 229786
rect 569788 229774 570012 229780
rect 569788 229758 570000 229774
rect 569788 225808 569816 229758
rect 570064 229702 570092 246502
rect 570156 239494 570184 251738
rect 570144 239488 570196 239494
rect 570144 239430 570196 239436
rect 570144 233572 570196 233578
rect 570144 233514 570196 233520
rect 570156 230042 570184 233514
rect 570144 230036 570196 230042
rect 570144 229978 570196 229984
rect 570144 229764 570196 229770
rect 570144 229706 570196 229712
rect 570052 229696 570104 229702
rect 570052 229638 570104 229644
rect 569960 229288 570012 229294
rect 569960 229230 570012 229236
rect 569972 228426 570000 229230
rect 569880 228398 570000 228426
rect 569880 227066 569908 228398
rect 569880 227038 570000 227066
rect 569972 226030 570000 227038
rect 570052 227044 570104 227050
rect 570052 226986 570104 226992
rect 569960 226024 570012 226030
rect 569960 225966 570012 225972
rect 569960 225820 570012 225826
rect 569788 225780 569960 225808
rect 569960 225762 570012 225768
rect 569604 224318 569724 224346
rect 569604 224074 569632 224318
rect 569604 224046 570000 224074
rect 569512 223910 569908 223938
rect 568960 218742 569356 218770
rect 568960 209658 568988 218742
rect 569880 216050 569908 223910
rect 569144 216022 569908 216050
rect 569144 209794 569172 216022
rect 569972 215694 570000 224046
rect 569960 215688 570012 215694
rect 569960 215630 570012 215636
rect 569960 215416 570012 215422
rect 569512 215376 569960 215404
rect 569144 209766 569448 209794
rect 568960 209630 569172 209658
rect 568868 209494 568988 209522
rect 568960 209386 568988 209494
rect 568960 209358 569080 209386
rect 569052 208570 569080 209358
rect 568776 208542 569080 208570
rect 568776 208400 568804 208542
rect 3160 182974 3280 183002
rect 3528 189094 3648 189122
rect 3712 195350 3832 195378
rect 568224 208372 568804 208400
rect 3160 180146 3188 182974
rect 3528 180282 3556 189094
rect 3712 184906 3740 195350
rect 568224 193474 568252 208372
rect 568316 203028 568344 208372
rect 568684 208298 568712 208372
rect 568684 208270 568804 208298
rect 568776 208026 568804 208270
rect 568684 207998 568804 208026
rect 568684 205578 568712 207998
rect 569144 205578 569172 209630
rect 568500 205550 569172 205578
rect 568500 203402 568528 205550
rect 568684 205442 568712 205550
rect 568592 205414 568712 205442
rect 568592 205170 568620 205414
rect 569420 205306 569448 209766
rect 568960 205278 569448 205306
rect 568592 205142 568712 205170
rect 568684 203402 568712 205142
rect 568960 203946 568988 205278
rect 569512 205034 569540 215376
rect 569960 215358 570012 215364
rect 569960 214668 570012 214674
rect 569960 214610 570012 214616
rect 569972 214146 570000 214610
rect 569696 214118 570000 214146
rect 569696 210202 569724 214118
rect 569960 214056 570012 214062
rect 569788 214004 569960 214010
rect 569788 213998 570012 214004
rect 569788 213982 570000 213998
rect 569788 212922 569816 213982
rect 569788 212894 569908 212922
rect 569880 211154 569908 212894
rect 569880 211126 570000 211154
rect 568868 203918 568988 203946
rect 569052 205006 569540 205034
rect 569604 210174 569724 210202
rect 568868 203402 568896 203918
rect 569052 203674 569080 205006
rect 569604 204898 569632 210174
rect 569972 209794 570000 211126
rect 569696 209766 570000 209794
rect 569696 205068 569724 209766
rect 569960 205080 570012 205086
rect 569696 205040 569960 205068
rect 569960 205022 570012 205028
rect 569236 204870 569632 204898
rect 569236 204320 569264 204870
rect 569960 204808 570012 204814
rect 568960 203646 569080 203674
rect 569144 204292 569264 204320
rect 569328 204768 569960 204796
rect 568960 203402 568988 203646
rect 568500 203374 568620 203402
rect 568684 203374 568804 203402
rect 568868 203374 569080 203402
rect 568592 203028 568620 203374
rect 568776 203130 568804 203374
rect 568776 203102 568896 203130
rect 568316 203000 568804 203028
rect 568592 193633 568620 203000
rect 568578 193624 568634 193633
rect 568578 193559 568634 193568
rect 568302 193488 568358 193497
rect 568224 193446 568302 193474
rect 568302 193423 568358 193432
rect 568776 191842 568804 203000
rect 568684 191814 568804 191842
rect 568684 188306 568712 191814
rect 568868 188408 568896 203102
rect 568592 188278 568712 188306
rect 568776 188380 568896 188408
rect 568592 188034 568620 188278
rect 568776 188034 568804 188380
rect 568960 188306 568988 203374
rect 569052 188408 569080 203374
rect 569144 191740 569172 204292
rect 569328 203708 569356 204768
rect 569960 204750 570012 204756
rect 570064 204626 570092 226986
rect 570156 214606 570184 229706
rect 570248 226914 570276 256498
rect 574744 251252 574796 251258
rect 574744 251194 574796 251200
rect 570328 250844 570380 250850
rect 570328 250786 570380 250792
rect 570340 229838 570368 250786
rect 570420 229900 570472 229906
rect 570420 229842 570472 229848
rect 570328 229832 570380 229838
rect 570328 229774 570380 229780
rect 570236 226908 570288 226914
rect 570236 226850 570288 226856
rect 570236 226024 570288 226030
rect 570236 225966 570288 225972
rect 570144 214600 570196 214606
rect 570144 214542 570196 214548
rect 570248 214062 570276 225966
rect 570236 214056 570288 214062
rect 570236 213998 570288 214004
rect 570432 208418 570460 229842
rect 570144 208412 570196 208418
rect 570144 208354 570196 208360
rect 570420 208412 570472 208418
rect 570420 208354 570472 208360
rect 569972 204598 570092 204626
rect 569972 203726 570000 204598
rect 570052 204468 570104 204474
rect 570052 204410 570104 204416
rect 569236 203680 569356 203708
rect 569960 203720 570012 203726
rect 569236 191842 569264 203680
rect 569960 203662 570012 203668
rect 569960 203584 570012 203590
rect 569328 203544 569960 203572
rect 569328 192114 569356 203544
rect 569960 203526 570012 203532
rect 569960 203448 570012 203454
rect 569420 203396 569960 203402
rect 569420 203390 570012 203396
rect 569420 203374 570000 203390
rect 569420 192250 569448 203374
rect 569960 203176 570012 203182
rect 569512 203124 569960 203130
rect 569512 203118 570012 203124
rect 569512 203102 570000 203118
rect 569512 192386 569540 203102
rect 569960 203040 570012 203046
rect 569604 202988 569960 202994
rect 569604 202982 570012 202988
rect 569604 202966 570000 202982
rect 569604 192488 569632 202966
rect 569960 202632 570012 202638
rect 569696 202580 569960 202586
rect 569696 202574 570012 202580
rect 569696 202558 570000 202574
rect 569696 192794 569724 202558
rect 570064 198914 570092 204410
rect 569788 198886 570092 198914
rect 569788 192930 569816 198886
rect 570156 198778 570184 208354
rect 570236 205080 570288 205086
rect 570236 205022 570288 205028
rect 570248 203454 570276 205022
rect 570236 203448 570288 203454
rect 570236 203390 570288 203396
rect 569880 198750 570184 198778
rect 569880 196602 569908 198750
rect 569880 196574 570000 196602
rect 569972 193934 570000 196574
rect 569960 193928 570012 193934
rect 569960 193870 570012 193876
rect 570326 193624 570382 193633
rect 570326 193559 570382 193568
rect 569788 192902 570000 192930
rect 569696 192766 569816 192794
rect 569972 192778 570000 192902
rect 569788 192658 569816 192766
rect 569960 192772 570012 192778
rect 569960 192714 570012 192720
rect 569788 192630 570000 192658
rect 569972 192506 570000 192630
rect 569960 192500 570012 192506
rect 569604 192460 569908 192488
rect 569880 192386 569908 192460
rect 569960 192442 570012 192448
rect 569512 192358 569632 192386
rect 569880 192358 570092 192386
rect 569420 192222 569540 192250
rect 569512 192114 569540 192222
rect 569604 192216 569632 192358
rect 569960 192228 570012 192234
rect 569604 192188 569960 192216
rect 569960 192170 570012 192176
rect 569328 192086 569448 192114
rect 569512 192098 570000 192114
rect 569512 192092 570012 192098
rect 569512 192086 569960 192092
rect 569420 191978 569448 192086
rect 569960 192034 570012 192040
rect 570064 192030 570092 192358
rect 570052 192024 570104 192030
rect 569420 191962 570000 191978
rect 570052 191966 570104 191972
rect 569420 191956 570012 191962
rect 569420 191950 569960 191956
rect 569960 191898 570012 191904
rect 569236 191814 570276 191842
rect 569960 191752 570012 191758
rect 569144 191712 569960 191740
rect 569960 191694 570012 191700
rect 570052 191752 570104 191758
rect 570052 191694 570104 191700
rect 569960 191616 570012 191622
rect 569328 191564 569960 191570
rect 569328 191558 570012 191564
rect 569328 191542 570000 191558
rect 569328 188408 569356 191542
rect 569960 191480 570012 191486
rect 569960 191422 570012 191428
rect 569972 191298 570000 191422
rect 569880 191270 570000 191298
rect 569880 188714 569908 191270
rect 569696 188686 569908 188714
rect 569052 188380 569632 188408
rect 568960 188278 569172 188306
rect 568224 188006 568804 188034
rect 3712 184878 3832 184906
rect 3528 180254 3740 180282
rect 3160 180118 3280 180146
rect 3252 180010 3280 180118
rect 3252 179982 3464 180010
rect 3436 179602 3464 179982
rect 3436 179574 3556 179602
rect 3160 179302 3464 179330
rect 3160 173074 3188 179302
rect 3436 178922 3464 179302
rect 3528 179058 3556 179574
rect 3528 179030 3648 179058
rect 3620 178922 3648 179030
rect 3712 178922 3740 180254
rect 3436 178894 3740 178922
rect 3620 178786 3648 178894
rect 3252 178758 3648 178786
rect 3252 174298 3280 178758
rect 3804 177018 3832 184878
rect 3620 176990 3832 177018
rect 3620 174298 3648 176990
rect 3252 174270 3832 174298
rect 3620 173074 3648 174270
rect 3160 173046 3740 173074
rect 3068 172774 3372 172802
rect 3344 172666 3372 172774
rect 2976 172638 3556 172666
rect 3344 172394 3372 172638
rect 2004 165996 2176 166002
rect 1952 165990 2176 165996
rect 1964 165974 2176 165990
rect 2332 165974 2912 166002
rect 2976 172366 3372 172394
rect 1952 165912 2004 165918
rect 1952 165854 2004 165860
rect 1964 165594 1992 165854
rect 2148 165730 2176 165974
rect 2148 165702 2820 165730
rect 1964 165566 2728 165594
rect 1952 165504 2004 165510
rect 1952 165446 2004 165452
rect 1964 160002 1992 165446
rect 2700 160290 2728 165566
rect 2424 160262 2728 160290
rect 1952 159996 2004 160002
rect 1952 159938 2004 159944
rect 1952 159860 2004 159866
rect 2004 159820 2084 159848
rect 1952 159802 2004 159808
rect 1952 159724 2004 159730
rect 1952 159666 2004 159672
rect 1964 159474 1992 159666
rect 2056 159576 2084 159820
rect 2056 159548 2268 159576
rect 1964 159446 2176 159474
rect 1952 159316 2004 159322
rect 2004 159276 2084 159304
rect 1952 159258 2004 159264
rect 1952 159180 2004 159186
rect 1952 159122 2004 159128
rect 1964 154086 1992 159122
rect 1952 154080 2004 154086
rect 1952 154022 2004 154028
rect 1860 153808 1912 153814
rect 1860 153750 1912 153756
rect 2056 151178 2084 159276
rect 1872 151150 2084 151178
rect 1872 145926 1900 151150
rect 2148 151042 2176 159446
rect 1964 151014 2176 151042
rect 1964 147150 1992 151014
rect 2240 150906 2268 159548
rect 2424 153218 2452 160262
rect 2792 160120 2820 165702
rect 2056 150878 2268 150906
rect 2332 153190 2452 153218
rect 2608 160092 2820 160120
rect 1952 147144 2004 147150
rect 1952 147086 2004 147092
rect 1952 147008 2004 147014
rect 1952 146950 2004 146956
rect 1860 145920 1912 145926
rect 1860 145862 1912 145868
rect 1964 145858 1992 146950
rect 1952 145852 2004 145858
rect 1952 145794 2004 145800
rect 2056 145738 2084 150878
rect 2332 148322 2360 153190
rect 1872 145722 2084 145738
rect 1860 145716 2084 145722
rect 1912 145710 2084 145716
rect 2240 148294 2360 148322
rect 1860 145658 1912 145664
rect 1952 145648 2004 145654
rect 1952 145590 2004 145596
rect 1860 143132 1912 143138
rect 1860 143074 1912 143080
rect 1872 141302 1900 143074
rect 1964 141370 1992 145590
rect 1952 141364 2004 141370
rect 1952 141306 2004 141312
rect 1860 141296 1912 141302
rect 2240 141250 2268 148294
rect 2608 146690 2636 160092
rect 2976 160018 3004 172366
rect 2700 159990 3004 160018
rect 3068 172230 3372 172258
rect 2700 148050 2728 159990
rect 3068 158794 3096 172230
rect 3344 171850 3372 172230
rect 3528 171850 3556 172638
rect 3620 171850 3648 173046
rect 3344 171822 3648 171850
rect 3528 171714 3556 171822
rect 3528 171686 3648 171714
rect 3068 158766 3280 158794
rect 3252 151178 3280 158766
rect 3068 151150 3280 151178
rect 2700 148022 2912 148050
rect 2608 146662 2728 146690
rect 1860 141238 1912 141244
rect 1964 141234 2268 141250
rect 1952 141228 2268 141234
rect 2004 141222 2268 141228
rect 1952 141170 2004 141176
rect 1860 141160 1912 141166
rect 1860 141102 1912 141108
rect 1872 134638 1900 141102
rect 1952 140004 2004 140010
rect 2700 139992 2728 146662
rect 2780 143676 2832 143682
rect 2780 143618 2832 143624
rect 2004 139964 2728 139992
rect 1952 139946 2004 139952
rect 2792 139856 2820 143618
rect 2516 139828 2820 139856
rect 1952 139120 2004 139126
rect 2004 139068 2452 139074
rect 1952 139062 2452 139068
rect 1964 139046 2452 139062
rect 1952 138916 2004 138922
rect 2004 138876 2360 138904
rect 1952 138858 2004 138864
rect 1952 138644 2004 138650
rect 2004 138604 2268 138632
rect 1952 138586 2004 138592
rect 1952 138304 2004 138310
rect 2004 138252 2084 138258
rect 1952 138246 2084 138252
rect 1964 138230 2084 138246
rect 1952 137964 2004 137970
rect 1952 137906 2004 137912
rect 1860 134632 1912 134638
rect 1860 134574 1912 134580
rect 1964 134502 1992 137906
rect 1952 134496 2004 134502
rect 1952 134438 2004 134444
rect 1768 133476 1820 133482
rect 1768 133418 1820 133424
rect 2056 133362 2084 138230
rect 1504 132382 1716 132410
rect 1780 133334 2084 133362
rect 1400 124772 1452 124778
rect 1400 124714 1452 124720
rect 1400 124636 1452 124642
rect 1400 124578 1452 124584
rect 1306 122088 1362 122097
rect 1306 122023 1362 122032
rect 1216 121100 1268 121106
rect 1216 121042 1268 121048
rect 1216 117564 1268 117570
rect 1216 117506 1268 117512
rect 1228 115122 1256 117506
rect 1308 116476 1360 116482
rect 1308 116418 1360 116424
rect 1216 115116 1268 115122
rect 1216 115058 1268 115064
rect 1216 110084 1268 110090
rect 1216 110026 1268 110032
rect 1228 108225 1256 110026
rect 1214 108216 1270 108225
rect 1214 108151 1270 108160
rect 1216 108112 1268 108118
rect 1216 108054 1268 108060
rect 1228 107137 1256 108054
rect 1320 107370 1348 116418
rect 1308 107364 1360 107370
rect 1308 107306 1360 107312
rect 1214 107128 1270 107137
rect 1214 107063 1270 107072
rect 1216 102604 1268 102610
rect 1216 102546 1268 102552
rect 1228 80889 1256 102546
rect 1306 99648 1362 99657
rect 1306 99583 1362 99592
rect 1320 98326 1348 99583
rect 1308 98320 1360 98326
rect 1308 98262 1360 98268
rect 1308 98184 1360 98190
rect 1308 98126 1360 98132
rect 1320 83502 1348 98126
rect 1308 83496 1360 83502
rect 1308 83438 1360 83444
rect 1214 80880 1270 80889
rect 1214 80815 1270 80824
rect 1308 72208 1360 72214
rect 1308 72150 1360 72156
rect 1216 71052 1268 71058
rect 1216 70994 1268 71000
rect 1228 65482 1256 70994
rect 1320 69358 1348 72150
rect 1308 69352 1360 69358
rect 1308 69294 1360 69300
rect 1308 67380 1360 67386
rect 1308 67322 1360 67328
rect 1216 65476 1268 65482
rect 1216 65418 1268 65424
rect 1320 65362 1348 67322
rect 1228 65334 1348 65362
rect 1228 63374 1256 65334
rect 1308 65272 1360 65278
rect 1308 65214 1360 65220
rect 1216 63368 1268 63374
rect 1216 63310 1268 63316
rect 1320 58041 1348 65214
rect 1306 58032 1362 58041
rect 1306 57967 1362 57976
rect 1308 57928 1360 57934
rect 1308 57870 1360 57876
rect 1320 45937 1348 57870
rect 1306 45928 1362 45937
rect 1306 45863 1362 45872
rect 1308 38548 1360 38554
rect 1308 38490 1360 38496
rect 1214 33280 1270 33289
rect 1214 33215 1270 33224
rect 1228 27130 1256 33215
rect 1216 27124 1268 27130
rect 1216 27066 1268 27072
rect 1214 27024 1270 27033
rect 1214 26959 1216 26968
rect 1268 26959 1270 26968
rect 1216 26930 1268 26936
rect 1214 26888 1270 26897
rect 1214 26823 1270 26832
rect 1124 16720 1176 16726
rect 1124 16662 1176 16668
rect 1124 15632 1176 15638
rect 1124 15574 1176 15580
rect 1136 14822 1164 15574
rect 1124 14816 1176 14822
rect 1124 14758 1176 14764
rect 1124 14680 1176 14686
rect 1124 14622 1176 14628
rect 1136 13054 1164 14622
rect 1124 13048 1176 13054
rect 1124 12990 1176 12996
rect 1122 12880 1178 12889
rect 1122 12815 1124 12824
rect 1176 12815 1178 12824
rect 1124 12786 1176 12792
rect 1124 12368 1176 12374
rect 1124 12310 1176 12316
rect 1136 12209 1164 12310
rect 1122 12200 1178 12209
rect 1122 12135 1178 12144
rect 1228 10418 1256 26823
rect 1320 21622 1348 38490
rect 1412 35465 1440 124578
rect 1504 39370 1532 132382
rect 1780 132002 1808 133334
rect 2240 132138 2268 138604
rect 1964 132122 2268 132138
rect 1952 132116 2268 132122
rect 2004 132110 2268 132116
rect 1952 132058 2004 132064
rect 1596 131974 1808 132002
rect 1596 126449 1624 131974
rect 2332 131866 2360 138876
rect 1688 131838 2360 131866
rect 1582 126440 1638 126449
rect 1582 126375 1638 126384
rect 1584 126268 1636 126274
rect 1584 126210 1636 126216
rect 1492 39364 1544 39370
rect 1492 39306 1544 39312
rect 1398 35456 1454 35465
rect 1398 35391 1454 35400
rect 1490 30288 1546 30297
rect 1490 30223 1546 30232
rect 1398 29744 1454 29753
rect 1398 29679 1454 29688
rect 1308 21616 1360 21622
rect 1308 21558 1360 21564
rect 1412 20194 1440 29679
rect 1504 29510 1532 30223
rect 1492 29504 1544 29510
rect 1492 29446 1544 29452
rect 1492 28008 1544 28014
rect 1492 27950 1544 27956
rect 1504 26858 1532 27950
rect 1492 26852 1544 26858
rect 1492 26794 1544 26800
rect 1490 25800 1546 25809
rect 1490 25735 1546 25744
rect 1504 24070 1532 25735
rect 1492 24064 1544 24070
rect 1492 24006 1544 24012
rect 1492 23792 1544 23798
rect 1492 23734 1544 23740
rect 1400 20188 1452 20194
rect 1400 20130 1452 20136
rect 1398 20088 1454 20097
rect 1398 20023 1454 20032
rect 1412 19990 1440 20023
rect 1400 19984 1452 19990
rect 1400 19926 1452 19932
rect 1398 19816 1454 19825
rect 1398 19751 1454 19760
rect 1308 18896 1360 18902
rect 1308 18838 1360 18844
rect 1320 12238 1348 18838
rect 1412 18766 1440 19751
rect 1400 18760 1452 18766
rect 1400 18702 1452 18708
rect 1400 18624 1452 18630
rect 1400 18566 1452 18572
rect 1412 15978 1440 18566
rect 1400 15972 1452 15978
rect 1400 15914 1452 15920
rect 1504 15858 1532 23734
rect 1412 15830 1532 15858
rect 1308 12232 1360 12238
rect 1308 12174 1360 12180
rect 1308 12096 1360 12102
rect 1308 12038 1360 12044
rect 1032 10396 1084 10402
rect 1032 10338 1084 10344
rect 1136 10390 1256 10418
rect 940 10260 992 10266
rect 940 10202 992 10208
rect 860 10118 980 10146
rect 848 7540 900 7546
rect 848 7482 900 7488
rect 756 4752 808 4758
rect 756 4694 808 4700
rect 756 3732 808 3738
rect 756 3674 808 3680
rect 768 1329 796 3674
rect 754 1320 810 1329
rect 754 1255 810 1264
rect 662 776 718 785
rect 860 746 888 7482
rect 952 1426 980 10118
rect 1032 10124 1084 10130
rect 1032 10066 1084 10072
rect 940 1420 992 1426
rect 940 1362 992 1368
rect 662 711 718 720
rect 848 740 900 746
rect 848 682 900 688
rect 386 439 442 448
rect 294 368 350 377
rect 294 303 350 312
rect 542 -960 654 480
rect 1044 474 1072 10066
rect 1136 882 1164 10390
rect 1320 10282 1348 12038
rect 1228 10254 1348 10282
rect 1228 4457 1256 10254
rect 1308 9444 1360 9450
rect 1308 9386 1360 9392
rect 1214 4448 1270 4457
rect 1214 4383 1270 4392
rect 1216 3324 1268 3330
rect 1216 3266 1268 3272
rect 1228 1057 1256 3266
rect 1214 1048 1270 1057
rect 1214 983 1270 992
rect 1124 876 1176 882
rect 1124 818 1176 824
rect 1320 678 1348 9386
rect 1308 672 1360 678
rect 1308 614 1360 620
rect 1032 468 1084 474
rect 1032 410 1084 416
rect 1412 270 1440 15830
rect 1492 15768 1544 15774
rect 1492 15710 1544 15716
rect 1504 15162 1532 15710
rect 1492 15156 1544 15162
rect 1492 15098 1544 15104
rect 1492 15020 1544 15026
rect 1492 14962 1544 14968
rect 1504 12510 1532 14962
rect 1492 12504 1544 12510
rect 1492 12446 1544 12452
rect 1596 10418 1624 126210
rect 1688 126070 1716 131838
rect 2424 131730 2452 139046
rect 1780 131702 2452 131730
rect 1780 128466 1808 131702
rect 2516 131594 2544 139828
rect 1872 131566 2544 131594
rect 1872 129282 1900 131566
rect 1952 130892 2004 130898
rect 2884 130880 2912 148022
rect 3068 142202 3096 151150
rect 3620 150770 3648 171686
rect 3436 150742 3648 150770
rect 3436 150634 3464 150742
rect 3712 150634 3740 173046
rect 3160 150606 3464 150634
rect 3528 150606 3740 150634
rect 3160 143682 3188 150606
rect 3528 150362 3556 150606
rect 3804 150362 3832 174270
rect 3252 150334 3832 150362
rect 3148 143676 3200 143682
rect 3148 143618 3200 143624
rect 3252 143534 3280 150334
rect 3528 150226 3556 150334
rect 3528 150198 3648 150226
rect 3620 143562 3648 150198
rect 3528 143534 3648 143562
rect 3252 143506 3372 143534
rect 3344 142202 3372 143506
rect 2004 130852 2912 130880
rect 2976 142174 3372 142202
rect 1952 130834 2004 130840
rect 2976 130778 3004 142174
rect 3068 138938 3096 142174
rect 3528 139754 3556 143534
rect 3344 139726 3556 139754
rect 3344 139210 3372 139726
rect 3344 139182 3464 139210
rect 3436 138938 3464 139182
rect 3068 138910 3832 138938
rect 3436 138836 3464 138910
rect 3436 138808 3556 138836
rect 3528 138530 3556 138808
rect 3528 138502 3648 138530
rect 1964 130750 3004 130778
rect 1964 130626 1992 130750
rect 1952 130620 2004 130626
rect 1952 130562 2004 130568
rect 1952 129464 2004 129470
rect 2004 129412 2912 129418
rect 1952 129406 2912 129412
rect 1964 129390 2912 129406
rect 1872 129254 2176 129282
rect 1952 129192 2004 129198
rect 2148 129180 2176 129254
rect 2884 129180 2912 129390
rect 2004 129152 2084 129180
rect 2148 129152 2820 129180
rect 2884 129152 3096 129180
rect 1952 129134 2004 129140
rect 1780 128438 1992 128466
rect 1860 128376 1912 128382
rect 1860 128318 1912 128324
rect 1768 126676 1820 126682
rect 1768 126618 1820 126624
rect 1676 126064 1728 126070
rect 1676 126006 1728 126012
rect 1780 126018 1808 126618
rect 1872 126410 1900 128318
rect 1860 126404 1912 126410
rect 1860 126346 1912 126352
rect 1964 126138 1992 128438
rect 2056 128058 2084 129152
rect 2056 128030 2360 128058
rect 1952 126132 2004 126138
rect 1952 126074 2004 126080
rect 1780 125990 2084 126018
rect 1860 124976 1912 124982
rect 1860 124918 1912 124924
rect 1952 124976 2004 124982
rect 1952 124918 2004 124924
rect 1676 124908 1728 124914
rect 1676 124850 1728 124856
rect 1688 65890 1716 124850
rect 1768 124772 1820 124778
rect 1768 124714 1820 124720
rect 1676 65884 1728 65890
rect 1676 65826 1728 65832
rect 1676 64796 1728 64802
rect 1676 64738 1728 64744
rect 1504 10390 1624 10418
rect 1504 1834 1532 10390
rect 1582 8800 1638 8809
rect 1582 8735 1584 8744
rect 1636 8735 1638 8744
rect 1584 8706 1636 8712
rect 1688 5114 1716 64738
rect 1780 29714 1808 124714
rect 1872 94790 1900 124918
rect 1964 118046 1992 124918
rect 1952 118040 2004 118046
rect 1952 117982 2004 117988
rect 2056 117858 2084 125990
rect 2332 120306 2360 128030
rect 2792 124896 2820 129152
rect 2792 124868 2912 124896
rect 2332 120278 2820 120306
rect 1964 117842 2084 117858
rect 1952 117836 2084 117842
rect 2004 117830 2084 117836
rect 1952 117778 2004 117784
rect 1952 117564 2004 117570
rect 2792 117552 2820 120278
rect 2004 117524 2820 117552
rect 1952 117506 2004 117512
rect 1952 117428 2004 117434
rect 1952 117370 2004 117376
rect 1964 111042 1992 117370
rect 1952 111036 2004 111042
rect 1952 110978 2004 110984
rect 2884 110378 2912 124868
rect 3068 124658 3096 129152
rect 3620 124964 3648 138502
rect 3528 124936 3648 124964
rect 3068 124630 3464 124658
rect 3436 117824 3464 124630
rect 2240 110350 2912 110378
rect 3252 117796 3464 117824
rect 2240 110242 2268 110350
rect 3252 110242 3280 117796
rect 3528 116906 3556 124936
rect 3804 124114 3832 138910
rect 568224 135810 568252 188006
rect 568592 187762 568620 188006
rect 568408 187734 568620 187762
rect 568408 179874 568436 187734
rect 569144 187490 569172 188278
rect 568500 187462 569172 187490
rect 568500 180010 568528 187462
rect 569328 187218 569356 188380
rect 569052 187190 569356 187218
rect 569052 180146 569080 187190
rect 569052 180118 569172 180146
rect 568500 179982 568620 180010
rect 568592 179874 568620 179982
rect 568408 179846 568528 179874
rect 568592 179846 568712 179874
rect 568500 178786 568528 179846
rect 568316 178758 568528 178786
rect 568316 163282 568344 178758
rect 568500 178486 568620 178514
rect 568500 174593 568528 178486
rect 568486 174584 568542 174593
rect 568486 174519 568542 174528
rect 568592 163282 568620 178486
rect 568684 174026 568712 179846
rect 568684 173998 569080 174026
rect 569052 166274 569080 173998
rect 569144 171986 569172 180118
rect 569222 178528 569278 178537
rect 569222 178463 569278 178472
rect 569236 172122 569264 178463
rect 569604 173482 569632 188380
rect 569696 187082 569724 188686
rect 569960 188624 570012 188630
rect 569788 188572 569960 188578
rect 569788 188566 570012 188572
rect 569788 188550 570000 188566
rect 569788 187218 569816 188550
rect 569960 188420 570012 188426
rect 569960 188362 570012 188368
rect 569788 187190 569908 187218
rect 569696 187054 569816 187082
rect 569788 174570 569816 187054
rect 569880 174978 569908 187190
rect 569972 180470 570000 188362
rect 569960 180464 570012 180470
rect 569960 180406 570012 180412
rect 569960 179852 570012 179858
rect 569960 179794 570012 179800
rect 569972 177750 570000 179794
rect 569960 177744 570012 177750
rect 569960 177686 570012 177692
rect 569960 176860 570012 176866
rect 569960 176802 570012 176808
rect 569972 175234 570000 176802
rect 569960 175228 570012 175234
rect 569960 175170 570012 175176
rect 569880 174962 570000 174978
rect 569880 174956 570012 174962
rect 569880 174950 569960 174956
rect 569960 174898 570012 174904
rect 569788 174542 570000 174570
rect 569972 173670 570000 174542
rect 569960 173664 570012 173670
rect 569960 173606 570012 173612
rect 569604 173454 569724 173482
rect 569696 172122 569724 173454
rect 569880 172230 570000 172258
rect 569880 172122 569908 172230
rect 569236 172094 569540 172122
rect 569696 172094 569908 172122
rect 569144 171958 569356 171986
rect 569328 171850 569356 171958
rect 569328 171822 569448 171850
rect 569420 170354 569448 171822
rect 569144 170326 569448 170354
rect 569144 169538 569172 170326
rect 569144 169510 569448 169538
rect 569052 166246 569356 166274
rect 568316 163254 568712 163282
rect 568592 163146 568620 163254
rect 568316 163118 568620 163146
rect 568316 153898 568344 163118
rect 568684 162330 568712 163254
rect 568592 162302 568712 162330
rect 568592 162058 568620 162302
rect 568592 162030 568896 162058
rect 568868 160970 568896 162030
rect 568776 160942 568896 160970
rect 568316 153870 568436 153898
rect 568408 147676 568436 153870
rect 568776 151722 568804 160942
rect 569328 155224 569356 166246
rect 569420 155802 569448 169510
rect 569512 169266 569540 172094
rect 569972 169386 570000 172230
rect 570064 171970 570092 191694
rect 570144 191548 570196 191554
rect 570144 191490 570196 191496
rect 570156 177342 570184 191490
rect 570248 188630 570276 191814
rect 570340 191622 570368 193559
rect 570328 191616 570380 191622
rect 570328 191558 570380 191564
rect 570236 188624 570288 188630
rect 570236 188566 570288 188572
rect 570328 177744 570380 177750
rect 570328 177686 570380 177692
rect 570144 177336 570196 177342
rect 570144 177278 570196 177284
rect 570144 173664 570196 173670
rect 570144 173606 570196 173612
rect 570052 171964 570104 171970
rect 570052 171906 570104 171912
rect 569960 169380 570012 169386
rect 569960 169322 570012 169328
rect 569512 169238 570092 169266
rect 569960 169176 570012 169182
rect 569512 169136 569960 169164
rect 569512 156210 569540 169136
rect 569960 169118 570012 169124
rect 569960 169040 570012 169046
rect 569960 168982 570012 168988
rect 569972 163962 570000 168982
rect 570064 168858 570092 169238
rect 570156 169046 570184 173606
rect 570144 169040 570196 169046
rect 570144 168982 570196 168988
rect 570064 168830 570184 168858
rect 569788 163934 570000 163962
rect 569788 157400 569816 163934
rect 569960 163736 570012 163742
rect 569880 163684 569960 163690
rect 569880 163678 570012 163684
rect 569880 163662 570000 163678
rect 569880 157536 569908 163662
rect 569960 163532 570012 163538
rect 569960 163474 570012 163480
rect 569972 157894 570000 163474
rect 570052 162036 570104 162042
rect 570052 161978 570104 161984
rect 569960 157888 570012 157894
rect 569960 157830 570012 157836
rect 569960 157548 570012 157554
rect 569880 157508 569960 157536
rect 569960 157490 570012 157496
rect 569960 157412 570012 157418
rect 569788 157372 569960 157400
rect 569960 157354 570012 157360
rect 569512 156182 570000 156210
rect 569972 155922 570000 156182
rect 569960 155916 570012 155922
rect 569960 155858 570012 155864
rect 569420 155774 570000 155802
rect 569972 155242 570000 155774
rect 570064 155650 570092 161978
rect 570156 157690 570184 168830
rect 570144 157684 570196 157690
rect 570144 157626 570196 157632
rect 570144 157548 570196 157554
rect 570144 157490 570196 157496
rect 570052 155644 570104 155650
rect 570052 155586 570104 155592
rect 569960 155236 570012 155242
rect 569328 155196 569816 155224
rect 569788 155156 569816 155196
rect 569960 155178 570012 155184
rect 569868 155168 569920 155174
rect 569788 155128 569868 155156
rect 569420 155094 569632 155122
rect 569868 155110 569920 155116
rect 569420 151722 569448 155094
rect 569604 155020 569632 155094
rect 570052 155100 570104 155106
rect 570052 155042 570104 155048
rect 569960 155032 570012 155038
rect 569604 154992 569960 155020
rect 569960 154974 570012 154980
rect 569960 154896 570012 154902
rect 568684 151694 568804 151722
rect 568868 151694 569448 151722
rect 569512 154856 569960 154884
rect 568408 147648 568620 147676
rect 568592 146554 568620 147648
rect 568500 146526 568620 146554
rect 568500 143426 568528 146526
rect 568684 143970 568712 151694
rect 568868 151586 568896 151694
rect 568408 143398 568528 143426
rect 568592 143942 568712 143970
rect 568776 151558 568896 151586
rect 568408 139482 568436 143398
rect 568592 139618 568620 143942
rect 568592 139590 568712 139618
rect 568408 139454 568620 139482
rect 568224 135782 568436 135810
rect 2056 110214 2268 110242
rect 2332 110214 3280 110242
rect 3344 116878 3556 116906
rect 3620 124086 3832 124114
rect 2056 110106 2084 110214
rect 1964 110090 2084 110106
rect 1952 110084 2084 110090
rect 2004 110078 2084 110084
rect 1952 110026 2004 110032
rect 1952 109744 2004 109750
rect 2332 109732 2360 110214
rect 3344 109970 3372 116878
rect 3620 114594 3648 124086
rect 568408 121530 568436 135782
rect 568316 121502 568436 121530
rect 3620 114566 3740 114594
rect 3068 109942 3372 109970
rect 2004 109704 2360 109732
rect 2424 109772 2728 109800
rect 1952 109686 2004 109692
rect 2424 109562 2452 109772
rect 1964 109534 2452 109562
rect 2700 109562 2728 109772
rect 3068 109562 3096 109942
rect 3712 109800 3740 114566
rect 3712 109772 3832 109800
rect 2700 109534 3096 109562
rect 1964 109478 1992 109534
rect 1952 109472 2004 109478
rect 1952 109414 2004 109420
rect 2516 109398 3740 109426
rect 1952 109336 2004 109342
rect 2516 109324 2544 109398
rect 2004 109296 2544 109324
rect 1952 109278 2004 109284
rect 2700 109262 3372 109290
rect 1952 109200 2004 109206
rect 2700 109154 2728 109262
rect 2004 109148 2728 109154
rect 1952 109142 2728 109148
rect 1964 109126 2728 109142
rect 1952 108928 2004 108934
rect 3344 108882 3372 109262
rect 2004 108876 3280 108882
rect 1952 108870 3280 108876
rect 1964 108854 3280 108870
rect 3344 108854 3464 108882
rect 1952 108792 2004 108798
rect 3252 108746 3280 108854
rect 2004 108740 3096 108746
rect 1952 108734 3096 108740
rect 1964 108718 3096 108734
rect 3252 108718 3372 108746
rect 1952 108656 2004 108662
rect 2004 108604 2912 108610
rect 1952 108598 2912 108604
rect 1964 108582 2912 108598
rect 1952 108520 2004 108526
rect 2004 108468 2820 108474
rect 1952 108462 2820 108468
rect 1964 108446 2820 108462
rect 1952 108384 2004 108390
rect 2004 108344 2728 108372
rect 1952 108326 2004 108332
rect 1952 108112 2004 108118
rect 2004 108060 2636 108066
rect 1952 108054 2636 108060
rect 1964 108038 2636 108054
rect 1952 107704 2004 107710
rect 2004 107664 2360 107692
rect 1952 107646 2004 107652
rect 1952 107364 2004 107370
rect 2004 107324 2268 107352
rect 1952 107306 2004 107312
rect 1952 107228 2004 107234
rect 2004 107188 2176 107216
rect 1952 107170 2004 107176
rect 1952 107092 2004 107098
rect 1952 107034 2004 107040
rect 1964 98462 1992 107034
rect 2148 103578 2176 107188
rect 2056 103550 2176 103578
rect 1952 98456 2004 98462
rect 1952 98398 2004 98404
rect 1952 98320 2004 98326
rect 2056 98308 2084 103550
rect 2240 103442 2268 107324
rect 2004 98280 2084 98308
rect 2148 103414 2268 103442
rect 1952 98262 2004 98268
rect 1952 98184 2004 98190
rect 2148 98172 2176 103414
rect 2004 98144 2176 98172
rect 1952 98126 2004 98132
rect 1860 94784 1912 94790
rect 1860 94726 1912 94732
rect 1952 94716 2004 94722
rect 2332 94704 2360 107664
rect 2004 94676 2360 94704
rect 1952 94658 2004 94664
rect 1952 94036 2004 94042
rect 2608 94024 2636 108038
rect 2004 93996 2636 94024
rect 1952 93978 2004 93984
rect 1952 93628 2004 93634
rect 2700 93616 2728 108344
rect 2004 93588 2728 93616
rect 1952 93570 2004 93576
rect 2792 93514 2820 108446
rect 1872 93498 2820 93514
rect 1860 93492 2820 93498
rect 1912 93486 2820 93492
rect 1860 93434 1912 93440
rect 1952 93424 2004 93430
rect 2884 93412 2912 108582
rect 3068 105618 3096 108718
rect 3068 105590 3280 105618
rect 3252 100722 3280 105590
rect 2004 93384 2912 93412
rect 3068 100694 3280 100722
rect 1952 93366 2004 93372
rect 1860 93288 1912 93294
rect 1860 93230 1912 93236
rect 1952 93288 2004 93294
rect 2004 93248 2820 93276
rect 1952 93230 2004 93236
rect 1872 86358 1900 93230
rect 1952 92200 2004 92206
rect 2792 92188 2820 93248
rect 2004 92160 2820 92188
rect 1952 92142 2004 92148
rect 1952 92064 2004 92070
rect 3068 92018 3096 100694
rect 2004 92012 3096 92018
rect 1952 92006 3096 92012
rect 1964 91990 3096 92006
rect 1952 91928 2004 91934
rect 2004 91876 2820 91882
rect 1952 91870 2820 91876
rect 1964 91854 2820 91870
rect 1952 91792 2004 91798
rect 2004 91752 2728 91780
rect 1952 91734 2004 91740
rect 1952 91656 2004 91662
rect 2004 91616 2636 91644
rect 1952 91598 2004 91604
rect 1952 91520 2004 91526
rect 2004 91480 2360 91508
rect 1952 91462 2004 91468
rect 1952 91384 2004 91390
rect 2004 91332 2084 91338
rect 1952 91326 2084 91332
rect 1964 91310 2084 91326
rect 1952 91248 2004 91254
rect 1952 91190 2004 91196
rect 1964 86426 1992 91190
rect 1952 86420 2004 86426
rect 1952 86362 2004 86368
rect 1860 86352 1912 86358
rect 2056 86306 2084 91310
rect 1860 86294 1912 86300
rect 1964 86278 2084 86306
rect 1964 86222 1992 86278
rect 1952 86216 2004 86222
rect 1952 86158 2004 86164
rect 1860 86148 1912 86154
rect 1860 86090 1912 86096
rect 1872 83722 1900 86090
rect 2332 84946 2360 91480
rect 1964 84918 2360 84946
rect 1964 84794 1992 84918
rect 1952 84788 2004 84794
rect 1952 84730 2004 84736
rect 2608 84674 2636 91616
rect 1964 84658 2636 84674
rect 1952 84652 2636 84658
rect 2004 84646 2636 84652
rect 1952 84594 2004 84600
rect 1952 83836 2004 83842
rect 2700 83824 2728 91752
rect 2792 83994 2820 91854
rect 3344 89706 3372 108718
rect 2976 89678 3372 89706
rect 2976 84130 3004 89678
rect 3436 88210 3464 108854
rect 3514 96112 3570 96121
rect 3514 96047 3570 96056
rect 3068 88182 3464 88210
rect 3068 84266 3096 88182
rect 3528 87802 3556 96047
rect 3712 94874 3740 109398
rect 3804 94874 3832 109772
rect 568316 98682 568344 121502
rect 568224 98654 568344 98682
rect 568224 96370 568252 98654
rect 568592 97050 568620 139454
rect 568408 97022 568620 97050
rect 568224 96342 568344 96370
rect 3436 87774 3556 87802
rect 3620 94846 3832 94874
rect 3068 84238 3280 84266
rect 2976 84102 3188 84130
rect 2792 83966 3004 83994
rect 2004 83796 2728 83824
rect 1952 83778 2004 83784
rect 1872 83694 2912 83722
rect 1952 83632 2004 83638
rect 2004 83580 2820 83586
rect 1952 83574 2820 83580
rect 1964 83558 2820 83574
rect 1860 83496 1912 83502
rect 1860 83438 1912 83444
rect 1872 72622 1900 83438
rect 2792 82634 2820 83558
rect 2332 82606 2820 82634
rect 1952 82136 2004 82142
rect 2004 82084 2084 82090
rect 1952 82078 2084 82084
rect 1964 82062 2084 82078
rect 1952 80776 2004 80782
rect 1952 80718 2004 80724
rect 1860 72616 1912 72622
rect 1860 72558 1912 72564
rect 1860 72480 1912 72486
rect 1860 72422 1912 72428
rect 1872 38554 1900 72422
rect 1964 72214 1992 80718
rect 1952 72208 2004 72214
rect 1952 72150 2004 72156
rect 2056 72026 2084 82062
rect 1964 72010 2084 72026
rect 1952 72004 2084 72010
rect 2004 71998 2084 72004
rect 1952 71946 2004 71952
rect 2332 71074 2360 82606
rect 2884 82498 2912 83694
rect 1964 71058 2360 71074
rect 1952 71052 2360 71058
rect 2004 71046 2360 71052
rect 2516 82470 2912 82498
rect 1952 70994 2004 71000
rect 2516 67674 2544 82470
rect 2976 78826 3004 83966
rect 3160 83858 3188 84102
rect 3252 83994 3280 84238
rect 3252 83966 3372 83994
rect 3160 83830 3280 83858
rect 2608 78798 3004 78826
rect 2608 76106 2636 78798
rect 3252 77466 3280 83830
rect 3344 83042 3372 83966
rect 3436 83586 3464 87774
rect 3620 84946 3648 94846
rect 3712 90386 3740 94846
rect 3712 90358 3832 90386
rect 3528 84918 3648 84946
rect 3528 83586 3556 84918
rect 3436 83558 3648 83586
rect 3344 83014 3464 83042
rect 2976 77438 3280 77466
rect 2608 76078 2912 76106
rect 2884 75562 2912 76078
rect 2976 75562 3004 77438
rect 3436 77058 3464 83014
rect 2700 75534 3004 75562
rect 3068 77030 3464 77058
rect 2700 71992 2728 75534
rect 2056 67646 2544 67674
rect 2608 71964 2728 71992
rect 2056 67538 2084 67646
rect 1964 67522 2084 67538
rect 1952 67516 2084 67522
rect 2004 67510 2084 67516
rect 1952 67458 2004 67464
rect 2608 67402 2636 71964
rect 2884 71890 2912 75534
rect 1964 67386 2636 67402
rect 1952 67380 2636 67386
rect 2004 67374 2636 67380
rect 2700 71862 2912 71890
rect 1952 67322 2004 67328
rect 2700 67266 2728 71862
rect 1964 67250 2728 67266
rect 1952 67244 2728 67250
rect 2004 67238 2728 67244
rect 1952 67186 2004 67192
rect 1952 66768 2004 66774
rect 2004 66728 2728 66756
rect 1952 66710 2004 66716
rect 1952 66632 2004 66638
rect 2004 66580 2636 66586
rect 1952 66574 2636 66580
rect 1964 66558 2636 66574
rect 1952 66496 2004 66502
rect 1952 66438 2004 66444
rect 1964 64802 1992 66438
rect 2608 66314 2636 66558
rect 2700 66450 2728 66728
rect 3068 66722 3096 77030
rect 3528 73114 3556 83558
rect 3436 73086 3556 73114
rect 3436 69034 3464 73086
rect 2976 66694 3096 66722
rect 3344 69006 3464 69034
rect 2976 66450 3004 66694
rect 2700 66422 3004 66450
rect 3344 66314 3372 69006
rect 2608 66286 3372 66314
rect 2044 65476 2096 65482
rect 2044 65418 2096 65424
rect 2056 64954 2084 65418
rect 3620 64954 3648 83558
rect 3804 75426 3832 90358
rect 568316 77194 568344 96342
rect 568408 93922 568436 97022
rect 568684 96642 568712 139590
rect 568592 96614 568712 96642
rect 568592 96098 568620 96614
rect 568776 96540 568804 151558
rect 569512 151314 569540 154856
rect 569960 154838 570012 154844
rect 570064 154204 570092 155042
rect 568500 96070 568620 96098
rect 568684 96512 568804 96540
rect 568868 151286 569540 151314
rect 569880 154176 570092 154204
rect 568500 95146 568528 96070
rect 568500 95118 568620 95146
rect 568408 93894 568528 93922
rect 568500 85626 568528 93894
rect 568592 87530 568620 95118
rect 568684 87802 568712 96512
rect 568684 87774 568804 87802
rect 568592 87502 568712 87530
rect 568500 85598 568620 85626
rect 568316 77166 568528 77194
rect 3712 75398 3832 75426
rect 3712 74882 3740 75398
rect 3712 74854 3832 74882
rect 2056 64926 3648 64954
rect 3804 64818 3832 74854
rect 568500 73148 568528 77166
rect 1952 64796 2004 64802
rect 1952 64738 2004 64744
rect 3620 64790 3832 64818
rect 568316 73120 568528 73148
rect 1952 64660 2004 64666
rect 2004 64620 3004 64648
rect 1952 64602 2004 64608
rect 1952 63368 2004 63374
rect 2004 63316 2820 63322
rect 1952 63310 2820 63316
rect 1964 63294 2820 63310
rect 1952 63164 2004 63170
rect 2004 63124 2728 63152
rect 1952 63106 2004 63112
rect 1952 63028 2004 63034
rect 2004 62988 2452 63016
rect 1952 62970 2004 62976
rect 1952 62892 2004 62898
rect 1952 62834 2004 62840
rect 1964 62778 1992 62834
rect 1964 62750 2268 62778
rect 1952 62280 2004 62286
rect 2004 62240 2176 62268
rect 1952 62222 2004 62228
rect 1952 57112 2004 57118
rect 2148 57100 2176 62240
rect 2004 57072 2176 57100
rect 1952 57054 2004 57060
rect 1952 56908 2004 56914
rect 2240 56896 2268 62750
rect 2004 56868 2268 56896
rect 1952 56850 2004 56856
rect 1952 56772 2004 56778
rect 2004 56732 2084 56760
rect 1952 56714 2004 56720
rect 2056 56658 2084 56732
rect 2424 56658 2452 62988
rect 1952 56636 2004 56642
rect 2056 56630 2452 56658
rect 1952 56578 2004 56584
rect 1964 55978 1992 56578
rect 1964 55950 2636 55978
rect 1952 55888 2004 55894
rect 2004 55848 2544 55876
rect 1952 55830 2004 55836
rect 1952 55208 2004 55214
rect 2004 55156 2452 55162
rect 1952 55150 2452 55156
rect 1964 55134 2452 55150
rect 1952 52760 2004 52766
rect 2004 52720 2084 52748
rect 1952 52702 2004 52708
rect 1952 52624 2004 52630
rect 1952 52566 2004 52572
rect 1964 43194 1992 52566
rect 2056 51490 2084 52720
rect 2056 51462 2176 51490
rect 2148 43466 2176 51462
rect 2424 43466 2452 55134
rect 2516 43602 2544 55848
rect 2608 43738 2636 55950
rect 2700 44554 2728 63124
rect 2792 63016 2820 63294
rect 2976 63152 3004 64620
rect 2976 63124 3556 63152
rect 2792 62988 3188 63016
rect 3160 51082 3188 62988
rect 3528 51082 3556 63124
rect 3620 56522 3648 64790
rect 3620 56494 3740 56522
rect 2792 51054 3188 51082
rect 3344 51054 3556 51082
rect 2792 44826 2820 51054
rect 3344 50810 3372 51054
rect 3712 50946 3740 56494
rect 3712 50918 3832 50946
rect 3344 50782 3556 50810
rect 2792 44798 3280 44826
rect 2700 44526 3096 44554
rect 2608 43710 2820 43738
rect 2792 43602 2820 43710
rect 2516 43574 2636 43602
rect 2792 43574 2912 43602
rect 2608 43466 2636 43574
rect 2148 43438 2360 43466
rect 2424 43438 2544 43466
rect 2608 43438 2820 43466
rect 2332 43194 2360 43438
rect 2516 43330 2544 43438
rect 2516 43302 2728 43330
rect 1964 43166 2176 43194
rect 2332 43166 2636 43194
rect 1952 43104 2004 43110
rect 1952 43046 2004 43052
rect 2148 43058 2176 43166
rect 1964 42922 1992 43046
rect 2148 43030 2544 43058
rect 1964 42894 2176 42922
rect 1952 42832 2004 42838
rect 2004 42780 2084 42786
rect 1952 42774 2084 42780
rect 1964 42758 2084 42774
rect 2056 39522 2084 42758
rect 1964 39506 2084 39522
rect 1952 39500 2084 39506
rect 2004 39494 2084 39500
rect 1952 39442 2004 39448
rect 2148 39386 2176 42894
rect 1964 39370 2176 39386
rect 1952 39364 2176 39370
rect 2004 39358 2176 39364
rect 1952 39306 2004 39312
rect 1952 39228 2004 39234
rect 1952 39170 2004 39176
rect 1964 39114 1992 39170
rect 1964 39086 2452 39114
rect 1860 38548 1912 38554
rect 1860 38490 1912 38496
rect 2424 35714 2452 39086
rect 1964 35698 2452 35714
rect 1952 35692 2452 35698
rect 2004 35686 2452 35692
rect 1952 35634 2004 35640
rect 2516 35578 2544 43030
rect 1964 35562 2544 35578
rect 1952 35556 2544 35562
rect 2004 35550 2544 35556
rect 1952 35498 2004 35504
rect 2608 35442 2636 43166
rect 1964 35426 2636 35442
rect 1952 35420 2636 35426
rect 2004 35414 2636 35420
rect 1952 35362 2004 35368
rect 2700 35306 2728 43302
rect 1964 35290 2728 35306
rect 1952 35284 2728 35290
rect 2004 35278 2728 35284
rect 1952 35226 2004 35232
rect 2792 34626 2820 43438
rect 1872 34598 2820 34626
rect 1872 29782 1900 34598
rect 2884 29866 2912 43574
rect 3068 40474 3096 44526
rect 3252 40610 3280 44798
rect 3528 42786 3556 50782
rect 3528 42758 3648 42786
rect 3620 40746 3648 42758
rect 3804 40746 3832 50918
rect 3436 40718 3832 40746
rect 3436 40610 3464 40718
rect 3620 40610 3648 40718
rect 3252 40582 3740 40610
rect 3068 40446 3372 40474
rect 3344 35680 3372 40446
rect 2056 29838 2912 29866
rect 3068 35652 3372 35680
rect 1860 29776 1912 29782
rect 1860 29718 1912 29724
rect 1768 29708 1820 29714
rect 1768 29650 1820 29656
rect 1768 29572 1820 29578
rect 1768 29514 1820 29520
rect 1780 15026 1808 29514
rect 2056 28370 2084 29838
rect 1964 28354 2084 28370
rect 1952 28348 2084 28354
rect 2004 28342 2084 28348
rect 1952 28290 2004 28296
rect 3068 28098 3096 35652
rect 3436 35544 3464 40582
rect 3620 40066 3648 40582
rect 3528 40038 3648 40066
rect 3528 37210 3556 40038
rect 3528 37182 3648 37210
rect 1964 28070 3096 28098
rect 3252 35516 3464 35544
rect 1964 28014 1992 28070
rect 1952 28008 2004 28014
rect 1952 27950 2004 27956
rect 3252 27826 3280 35516
rect 3620 35408 3648 37182
rect 1872 27798 3280 27826
rect 3436 35380 3648 35408
rect 1872 23746 1900 27798
rect 3436 27690 3464 35380
rect 3712 33810 3740 40582
rect 3790 40352 3846 40361
rect 3790 40287 3846 40296
rect 3344 27662 3464 27690
rect 3620 33782 3740 33810
rect 3344 27282 3372 27662
rect 1964 27266 3372 27282
rect 1952 27260 3372 27266
rect 2004 27254 3372 27260
rect 1952 27202 2004 27208
rect 1952 27124 2004 27130
rect 2004 27084 3096 27112
rect 1952 27066 2004 27072
rect 1952 26988 2004 26994
rect 2004 26948 2820 26976
rect 1952 26930 2004 26936
rect 2792 26874 2820 26948
rect 1952 26852 2004 26858
rect 2792 26846 2912 26874
rect 1952 26794 2004 26800
rect 1964 26738 1992 26794
rect 1964 26710 2820 26738
rect 1872 23718 2544 23746
rect 1952 22228 2004 22234
rect 2004 22188 2268 22216
rect 1952 22170 2004 22176
rect 1952 22092 2004 22098
rect 1952 22034 2004 22040
rect 1964 19666 1992 22034
rect 1964 19638 2084 19666
rect 2056 18578 2084 19638
rect 1964 18550 2084 18578
rect 1964 18494 1992 18550
rect 1952 18488 2004 18494
rect 1952 18430 2004 18436
rect 2240 18034 2268 22188
rect 1872 18006 2268 18034
rect 1872 17950 1900 18006
rect 1860 17944 1912 17950
rect 1860 17886 1912 17892
rect 1860 16584 1912 16590
rect 2516 16538 2544 23718
rect 2792 21570 2820 26710
rect 2700 21542 2820 21570
rect 2700 17626 2728 21542
rect 2700 17598 2820 17626
rect 1912 16532 2544 16538
rect 1860 16526 2544 16532
rect 1872 16510 2544 16526
rect 1860 16448 1912 16454
rect 1912 16396 2084 16402
rect 1860 16390 2084 16396
rect 1872 16374 2084 16390
rect 1952 16312 2004 16318
rect 1952 16254 2004 16260
rect 2056 16266 2084 16374
rect 2792 16266 2820 17598
rect 1860 16108 1912 16114
rect 1860 16050 1912 16056
rect 1768 15020 1820 15026
rect 1768 14962 1820 14968
rect 1872 14906 1900 16050
rect 1964 15774 1992 16254
rect 2056 16238 2820 16266
rect 2884 16096 2912 26846
rect 3068 16674 3096 27084
rect 3620 16674 3648 33782
rect 2608 16068 2912 16096
rect 2976 16646 3648 16674
rect 2608 15960 2636 16068
rect 2976 15960 3004 16646
rect 3068 16572 3096 16646
rect 3068 16544 3740 16572
rect 2056 15932 3004 15960
rect 1952 15768 2004 15774
rect 1952 15710 2004 15716
rect 1952 15632 2004 15638
rect 2056 15620 2084 15932
rect 2608 15858 2636 15932
rect 2608 15830 3648 15858
rect 2004 15592 2084 15620
rect 1952 15574 2004 15580
rect 1952 15496 2004 15502
rect 2004 15456 2360 15484
rect 1952 15438 2004 15444
rect 1952 15360 2004 15366
rect 2004 15320 2176 15348
rect 1952 15302 2004 15308
rect 1952 15156 2004 15162
rect 1952 15098 2004 15104
rect 1596 5086 1716 5114
rect 1780 14878 1900 14906
rect 1492 1828 1544 1834
rect 1492 1770 1544 1776
rect 1492 1692 1544 1698
rect 1492 1634 1544 1640
rect 1504 1465 1532 1634
rect 1596 1494 1624 5086
rect 1676 1760 1728 1766
rect 1676 1702 1728 1708
rect 1584 1488 1636 1494
rect 1490 1456 1546 1465
rect 1584 1430 1636 1436
rect 1490 1391 1546 1400
rect 1688 480 1716 1702
rect 1780 921 1808 14878
rect 1860 14816 1912 14822
rect 1860 14758 1912 14764
rect 1872 12594 1900 14758
rect 1964 13530 1992 15098
rect 2148 15008 2176 15320
rect 2332 15144 2360 15456
rect 2332 15116 3556 15144
rect 2148 14980 3464 15008
rect 1952 13524 2004 13530
rect 1952 13466 2004 13472
rect 1952 13388 2004 13394
rect 2004 13348 3372 13376
rect 1952 13330 2004 13336
rect 1952 13048 2004 13054
rect 2004 13008 3280 13036
rect 1952 12990 2004 12996
rect 1952 12844 2004 12850
rect 2004 12804 3188 12832
rect 1952 12786 2004 12792
rect 1872 12566 3096 12594
rect 1952 12504 2004 12510
rect 2004 12464 3004 12492
rect 1952 12446 2004 12452
rect 1952 4752 2004 4758
rect 1952 4694 2004 4700
rect 1860 3732 1912 3738
rect 1860 3674 1912 3680
rect 1872 1601 1900 3674
rect 1858 1592 1914 1601
rect 1858 1527 1914 1536
rect 1766 912 1822 921
rect 1766 847 1822 856
rect 1400 264 1452 270
rect 1400 206 1452 212
rect 1646 -960 1758 480
rect 1964 377 1992 4694
rect 2976 1698 3004 12464
rect 2964 1692 3016 1698
rect 2964 1634 3016 1640
rect 3068 814 3096 12566
rect 3160 1290 3188 12804
rect 3148 1284 3200 1290
rect 3148 1226 3200 1232
rect 3252 1018 3280 13008
rect 3240 1012 3292 1018
rect 3240 954 3292 960
rect 3344 950 3372 13348
rect 3332 944 3384 950
rect 3332 886 3384 892
rect 3056 808 3108 814
rect 3056 750 3108 756
rect 2884 564 3096 592
rect 2884 480 2912 564
rect 1950 368 2006 377
rect 1950 303 2006 312
rect 2842 -960 2954 480
rect 3068 202 3096 564
rect 3436 241 3464 14980
rect 3528 1494 3556 15116
rect 3516 1488 3568 1494
rect 3516 1430 3568 1436
rect 3620 542 3648 15830
rect 3712 1465 3740 16544
rect 3804 1766 3832 40287
rect 568316 40032 568344 73120
rect 568592 55298 568620 85598
rect 568684 64410 568712 87502
rect 568776 64546 568804 87774
rect 568868 73522 568896 151286
rect 569880 151178 569908 154176
rect 570052 153944 570104 153950
rect 570052 153886 570104 153892
rect 569960 153876 570012 153882
rect 569960 153818 570012 153824
rect 569144 151150 569908 151178
rect 569144 146996 569172 151150
rect 569972 149444 570000 153818
rect 570064 149598 570092 153886
rect 570052 149592 570104 149598
rect 570052 149534 570104 149540
rect 568960 146968 569172 146996
rect 569236 149416 570000 149444
rect 570052 149456 570104 149462
rect 568960 73658 568988 146968
rect 569236 142100 569264 149416
rect 570052 149398 570104 149404
rect 569960 149320 570012 149326
rect 569960 149262 570012 149268
rect 569972 148510 570000 149262
rect 569960 148504 570012 148510
rect 569960 148446 570012 148452
rect 570064 148374 570092 149398
rect 570052 148368 570104 148374
rect 570052 148310 570104 148316
rect 569960 147960 570012 147966
rect 569512 147920 569960 147948
rect 569512 142746 569540 147920
rect 569960 147902 570012 147908
rect 570156 147830 570184 157490
rect 570236 155780 570288 155786
rect 570236 155722 570288 155728
rect 570248 153882 570276 155722
rect 570236 153876 570288 153882
rect 570236 153818 570288 153824
rect 570236 153468 570288 153474
rect 570236 153410 570288 153416
rect 570248 149308 570276 153410
rect 570340 149462 570368 177686
rect 570420 162240 570472 162246
rect 570420 162182 570472 162188
rect 570328 149456 570380 149462
rect 570328 149398 570380 149404
rect 570248 149280 570368 149308
rect 570236 149116 570288 149122
rect 570236 149058 570288 149064
rect 569960 147824 570012 147830
rect 569420 142718 569540 142746
rect 569604 147784 569960 147812
rect 569420 142338 569448 142718
rect 569052 142072 569264 142100
rect 569328 142310 569448 142338
rect 569052 74066 569080 142072
rect 569328 138802 569356 142310
rect 569604 142236 569632 147784
rect 569960 147766 570012 147772
rect 570144 147824 570196 147830
rect 570144 147766 570196 147772
rect 569960 147688 570012 147694
rect 569144 138774 569356 138802
rect 569420 142208 569632 142236
rect 569696 147648 569960 147676
rect 569144 76106 569172 138774
rect 569420 138666 569448 142208
rect 569696 142100 569724 147648
rect 569960 147630 570012 147636
rect 569960 147008 570012 147014
rect 569236 138638 569448 138666
rect 569604 142072 569724 142100
rect 569788 146968 569960 146996
rect 569236 76242 569264 138638
rect 569604 138258 569632 142072
rect 569788 139482 569816 146968
rect 569960 146950 570012 146956
rect 569960 144288 570012 144294
rect 569328 138230 569632 138258
rect 569696 139454 569816 139482
rect 569880 144236 569960 144242
rect 569880 144230 570012 144236
rect 569880 144214 570000 144230
rect 569328 76344 569356 138230
rect 569696 135640 569724 139454
rect 569880 135810 569908 144214
rect 569880 135782 570092 135810
rect 569696 135612 569908 135640
rect 569880 134994 569908 135612
rect 569880 134978 570000 134994
rect 569880 134972 570012 134978
rect 569880 134966 569960 134972
rect 569960 134914 570012 134920
rect 570064 134858 570092 135782
rect 569788 134830 570092 134858
rect 569788 134722 569816 134830
rect 569420 134694 569816 134722
rect 569960 134768 570012 134774
rect 569960 134710 570012 134716
rect 569420 76480 569448 134694
rect 569972 134450 570000 134710
rect 570052 134564 570104 134570
rect 570052 134506 570104 134512
rect 569512 134422 570000 134450
rect 569512 76616 569540 134422
rect 569960 134360 570012 134366
rect 569604 134308 569960 134314
rect 569604 134302 570012 134308
rect 569604 134286 570000 134302
rect 569604 76752 569632 134286
rect 569960 134224 570012 134230
rect 569696 134184 569960 134212
rect 569696 77058 569724 134184
rect 569960 134166 570012 134172
rect 569960 133136 570012 133142
rect 569788 133084 569960 133090
rect 569788 133078 570012 133084
rect 569788 133062 570000 133078
rect 569788 77194 569816 133062
rect 570064 104258 570092 134506
rect 570248 134366 570276 149058
rect 570340 144294 570368 149280
rect 570432 149122 570460 162182
rect 574756 150657 574784 251194
rect 574848 232257 574876 391954
rect 580170 346080 580226 346089
rect 580170 346015 580226 346024
rect 580184 345098 580212 346015
rect 574928 345092 574980 345098
rect 574928 345034 574980 345040
rect 580172 345092 580224 345098
rect 580172 345034 580224 345040
rect 574834 232248 574890 232257
rect 574834 232183 574890 232192
rect 574940 205057 574968 345034
rect 580170 299160 580226 299169
rect 580170 299095 580226 299104
rect 580184 298178 580212 299095
rect 575020 298172 575072 298178
rect 575020 298114 575072 298120
rect 580172 298172 580224 298178
rect 580172 298114 580224 298120
rect 574926 205048 574982 205057
rect 574926 204983 574982 204992
rect 574836 204332 574888 204338
rect 574836 204274 574888 204280
rect 574742 150648 574798 150657
rect 574742 150583 574798 150592
rect 570420 149116 570472 149122
rect 570420 149058 570472 149064
rect 570328 144288 570380 144294
rect 570328 144230 570380 144236
rect 570236 134360 570288 134366
rect 570236 134302 570288 134308
rect 574848 124098 574876 204274
rect 575032 177857 575060 298114
rect 580170 252240 580226 252249
rect 580170 252175 580226 252184
rect 580184 251258 580212 252175
rect 580172 251252 580224 251258
rect 580172 251194 580224 251200
rect 580170 205320 580226 205329
rect 580170 205255 580226 205264
rect 580184 204338 580212 205255
rect 580172 204332 580224 204338
rect 580172 204274 580224 204280
rect 575018 177848 575074 177857
rect 575018 177783 575074 177792
rect 580170 158400 580226 158409
rect 580170 158335 580226 158344
rect 580184 157418 580212 158335
rect 574928 157412 574980 157418
rect 574928 157354 574980 157360
rect 580172 157412 580224 157418
rect 580172 157354 580224 157360
rect 572720 124092 572772 124098
rect 572720 124034 572772 124040
rect 574836 124092 574888 124098
rect 574836 124034 574888 124040
rect 572732 123457 572760 124034
rect 572718 123448 572774 123457
rect 572718 123383 572774 123392
rect 574744 110492 574796 110498
rect 574744 110434 574796 110440
rect 569880 104230 570092 104258
rect 569880 77296 569908 104230
rect 570326 99376 570382 99385
rect 570326 99311 570382 99320
rect 570340 90137 570368 99311
rect 572720 96552 572772 96558
rect 572720 96494 572772 96500
rect 572732 96257 572760 96494
rect 572718 96248 572774 96257
rect 572718 96183 572774 96192
rect 570326 90128 570382 90137
rect 570326 90063 570382 90072
rect 569960 77308 570012 77314
rect 569880 77268 569960 77296
rect 569960 77250 570012 77256
rect 569788 77166 570092 77194
rect 569696 77030 569816 77058
rect 569788 76786 569816 77030
rect 569788 76770 570000 76786
rect 569788 76764 570012 76770
rect 569788 76758 569960 76764
rect 569604 76724 569724 76752
rect 569696 76616 569724 76724
rect 569960 76706 570012 76712
rect 569880 76634 570000 76650
rect 569880 76628 570012 76634
rect 569880 76622 569960 76628
rect 569880 76616 569908 76622
rect 569512 76588 569632 76616
rect 569696 76588 569908 76616
rect 569604 76514 569632 76588
rect 569960 76570 570012 76576
rect 569604 76498 570000 76514
rect 569604 76492 570012 76498
rect 569604 76486 569960 76492
rect 569420 76452 569540 76480
rect 569512 76344 569540 76452
rect 569960 76434 570012 76440
rect 569788 76362 570000 76378
rect 569788 76356 570012 76362
rect 569788 76350 569960 76356
rect 569788 76344 569816 76350
rect 569328 76316 569448 76344
rect 569512 76316 569816 76344
rect 569420 76242 569448 76316
rect 569960 76298 570012 76304
rect 569236 76214 569356 76242
rect 569420 76226 570000 76242
rect 569420 76220 570012 76226
rect 569420 76214 569960 76220
rect 569328 76106 569356 76214
rect 569960 76162 570012 76168
rect 569144 76078 569264 76106
rect 569328 76078 569448 76106
rect 569236 75970 569264 76078
rect 569236 75942 569356 75970
rect 569328 74712 569356 75942
rect 569420 74848 569448 76078
rect 569960 74860 570012 74866
rect 569420 74820 569960 74848
rect 569960 74802 570012 74808
rect 569960 74724 570012 74730
rect 569328 74684 569960 74712
rect 569960 74666 570012 74672
rect 569052 74038 570000 74066
rect 569972 73778 570000 74038
rect 569960 73772 570012 73778
rect 569960 73714 570012 73720
rect 568960 73642 570000 73658
rect 568960 73636 570012 73642
rect 568960 73630 569960 73636
rect 569960 73578 570012 73584
rect 568868 73494 570000 73522
rect 569972 73438 570000 73494
rect 569960 73432 570012 73438
rect 568960 73358 569724 73386
rect 569960 73374 570012 73380
rect 568960 64682 568988 73358
rect 569696 73284 569724 73358
rect 569960 73296 570012 73302
rect 569696 73256 569960 73284
rect 569052 73222 569448 73250
rect 569960 73238 570012 73244
rect 569052 64818 569080 73222
rect 569420 73148 569448 73222
rect 569960 73160 570012 73166
rect 569420 73120 569960 73148
rect 569960 73102 570012 73108
rect 569960 73024 570012 73030
rect 569604 72984 569960 73012
rect 569604 68082 569632 72984
rect 569960 72966 570012 72972
rect 569960 72480 570012 72486
rect 569696 72440 569960 72468
rect 569696 68388 569724 72440
rect 569960 72422 570012 72428
rect 569960 68400 570012 68406
rect 569696 68360 569960 68388
rect 569960 68342 570012 68348
rect 569604 68066 570000 68082
rect 569604 68060 570012 68066
rect 569604 68054 569960 68060
rect 569960 68002 570012 68008
rect 569960 67924 570012 67930
rect 569960 67866 570012 67872
rect 569972 65006 570000 67866
rect 570064 66026 570092 77166
rect 570144 76492 570196 76498
rect 570144 76434 570196 76440
rect 570156 67930 570184 76434
rect 570236 74724 570288 74730
rect 570236 74666 570288 74672
rect 570248 73302 570276 74666
rect 570236 73296 570288 73302
rect 570236 73238 570288 73244
rect 574756 69057 574784 110434
rect 574940 96558 574968 157354
rect 580170 111480 580226 111489
rect 580170 111415 580226 111424
rect 580184 110498 580212 111415
rect 580172 110492 580224 110498
rect 580172 110434 580224 110440
rect 574928 96552 574980 96558
rect 574928 96494 574980 96500
rect 574742 69048 574798 69057
rect 574742 68983 574798 68992
rect 570236 68400 570288 68406
rect 570236 68342 570288 68348
rect 570144 67924 570196 67930
rect 570144 67866 570196 67872
rect 570144 66156 570196 66162
rect 570144 66098 570196 66104
rect 570052 66020 570104 66026
rect 570052 65962 570104 65968
rect 569960 65000 570012 65006
rect 569960 64942 570012 64948
rect 569052 64790 570000 64818
rect 568960 64654 569448 64682
rect 568776 64518 569356 64546
rect 568684 64382 568988 64410
rect 568960 64002 568988 64382
rect 568960 63974 569172 64002
rect 569144 63186 569172 63974
rect 568408 55270 568620 55298
rect 568684 63158 569172 63186
rect 568408 54346 568436 55270
rect 568408 54318 568528 54346
rect 568500 49042 568528 54318
rect 568684 49722 568712 63158
rect 569328 63050 569356 64518
rect 568224 40004 568344 40032
rect 568408 49014 568528 49042
rect 568592 49694 568712 49722
rect 568776 63022 569356 63050
rect 20074 13288 20130 13297
rect 19996 13246 20074 13274
rect 19996 7993 20024 13246
rect 20074 13223 20130 13232
rect 19982 7984 20038 7993
rect 19982 7919 20038 7928
rect 225694 6488 225750 6497
rect 225750 6446 225828 6474
rect 225694 6423 225750 6432
rect 225800 5137 225828 6446
rect 225786 5128 225842 5137
rect 225786 5063 225842 5072
rect 124310 3768 124366 3777
rect 124310 3703 124366 3712
rect 177946 3768 178002 3777
rect 177946 3703 178002 3712
rect 268382 3768 268438 3777
rect 268382 3703 268438 3712
rect 124324 3126 124352 3703
rect 177960 3126 177988 3703
rect 268396 3126 268424 3703
rect 124312 3120 124364 3126
rect 124312 3062 124364 3068
rect 177948 3120 178000 3126
rect 177948 3062 178000 3068
rect 268384 3120 268436 3126
rect 268384 3062 268436 3068
rect 3792 1760 3844 1766
rect 7656 1760 7708 1766
rect 6090 1728 6146 1737
rect 3792 1702 3844 1708
rect 5460 1698 5750 1714
rect 4068 1692 4120 1698
rect 4068 1634 4120 1640
rect 5448 1692 5750 1698
rect 5500 1686 5750 1692
rect 6090 1663 6146 1672
rect 6826 1728 6882 1737
rect 22100 1760 22152 1766
rect 7656 1702 7708 1708
rect 11242 1728 11298 1737
rect 6826 1663 6882 1672
rect 5448 1634 5500 1640
rect 3698 1456 3754 1465
rect 3698 1391 3754 1400
rect 3608 536 3660 542
rect 3608 478 3660 484
rect 4080 480 4108 1634
rect 6104 1465 6132 1663
rect 6840 1494 6868 1663
rect 6828 1488 6880 1494
rect 5906 1456 5962 1465
rect 4908 1426 5304 1442
rect 4908 1420 5316 1426
rect 4908 1414 5264 1420
rect 4908 610 4936 1414
rect 5906 1391 5908 1400
rect 5264 1362 5316 1368
rect 5960 1391 5962 1400
rect 6090 1456 6146 1465
rect 6828 1430 6880 1436
rect 6090 1391 6146 1400
rect 6460 1420 6512 1426
rect 5908 1362 5960 1368
rect 6460 1362 6512 1368
rect 4988 1352 5040 1358
rect 5356 1352 5408 1358
rect 5040 1300 5356 1306
rect 4988 1294 5408 1300
rect 5000 1278 5396 1294
rect 5000 1154 5672 1170
rect 4988 1148 5672 1154
rect 5040 1142 5672 1148
rect 4988 1090 5040 1096
rect 5080 1080 5132 1086
rect 5540 1080 5592 1086
rect 5132 1028 5540 1034
rect 5080 1022 5592 1028
rect 5092 1006 5580 1022
rect 5644 898 5672 1142
rect 4988 876 5040 882
rect 4988 818 5040 824
rect 5552 870 5672 898
rect 5000 762 5028 818
rect 5000 734 5304 762
rect 4986 640 5042 649
rect 4896 604 4948 610
rect 4986 575 5042 584
rect 4896 546 4948 552
rect 5000 542 5028 575
rect 4988 536 5040 542
rect 3422 232 3478 241
rect 3056 196 3108 202
rect 3422 167 3478 176
rect 3056 138 3108 144
rect 4038 -960 4150 480
rect 4988 478 5040 484
rect 5276 480 5304 734
rect 5552 626 5580 870
rect 5630 640 5686 649
rect 5552 598 5630 626
rect 5630 575 5686 584
rect 6472 480 6500 1362
rect 7380 672 7432 678
rect 7380 614 7432 620
rect 7392 513 7420 614
rect 7378 504 7434 513
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7668 480 7696 1702
rect 11242 1663 11298 1672
rect 14462 1728 14518 1737
rect 22100 1702 22152 1708
rect 22192 1760 22244 1766
rect 22192 1702 22244 1708
rect 26424 1760 26476 1766
rect 48688 1760 48740 1766
rect 26424 1702 26476 1708
rect 37370 1728 37426 1737
rect 14462 1663 14518 1672
rect 18328 1692 18380 1698
rect 10416 1624 10468 1630
rect 10416 1566 10468 1572
rect 8852 1284 8904 1290
rect 8852 1226 8904 1232
rect 8864 480 8892 1226
rect 10428 1193 10456 1566
rect 10692 1420 10744 1426
rect 10692 1362 10744 1368
rect 10600 1352 10652 1358
rect 10520 1312 10600 1340
rect 10414 1184 10470 1193
rect 10414 1119 10470 1128
rect 10520 898 10548 1312
rect 10600 1294 10652 1300
rect 10244 870 10548 898
rect 10244 785 10272 870
rect 10230 776 10286 785
rect 10230 711 10286 720
rect 10060 598 10272 626
rect 10060 480 10088 598
rect 7378 439 7434 448
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 9864 128 9916 134
rect 9862 96 9864 105
rect 9916 96 9918 105
rect 9862 31 9918 40
rect 10018 -960 10130 480
rect 10244 105 10272 598
rect 10508 604 10560 610
rect 10508 546 10560 552
rect 10520 354 10548 546
rect 10704 377 10732 1362
rect 11256 480 11284 1663
rect 14476 1465 14504 1663
rect 18328 1634 18380 1640
rect 19340 1692 19392 1698
rect 19340 1634 19392 1640
rect 17960 1556 18012 1562
rect 17960 1498 18012 1504
rect 18052 1556 18104 1562
rect 18052 1498 18104 1504
rect 14462 1456 14518 1465
rect 14462 1391 14518 1400
rect 14646 1456 14702 1465
rect 14646 1391 14702 1400
rect 14464 1352 14516 1358
rect 14464 1294 14516 1300
rect 14556 1352 14608 1358
rect 14556 1294 14608 1300
rect 14476 921 14504 1294
rect 13634 912 13690 921
rect 13634 847 13690 856
rect 14462 912 14518 921
rect 14462 847 14518 856
rect 13268 740 13320 746
rect 13268 682 13320 688
rect 13280 649 13308 682
rect 13266 640 13322 649
rect 12452 598 12664 626
rect 12452 480 12480 598
rect 10428 326 10548 354
rect 10690 368 10746 377
rect 10428 270 10456 326
rect 10690 303 10746 312
rect 10416 264 10468 270
rect 10416 206 10468 212
rect 10230 96 10286 105
rect 10230 31 10286 40
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 12636 377 12664 598
rect 13266 575 13322 584
rect 13450 640 13506 649
rect 13450 575 13452 584
rect 13504 575 13506 584
rect 13452 546 13504 552
rect 13648 480 13676 847
rect 12622 368 12678 377
rect 12622 303 12678 312
rect 13082 232 13138 241
rect 13082 167 13138 176
rect 13096 66 13124 167
rect 13084 60 13136 66
rect 13084 2 13136 8
rect 13606 -960 13718 480
rect 14568 241 14596 1294
rect 14660 377 14688 1391
rect 15212 746 15240 1020
rect 17972 746 18000 1498
rect 18064 1358 18092 1498
rect 18052 1352 18104 1358
rect 18052 1294 18104 1300
rect 15200 740 15252 746
rect 15200 682 15252 688
rect 17960 740 18012 746
rect 17960 682 18012 688
rect 14844 598 15056 626
rect 14844 480 14872 598
rect 14646 368 14702 377
rect 14646 303 14702 312
rect 14554 232 14610 241
rect 14554 167 14610 176
rect 14802 -960 14914 480
rect 15028 241 15056 598
rect 17236 598 17448 626
rect 15856 564 16068 592
rect 15856 377 15884 564
rect 16040 480 16068 564
rect 17236 480 17264 598
rect 15842 368 15898 377
rect 15842 303 15898 312
rect 15014 232 15070 241
rect 15014 167 15070 176
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 17420 66 17448 598
rect 18340 480 18368 1634
rect 17408 60 17460 66
rect 17408 2 17460 8
rect 18298 -960 18410 480
rect 19352 241 19380 1634
rect 22112 921 22140 1702
rect 22098 912 22154 921
rect 22098 847 22154 856
rect 19432 808 19484 814
rect 19484 768 19840 796
rect 19432 750 19484 756
rect 19536 564 19748 592
rect 19536 480 19564 564
rect 19338 232 19394 241
rect 19338 167 19394 176
rect 19494 -960 19606 480
rect 19720 241 19748 564
rect 19812 377 19840 768
rect 20718 640 20774 649
rect 20718 575 20774 584
rect 21914 640 21970 649
rect 22204 610 22232 1702
rect 26436 1601 26464 1702
rect 26608 1692 26660 1698
rect 37370 1663 37426 1672
rect 37738 1728 37794 1737
rect 40958 1728 41014 1737
rect 39040 1698 39620 1714
rect 37738 1663 37740 1672
rect 26608 1634 26660 1640
rect 26620 1601 26648 1634
rect 26422 1592 26478 1601
rect 26422 1527 26478 1536
rect 26606 1592 26662 1601
rect 29734 1592 29790 1601
rect 26606 1527 26662 1536
rect 28356 1556 28408 1562
rect 29734 1527 29790 1536
rect 32678 1592 32734 1601
rect 32678 1527 32734 1536
rect 36176 1556 36228 1562
rect 28356 1498 28408 1504
rect 28262 1456 28318 1465
rect 28262 1391 28318 1400
rect 27896 1284 27948 1290
rect 27896 1226 27948 1232
rect 24308 1216 24360 1222
rect 24360 1164 24702 1170
rect 24308 1158 24702 1164
rect 24320 1142 24702 1158
rect 27908 1057 27936 1226
rect 26882 1048 26938 1057
rect 26882 983 26938 992
rect 27894 1048 27950 1057
rect 27894 983 27950 992
rect 23110 776 23166 785
rect 23110 711 23166 720
rect 24306 776 24362 785
rect 24306 711 24362 720
rect 21914 575 21970 584
rect 22192 604 22244 610
rect 20732 480 20760 575
rect 21928 480 21956 575
rect 22192 546 22244 552
rect 23124 480 23152 711
rect 24320 480 24348 711
rect 26700 672 26752 678
rect 25332 598 25544 626
rect 26700 614 26752 620
rect 19798 368 19854 377
rect 19798 303 19854 312
rect 19706 232 19762 241
rect 19706 167 19762 176
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25332 270 25360 598
rect 25516 480 25544 598
rect 26712 480 26740 614
rect 25320 264 25372 270
rect 25320 206 25372 212
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 26896 338 26924 983
rect 27894 912 27950 921
rect 28276 882 28304 1391
rect 27894 847 27950 856
rect 28264 876 28316 882
rect 27908 480 27936 847
rect 28264 818 28316 824
rect 26884 332 26936 338
rect 26884 274 26936 280
rect 27866 -960 27978 480
rect 28368 377 28396 1498
rect 29092 1420 29144 1426
rect 29092 1362 29144 1368
rect 29104 480 29132 1362
rect 29748 814 29776 1527
rect 31482 1456 31538 1465
rect 31482 1391 31538 1400
rect 29736 808 29788 814
rect 29736 750 29788 756
rect 30300 598 30512 626
rect 30300 480 30328 598
rect 28354 368 28410 377
rect 28354 303 28410 312
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 30484 377 30512 598
rect 31496 480 31524 1391
rect 32692 480 32720 1527
rect 36176 1498 36228 1504
rect 33888 1154 34178 1170
rect 33876 1148 34178 1154
rect 33928 1142 34178 1148
rect 33876 1090 33928 1096
rect 34978 912 35034 921
rect 34978 847 35034 856
rect 33704 598 33916 626
rect 33704 513 33732 598
rect 33690 504 33746 513
rect 30470 368 30526 377
rect 30470 303 30526 312
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33888 480 33916 598
rect 34992 480 35020 847
rect 35162 504 35218 513
rect 33690 439 33746 448
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36188 480 36216 1498
rect 37384 480 37412 1663
rect 37792 1663 37794 1672
rect 39028 1692 39620 1698
rect 37740 1634 37792 1640
rect 39080 1686 39620 1692
rect 39028 1634 39080 1640
rect 39394 1592 39450 1601
rect 39592 1562 39620 1686
rect 40958 1663 41014 1672
rect 41142 1728 41198 1737
rect 48686 1728 48688 1737
rect 48872 1760 48924 1766
rect 48740 1728 48742 1737
rect 41142 1663 41198 1672
rect 42708 1692 42760 1698
rect 39762 1592 39818 1601
rect 39394 1527 39450 1536
rect 39580 1556 39632 1562
rect 39302 1456 39358 1465
rect 39302 1391 39358 1400
rect 39316 1193 39344 1391
rect 39408 1222 39436 1527
rect 39762 1527 39818 1536
rect 39580 1498 39632 1504
rect 39396 1216 39448 1222
rect 39302 1184 39358 1193
rect 39396 1158 39448 1164
rect 39302 1119 39358 1128
rect 38566 912 38622 921
rect 38566 847 38622 856
rect 38200 808 38252 814
rect 38198 776 38200 785
rect 38252 776 38254 785
rect 38198 711 38254 720
rect 38382 776 38438 785
rect 38382 711 38438 720
rect 35162 439 35218 448
rect 35176 338 35204 439
rect 35164 332 35216 338
rect 35164 274 35216 280
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38396 270 38424 711
rect 38580 480 38608 847
rect 39776 480 39804 1527
rect 40972 480 41000 1663
rect 41156 1562 41184 1663
rect 42708 1634 42760 1640
rect 45560 1692 45612 1698
rect 50620 1760 50672 1766
rect 48924 1708 49096 1714
rect 48872 1702 49096 1708
rect 50620 1702 50672 1708
rect 50804 1760 50856 1766
rect 56416 1760 56468 1766
rect 50804 1702 50856 1708
rect 55034 1728 55090 1737
rect 48884 1686 49096 1702
rect 48686 1663 48742 1672
rect 45560 1634 45612 1640
rect 42524 1624 42576 1630
rect 42522 1592 42524 1601
rect 42720 1601 42748 1634
rect 42576 1592 42578 1601
rect 41144 1556 41196 1562
rect 42522 1527 42578 1536
rect 42706 1592 42762 1601
rect 42706 1527 42762 1536
rect 45468 1556 45520 1562
rect 41144 1498 41196 1504
rect 45468 1498 45520 1504
rect 45480 1465 45508 1498
rect 42246 1456 42302 1465
rect 44086 1456 44142 1465
rect 43746 1414 44086 1442
rect 42246 1391 42302 1400
rect 44086 1391 44142 1400
rect 45466 1456 45522 1465
rect 45572 1442 45600 1634
rect 48042 1592 48098 1601
rect 48042 1527 48098 1536
rect 48686 1592 48742 1601
rect 49068 1578 49096 1686
rect 49330 1592 49386 1601
rect 49068 1550 49330 1578
rect 48686 1527 48742 1536
rect 49330 1527 49386 1536
rect 45650 1456 45706 1465
rect 45572 1414 45650 1442
rect 45466 1391 45522 1400
rect 45650 1391 45706 1400
rect 42260 1193 42288 1391
rect 47032 1352 47084 1358
rect 47032 1294 47084 1300
rect 42062 1184 42118 1193
rect 42062 1119 42118 1128
rect 42246 1184 42302 1193
rect 42246 1119 42302 1128
rect 42076 814 42104 1119
rect 47044 1057 47072 1294
rect 47952 1284 48004 1290
rect 47952 1226 48004 1232
rect 46570 1048 46626 1057
rect 46570 983 46626 992
rect 46754 1048 46810 1057
rect 46754 983 46810 992
rect 47030 1048 47086 1057
rect 47030 983 47086 992
rect 42156 876 42208 882
rect 42156 818 42208 824
rect 42064 808 42116 814
rect 42064 750 42116 756
rect 42168 480 42196 818
rect 43352 808 43404 814
rect 46584 785 46612 983
rect 46664 876 46716 882
rect 46664 818 46716 824
rect 43352 750 43404 756
rect 46294 776 46350 785
rect 43364 480 43392 750
rect 46294 711 46350 720
rect 46570 776 46626 785
rect 46570 711 46626 720
rect 44376 598 44588 626
rect 38384 264 38436 270
rect 38384 206 38436 212
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44376 134 44404 598
rect 44560 480 44588 598
rect 45572 598 45784 626
rect 45572 513 45600 598
rect 45558 504 45614 513
rect 44364 128 44416 134
rect 44364 70 44416 76
rect 44518 -960 44630 480
rect 45756 480 45784 598
rect 45558 439 45614 448
rect 45714 -960 45826 480
rect 46308 134 46336 711
rect 46676 513 46704 818
rect 46768 678 46796 983
rect 47964 921 47992 1226
rect 47950 912 48006 921
rect 47950 847 48006 856
rect 48056 814 48084 1527
rect 48700 1290 48728 1527
rect 48964 1488 49016 1494
rect 50632 1476 50660 1702
rect 50816 1601 50844 1702
rect 55034 1663 55090 1672
rect 55218 1728 55274 1737
rect 56416 1702 56468 1708
rect 56692 1760 56744 1766
rect 111984 1760 112036 1766
rect 56692 1702 56744 1708
rect 59082 1728 59138 1737
rect 55218 1663 55274 1672
rect 50802 1592 50858 1601
rect 50986 1592 51042 1601
rect 50802 1527 50858 1536
rect 50908 1550 50986 1578
rect 50908 1476 50936 1550
rect 50986 1527 51042 1536
rect 50632 1448 50936 1476
rect 55048 1465 55076 1663
rect 55034 1456 55090 1465
rect 48964 1430 49016 1436
rect 48688 1284 48740 1290
rect 48688 1226 48740 1232
rect 48134 912 48190 921
rect 48134 847 48190 856
rect 48044 808 48096 814
rect 48044 750 48096 756
rect 46756 672 46808 678
rect 46756 614 46808 620
rect 46940 672 46992 678
rect 46940 614 46992 620
rect 46662 504 46718 513
rect 46952 480 46980 614
rect 48148 480 48176 847
rect 48976 785 49004 1430
rect 55034 1391 55090 1400
rect 55036 1352 55088 1358
rect 54036 1312 55036 1340
rect 48962 776 49018 785
rect 48962 711 49018 720
rect 49514 776 49570 785
rect 49514 711 49570 720
rect 49160 598 49372 626
rect 46662 439 46718 448
rect 46296 128 46348 134
rect 46296 70 46348 76
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49160 338 49188 598
rect 49344 480 49372 598
rect 49148 332 49200 338
rect 49148 274 49200 280
rect 49302 -960 49414 480
rect 49528 241 49556 711
rect 50540 598 50752 626
rect 49882 504 49938 513
rect 50540 480 50568 598
rect 50724 513 50752 598
rect 51644 598 51856 626
rect 50710 504 50766 513
rect 49882 439 49938 448
rect 49514 232 49570 241
rect 49896 202 49924 439
rect 49514 167 49570 176
rect 49884 196 49936 202
rect 49884 138 49936 144
rect 50498 -960 50610 480
rect 51644 480 51672 598
rect 50710 439 50766 448
rect 51602 -960 51714 480
rect 51828 241 51856 598
rect 52828 604 52880 610
rect 52828 546 52880 552
rect 52840 480 52868 546
rect 51814 232 51870 241
rect 51814 167 51870 176
rect 52798 -960 52910 480
rect 53208 270 53236 1020
rect 54036 480 54064 1312
rect 55036 1294 55088 1300
rect 55232 814 55260 1663
rect 55954 912 56010 921
rect 55954 847 56010 856
rect 55220 808 55272 814
rect 55220 750 55272 756
rect 55678 776 55734 785
rect 55678 711 55734 720
rect 55232 598 55444 626
rect 55232 480 55260 598
rect 53196 264 53248 270
rect 53196 206 53248 212
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 55416 134 55444 598
rect 55692 270 55720 711
rect 55588 264 55640 270
rect 55588 206 55640 212
rect 55680 264 55732 270
rect 55968 241 55996 847
rect 56428 480 56456 1702
rect 56600 1556 56652 1562
rect 56600 1498 56652 1504
rect 56612 1465 56640 1498
rect 56598 1456 56654 1465
rect 56598 1391 56654 1400
rect 56704 1222 56732 1702
rect 56784 1692 56836 1698
rect 56784 1634 56836 1640
rect 57888 1692 57940 1698
rect 59082 1663 59138 1672
rect 59266 1728 59322 1737
rect 64878 1728 64934 1737
rect 59266 1663 59322 1672
rect 57888 1634 57940 1640
rect 56692 1216 56744 1222
rect 56692 1158 56744 1164
rect 56796 950 56824 1634
rect 57900 1601 57928 1634
rect 57886 1592 57942 1601
rect 58438 1592 58494 1601
rect 57886 1527 57942 1536
rect 58072 1556 58124 1562
rect 58494 1550 58572 1578
rect 58438 1527 58494 1536
rect 58072 1498 58124 1504
rect 57980 1488 58032 1494
rect 57980 1430 58032 1436
rect 57992 1222 58020 1430
rect 57980 1216 58032 1222
rect 57980 1158 58032 1164
rect 58084 950 58112 1498
rect 58544 1465 58572 1550
rect 58530 1456 58586 1465
rect 58530 1391 58586 1400
rect 58256 1352 58308 1358
rect 59096 1340 59124 1663
rect 59280 1562 59308 1663
rect 64432 1652 64644 1680
rect 68834 1728 68890 1737
rect 64934 1686 65288 1714
rect 64878 1663 64934 1672
rect 61014 1592 61070 1601
rect 59268 1556 59320 1562
rect 59268 1498 59320 1504
rect 59360 1556 59412 1562
rect 61014 1527 61070 1536
rect 61198 1592 61254 1601
rect 61198 1527 61254 1536
rect 59360 1498 59412 1504
rect 59176 1352 59228 1358
rect 59096 1312 59176 1340
rect 58256 1294 58308 1300
rect 59176 1294 59228 1300
rect 58162 1184 58218 1193
rect 58268 1170 58296 1294
rect 58218 1142 58296 1170
rect 58346 1184 58402 1193
rect 58162 1119 58218 1128
rect 58346 1119 58402 1128
rect 56784 944 56836 950
rect 56784 886 56836 892
rect 58072 944 58124 950
rect 58072 886 58124 892
rect 58360 796 58388 1119
rect 57440 768 58388 796
rect 55680 206 55732 212
rect 55954 232 56010 241
rect 55404 128 55456 134
rect 55600 116 55628 206
rect 56138 232 56194 241
rect 55954 167 56010 176
rect 56060 190 56138 218
rect 56060 116 56088 190
rect 56138 167 56194 176
rect 55600 88 56088 116
rect 55404 70 55456 76
rect 56386 -960 56498 480
rect 57440 241 57468 768
rect 59372 678 59400 1498
rect 60740 1488 60792 1494
rect 60740 1430 60792 1436
rect 60278 1320 60334 1329
rect 60278 1255 60334 1264
rect 60292 1068 60320 1255
rect 60752 1193 60780 1430
rect 60830 1320 60886 1329
rect 60830 1255 60886 1264
rect 60738 1184 60794 1193
rect 60738 1119 60794 1128
rect 60844 1068 60872 1255
rect 60292 1040 60872 1068
rect 59360 672 59412 678
rect 57624 598 57836 626
rect 57624 480 57652 598
rect 57426 232 57482 241
rect 57426 167 57482 176
rect 57582 -960 57694 480
rect 57808 241 57836 598
rect 58636 598 58848 626
rect 59360 614 59412 620
rect 60004 672 60056 678
rect 60004 614 60056 620
rect 57794 232 57850 241
rect 58636 202 58664 598
rect 58820 480 58848 598
rect 60016 480 60044 614
rect 57794 167 57850 176
rect 58624 196 58676 202
rect 58624 138 58676 144
rect 58778 -960 58890 480
rect 58992 332 59044 338
rect 58992 274 59044 280
rect 59004 202 59032 274
rect 58992 196 59044 202
rect 58992 138 59044 144
rect 59974 -960 60086 480
rect 61028 270 61056 1527
rect 61212 950 61240 1527
rect 62394 1456 62450 1465
rect 62304 1420 62356 1426
rect 62946 1456 63002 1465
rect 62450 1414 62698 1442
rect 62394 1391 62450 1400
rect 62946 1391 63002 1400
rect 62304 1362 62356 1368
rect 62316 1086 62344 1362
rect 62304 1080 62356 1086
rect 62304 1022 62356 1028
rect 62396 1080 62448 1086
rect 62396 1022 62448 1028
rect 61200 944 61252 950
rect 61200 886 61252 892
rect 61212 598 61424 626
rect 61212 480 61240 598
rect 61016 264 61068 270
rect 61016 206 61068 212
rect 61170 -960 61282 480
rect 61396 241 61424 598
rect 62408 480 62436 1022
rect 62960 950 62988 1391
rect 63052 1380 63816 1408
rect 63052 1329 63080 1380
rect 63788 1329 63816 1380
rect 63038 1320 63094 1329
rect 63774 1320 63830 1329
rect 63038 1255 63094 1264
rect 63512 1290 63724 1306
rect 63512 1284 63736 1290
rect 63512 1278 63684 1284
rect 63314 1184 63370 1193
rect 63314 1119 63370 1128
rect 62948 944 63000 950
rect 63328 932 63356 1119
rect 63512 1057 63540 1278
rect 63774 1255 63830 1264
rect 63684 1226 63736 1232
rect 63592 1216 63644 1222
rect 63866 1184 63922 1193
rect 63592 1158 63644 1164
rect 63498 1048 63554 1057
rect 63498 983 63554 992
rect 63604 932 63632 1158
rect 63328 904 63632 932
rect 63788 1142 63866 1170
rect 62948 886 63000 892
rect 63788 882 63816 1142
rect 63866 1119 63922 1128
rect 63776 876 63828 882
rect 63776 818 63828 824
rect 63868 876 63920 882
rect 63868 818 63920 824
rect 63880 762 63908 818
rect 63604 734 63908 762
rect 63604 480 63632 734
rect 61382 232 61438 241
rect 61382 167 61438 176
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64432 241 64460 1652
rect 64510 1592 64566 1601
rect 64510 1527 64566 1536
rect 64524 1340 64552 1527
rect 64616 1442 64644 1652
rect 65260 1578 65288 1686
rect 65536 1686 68834 1714
rect 65338 1592 65394 1601
rect 65260 1550 65338 1578
rect 65338 1527 65394 1536
rect 65536 1442 65564 1686
rect 72422 1728 72478 1737
rect 71792 1698 72174 1714
rect 68834 1663 68890 1672
rect 71780 1692 72174 1698
rect 71832 1686 72174 1692
rect 73710 1728 73766 1737
rect 72478 1672 73200 1680
rect 72422 1663 73200 1672
rect 82634 1728 82690 1737
rect 75656 1686 76420 1714
rect 73766 1672 75500 1680
rect 73710 1663 75500 1672
rect 72436 1652 73200 1663
rect 73724 1652 75500 1663
rect 71780 1634 71832 1640
rect 66902 1592 66958 1601
rect 73172 1578 73200 1652
rect 74078 1592 74134 1601
rect 73172 1550 73752 1578
rect 66902 1527 66904 1536
rect 66956 1527 66958 1536
rect 66904 1498 66956 1504
rect 68848 1516 72096 1544
rect 64616 1414 65564 1442
rect 66902 1456 66958 1465
rect 67086 1456 67142 1465
rect 66902 1391 66958 1400
rect 67008 1414 67086 1442
rect 64524 1312 64736 1340
rect 64708 1272 64736 1312
rect 64708 1244 65104 1272
rect 64786 1184 64842 1193
rect 64786 1119 64842 1128
rect 64800 480 64828 1119
rect 64880 944 64932 950
rect 64932 892 65012 898
rect 64880 886 65012 892
rect 64892 870 65012 886
rect 64984 490 65012 870
rect 65076 864 65104 1244
rect 66916 1222 66944 1391
rect 66904 1216 66956 1222
rect 66718 1184 66774 1193
rect 66904 1158 66956 1164
rect 66718 1119 66774 1128
rect 66732 1086 66760 1119
rect 66628 1080 66680 1086
rect 66628 1022 66680 1028
rect 66720 1080 66772 1086
rect 66720 1022 66772 1028
rect 66640 898 66668 1022
rect 67008 898 67036 1414
rect 68848 1426 68876 1516
rect 67086 1391 67142 1400
rect 68836 1420 68888 1426
rect 68836 1362 68888 1368
rect 68928 1420 68980 1426
rect 68928 1362 68980 1368
rect 71872 1420 71924 1426
rect 71872 1362 71924 1368
rect 68940 1170 68968 1362
rect 66640 870 67036 898
rect 68112 1142 68968 1170
rect 65076 836 66024 864
rect 65338 504 65394 513
rect 64418 232 64474 241
rect 64418 167 64474 176
rect 64758 -960 64870 480
rect 64984 462 65338 490
rect 65996 480 66024 836
rect 67192 598 67404 626
rect 67192 480 67220 598
rect 65338 439 65394 448
rect 65062 368 65118 377
rect 65338 368 65394 377
rect 65118 326 65338 354
rect 65062 303 65118 312
rect 65338 303 65394 312
rect 65954 -960 66066 480
rect 66732 326 67036 354
rect 66732 241 66760 326
rect 67008 270 67036 326
rect 66904 264 66956 270
rect 66718 232 66774 241
rect 66718 167 66774 176
rect 66902 232 66904 241
rect 66996 264 67048 270
rect 66956 232 66958 241
rect 66996 206 67048 212
rect 66902 167 66958 176
rect 67150 -960 67262 480
rect 67376 270 67404 598
rect 68112 513 68140 1142
rect 68836 1080 68888 1086
rect 68888 1028 68968 1034
rect 68836 1022 68968 1028
rect 68848 1006 68968 1022
rect 68940 950 68968 1006
rect 68928 944 68980 950
rect 68928 886 68980 892
rect 70676 944 70728 950
rect 70676 886 70728 892
rect 68296 598 68508 626
rect 68098 504 68154 513
rect 68296 480 68324 598
rect 68480 513 68508 598
rect 69308 598 69520 626
rect 68466 504 68522 513
rect 68098 439 68154 448
rect 67364 264 67416 270
rect 67364 206 67416 212
rect 68254 -960 68366 480
rect 68466 439 68522 448
rect 69308 202 69336 598
rect 69492 480 69520 598
rect 70688 480 70716 886
rect 71884 480 71912 1362
rect 69296 196 69348 202
rect 69296 138 69348 144
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 72068 354 72096 1516
rect 73724 1442 73752 1550
rect 75366 1592 75422 1601
rect 74078 1527 74134 1536
rect 73986 1456 74042 1465
rect 73724 1414 73986 1442
rect 73986 1391 74042 1400
rect 74092 1306 74120 1527
rect 73172 1278 74120 1306
rect 74276 1516 74580 1544
rect 75472 1578 75500 1652
rect 75656 1578 75684 1686
rect 76392 1680 76420 1686
rect 82372 1686 82634 1714
rect 76392 1652 77248 1680
rect 75472 1550 75684 1578
rect 76194 1592 76250 1601
rect 75366 1527 75422 1536
rect 77114 1592 77170 1601
rect 76194 1527 76250 1536
rect 76392 1550 77114 1578
rect 73172 762 73200 1278
rect 72620 734 73200 762
rect 73264 1142 73660 1170
rect 72620 513 72648 734
rect 73264 626 73292 1142
rect 73342 1048 73398 1057
rect 73342 983 73398 992
rect 73080 598 73292 626
rect 73356 626 73384 983
rect 73632 932 73660 1142
rect 74276 1057 74304 1516
rect 74552 1426 74580 1516
rect 74448 1420 74500 1426
rect 74448 1362 74500 1368
rect 74540 1420 74592 1426
rect 74540 1362 74592 1368
rect 74460 1057 74488 1362
rect 74262 1048 74318 1057
rect 74262 983 74318 992
rect 74446 1048 74502 1057
rect 74446 983 74502 992
rect 75380 932 75408 1527
rect 73632 904 74580 932
rect 75380 904 75960 932
rect 73356 598 74304 626
rect 72606 504 72662 513
rect 72790 504 72846 513
rect 72606 439 72662 448
rect 72712 462 72790 490
rect 72712 354 72740 462
rect 73080 480 73108 598
rect 73252 536 73304 542
rect 74078 504 74134 513
rect 73304 484 73936 490
rect 72790 439 72846 448
rect 72068 326 72740 354
rect 73038 -960 73150 480
rect 73252 478 73936 484
rect 73264 462 73936 478
rect 73342 368 73398 377
rect 73802 368 73858 377
rect 73398 326 73660 354
rect 73342 303 73398 312
rect 73528 264 73580 270
rect 73526 232 73528 241
rect 73632 252 73660 326
rect 73802 303 73858 312
rect 73816 252 73844 303
rect 73580 232 73582 241
rect 73632 224 73844 252
rect 73526 167 73582 176
rect 73908 105 73936 462
rect 74276 480 74304 598
rect 74078 439 74134 448
rect 74092 241 74120 439
rect 74078 232 74134 241
rect 74078 167 74134 176
rect 73894 96 73950 105
rect 73894 31 73950 40
rect 74234 -960 74346 480
rect 74552 105 74580 904
rect 75644 672 75696 678
rect 75472 620 75644 626
rect 75472 614 75696 620
rect 75472 598 75684 614
rect 75472 480 75500 598
rect 75932 513 75960 904
rect 76208 513 76236 1527
rect 75734 504 75790 513
rect 74538 96 74594 105
rect 74538 31 74594 40
rect 75430 -960 75542 480
rect 75734 439 75790 448
rect 75918 504 75974 513
rect 75918 439 75974 448
rect 76194 504 76250 513
rect 76194 439 76250 448
rect 75748 354 75776 439
rect 76392 354 76420 1550
rect 77114 1527 77170 1536
rect 77220 1442 77248 1652
rect 78416 1652 78720 1680
rect 78416 1601 78444 1652
rect 78402 1592 78458 1601
rect 78402 1527 78458 1536
rect 78586 1592 78642 1601
rect 78586 1527 78642 1536
rect 78600 1494 78628 1527
rect 76576 1414 77248 1442
rect 78588 1488 78640 1494
rect 78588 1430 78640 1436
rect 76472 944 76524 950
rect 76472 886 76524 892
rect 76484 762 76512 886
rect 76576 864 76604 1414
rect 78692 1408 78720 1652
rect 82266 1592 82322 1601
rect 82266 1527 82322 1536
rect 81360 1426 81742 1442
rect 78864 1420 78916 1426
rect 78692 1380 78864 1408
rect 78864 1362 78916 1368
rect 81348 1420 81742 1426
rect 81400 1414 81742 1420
rect 81808 1420 81860 1426
rect 81348 1362 81400 1368
rect 81808 1362 81860 1368
rect 76656 1352 76708 1358
rect 76708 1300 78260 1306
rect 76656 1294 78260 1300
rect 76668 1278 78260 1294
rect 76840 876 76892 882
rect 76576 836 76840 864
rect 76840 818 76892 824
rect 76484 734 76696 762
rect 76668 480 76696 734
rect 77680 598 77892 626
rect 75748 326 76420 354
rect 76626 -960 76738 480
rect 77680 241 77708 598
rect 77864 480 77892 598
rect 77666 232 77722 241
rect 77666 167 77722 176
rect 77822 -960 77934 480
rect 78232 241 78260 1278
rect 78772 1284 78824 1290
rect 78508 1244 78772 1272
rect 78508 513 78536 1244
rect 78772 1226 78824 1232
rect 78864 1148 78916 1154
rect 78864 1090 78916 1096
rect 78494 504 78550 513
rect 78494 439 78550 448
rect 78218 232 78274 241
rect 78218 167 78274 176
rect 78876 105 78904 1090
rect 79048 808 79100 814
rect 81820 762 81848 1362
rect 82174 1184 82230 1193
rect 82280 1170 82308 1527
rect 82372 1290 82400 1686
rect 83738 1728 83794 1737
rect 82634 1663 82690 1672
rect 82740 1686 83412 1714
rect 82740 1306 82768 1686
rect 83384 1578 83412 1686
rect 83738 1663 83794 1672
rect 85670 1728 85726 1737
rect 100482 1728 100538 1737
rect 85726 1686 86172 1714
rect 85670 1663 85726 1672
rect 83384 1550 83596 1578
rect 83186 1456 83242 1465
rect 83370 1456 83426 1465
rect 83242 1414 83320 1442
rect 83186 1391 83242 1400
rect 82360 1284 82412 1290
rect 82360 1226 82412 1232
rect 82464 1278 82768 1306
rect 82464 1170 82492 1278
rect 82280 1142 82492 1170
rect 82556 1142 83044 1170
rect 82174 1119 82230 1128
rect 82188 1068 82216 1119
rect 82556 1068 82584 1142
rect 83016 1086 83044 1142
rect 83188 1148 83240 1154
rect 83292 1136 83320 1414
rect 83568 1442 83596 1550
rect 83646 1456 83702 1465
rect 83568 1414 83646 1442
rect 83370 1391 83426 1400
rect 83646 1391 83702 1400
rect 83384 1154 83412 1391
rect 83240 1108 83320 1136
rect 83372 1148 83424 1154
rect 83188 1090 83240 1096
rect 83556 1148 83608 1154
rect 83372 1090 83424 1096
rect 83476 1108 83556 1136
rect 82188 1040 82584 1068
rect 83004 1080 83056 1086
rect 82648 1006 82860 1034
rect 83004 1022 83056 1028
rect 82450 912 82506 921
rect 79048 750 79100 756
rect 79060 480 79088 750
rect 79244 734 81848 762
rect 82188 870 82450 898
rect 79244 513 79272 734
rect 80256 598 80468 626
rect 79230 504 79286 513
rect 78862 96 78918 105
rect 78862 31 78918 40
rect 79018 -960 79130 480
rect 80256 480 80284 598
rect 80440 513 80468 598
rect 81452 598 81664 626
rect 80426 504 80482 513
rect 79230 439 79286 448
rect 80214 -960 80326 480
rect 81452 480 81480 598
rect 80426 439 80482 448
rect 81410 -960 81522 480
rect 81636 105 81664 598
rect 82188 241 82216 870
rect 82648 898 82676 1006
rect 82832 932 82860 1006
rect 83476 932 83504 1108
rect 83556 1090 83608 1096
rect 82832 904 83504 932
rect 82556 882 82676 898
rect 82450 847 82506 856
rect 82544 876 82676 882
rect 82596 870 82676 876
rect 82728 876 82780 882
rect 82544 818 82596 824
rect 82728 818 82780 824
rect 82740 728 82768 818
rect 83648 808 83700 814
rect 83752 796 83780 1663
rect 85672 1420 85724 1426
rect 85672 1362 85724 1368
rect 85856 1420 85908 1426
rect 85856 1362 85908 1368
rect 84764 1278 85068 1306
rect 83844 882 84240 898
rect 84764 882 84792 1278
rect 84936 1216 84988 1222
rect 84936 1158 84988 1164
rect 83832 876 84240 882
rect 83884 870 84240 876
rect 83832 818 83884 824
rect 83700 768 83780 796
rect 83648 750 83700 756
rect 82648 700 82768 728
rect 83832 740 83884 746
rect 82648 480 82676 700
rect 83832 682 83884 688
rect 83844 480 83872 682
rect 84212 626 84240 870
rect 84752 876 84804 882
rect 84752 818 84804 824
rect 84212 598 84700 626
rect 82174 232 82230 241
rect 82174 167 82230 176
rect 81622 96 81678 105
rect 81622 31 81678 40
rect 82606 -960 82718 480
rect 83464 196 83516 202
rect 83464 138 83516 144
rect 82910 96 82966 105
rect 83476 82 83504 138
rect 82966 54 83504 82
rect 82910 31 82966 40
rect 83802 -960 83914 480
rect 84212 326 84516 354
rect 84212 241 84240 326
rect 84198 232 84254 241
rect 84198 167 84254 176
rect 84382 232 84438 241
rect 84488 202 84516 326
rect 84672 202 84700 598
rect 84948 480 84976 1158
rect 85040 1034 85068 1278
rect 85684 1204 85712 1362
rect 85868 1329 85896 1362
rect 86144 1340 86172 1686
rect 92584 1686 96936 1714
rect 92584 1601 92612 1686
rect 92570 1592 92626 1601
rect 92570 1527 92626 1536
rect 92754 1592 92810 1601
rect 96434 1592 96490 1601
rect 92754 1527 92810 1536
rect 92860 1550 96434 1578
rect 91926 1456 91982 1465
rect 86880 1414 87184 1442
rect 86880 1358 86908 1414
rect 87156 1408 87184 1414
rect 87156 1380 91324 1408
rect 91982 1414 92060 1442
rect 91926 1391 91982 1400
rect 86316 1352 86368 1358
rect 85854 1320 85910 1329
rect 86038 1320 86094 1329
rect 85854 1255 85910 1264
rect 85960 1278 86038 1306
rect 85960 1204 85988 1278
rect 86144 1312 86316 1340
rect 86316 1294 86368 1300
rect 86868 1352 86920 1358
rect 86868 1294 86920 1300
rect 86038 1255 86094 1264
rect 88536 1278 88748 1306
rect 88536 1222 88564 1278
rect 87880 1216 87932 1222
rect 85684 1176 85988 1204
rect 86420 1176 87880 1204
rect 86420 1034 86448 1176
rect 88156 1216 88208 1222
rect 87880 1158 87932 1164
rect 88076 1176 88156 1204
rect 88076 1034 88104 1176
rect 88156 1158 88208 1164
rect 88524 1216 88576 1222
rect 88524 1158 88576 1164
rect 88616 1216 88668 1222
rect 88616 1158 88668 1164
rect 88720 1170 88748 1278
rect 91296 1272 91324 1380
rect 92032 1306 92060 1414
rect 92768 1408 92796 1527
rect 92584 1380 92796 1408
rect 92202 1320 92258 1329
rect 91928 1284 91980 1290
rect 91296 1244 91928 1272
rect 92032 1278 92202 1306
rect 92584 1290 92612 1380
rect 92202 1255 92258 1264
rect 92572 1284 92624 1290
rect 91928 1226 91980 1232
rect 92572 1226 92624 1232
rect 92664 1284 92716 1290
rect 92860 1272 92888 1550
rect 96434 1527 96490 1536
rect 96618 1592 96674 1601
rect 96908 1578 96936 1686
rect 97092 1686 100482 1714
rect 96986 1592 97042 1601
rect 96908 1550 96986 1578
rect 96618 1527 96674 1536
rect 96986 1527 97042 1536
rect 96632 1442 96660 1527
rect 97092 1442 97120 1686
rect 100956 1720 107608 1748
rect 100956 1714 100984 1720
rect 100482 1663 100538 1672
rect 100864 1686 100984 1714
rect 100864 1544 100892 1686
rect 101968 1652 103652 1680
rect 101678 1592 101734 1601
rect 96632 1414 97120 1442
rect 100220 1516 100892 1544
rect 100956 1516 101260 1544
rect 101678 1527 101680 1536
rect 100220 1329 100248 1516
rect 100956 1465 100984 1516
rect 100942 1456 100998 1465
rect 100942 1391 100998 1400
rect 101126 1456 101182 1465
rect 101232 1442 101260 1516
rect 101732 1527 101734 1536
rect 101680 1498 101732 1504
rect 101310 1456 101366 1465
rect 101232 1414 101310 1442
rect 101126 1391 101182 1400
rect 101310 1391 101366 1400
rect 101140 1340 101168 1391
rect 101140 1329 101444 1340
rect 96618 1320 96674 1329
rect 92716 1244 92888 1272
rect 93136 1278 96618 1306
rect 92664 1226 92716 1232
rect 93136 1222 93164 1278
rect 97906 1320 97962 1329
rect 96618 1255 96674 1264
rect 97828 1278 97906 1306
rect 92204 1216 92256 1222
rect 90730 1184 90786 1193
rect 85040 1006 86448 1034
rect 87800 1006 88104 1034
rect 86144 734 87552 762
rect 86144 480 86172 734
rect 87524 728 87552 734
rect 87800 728 87828 1006
rect 87880 876 87932 882
rect 87880 818 87932 824
rect 87524 700 87828 728
rect 87340 598 87552 626
rect 87340 480 87368 598
rect 84382 167 84438 176
rect 84476 196 84528 202
rect 84198 96 84254 105
rect 84396 82 84424 167
rect 84476 138 84528 144
rect 84660 196 84712 202
rect 84660 138 84712 144
rect 84254 54 84424 82
rect 84198 31 84254 40
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 87524 241 87552 598
rect 87510 232 87566 241
rect 87892 218 87920 818
rect 88628 592 88656 1158
rect 88720 1142 90730 1170
rect 90730 1119 90786 1128
rect 92202 1184 92204 1193
rect 93124 1216 93176 1222
rect 92256 1184 92258 1193
rect 92202 1119 92258 1128
rect 92308 1142 92980 1170
rect 93124 1158 93176 1164
rect 92020 1080 92072 1086
rect 88536 564 88656 592
rect 89548 1006 91218 1034
rect 92308 1034 92336 1142
rect 92072 1028 92336 1034
rect 92020 1022 92336 1028
rect 92756 1080 92808 1086
rect 92756 1022 92808 1028
rect 92848 1080 92900 1086
rect 92848 1022 92900 1028
rect 92032 1006 92336 1022
rect 88536 480 88564 564
rect 87708 202 87920 218
rect 87510 167 87566 176
rect 87696 196 87920 202
rect 87748 190 87920 196
rect 87696 138 87748 144
rect 88494 -960 88606 480
rect 89548 406 89576 1006
rect 91466 912 91522 921
rect 91466 847 91522 856
rect 92110 912 92166 921
rect 92166 870 92336 898
rect 92110 847 92166 856
rect 91480 728 91508 847
rect 89732 700 91508 728
rect 91742 776 91798 785
rect 92018 776 92074 785
rect 91798 734 92018 762
rect 91742 711 91798 720
rect 92018 711 92074 720
rect 89732 480 89760 700
rect 90744 632 92152 660
rect 89536 400 89588 406
rect 89536 342 89588 348
rect 89690 -960 89802 480
rect 90744 406 90772 632
rect 90928 564 91140 592
rect 90928 480 90956 564
rect 90732 400 90784 406
rect 90732 342 90784 348
rect 90886 -960 90998 480
rect 91112 406 91140 564
rect 92124 480 92152 632
rect 91100 400 91152 406
rect 91100 342 91152 348
rect 92082 -960 92194 480
rect 92308 218 92336 870
rect 92664 808 92716 814
rect 92664 750 92716 756
rect 92572 468 92624 474
rect 92676 456 92704 750
rect 92768 474 92796 1022
rect 92860 814 92888 1022
rect 92848 808 92900 814
rect 92848 750 92900 756
rect 92952 660 92980 1142
rect 97078 1048 97134 1057
rect 93044 1006 94176 1034
rect 93044 814 93072 1006
rect 93492 876 93544 882
rect 93136 836 93492 864
rect 93032 808 93084 814
rect 93032 750 93084 756
rect 93136 660 93164 836
rect 94044 876 94096 882
rect 93492 818 93544 824
rect 93596 836 94044 864
rect 92952 632 93164 660
rect 93228 700 93532 728
rect 93228 592 93256 700
rect 93400 604 93452 610
rect 92860 564 93256 592
rect 93320 564 93400 592
rect 92624 428 92704 456
rect 92756 468 92808 474
rect 92572 410 92624 416
rect 92756 410 92808 416
rect 92478 368 92534 377
rect 92662 368 92718 377
rect 92534 326 92662 354
rect 92478 303 92534 312
rect 92662 303 92718 312
rect 92860 218 92888 564
rect 93320 480 93348 564
rect 93400 546 93452 552
rect 92308 190 92888 218
rect 93278 -960 93390 480
rect 93504 82 93532 700
rect 93596 241 93624 836
rect 94044 818 94096 824
rect 93860 604 93912 610
rect 93860 546 93912 552
rect 93582 232 93638 241
rect 93766 232 93822 241
rect 93582 167 93638 176
rect 93688 190 93766 218
rect 93688 82 93716 190
rect 93766 167 93822 176
rect 93872 105 93900 546
rect 94148 105 94176 1006
rect 97078 983 97134 992
rect 97262 1048 97318 1057
rect 97262 983 97318 992
rect 97092 882 97120 983
rect 97276 950 97304 983
rect 97264 944 97316 950
rect 97264 886 97316 892
rect 97080 876 97132 882
rect 97080 818 97132 824
rect 94240 564 94544 592
rect 94240 406 94268 564
rect 94516 480 94544 564
rect 95712 564 95924 592
rect 95712 480 95740 564
rect 94228 400 94280 406
rect 94228 342 94280 348
rect 93504 54 93716 82
rect 93858 96 93914 105
rect 93858 31 93914 40
rect 94134 96 94190 105
rect 94134 31 94190 40
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 95896 406 95924 564
rect 96908 564 97120 592
rect 96908 480 96936 564
rect 95884 400 95936 406
rect 95884 342 95936 348
rect 96866 -960 96978 480
rect 97092 82 97120 564
rect 97828 241 97856 1278
rect 97906 1255 97962 1264
rect 100206 1320 100262 1329
rect 101140 1320 101458 1329
rect 101140 1312 101402 1320
rect 100312 1290 100694 1306
rect 100206 1255 100262 1264
rect 100300 1284 100694 1290
rect 100352 1278 100694 1284
rect 101968 1290 101996 1652
rect 102336 1584 103192 1612
rect 102232 1556 102284 1562
rect 102336 1544 102364 1584
rect 102284 1516 102364 1544
rect 102232 1498 102284 1504
rect 102782 1456 102838 1465
rect 103058 1456 103114 1465
rect 102838 1414 103058 1442
rect 102782 1391 102838 1400
rect 103058 1391 103114 1400
rect 102232 1352 102284 1358
rect 102322 1320 102378 1329
rect 102284 1300 102322 1306
rect 102232 1294 102322 1300
rect 101402 1255 101458 1264
rect 101956 1284 102008 1290
rect 100300 1226 100352 1232
rect 102244 1278 102322 1294
rect 102598 1320 102654 1329
rect 102322 1255 102378 1264
rect 102428 1278 102598 1306
rect 101956 1226 102008 1232
rect 101402 1184 101458 1193
rect 100864 1128 101402 1136
rect 100864 1119 101458 1128
rect 100864 1108 101444 1119
rect 100864 1068 100892 1108
rect 100772 1040 100892 1068
rect 100772 932 100800 1040
rect 102428 1034 102456 1278
rect 103058 1320 103114 1329
rect 102784 1284 102836 1290
rect 102598 1255 102654 1264
rect 97920 904 100800 932
rect 100956 1006 102456 1034
rect 102704 1244 102784 1272
rect 97814 232 97870 241
rect 97814 167 97870 176
rect 97920 82 97948 904
rect 100956 864 100984 1006
rect 101680 944 101732 950
rect 99300 836 100984 864
rect 101140 904 101680 932
rect 98104 564 98316 592
rect 98104 480 98132 564
rect 97092 54 97948 82
rect 98062 -960 98174 480
rect 98288 241 98316 564
rect 99300 480 99328 836
rect 100760 740 100812 746
rect 100496 700 100760 728
rect 100496 480 100524 700
rect 100760 682 100812 688
rect 98274 232 98330 241
rect 98274 167 98330 176
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101140 354 101168 904
rect 102704 932 102732 1244
rect 103058 1255 103114 1264
rect 102784 1226 102836 1232
rect 101680 886 101732 892
rect 101784 904 102732 932
rect 101404 808 101456 814
rect 101404 750 101456 756
rect 101416 592 101444 750
rect 101416 564 101628 592
rect 101600 480 101628 564
rect 101048 326 101168 354
rect 101048 105 101076 326
rect 101034 96 101090 105
rect 101034 31 101090 40
rect 101558 -960 101670 480
rect 101784 105 101812 904
rect 101956 808 102008 814
rect 101956 750 102008 756
rect 102230 776 102286 785
rect 101968 105 101996 750
rect 102690 776 102746 785
rect 102416 740 102468 746
rect 102286 720 102416 728
rect 102230 711 102416 720
rect 102244 700 102416 711
rect 102690 711 102692 720
rect 102416 682 102468 688
rect 102744 711 102746 720
rect 102692 682 102744 688
rect 103072 610 103100 1255
rect 103164 1170 103192 1584
rect 103426 1592 103482 1601
rect 103336 1556 103388 1562
rect 103426 1527 103482 1536
rect 103336 1498 103388 1504
rect 103348 1290 103376 1498
rect 103336 1284 103388 1290
rect 103336 1226 103388 1232
rect 103440 1170 103468 1527
rect 103624 1408 103652 1652
rect 103716 1652 107148 1680
rect 103716 1562 103744 1652
rect 103704 1556 103756 1562
rect 103704 1498 103756 1504
rect 106924 1488 106976 1494
rect 106924 1430 106976 1436
rect 103624 1380 106872 1408
rect 103518 1320 103574 1329
rect 106738 1320 106794 1329
rect 103518 1255 103574 1264
rect 103808 1278 106320 1306
rect 103164 1142 103468 1170
rect 103532 1000 103560 1255
rect 103164 972 103560 1000
rect 103060 604 103112 610
rect 102796 564 103008 592
rect 102796 480 102824 564
rect 102980 490 103008 564
rect 103060 546 103112 552
rect 103164 490 103192 972
rect 103428 876 103480 882
rect 103428 818 103480 824
rect 103440 626 103468 818
rect 103808 785 103836 1278
rect 104624 1216 104676 1222
rect 104622 1184 104624 1193
rect 106292 1204 106320 1278
rect 106648 1284 106700 1290
rect 106844 1290 106872 1380
rect 106738 1255 106794 1264
rect 106832 1284 106884 1290
rect 106648 1226 106700 1232
rect 106556 1216 106608 1222
rect 104676 1184 104678 1193
rect 103980 1148 104032 1154
rect 104622 1119 104678 1128
rect 104806 1184 104862 1193
rect 106292 1176 106556 1204
rect 106556 1158 106608 1164
rect 104806 1119 104808 1128
rect 103980 1090 104032 1096
rect 104860 1119 104862 1128
rect 105820 1148 105872 1154
rect 104808 1090 104860 1096
rect 105872 1108 106504 1136
rect 105820 1090 105872 1096
rect 103992 1034 104020 1090
rect 103992 1006 106412 1034
rect 103900 836 105216 864
rect 103794 776 103850 785
rect 103794 711 103850 720
rect 103900 626 103928 836
rect 103978 776 104034 785
rect 103978 711 104034 720
rect 103440 598 103928 626
rect 101770 96 101826 105
rect 101770 31 101826 40
rect 101954 96 102010 105
rect 101954 31 102010 40
rect 102754 -960 102866 480
rect 102980 462 103192 490
rect 103992 480 104020 711
rect 105188 480 105216 836
rect 106384 480 106412 1006
rect 106476 882 106504 1108
rect 106660 1000 106688 1226
rect 106752 1068 106780 1255
rect 106832 1226 106884 1232
rect 106830 1184 106886 1193
rect 106936 1170 106964 1430
rect 106886 1142 106964 1170
rect 106830 1119 106886 1128
rect 106752 1040 107056 1068
rect 107120 1057 107148 1652
rect 107580 1578 107608 1720
rect 111430 1728 111486 1737
rect 110800 1686 111380 1714
rect 107580 1550 109080 1578
rect 109052 1544 109080 1550
rect 109052 1516 109356 1544
rect 107304 1244 107516 1272
rect 106660 972 106780 1000
rect 106464 876 106516 882
rect 106464 818 106516 824
rect 106752 490 106780 972
rect 107028 814 107056 1040
rect 107106 1048 107162 1057
rect 107106 983 107162 992
rect 106924 808 106976 814
rect 106924 750 106976 756
rect 107016 808 107068 814
rect 107016 750 107068 756
rect 106936 592 106964 750
rect 107304 592 107332 1244
rect 107488 1204 107516 1244
rect 107382 1184 107438 1193
rect 107488 1176 109264 1204
rect 107438 1128 109172 1136
rect 107382 1119 109172 1128
rect 107396 1108 109172 1119
rect 109038 1048 109094 1057
rect 109038 983 109094 992
rect 108856 876 108908 882
rect 109052 864 109080 983
rect 109144 932 109172 1108
rect 109236 1057 109264 1176
rect 109328 1170 109356 1516
rect 110800 1465 110828 1686
rect 111352 1630 111380 1686
rect 111430 1663 111486 1672
rect 111628 1720 111984 1748
rect 111340 1624 111392 1630
rect 111246 1592 111302 1601
rect 111168 1550 111246 1578
rect 110786 1456 110842 1465
rect 109880 1426 110170 1442
rect 109868 1420 110170 1426
rect 109920 1414 110170 1420
rect 109868 1362 109920 1368
rect 110248 1380 110644 1408
rect 110786 1391 110842 1400
rect 110248 1170 110276 1380
rect 110616 1290 110644 1380
rect 111168 1290 111196 1550
rect 111340 1566 111392 1572
rect 111444 1578 111472 1663
rect 111628 1578 111656 1720
rect 128268 1760 128320 1766
rect 111984 1702 112036 1708
rect 112732 1720 117084 1748
rect 112168 1624 112220 1630
rect 111444 1550 111656 1578
rect 112166 1592 112168 1601
rect 112220 1592 112222 1601
rect 111246 1527 111302 1536
rect 111720 1516 112116 1544
rect 112166 1527 112222 1536
rect 111248 1488 111300 1494
rect 111246 1456 111248 1465
rect 111300 1456 111302 1465
rect 111246 1391 111302 1400
rect 111430 1456 111486 1465
rect 111430 1391 111432 1400
rect 111484 1391 111486 1400
rect 111432 1362 111484 1368
rect 111720 1306 111748 1516
rect 111982 1456 112038 1465
rect 111982 1391 112038 1400
rect 110420 1284 110472 1290
rect 110420 1226 110472 1232
rect 110604 1284 110656 1290
rect 110604 1226 110656 1232
rect 111156 1284 111208 1290
rect 111156 1226 111208 1232
rect 111260 1278 111748 1306
rect 111892 1284 111944 1290
rect 109328 1142 110276 1170
rect 110326 1184 110382 1193
rect 110326 1119 110382 1128
rect 109222 1048 109278 1057
rect 110340 1000 110368 1119
rect 110432 1068 110460 1226
rect 110512 1216 110564 1222
rect 110510 1184 110512 1193
rect 110564 1184 110566 1193
rect 110510 1119 110566 1128
rect 111260 1068 111288 1278
rect 111892 1226 111944 1232
rect 111614 1184 111670 1193
rect 111614 1119 111670 1128
rect 110432 1040 111288 1068
rect 111628 1000 111656 1119
rect 109222 983 109278 992
rect 109328 972 110092 1000
rect 110340 972 111656 1000
rect 109328 932 109356 972
rect 109144 904 109356 932
rect 110064 882 110092 972
rect 111904 932 111932 1226
rect 111996 1222 112024 1391
rect 111984 1216 112036 1222
rect 111984 1158 112036 1164
rect 112088 1170 112116 1516
rect 112626 1184 112682 1193
rect 112088 1142 112626 1170
rect 112626 1119 112682 1128
rect 112732 1068 112760 1720
rect 115204 1624 115256 1630
rect 115204 1566 115256 1572
rect 115216 1426 115244 1566
rect 115492 1550 116164 1578
rect 115204 1420 115256 1426
rect 115204 1362 115256 1368
rect 111168 904 111932 932
rect 111996 1040 112760 1068
rect 109408 876 109460 882
rect 108908 836 108988 864
rect 109052 836 109408 864
rect 108856 818 108908 824
rect 108028 808 108080 814
rect 107382 776 107438 785
rect 107382 711 107438 720
rect 107842 776 107898 785
rect 107842 711 107844 720
rect 106936 564 107332 592
rect 107396 490 107424 711
rect 107896 711 107898 720
rect 107948 768 108028 796
rect 107844 682 107896 688
rect 107948 626 107976 768
rect 108028 750 108080 756
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 106752 462 107424 490
rect 107580 598 107976 626
rect 108592 598 108804 626
rect 107580 480 107608 598
rect 107538 -960 107650 480
rect 108592 105 108620 598
rect 108776 480 108804 598
rect 108578 96 108634 105
rect 108578 31 108634 40
rect 108734 -960 108846 480
rect 108960 241 108988 836
rect 109408 818 109460 824
rect 109960 876 110012 882
rect 109960 818 110012 824
rect 110052 876 110104 882
rect 110052 818 110104 824
rect 109972 480 110000 818
rect 111168 480 111196 904
rect 111536 836 111840 864
rect 111536 746 111564 836
rect 111524 740 111576 746
rect 111524 682 111576 688
rect 111616 740 111668 746
rect 111616 682 111668 688
rect 111628 649 111656 682
rect 111812 649 111840 836
rect 111614 640 111670 649
rect 111614 575 111670 584
rect 111798 640 111854 649
rect 111798 575 111854 584
rect 111890 504 111946 513
rect 108946 232 109002 241
rect 108946 167 109002 176
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 111890 439 111946 448
rect 111904 406 111932 439
rect 111892 400 111944 406
rect 111892 342 111944 348
rect 111706 232 111762 241
rect 111996 218 112024 1040
rect 115492 1000 115520 1550
rect 116136 1476 116164 1550
rect 116136 1448 116256 1476
rect 112272 972 115520 1000
rect 115584 1414 115980 1442
rect 112076 740 112128 746
rect 112076 682 112128 688
rect 112088 649 112116 682
rect 112074 640 112130 649
rect 112272 592 112300 972
rect 112824 870 113680 898
rect 112824 814 112852 870
rect 112352 808 112404 814
rect 112812 808 112864 814
rect 112404 768 112668 796
rect 112352 750 112404 756
rect 112074 575 112130 584
rect 112180 564 112300 592
rect 112350 640 112406 649
rect 112350 575 112406 584
rect 112074 504 112130 513
rect 112074 439 112130 448
rect 112088 406 112116 439
rect 112076 400 112128 406
rect 112076 342 112128 348
rect 111762 190 112024 218
rect 112180 202 112208 564
rect 112364 480 112392 575
rect 112168 196 112220 202
rect 111706 167 111762 176
rect 112168 138 112220 144
rect 112322 -960 112434 480
rect 112640 105 112668 768
rect 112812 750 112864 756
rect 113548 808 113600 814
rect 113548 750 113600 756
rect 113560 480 113588 750
rect 113652 626 113680 870
rect 113732 808 113784 814
rect 113730 776 113732 785
rect 113784 776 113786 785
rect 113730 711 113786 720
rect 114098 640 114154 649
rect 113652 598 114098 626
rect 115584 626 115612 1414
rect 115952 1154 115980 1414
rect 115940 1148 115992 1154
rect 115940 1090 115992 1096
rect 116228 1018 116256 1448
rect 117056 1329 117084 1720
rect 120630 1728 120686 1737
rect 120092 1652 120304 1680
rect 122286 1728 122342 1737
rect 120686 1686 121408 1714
rect 120630 1663 120686 1672
rect 119448 1426 119738 1442
rect 119436 1420 119738 1426
rect 119488 1414 119738 1420
rect 119804 1420 119856 1426
rect 119436 1362 119488 1368
rect 119804 1362 119856 1368
rect 116858 1320 116914 1329
rect 116504 1290 116716 1306
rect 116492 1284 116728 1290
rect 116544 1278 116676 1284
rect 116492 1226 116544 1232
rect 116676 1226 116728 1232
rect 116768 1284 116820 1290
rect 116858 1255 116914 1264
rect 117042 1320 117098 1329
rect 117042 1255 117098 1264
rect 116768 1226 116820 1232
rect 116780 1170 116808 1226
rect 116872 1204 116900 1255
rect 119344 1216 119396 1222
rect 116872 1176 119344 1204
rect 116412 1142 116808 1170
rect 119816 1170 119844 1362
rect 119344 1158 119396 1164
rect 119448 1142 119844 1170
rect 116216 1012 116268 1018
rect 116216 954 116268 960
rect 116412 785 116440 1142
rect 119448 1034 119476 1142
rect 116504 1006 119476 1034
rect 120092 1018 120120 1652
rect 120170 1592 120226 1601
rect 120276 1578 120304 1652
rect 120276 1550 121316 1578
rect 120170 1527 120226 1536
rect 120184 1068 120212 1527
rect 120630 1456 120686 1465
rect 120356 1420 120408 1426
rect 120906 1456 120962 1465
rect 120686 1414 120906 1442
rect 120630 1391 120686 1400
rect 120906 1391 120962 1400
rect 121000 1420 121052 1426
rect 120356 1362 120408 1368
rect 121000 1362 121052 1368
rect 120368 1193 120396 1362
rect 120354 1184 120410 1193
rect 120354 1119 120410 1128
rect 120184 1040 120856 1068
rect 120080 1012 120132 1018
rect 116398 776 116454 785
rect 115768 700 116072 728
rect 116398 711 116454 720
rect 115768 649 115796 700
rect 116044 660 116072 700
rect 116504 660 116532 1006
rect 120080 954 120132 960
rect 116584 944 116636 950
rect 116584 886 116636 892
rect 117136 944 117188 950
rect 117136 886 117188 892
rect 116596 785 116624 886
rect 116582 776 116638 785
rect 116582 711 116638 720
rect 114098 575 114154 584
rect 114756 598 115612 626
rect 115754 640 115810 649
rect 114756 480 114784 598
rect 115754 575 115810 584
rect 115938 640 115994 649
rect 116044 632 116532 660
rect 115938 575 115994 584
rect 115952 480 115980 575
rect 117148 480 117176 886
rect 118252 870 120764 898
rect 118252 480 118280 870
rect 120736 814 120764 870
rect 120540 808 120592 814
rect 120724 808 120776 814
rect 120592 768 120672 796
rect 120540 750 120592 756
rect 119448 564 119660 592
rect 119448 480 119476 564
rect 112626 96 112682 105
rect 112626 31 112682 40
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 116582 232 116638 241
rect 116858 232 116914 241
rect 116638 190 116858 218
rect 116582 167 116638 176
rect 116858 167 116914 176
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 119632 105 119660 564
rect 120644 480 120672 768
rect 120724 750 120776 756
rect 120828 490 120856 1040
rect 121012 660 121040 1362
rect 121288 1170 121316 1550
rect 121380 1290 121408 1686
rect 121840 1686 122286 1714
rect 121840 1329 121868 1686
rect 122286 1663 122342 1672
rect 124310 1728 124366 1737
rect 125782 1728 125838 1737
rect 124366 1686 124444 1714
rect 124310 1663 124366 1672
rect 121918 1592 121974 1601
rect 121918 1527 121974 1536
rect 121932 1408 121960 1527
rect 122748 1488 122800 1494
rect 122116 1448 122748 1476
rect 122012 1420 122064 1426
rect 121932 1380 122012 1408
rect 122012 1362 122064 1368
rect 121826 1320 121882 1329
rect 121368 1284 121420 1290
rect 122010 1320 122066 1329
rect 121826 1255 121882 1264
rect 121932 1278 122010 1306
rect 121368 1226 121420 1232
rect 121932 1170 121960 1278
rect 122010 1255 122066 1264
rect 121288 1142 121960 1170
rect 121184 1080 121236 1086
rect 121184 1022 121236 1028
rect 120920 649 121040 660
rect 121196 649 121224 1022
rect 122116 864 122144 1448
rect 122748 1430 122800 1436
rect 124416 1340 124444 1686
rect 124588 1692 124640 1698
rect 128266 1728 128268 1737
rect 138940 1760 138992 1766
rect 128320 1728 128322 1737
rect 129002 1728 129058 1737
rect 125782 1663 125838 1672
rect 124588 1634 124640 1640
rect 124600 1476 124628 1634
rect 125796 1630 125824 1663
rect 125888 1652 127940 1680
rect 128266 1663 128322 1672
rect 128924 1686 129002 1714
rect 125784 1624 125836 1630
rect 125784 1566 125836 1572
rect 125888 1476 125916 1652
rect 127806 1592 127862 1601
rect 127806 1527 127862 1536
rect 124600 1448 125916 1476
rect 125968 1488 126020 1494
rect 125968 1430 126020 1436
rect 127714 1456 127770 1465
rect 125980 1340 126008 1430
rect 127714 1391 127770 1400
rect 124416 1312 126008 1340
rect 126152 1284 126204 1290
rect 122852 1244 126152 1272
rect 122852 1154 122880 1244
rect 127728 1272 127756 1391
rect 127820 1340 127848 1527
rect 127912 1465 127940 1652
rect 128820 1624 128872 1630
rect 127990 1592 128046 1601
rect 127990 1527 128046 1536
rect 128648 1584 128820 1612
rect 128004 1494 128032 1527
rect 127992 1488 128044 1494
rect 127898 1456 127954 1465
rect 127992 1430 128044 1436
rect 128452 1488 128504 1494
rect 128452 1430 128504 1436
rect 127898 1391 127954 1400
rect 128464 1340 128492 1430
rect 128648 1358 128676 1584
rect 128820 1566 128872 1572
rect 128924 1358 128952 1686
rect 135166 1728 135222 1737
rect 129002 1663 129058 1672
rect 134524 1692 134576 1698
rect 134576 1652 135024 1680
rect 135166 1663 135168 1672
rect 134524 1634 134576 1640
rect 134890 1592 134946 1601
rect 134996 1578 135024 1652
rect 135220 1663 135222 1672
rect 135350 1728 135406 1737
rect 135350 1663 135406 1672
rect 135626 1728 135682 1737
rect 135626 1663 135682 1672
rect 136270 1728 136326 1737
rect 138386 1728 138442 1737
rect 136326 1686 137048 1714
rect 136270 1663 136326 1672
rect 135168 1634 135220 1640
rect 135364 1612 135392 1663
rect 135640 1612 135668 1663
rect 135074 1592 135130 1601
rect 134996 1550 135074 1578
rect 134890 1527 134946 1536
rect 135364 1584 135576 1612
rect 135640 1584 136496 1612
rect 135074 1527 135130 1536
rect 129002 1456 129058 1465
rect 129002 1391 129058 1400
rect 129476 1448 131988 1476
rect 127820 1312 128492 1340
rect 128636 1352 128688 1358
rect 128636 1294 128688 1300
rect 128912 1352 128964 1358
rect 128912 1294 128964 1300
rect 128544 1284 128596 1290
rect 127728 1244 128544 1272
rect 126152 1226 126204 1232
rect 128544 1226 128596 1232
rect 125506 1184 125562 1193
rect 122840 1148 122892 1154
rect 123208 1148 123260 1154
rect 122840 1090 122892 1096
rect 122944 1108 123208 1136
rect 122944 1034 122972 1108
rect 123208 1090 123260 1096
rect 123404 1142 125506 1170
rect 122472 1012 122524 1018
rect 122472 954 122524 960
rect 122760 1006 122972 1034
rect 121288 836 122144 864
rect 120906 640 121040 649
rect 120962 632 121040 640
rect 121182 640 121238 649
rect 120906 575 120962 584
rect 121182 575 121238 584
rect 121288 490 121316 836
rect 122484 814 122512 954
rect 122564 944 122616 950
rect 122564 886 122616 892
rect 122576 814 122604 886
rect 122472 808 122524 814
rect 122472 750 122524 756
rect 122564 808 122616 814
rect 122760 785 122788 1006
rect 122564 750 122616 756
rect 122746 776 122802 785
rect 122746 711 122802 720
rect 122852 734 123340 762
rect 122196 672 122248 678
rect 119618 96 119674 105
rect 119618 31 119674 40
rect 120602 -960 120714 480
rect 120828 462 121316 490
rect 121840 632 122196 660
rect 121840 480 121868 632
rect 122196 614 122248 620
rect 122852 490 122880 734
rect 121798 -960 121910 480
rect 122668 462 122880 490
rect 123036 564 123248 592
rect 123036 480 123064 564
rect 122668 377 122696 462
rect 122654 368 122710 377
rect 122654 303 122710 312
rect 122994 -960 123106 480
rect 123220 218 123248 564
rect 123312 377 123340 734
rect 123298 368 123354 377
rect 123298 303 123354 312
rect 123404 218 123432 1142
rect 125506 1119 125562 1128
rect 126702 1184 126758 1193
rect 128450 1184 128506 1193
rect 126758 1142 128450 1170
rect 126702 1119 126758 1128
rect 128450 1119 128506 1128
rect 123574 1048 123630 1057
rect 123758 1048 123814 1057
rect 123574 983 123630 992
rect 123680 1006 123758 1034
rect 123588 950 123616 983
rect 123484 944 123536 950
rect 123484 886 123536 892
rect 123576 944 123628 950
rect 123576 886 123628 892
rect 123220 190 123432 218
rect 123496 218 123524 886
rect 123680 796 123708 1006
rect 128818 1048 128874 1057
rect 123758 983 123814 992
rect 123944 1012 123996 1018
rect 125600 1012 125652 1018
rect 123996 972 125600 1000
rect 123944 954 123996 960
rect 128818 983 128874 992
rect 125600 954 125652 960
rect 128832 898 128860 983
rect 124416 870 128860 898
rect 124416 864 124444 870
rect 129016 864 129044 1391
rect 129280 1352 129332 1358
rect 129280 1294 129332 1300
rect 129108 1006 129214 1034
rect 129108 950 129136 1006
rect 129096 944 129148 950
rect 129096 886 129148 892
rect 123588 768 123708 796
rect 123772 836 124444 864
rect 128924 836 129044 864
rect 123588 354 123616 768
rect 123772 649 123800 836
rect 128924 762 128952 836
rect 124048 734 128952 762
rect 129094 776 129150 785
rect 123758 640 123814 649
rect 123942 640 123998 649
rect 123758 575 123814 584
rect 123864 598 123942 626
rect 123864 354 123892 598
rect 123942 575 123998 584
rect 123588 326 123892 354
rect 124048 218 124076 734
rect 129292 762 129320 1294
rect 129476 950 129504 1448
rect 131960 1408 131988 1448
rect 134798 1456 134854 1465
rect 129752 1380 131804 1408
rect 131960 1380 134748 1408
rect 134798 1391 134800 1400
rect 129464 944 129516 950
rect 129464 886 129516 892
rect 129752 864 129780 1380
rect 131302 1320 131358 1329
rect 131486 1320 131542 1329
rect 131302 1255 131358 1264
rect 131408 1278 131486 1306
rect 129150 734 129320 762
rect 129568 836 129780 864
rect 129094 711 129150 720
rect 124218 640 124274 649
rect 129568 626 129596 836
rect 129646 776 129702 785
rect 131316 762 131344 1255
rect 131408 898 131436 1278
rect 131670 1320 131726 1329
rect 131486 1255 131542 1264
rect 131592 1278 131670 1306
rect 131486 1048 131542 1057
rect 131592 1034 131620 1278
rect 131670 1255 131726 1264
rect 131776 1170 131804 1380
rect 134720 1329 134748 1380
rect 134852 1391 134854 1400
rect 134800 1362 134852 1368
rect 134706 1320 134762 1329
rect 134616 1284 134668 1290
rect 132512 1244 134616 1272
rect 132512 1170 132540 1244
rect 134904 1306 134932 1527
rect 135548 1465 135576 1584
rect 135534 1456 135590 1465
rect 135534 1391 135590 1400
rect 135812 1420 135864 1426
rect 135812 1362 135864 1368
rect 135074 1320 135130 1329
rect 134706 1255 134762 1264
rect 134800 1284 134852 1290
rect 134616 1226 134668 1232
rect 134904 1278 135074 1306
rect 135074 1255 135130 1264
rect 134800 1226 134852 1232
rect 131776 1142 132540 1170
rect 134812 1154 134840 1226
rect 135824 1204 135852 1362
rect 135902 1320 135958 1329
rect 136362 1320 136418 1329
rect 135958 1278 136362 1306
rect 135902 1255 135958 1264
rect 136468 1306 136496 1584
rect 136546 1592 136602 1601
rect 136546 1527 136602 1536
rect 136560 1442 136588 1527
rect 136914 1456 136970 1465
rect 136560 1414 136914 1442
rect 136914 1391 136970 1400
rect 136914 1320 136970 1329
rect 136468 1278 136914 1306
rect 136362 1255 136418 1264
rect 136914 1255 136970 1264
rect 137020 1204 137048 1686
rect 137192 1692 137244 1698
rect 137192 1634 137244 1640
rect 138296 1692 138348 1698
rect 145564 1760 145616 1766
rect 139412 1720 140728 1748
rect 139412 1714 139440 1720
rect 138940 1702 138992 1708
rect 138386 1663 138388 1672
rect 138296 1634 138348 1640
rect 138440 1663 138442 1672
rect 138756 1692 138808 1698
rect 138388 1634 138440 1640
rect 138756 1634 138808 1640
rect 137204 1329 137232 1634
rect 138308 1578 138336 1634
rect 138308 1550 138690 1578
rect 138768 1426 138796 1634
rect 138756 1420 138808 1426
rect 138756 1362 138808 1368
rect 137190 1320 137246 1329
rect 137190 1255 137246 1264
rect 135534 1184 135590 1193
rect 134800 1148 134852 1154
rect 135824 1176 137048 1204
rect 135534 1119 135590 1128
rect 134800 1090 134852 1096
rect 131542 1006 131620 1034
rect 131670 1048 131726 1057
rect 131486 983 131542 992
rect 135548 1034 135576 1119
rect 135810 1048 135866 1057
rect 135548 1006 135810 1034
rect 131670 983 131672 992
rect 131724 983 131726 992
rect 135810 983 135866 992
rect 131672 954 131724 960
rect 132604 904 136404 932
rect 131408 870 132540 898
rect 132512 864 132540 870
rect 132604 864 132632 904
rect 136376 898 136404 904
rect 138386 912 138442 921
rect 136376 870 138386 898
rect 132512 836 132632 864
rect 135364 836 136220 864
rect 138386 847 138442 856
rect 131316 734 135208 762
rect 129646 711 129702 720
rect 129660 660 129688 711
rect 129660 632 135116 660
rect 124218 575 124274 584
rect 125428 598 129596 626
rect 124232 480 124260 575
rect 125428 480 125456 598
rect 129278 504 129334 513
rect 123496 190 124076 218
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 129922 504 129978 513
rect 129334 462 129922 490
rect 129278 439 129334 448
rect 129922 439 129978 448
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 135088 354 135116 632
rect 135180 456 135208 734
rect 135364 649 135392 836
rect 136086 776 136142 785
rect 136192 762 136220 836
rect 138952 762 138980 1702
rect 139320 1686 139440 1714
rect 139214 1456 139270 1465
rect 139124 1420 139176 1426
rect 139214 1391 139216 1400
rect 139124 1362 139176 1368
rect 139268 1391 139270 1400
rect 139216 1362 139268 1368
rect 139136 1306 139164 1362
rect 139320 1306 139348 1686
rect 139780 1584 140544 1612
rect 139582 1456 139638 1465
rect 139582 1391 139638 1400
rect 139136 1278 139348 1306
rect 139492 1216 139544 1222
rect 139596 1204 139624 1391
rect 139544 1176 139624 1204
rect 139780 1193 139808 1584
rect 139872 1516 140452 1544
rect 139766 1184 139822 1193
rect 139492 1158 139544 1164
rect 139766 1119 139822 1128
rect 139872 1068 139900 1516
rect 140042 1456 140098 1465
rect 140042 1391 140098 1400
rect 140226 1456 140282 1465
rect 140424 1426 140452 1516
rect 140226 1391 140282 1400
rect 140320 1420 140372 1426
rect 139030 1048 139086 1057
rect 139412 1040 139900 1068
rect 139412 1034 139440 1040
rect 139086 1006 139440 1034
rect 139030 983 139086 992
rect 139412 921 139624 932
rect 139398 912 139638 921
rect 139454 904 139582 912
rect 139398 847 139454 856
rect 139582 847 139638 856
rect 136192 734 138980 762
rect 139398 776 139454 785
rect 136086 711 136142 720
rect 139582 776 139638 785
rect 139454 720 139582 728
rect 139398 711 139638 720
rect 136100 660 136128 711
rect 139412 700 139624 711
rect 135350 640 135406 649
rect 136100 632 139992 660
rect 140056 649 140084 1391
rect 140240 1154 140268 1391
rect 140320 1362 140372 1368
rect 140412 1420 140464 1426
rect 140412 1362 140464 1368
rect 140228 1148 140280 1154
rect 140228 1090 140280 1096
rect 140332 1034 140360 1362
rect 140516 1170 140544 1584
rect 140700 1476 140728 1720
rect 141146 1728 141202 1737
rect 140792 1686 141146 1714
rect 140792 1601 140820 1686
rect 144366 1728 144422 1737
rect 141146 1663 141202 1672
rect 142632 1652 143028 1680
rect 144366 1663 144422 1672
rect 145102 1728 145158 1737
rect 145840 1760 145892 1766
rect 145564 1702 145616 1708
rect 145654 1728 145710 1737
rect 145102 1663 145158 1672
rect 140778 1592 140834 1601
rect 140962 1592 141018 1601
rect 140778 1527 140834 1536
rect 140884 1550 140962 1578
rect 140884 1476 140912 1550
rect 142528 1556 142580 1562
rect 140962 1527 141018 1536
rect 140700 1448 140912 1476
rect 141160 1516 142528 1544
rect 141160 1426 141188 1516
rect 142528 1498 142580 1504
rect 141238 1456 141294 1465
rect 141148 1420 141200 1426
rect 141514 1456 141570 1465
rect 141294 1414 141514 1442
rect 141238 1391 141294 1400
rect 141514 1391 141570 1400
rect 141148 1362 141200 1368
rect 140780 1284 140832 1290
rect 140832 1244 142476 1272
rect 140780 1226 140832 1232
rect 141330 1184 141386 1193
rect 140516 1142 141330 1170
rect 142344 1148 142396 1154
rect 141330 1119 141386 1128
rect 142080 1108 142344 1136
rect 142080 1034 142108 1108
rect 142344 1090 142396 1096
rect 140332 1006 142108 1034
rect 142448 950 142476 1244
rect 140504 944 140556 950
rect 140148 904 140504 932
rect 135350 575 135406 584
rect 135548 564 139900 592
rect 135444 468 135496 474
rect 135180 428 135444 456
rect 135444 410 135496 416
rect 135548 354 135576 564
rect 135088 326 135576 354
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 139872 354 139900 564
rect 139964 490 139992 632
rect 140042 640 140098 649
rect 140042 575 140098 584
rect 140148 490 140176 904
rect 140504 886 140556 892
rect 142436 944 142488 950
rect 142436 886 142488 892
rect 139964 462 140176 490
rect 140608 836 142384 864
rect 140608 354 140636 836
rect 142250 776 142306 785
rect 142356 762 142384 836
rect 142434 776 142490 785
rect 142356 734 142434 762
rect 142250 711 142306 720
rect 142434 711 142490 720
rect 142264 660 142292 711
rect 142264 632 142384 660
rect 139872 326 140636 354
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 142356 474 142384 632
rect 142252 468 142304 474
rect 142252 410 142304 416
rect 142344 468 142396 474
rect 142344 410 142396 416
rect 142264 354 142292 410
rect 142632 354 142660 1652
rect 142896 1556 142948 1562
rect 142896 1498 142948 1504
rect 142804 1284 142856 1290
rect 142804 1226 142856 1232
rect 142816 660 142844 1226
rect 142908 1000 142936 1498
rect 143000 1408 143028 1652
rect 144380 1544 144408 1663
rect 144736 1624 144788 1630
rect 144788 1584 144868 1612
rect 144736 1566 144788 1572
rect 144840 1578 144868 1584
rect 145010 1592 145066 1601
rect 144840 1550 145010 1578
rect 144380 1516 144500 1544
rect 145010 1527 145066 1536
rect 144472 1476 144500 1516
rect 144472 1448 145052 1476
rect 144184 1420 144236 1426
rect 143000 1380 144184 1408
rect 144184 1362 144236 1368
rect 145024 1306 145052 1448
rect 145116 1426 145144 1663
rect 145576 1494 145604 1702
rect 145654 1663 145710 1672
rect 145838 1728 145840 1737
rect 146208 1760 146260 1766
rect 145892 1728 145894 1737
rect 145838 1663 145894 1672
rect 146206 1728 146208 1737
rect 147036 1760 147088 1766
rect 146260 1728 146262 1737
rect 148324 1760 148376 1766
rect 147088 1720 147904 1748
rect 147036 1702 147088 1708
rect 146206 1663 146262 1672
rect 145564 1488 145616 1494
rect 145668 1476 145696 1663
rect 145838 1592 145894 1601
rect 147402 1592 147458 1601
rect 145894 1550 147402 1578
rect 145838 1527 145894 1536
rect 147402 1527 147458 1536
rect 145668 1448 147812 1476
rect 145564 1430 145616 1436
rect 145104 1420 145156 1426
rect 145104 1362 145156 1368
rect 145196 1420 145248 1426
rect 145196 1362 145248 1368
rect 145208 1306 145236 1362
rect 145024 1278 145236 1306
rect 145300 1312 147720 1340
rect 144828 1216 144880 1222
rect 144828 1158 144880 1164
rect 144920 1216 144972 1222
rect 145300 1193 145328 1312
rect 145392 1244 145788 1272
rect 144920 1158 144972 1164
rect 145286 1184 145342 1193
rect 144840 1068 144868 1158
rect 144932 1068 144960 1158
rect 145286 1119 145342 1128
rect 144840 1040 144960 1068
rect 145392 1000 145420 1244
rect 145470 1184 145526 1193
rect 145470 1119 145526 1128
rect 142908 972 145420 1000
rect 144182 776 144238 785
rect 145484 762 145512 1119
rect 145760 785 145788 1244
rect 146128 1142 146708 1170
rect 146128 1018 146156 1142
rect 146680 1068 146708 1142
rect 147588 1148 147640 1154
rect 147588 1090 147640 1096
rect 147496 1080 147548 1086
rect 146680 1040 147496 1068
rect 147496 1022 147548 1028
rect 146116 1012 146168 1018
rect 146116 954 146168 960
rect 147600 796 147628 1090
rect 147692 864 147720 1312
rect 147784 932 147812 1448
rect 147876 1329 147904 1720
rect 148046 1728 148102 1737
rect 148102 1686 148258 1714
rect 148324 1702 148376 1708
rect 148600 1760 148652 1766
rect 149244 1760 149296 1766
rect 148600 1702 148652 1708
rect 148966 1728 149022 1737
rect 148046 1663 148102 1672
rect 147862 1320 147918 1329
rect 147862 1255 147918 1264
rect 148336 932 148364 1702
rect 148612 1193 148640 1702
rect 149150 1728 149206 1737
rect 149022 1686 149100 1714
rect 148966 1663 149022 1672
rect 148968 1624 149020 1630
rect 148690 1592 148746 1601
rect 148968 1566 149020 1572
rect 148690 1527 148746 1536
rect 148704 1329 148732 1527
rect 148876 1420 148928 1426
rect 148876 1362 148928 1368
rect 148888 1329 148916 1362
rect 148690 1320 148746 1329
rect 148690 1255 148746 1264
rect 148874 1320 148930 1329
rect 148874 1255 148930 1264
rect 148598 1184 148654 1193
rect 148980 1170 149008 1566
rect 149072 1329 149100 1686
rect 149244 1702 149296 1708
rect 149336 1760 149388 1766
rect 149336 1702 149388 1708
rect 149980 1760 150032 1766
rect 156788 1760 156840 1766
rect 150032 1720 150112 1748
rect 154316 1737 156788 1748
rect 149980 1702 150032 1708
rect 149150 1663 149206 1672
rect 149058 1320 149114 1329
rect 149058 1255 149114 1264
rect 148598 1119 148654 1128
rect 148796 1142 149008 1170
rect 147784 904 148364 932
rect 148796 864 148824 1142
rect 148876 1080 148928 1086
rect 149164 1068 149192 1663
rect 149256 1494 149284 1702
rect 149244 1488 149296 1494
rect 149244 1430 149296 1436
rect 149242 1184 149298 1193
rect 149242 1119 149298 1128
rect 148928 1040 149192 1068
rect 148876 1022 148928 1028
rect 147692 836 148824 864
rect 149256 796 149284 1119
rect 144238 734 145512 762
rect 145746 776 145802 785
rect 144182 711 144238 720
rect 145746 711 145802 720
rect 146942 776 146998 785
rect 147600 768 149284 796
rect 149348 728 149376 1702
rect 150084 1578 150112 1720
rect 154302 1728 156788 1737
rect 150164 1692 150216 1698
rect 150624 1692 150676 1698
rect 150216 1652 150624 1680
rect 150164 1634 150216 1640
rect 150624 1634 150676 1640
rect 150728 1652 154252 1680
rect 154358 1720 156788 1728
rect 161572 1760 161624 1766
rect 158810 1728 158866 1737
rect 156788 1702 156840 1708
rect 154302 1663 154358 1672
rect 156892 1686 157196 1714
rect 150728 1578 150756 1652
rect 154224 1612 154252 1652
rect 156892 1612 156920 1686
rect 150084 1550 150756 1578
rect 152384 1601 153976 1612
rect 152384 1592 153990 1601
rect 152384 1584 153934 1592
rect 152004 1556 152056 1562
rect 150820 1516 152004 1544
rect 149428 1488 149480 1494
rect 150820 1442 150848 1516
rect 152004 1498 152056 1504
rect 149480 1436 150848 1442
rect 149428 1430 150848 1436
rect 149440 1414 150848 1430
rect 151542 1456 151598 1465
rect 151818 1456 151874 1465
rect 151598 1414 151818 1442
rect 151542 1391 151598 1400
rect 151818 1391 151874 1400
rect 150256 1352 150308 1358
rect 151912 1352 151964 1358
rect 150308 1312 151912 1340
rect 150256 1294 150308 1300
rect 152384 1329 152412 1584
rect 152660 1516 153056 1544
rect 154224 1584 156920 1612
rect 157064 1624 157116 1630
rect 157064 1566 157116 1572
rect 153934 1527 153990 1536
rect 152556 1488 152608 1494
rect 152556 1430 152608 1436
rect 152568 1329 152596 1430
rect 151912 1294 151964 1300
rect 152002 1320 152058 1329
rect 152370 1320 152426 1329
rect 152002 1255 152058 1264
rect 152096 1284 152148 1290
rect 149796 1216 149848 1222
rect 150898 1184 150954 1193
rect 149796 1158 149848 1164
rect 149520 944 149572 950
rect 149808 932 149836 1158
rect 149992 1154 150898 1170
rect 149980 1148 150898 1154
rect 150032 1142 150898 1148
rect 150898 1119 150954 1128
rect 149980 1090 150032 1096
rect 149808 904 150756 932
rect 149520 886 149572 892
rect 146998 720 149376 728
rect 146942 711 149376 720
rect 146956 700 149376 711
rect 149532 660 149560 886
rect 142816 632 143672 660
rect 143644 626 143672 632
rect 144748 632 149560 660
rect 149624 734 150664 762
rect 143644 598 144684 626
rect 142264 326 142660 354
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 144656 354 144684 598
rect 144748 474 144776 632
rect 149624 592 149652 734
rect 150256 672 150308 678
rect 144840 564 149652 592
rect 150254 640 150256 649
rect 150308 640 150310 649
rect 150254 575 150310 584
rect 144736 468 144788 474
rect 144736 410 144788 416
rect 144840 354 144868 564
rect 144656 326 144868 354
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 150636 354 150664 734
rect 150728 626 150756 904
rect 151174 912 151230 921
rect 152016 898 152044 1255
rect 152370 1255 152426 1264
rect 152554 1320 152610 1329
rect 152660 1290 152688 1516
rect 153028 1476 153056 1516
rect 154040 1516 156828 1544
rect 154040 1476 154068 1516
rect 153028 1448 154068 1476
rect 156800 1476 156828 1516
rect 157076 1476 157104 1566
rect 157168 1562 157196 1686
rect 158994 1728 159050 1737
rect 158810 1663 158866 1672
rect 158904 1692 158956 1698
rect 158824 1630 158852 1663
rect 158994 1663 159050 1672
rect 159652 1686 161428 1714
rect 169484 1760 169536 1766
rect 161624 1720 166396 1748
rect 161572 1702 161624 1708
rect 158904 1634 158956 1640
rect 158812 1624 158864 1630
rect 157352 1562 157734 1578
rect 158812 1566 158864 1572
rect 157156 1556 157208 1562
rect 157156 1498 157208 1504
rect 157340 1556 157734 1562
rect 157392 1550 157734 1556
rect 157984 1556 158036 1562
rect 157340 1498 157392 1504
rect 157904 1516 157984 1544
rect 156800 1448 157104 1476
rect 154118 1320 154174 1329
rect 152554 1255 152610 1264
rect 152648 1284 152700 1290
rect 152096 1226 152148 1232
rect 152648 1226 152700 1232
rect 152752 1278 153792 1306
rect 151230 870 152044 898
rect 151174 847 151230 856
rect 152108 814 152136 1226
rect 152464 1216 152516 1222
rect 152752 1170 152780 1278
rect 153764 1204 153792 1278
rect 157522 1320 157578 1329
rect 154118 1255 154174 1264
rect 156420 1284 156472 1290
rect 153844 1216 153896 1222
rect 152516 1164 152780 1170
rect 152464 1158 152780 1164
rect 152476 1142 152780 1158
rect 152844 1176 153700 1204
rect 153764 1176 153844 1204
rect 152372 944 152424 950
rect 152844 932 152872 1176
rect 152424 904 152872 932
rect 153028 1108 153608 1136
rect 152372 886 152424 892
rect 152096 808 152148 814
rect 152096 750 152148 756
rect 152188 740 152240 746
rect 151188 700 151860 728
rect 151082 640 151138 649
rect 150728 598 151082 626
rect 151082 575 151138 584
rect 150806 504 150862 513
rect 151188 490 151216 700
rect 151450 640 151506 649
rect 150862 462 151216 490
rect 151280 598 151450 626
rect 150806 439 150862 448
rect 151280 354 151308 598
rect 151832 626 151860 700
rect 153028 728 153056 1108
rect 153580 1057 153608 1108
rect 153382 1048 153438 1057
rect 153566 1048 153622 1057
rect 153438 1006 153516 1034
rect 153382 983 153438 992
rect 153488 814 153516 1006
rect 153566 983 153622 992
rect 153476 808 153528 814
rect 153672 796 153700 1176
rect 153844 1158 153896 1164
rect 154132 950 154160 1255
rect 157432 1284 157484 1290
rect 156472 1244 157432 1272
rect 156420 1226 156472 1232
rect 157522 1255 157578 1264
rect 157432 1226 157484 1232
rect 157536 1154 157564 1255
rect 157904 1193 157932 1516
rect 157984 1498 158036 1504
rect 157982 1456 158038 1465
rect 157982 1391 158038 1400
rect 158166 1456 158222 1465
rect 158166 1391 158222 1400
rect 157890 1184 157946 1193
rect 154212 1148 154264 1154
rect 157524 1148 157576 1154
rect 154264 1108 156644 1136
rect 154212 1090 154264 1096
rect 154316 1006 155264 1034
rect 154120 944 154172 950
rect 154120 886 154172 892
rect 154316 796 154344 1006
rect 154396 944 154448 950
rect 154396 886 154448 892
rect 155132 944 155184 950
rect 155132 886 155184 892
rect 153672 768 154344 796
rect 153476 750 153528 756
rect 152240 700 153056 728
rect 153568 740 153620 746
rect 152188 682 152240 688
rect 154408 728 154436 886
rect 153568 682 153620 688
rect 153672 700 154436 728
rect 153580 626 153608 682
rect 151832 598 153608 626
rect 151450 575 151506 584
rect 153672 490 153700 700
rect 155144 626 155172 886
rect 155236 728 155264 1006
rect 156616 932 156644 1108
rect 157076 1108 157380 1136
rect 157076 1057 157104 1108
rect 157062 1048 157118 1057
rect 157246 1048 157302 1057
rect 157062 983 157118 992
rect 157168 1006 157246 1034
rect 157168 932 157196 1006
rect 157246 983 157302 992
rect 156616 904 157196 932
rect 157352 932 157380 1108
rect 157996 1170 158024 1391
rect 158180 1290 158208 1391
rect 158168 1284 158220 1290
rect 158168 1226 158220 1232
rect 158628 1284 158680 1290
rect 158628 1226 158680 1232
rect 158812 1284 158864 1290
rect 158812 1226 158864 1232
rect 158640 1193 158668 1226
rect 158074 1184 158130 1193
rect 157996 1142 158074 1170
rect 157890 1119 157946 1128
rect 158074 1119 158130 1128
rect 158442 1184 158498 1193
rect 158442 1119 158444 1128
rect 157524 1090 157576 1096
rect 158496 1119 158498 1128
rect 158626 1184 158682 1193
rect 158626 1119 158682 1128
rect 158444 1090 158496 1096
rect 157352 904 157932 932
rect 156800 746 157840 762
rect 156604 740 156656 746
rect 155236 700 156604 728
rect 156604 682 156656 688
rect 156788 740 157840 746
rect 156840 734 157840 740
rect 156788 682 156840 688
rect 157812 678 157840 734
rect 157340 672 157392 678
rect 157154 640 157210 649
rect 150636 326 151308 354
rect 151360 264 151412 270
rect 150990 232 151046 241
rect 151046 212 151360 218
rect 151046 206 151412 212
rect 151046 190 151400 206
rect 150990 167 151046 176
rect 151514 -960 151626 480
rect 151728 264 151780 270
rect 151818 232 151874 241
rect 151780 212 151818 218
rect 151728 206 151818 212
rect 151740 190 151818 206
rect 151818 167 151874 176
rect 152710 -960 152822 480
rect 153120 462 153700 490
rect 153764 598 154160 626
rect 155144 598 157154 626
rect 153120 377 153148 462
rect 153764 406 153792 598
rect 153200 400 153252 406
rect 153106 368 153162 377
rect 153752 400 153804 406
rect 153290 368 153346 377
rect 153252 348 153290 354
rect 153200 342 153290 348
rect 153212 326 153290 342
rect 153106 303 153162 312
rect 153752 342 153804 348
rect 153290 303 153346 312
rect 153906 -960 154018 480
rect 154132 388 154160 598
rect 157616 672 157668 678
rect 157340 614 157392 620
rect 157614 640 157616 649
rect 157800 672 157852 678
rect 157668 640 157670 649
rect 157154 575 157210 584
rect 156878 504 156934 513
rect 154672 400 154724 406
rect 154132 360 154672 388
rect 154672 342 154724 348
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157154 504 157210 513
rect 156934 462 157154 490
rect 156878 439 156934 448
rect 157154 439 157210 448
rect 157248 400 157300 406
rect 156878 368 156934 377
rect 156934 348 157248 354
rect 157352 377 157380 614
rect 157904 649 157932 904
rect 158824 728 158852 1226
rect 158916 796 158944 1634
rect 159008 1465 159036 1663
rect 159364 1624 159416 1630
rect 159364 1566 159416 1572
rect 158994 1456 159050 1465
rect 158994 1391 159050 1400
rect 159376 1329 159404 1566
rect 159652 1465 159680 1686
rect 160282 1592 160338 1601
rect 161202 1592 161258 1601
rect 160940 1562 161202 1578
rect 160282 1527 160284 1536
rect 160336 1527 160338 1536
rect 160928 1556 161202 1562
rect 160284 1498 160336 1504
rect 160980 1550 161202 1556
rect 161202 1527 161258 1536
rect 160928 1498 160980 1504
rect 159638 1456 159694 1465
rect 159638 1391 159694 1400
rect 159362 1320 159418 1329
rect 159546 1320 159602 1329
rect 159362 1255 159418 1264
rect 159456 1284 159508 1290
rect 159546 1255 159602 1264
rect 159456 1226 159508 1232
rect 159468 1193 159496 1226
rect 159270 1184 159326 1193
rect 159270 1119 159326 1128
rect 159454 1184 159510 1193
rect 159454 1119 159510 1128
rect 159284 1068 159312 1119
rect 159560 1068 159588 1255
rect 161112 1216 161164 1222
rect 161296 1216 161348 1222
rect 161164 1164 161296 1170
rect 161112 1158 161348 1164
rect 161400 1170 161428 1686
rect 162044 1584 164004 1612
rect 161846 1320 161902 1329
rect 162044 1306 162072 1584
rect 161902 1278 162072 1306
rect 162320 1516 163820 1544
rect 162320 1290 162348 1516
rect 162860 1420 162912 1426
rect 162860 1362 162912 1368
rect 162308 1284 162360 1290
rect 161846 1255 161902 1264
rect 162872 1272 162900 1362
rect 163792 1329 163820 1516
rect 163976 1442 164004 1584
rect 164238 1456 164294 1465
rect 163976 1414 164238 1442
rect 164238 1391 164294 1400
rect 163778 1320 163834 1329
rect 163688 1284 163740 1290
rect 162872 1244 163688 1272
rect 162308 1226 162360 1232
rect 163778 1255 163834 1264
rect 163688 1226 163740 1232
rect 166368 1193 166396 1720
rect 166814 1728 166870 1737
rect 166814 1663 166870 1672
rect 169114 1728 169170 1737
rect 169484 1702 169536 1708
rect 170956 1760 171008 1766
rect 170956 1702 171008 1708
rect 171048 1760 171100 1766
rect 174268 1760 174320 1766
rect 171048 1702 171100 1708
rect 171520 1720 174268 1748
rect 169114 1663 169116 1672
rect 166460 1516 166764 1544
rect 166354 1184 166410 1193
rect 160560 1148 160612 1154
rect 161020 1148 161072 1154
rect 160612 1108 161020 1136
rect 160560 1090 160612 1096
rect 161124 1142 161336 1158
rect 161400 1142 163452 1170
rect 161020 1090 161072 1096
rect 159284 1040 159588 1068
rect 159284 972 161428 1000
rect 159284 796 159312 972
rect 158916 768 159312 796
rect 159376 870 160876 898
rect 159376 728 159404 870
rect 160848 814 160876 870
rect 160836 808 160888 814
rect 160836 750 160888 756
rect 160744 740 160796 746
rect 158824 700 159404 728
rect 159836 700 160744 728
rect 159456 672 159508 678
rect 157800 614 157852 620
rect 157890 640 157946 649
rect 157614 575 157670 584
rect 158074 640 158130 649
rect 157890 575 157946 584
rect 157996 598 158074 626
rect 156934 342 157300 348
rect 157338 368 157394 377
rect 156934 326 157288 342
rect 156878 303 156934 312
rect 157338 303 157394 312
rect 157494 -960 157606 480
rect 157996 388 158024 598
rect 159836 626 159864 700
rect 160744 682 160796 688
rect 159508 620 159864 626
rect 159456 614 159864 620
rect 160928 672 160980 678
rect 160980 620 161336 626
rect 160928 614 161336 620
rect 159468 598 159864 614
rect 160940 598 161336 614
rect 158074 575 158130 584
rect 157812 377 158024 388
rect 157798 368 158024 377
rect 157854 360 158024 368
rect 157798 303 157854 312
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 161308 218 161336 598
rect 161400 377 161428 972
rect 162584 944 162636 950
rect 163424 932 163452 1142
rect 166354 1119 166410 1128
rect 166460 1068 166488 1516
rect 163700 1057 166488 1068
rect 163686 1048 166488 1057
rect 163742 1040 166488 1048
rect 166630 1048 166686 1057
rect 163686 983 163742 992
rect 166736 1034 166764 1516
rect 166828 1426 166856 1663
rect 169168 1663 169170 1672
rect 169116 1634 169168 1640
rect 167288 1516 167500 1544
rect 167288 1426 167316 1516
rect 166816 1420 166868 1426
rect 166816 1362 166868 1368
rect 167276 1420 167328 1426
rect 167276 1362 167328 1368
rect 167368 1420 167420 1426
rect 167368 1362 167420 1368
rect 166920 1154 167210 1170
rect 166908 1148 167210 1154
rect 166960 1142 167210 1148
rect 166908 1090 166960 1096
rect 166814 1048 166870 1057
rect 166736 1006 166814 1034
rect 166630 983 166686 992
rect 166814 983 166870 992
rect 162636 904 163360 932
rect 163424 904 166304 932
rect 162584 886 162636 892
rect 161478 776 161534 785
rect 161754 776 161810 785
rect 161534 734 161754 762
rect 161478 711 161534 720
rect 161754 711 161810 720
rect 163134 776 163190 785
rect 163190 746 163268 762
rect 163190 740 163280 746
rect 163190 734 163228 740
rect 163134 711 163190 720
rect 163228 682 163280 688
rect 163136 672 163188 678
rect 161754 640 161810 649
rect 161492 598 161754 626
rect 161386 368 161442 377
rect 161386 303 161442 312
rect 161492 218 161520 598
rect 163136 614 163188 620
rect 161754 575 161810 584
rect 161308 190 161520 218
rect 162278 -960 162390 480
rect 163148 377 163176 614
rect 163332 377 163360 904
rect 163700 836 164004 864
rect 163700 785 163728 836
rect 163686 776 163742 785
rect 163686 711 163742 720
rect 163870 776 163926 785
rect 163976 746 164004 836
rect 163870 711 163872 720
rect 163924 711 163926 720
rect 163964 740 164016 746
rect 163872 682 163924 688
rect 163964 682 164016 688
rect 166172 672 166224 678
rect 163502 640 163558 649
rect 164068 632 166172 660
rect 164068 626 164096 632
rect 163558 598 164096 626
rect 166172 614 166224 620
rect 163502 575 163558 584
rect 166276 524 166304 904
rect 166644 678 166672 983
rect 166632 672 166684 678
rect 167380 660 167408 1362
rect 166632 614 166684 620
rect 166736 632 167408 660
rect 167472 660 167500 1516
rect 168944 1516 169340 1544
rect 168944 1329 168972 1516
rect 169022 1456 169078 1465
rect 169022 1391 169078 1400
rect 169206 1456 169262 1465
rect 169206 1391 169208 1400
rect 168930 1320 168986 1329
rect 168930 1255 168986 1264
rect 168654 1184 168710 1193
rect 169036 1154 169064 1391
rect 169260 1391 169262 1400
rect 169208 1362 169260 1368
rect 169114 1320 169170 1329
rect 169114 1255 169170 1264
rect 168654 1119 168710 1128
rect 169024 1148 169076 1154
rect 168668 1034 168696 1119
rect 169024 1090 169076 1096
rect 169128 1034 169156 1255
rect 169312 1068 169340 1516
rect 169392 1488 169444 1494
rect 169392 1430 169444 1436
rect 169496 1442 169524 1702
rect 169576 1692 169628 1698
rect 169576 1634 169628 1640
rect 169588 1544 169616 1634
rect 169852 1556 169904 1562
rect 169588 1516 169852 1544
rect 169852 1498 169904 1504
rect 169404 1193 169432 1430
rect 169496 1414 170904 1442
rect 170770 1320 170826 1329
rect 169944 1284 169996 1290
rect 170508 1278 170770 1306
rect 169996 1244 170444 1272
rect 169944 1226 169996 1232
rect 169390 1184 169446 1193
rect 169574 1184 169630 1193
rect 169390 1119 169446 1128
rect 169496 1142 169574 1170
rect 169496 1068 169524 1142
rect 169574 1119 169630 1128
rect 169312 1040 169524 1068
rect 168668 1006 169156 1034
rect 170416 898 170444 1244
rect 170508 1193 170536 1278
rect 170770 1255 170826 1264
rect 170494 1184 170550 1193
rect 170494 1119 170550 1128
rect 170876 1034 170904 1414
rect 170968 1306 170996 1702
rect 171060 1601 171088 1702
rect 171046 1592 171102 1601
rect 171046 1527 171102 1536
rect 171520 1494 171548 1720
rect 174268 1702 174320 1708
rect 175280 1760 175332 1766
rect 177856 1760 177908 1766
rect 175332 1720 175412 1748
rect 175280 1702 175332 1708
rect 171598 1592 171654 1601
rect 171598 1527 171654 1536
rect 175384 1544 175412 1720
rect 177500 1720 177856 1748
rect 171508 1488 171560 1494
rect 171508 1430 171560 1436
rect 171612 1442 171640 1527
rect 175384 1516 177252 1544
rect 173346 1456 173402 1465
rect 171612 1414 173346 1442
rect 173346 1391 173402 1400
rect 173624 1420 173676 1426
rect 173624 1362 173676 1368
rect 173636 1306 173664 1362
rect 170968 1278 173664 1306
rect 173806 1320 173862 1329
rect 176016 1284 176068 1290
rect 173862 1264 176016 1272
rect 173806 1255 176016 1264
rect 173820 1244 176016 1255
rect 176016 1226 176068 1232
rect 173254 1184 173310 1193
rect 176290 1184 176346 1193
rect 173310 1142 176290 1170
rect 173254 1119 173310 1128
rect 176290 1119 176346 1128
rect 177118 1184 177174 1193
rect 177118 1119 177174 1128
rect 170876 1006 176686 1034
rect 169496 870 169984 898
rect 170416 870 176148 898
rect 169496 814 169524 870
rect 169484 808 169536 814
rect 169484 750 169536 756
rect 169668 740 169720 746
rect 169668 682 169720 688
rect 167472 632 169616 660
rect 169680 649 169708 682
rect 166736 524 166764 632
rect 166276 496 166764 524
rect 169588 524 169616 632
rect 169666 640 169722 649
rect 169850 640 169906 649
rect 169666 575 169722 584
rect 169772 598 169850 626
rect 169772 524 169800 598
rect 169956 626 169984 870
rect 175648 808 175700 814
rect 175648 750 175700 756
rect 176014 776 176070 785
rect 170034 640 170090 649
rect 169956 598 170034 626
rect 169850 575 169906 584
rect 170034 575 170090 584
rect 169588 496 169800 524
rect 163134 368 163190 377
rect 163134 303 163190 312
rect 163318 368 163374 377
rect 163318 303 163374 312
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 175660 218 175688 750
rect 175924 740 175976 746
rect 176120 762 176148 870
rect 176198 776 176254 785
rect 176120 734 176198 762
rect 176014 711 176016 720
rect 175924 682 175976 688
rect 176068 711 176070 720
rect 176198 711 176254 720
rect 176016 682 176068 688
rect 175936 610 175964 682
rect 177132 678 177160 1119
rect 176108 672 176160 678
rect 176660 672 176712 678
rect 176160 632 176332 660
rect 176108 614 176160 620
rect 175924 604 175976 610
rect 175924 546 175976 552
rect 175740 536 175792 542
rect 176200 536 176252 542
rect 176028 496 176200 524
rect 176028 490 176056 496
rect 175792 484 176056 490
rect 175740 478 176056 484
rect 176200 478 176252 484
rect 175752 462 176056 478
rect 176304 406 176332 632
rect 176396 632 176660 660
rect 176292 400 176344 406
rect 176292 342 176344 348
rect 176396 218 176424 632
rect 176660 614 176712 620
rect 177120 672 177172 678
rect 177120 614 177172 620
rect 177224 626 177252 1516
rect 177500 1426 177528 1720
rect 183744 1760 183796 1766
rect 177856 1702 177908 1708
rect 178774 1728 178830 1737
rect 178774 1663 178830 1672
rect 179050 1728 179106 1737
rect 179616 1720 183744 1748
rect 179050 1663 179052 1672
rect 178788 1630 178816 1663
rect 179104 1663 179106 1672
rect 179144 1692 179196 1698
rect 179052 1634 179104 1640
rect 179144 1634 179196 1640
rect 179328 1692 179380 1698
rect 179512 1692 179564 1698
rect 179380 1652 179512 1680
rect 179328 1634 179380 1640
rect 179512 1634 179564 1640
rect 178684 1624 178736 1630
rect 177670 1592 177726 1601
rect 177726 1550 178448 1578
rect 178684 1566 178736 1572
rect 178776 1624 178828 1630
rect 178776 1566 178828 1572
rect 177670 1527 177726 1536
rect 177856 1488 177908 1494
rect 177908 1448 178172 1476
rect 177856 1430 177908 1436
rect 177488 1420 177540 1426
rect 177488 1362 177540 1368
rect 177762 1320 177818 1329
rect 177672 1284 177724 1290
rect 177762 1255 177818 1264
rect 178038 1320 178094 1329
rect 178144 1290 178172 1448
rect 178314 1456 178370 1465
rect 178314 1391 178370 1400
rect 178038 1255 178040 1264
rect 177672 1226 177724 1232
rect 177684 1193 177712 1226
rect 177670 1184 177726 1193
rect 177670 1119 177726 1128
rect 177776 882 177804 1255
rect 178092 1255 178094 1264
rect 178132 1284 178184 1290
rect 178040 1226 178092 1232
rect 178132 1226 178184 1232
rect 177580 876 177632 882
rect 177580 818 177632 824
rect 177764 876 177816 882
rect 177764 818 177816 824
rect 177592 762 177620 818
rect 177592 734 178080 762
rect 178328 746 178356 1391
rect 178420 1034 178448 1550
rect 178696 1465 178724 1566
rect 178682 1456 178738 1465
rect 178682 1391 178738 1400
rect 179156 1306 179184 1634
rect 178972 1278 179184 1306
rect 178972 1222 179000 1278
rect 178960 1216 179012 1222
rect 179236 1216 179288 1222
rect 179156 1193 179236 1204
rect 178960 1158 179012 1164
rect 179142 1184 179236 1193
rect 179198 1176 179236 1184
rect 179236 1158 179288 1164
rect 179326 1184 179382 1193
rect 179142 1119 179198 1128
rect 179326 1119 179382 1128
rect 179340 1034 179368 1119
rect 178420 1006 179368 1034
rect 179616 882 179644 1720
rect 190368 1760 190420 1766
rect 190012 1720 190368 1748
rect 183744 1702 183796 1708
rect 183848 1686 184244 1714
rect 179878 1592 179934 1601
rect 181718 1592 181774 1601
rect 179878 1527 179934 1536
rect 180076 1550 181116 1578
rect 179892 1426 179920 1527
rect 179788 1420 179840 1426
rect 179788 1362 179840 1368
rect 179880 1420 179932 1426
rect 179880 1362 179932 1368
rect 179694 1320 179750 1329
rect 179800 1306 179828 1362
rect 180076 1306 180104 1550
rect 181088 1476 181116 1550
rect 183848 1578 183876 1686
rect 184216 1630 184244 1686
rect 184308 1652 184796 1680
rect 181774 1550 183876 1578
rect 183928 1624 183980 1630
rect 183928 1566 183980 1572
rect 184204 1624 184256 1630
rect 184204 1566 184256 1572
rect 181718 1527 181774 1536
rect 182640 1488 182692 1494
rect 181088 1448 182640 1476
rect 183940 1476 183968 1566
rect 184308 1476 184336 1652
rect 184662 1592 184718 1601
rect 184662 1527 184718 1536
rect 182640 1430 182692 1436
rect 183742 1456 183798 1465
rect 179800 1278 180104 1306
rect 180168 1380 181024 1408
rect 183940 1448 184336 1476
rect 184386 1456 184442 1465
rect 183798 1400 184386 1408
rect 183742 1391 184442 1400
rect 183756 1380 184428 1391
rect 179694 1255 179750 1264
rect 179708 882 179736 1255
rect 179604 876 179656 882
rect 179604 818 179656 824
rect 179696 876 179748 882
rect 179696 818 179748 824
rect 180168 746 180196 1380
rect 180246 1320 180302 1329
rect 180246 1255 180302 1264
rect 180260 746 180288 1255
rect 180628 1244 180932 1272
rect 180628 882 180656 1244
rect 180798 1184 180854 1193
rect 180798 1119 180854 1128
rect 180616 876 180668 882
rect 180616 818 180668 824
rect 180708 876 180760 882
rect 180708 818 180760 824
rect 177948 672 178000 678
rect 177394 640 177450 649
rect 177224 598 177394 626
rect 177394 575 177450 584
rect 177946 640 177948 649
rect 178000 640 178002 649
rect 177946 575 178002 584
rect 178052 524 178080 734
rect 178316 740 178368 746
rect 178316 682 178368 688
rect 180156 740 180208 746
rect 180156 682 180208 688
rect 180248 740 180300 746
rect 180248 682 180300 688
rect 180720 592 180748 818
rect 180812 796 180840 1119
rect 180904 864 180932 1244
rect 180996 1170 181024 1380
rect 182638 1320 182694 1329
rect 182694 1278 184060 1306
rect 182638 1255 182694 1264
rect 183928 1216 183980 1222
rect 182914 1184 182970 1193
rect 180996 1142 182914 1170
rect 183928 1158 183980 1164
rect 184032 1170 184060 1278
rect 184202 1184 184258 1193
rect 182914 1119 182970 1128
rect 183940 1057 183968 1158
rect 184032 1142 184202 1170
rect 184202 1119 184258 1128
rect 183926 1048 183982 1057
rect 183926 983 183982 992
rect 184294 1048 184350 1057
rect 184350 1006 184520 1034
rect 184294 983 184350 992
rect 183572 870 184336 898
rect 183572 864 183600 870
rect 180904 836 183600 864
rect 183744 808 183796 814
rect 180812 768 183744 796
rect 183744 750 183796 756
rect 184202 776 184258 785
rect 184020 740 184072 746
rect 183940 700 184020 728
rect 183560 672 183612 678
rect 178420 564 180748 592
rect 183480 632 183560 660
rect 178420 524 178448 564
rect 178052 496 178448 524
rect 175660 190 176424 218
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183480 202 183508 632
rect 183560 614 183612 620
rect 183468 196 183520 202
rect 183468 138 183520 144
rect 183714 -960 183826 480
rect 183940 202 183968 700
rect 184308 762 184336 870
rect 184386 776 184442 785
rect 184308 734 184386 762
rect 184202 711 184258 720
rect 184492 762 184520 1006
rect 184676 898 184704 1527
rect 184768 1272 184796 1652
rect 190012 1562 190040 1720
rect 191012 1760 191064 1766
rect 190368 1702 190420 1708
rect 190642 1728 190698 1737
rect 190918 1728 190974 1737
rect 190698 1686 190776 1714
rect 190642 1663 190698 1672
rect 190642 1592 190698 1601
rect 190564 1562 190642 1578
rect 189908 1556 189960 1562
rect 189908 1498 189960 1504
rect 190000 1556 190052 1562
rect 190000 1498 190052 1504
rect 190092 1556 190144 1562
rect 190092 1498 190144 1504
rect 190552 1556 190642 1562
rect 190604 1550 190642 1556
rect 190642 1527 190698 1536
rect 190552 1498 190604 1504
rect 189920 1442 189948 1498
rect 190104 1442 190132 1498
rect 189920 1414 190132 1442
rect 190368 1488 190420 1494
rect 190368 1430 190420 1436
rect 190184 1352 190236 1358
rect 189630 1320 189686 1329
rect 184768 1244 186360 1272
rect 190012 1312 190184 1340
rect 190012 1306 190040 1312
rect 189686 1278 190040 1306
rect 190184 1294 190236 1300
rect 189630 1255 189686 1264
rect 185858 1184 185914 1193
rect 186332 1170 186360 1244
rect 189448 1216 189500 1222
rect 186502 1184 186558 1193
rect 185914 1142 186254 1170
rect 186332 1142 186502 1170
rect 185858 1119 185914 1128
rect 190380 1193 190408 1430
rect 190552 1216 190604 1222
rect 189448 1158 189500 1164
rect 190366 1184 190422 1193
rect 186502 1119 186558 1128
rect 189460 1034 189488 1158
rect 190366 1119 190422 1128
rect 190472 1176 190552 1204
rect 189906 1048 189962 1057
rect 189460 1006 189906 1034
rect 189906 983 189962 992
rect 190472 898 190500 1176
rect 190552 1158 190604 1164
rect 184676 870 190500 898
rect 190748 898 190776 1686
rect 191012 1702 191064 1708
rect 191196 1760 191248 1766
rect 191748 1760 191800 1766
rect 191248 1720 191748 1748
rect 191196 1702 191248 1708
rect 233516 1760 233568 1766
rect 191748 1702 191800 1708
rect 192206 1728 192262 1737
rect 190918 1663 190974 1672
rect 190932 1465 190960 1663
rect 191024 1578 191052 1702
rect 196438 1728 196494 1737
rect 192262 1686 192340 1714
rect 192206 1663 192262 1672
rect 192312 1578 192340 1686
rect 196438 1663 196494 1672
rect 196714 1728 196770 1737
rect 198738 1728 198794 1737
rect 196714 1663 196770 1672
rect 198476 1686 198738 1714
rect 195978 1592 196034 1601
rect 191024 1550 191788 1578
rect 191012 1488 191064 1494
rect 190918 1456 190974 1465
rect 191012 1430 191064 1436
rect 191288 1488 191340 1494
rect 191656 1488 191708 1494
rect 191340 1448 191656 1476
rect 191288 1430 191340 1436
rect 191760 1476 191788 1550
rect 191944 1550 192248 1578
rect 192312 1550 195730 1578
rect 195808 1550 195978 1578
rect 191840 1488 191892 1494
rect 191760 1448 191840 1476
rect 191656 1430 191708 1436
rect 191840 1430 191892 1436
rect 190918 1391 190974 1400
rect 190828 1352 190880 1358
rect 190828 1294 190880 1300
rect 190840 1193 190868 1294
rect 190920 1216 190972 1222
rect 190826 1184 190882 1193
rect 190920 1158 190972 1164
rect 191024 1170 191052 1430
rect 191472 1352 191524 1358
rect 191116 1329 191472 1340
rect 191102 1320 191472 1329
rect 191158 1312 191472 1320
rect 191472 1294 191524 1300
rect 191102 1255 191158 1264
rect 191562 1184 191618 1193
rect 190826 1119 190882 1128
rect 190932 1034 190960 1158
rect 191024 1142 191562 1170
rect 191562 1119 191618 1128
rect 191378 1048 191434 1057
rect 190932 1006 191378 1034
rect 191378 983 191434 992
rect 191944 898 191972 1550
rect 192116 1488 192168 1494
rect 192116 1430 192168 1436
rect 190748 870 191972 898
rect 192128 796 192156 1430
rect 190458 776 190514 785
rect 184492 734 190458 762
rect 184386 711 184442 720
rect 191576 768 192156 796
rect 192220 796 192248 1550
rect 195244 1352 195296 1358
rect 195244 1294 195296 1300
rect 195256 898 195284 1294
rect 195808 898 195836 1550
rect 195978 1527 196034 1536
rect 195256 870 195836 898
rect 196452 898 196480 1663
rect 196532 1488 196584 1494
rect 196532 1430 196584 1436
rect 196544 1034 196572 1430
rect 196728 1193 196756 1663
rect 197820 1556 197872 1562
rect 197872 1516 198320 1544
rect 197820 1498 197872 1504
rect 196992 1488 197044 1494
rect 196820 1448 196992 1476
rect 196714 1184 196770 1193
rect 196714 1119 196770 1128
rect 196820 1034 196848 1448
rect 196992 1430 197044 1436
rect 197268 1352 197320 1358
rect 197268 1294 197320 1300
rect 196544 1006 196848 1034
rect 197174 1048 197230 1057
rect 197280 1034 197308 1294
rect 198094 1184 198150 1193
rect 198292 1170 198320 1516
rect 198476 1358 198504 1686
rect 200026 1728 200082 1737
rect 198738 1663 198794 1672
rect 198844 1686 200026 1714
rect 198556 1556 198608 1562
rect 198844 1544 198872 1686
rect 207294 1728 207350 1737
rect 200026 1663 200082 1672
rect 200132 1652 204576 1680
rect 208122 1728 208178 1737
rect 207350 1686 208122 1714
rect 207294 1663 207350 1672
rect 216678 1728 216734 1737
rect 208122 1663 208178 1672
rect 198608 1516 198872 1544
rect 199106 1592 199162 1601
rect 199106 1527 199108 1536
rect 198556 1498 198608 1504
rect 199160 1527 199162 1536
rect 199750 1592 199806 1601
rect 200132 1578 200160 1652
rect 204442 1592 204498 1601
rect 199806 1550 200160 1578
rect 200224 1550 200344 1578
rect 199750 1527 199806 1536
rect 199108 1498 199160 1504
rect 200224 1494 200252 1550
rect 200316 1544 200344 1550
rect 200316 1536 204442 1544
rect 200316 1527 204498 1536
rect 200316 1516 204484 1527
rect 204548 1494 204576 1652
rect 208964 1652 211476 1680
rect 220450 1728 220506 1737
rect 216734 1698 216812 1714
rect 220188 1698 220450 1714
rect 216734 1692 216824 1698
rect 216734 1686 216772 1692
rect 216678 1663 216734 1672
rect 204810 1592 204866 1601
rect 204628 1556 204680 1562
rect 205454 1592 205510 1601
rect 204810 1527 204866 1536
rect 205284 1550 205454 1578
rect 204628 1498 204680 1504
rect 200212 1488 200264 1494
rect 204536 1488 204588 1494
rect 200212 1430 200264 1436
rect 200302 1456 200358 1465
rect 200358 1414 203196 1442
rect 204536 1430 204588 1436
rect 200302 1391 200358 1400
rect 198464 1352 198516 1358
rect 198464 1294 198516 1300
rect 199200 1352 199252 1358
rect 202972 1352 203024 1358
rect 199252 1312 202972 1340
rect 199200 1294 199252 1300
rect 202972 1294 203024 1300
rect 198292 1142 198504 1170
rect 198094 1119 198150 1128
rect 197230 1006 197308 1034
rect 198108 1034 198136 1119
rect 198370 1048 198426 1057
rect 198108 1006 198370 1034
rect 197174 983 197230 992
rect 198476 1034 198504 1142
rect 198476 1006 198780 1034
rect 198370 983 198426 992
rect 197726 912 197782 921
rect 196452 870 197032 898
rect 192220 768 193720 796
rect 191576 728 191604 768
rect 193692 762 193720 768
rect 193692 734 194640 762
rect 190458 711 190514 720
rect 184020 682 184072 688
rect 184216 626 184244 711
rect 190564 700 191144 728
rect 190564 660 190592 700
rect 187804 632 190592 660
rect 187804 626 187832 632
rect 184216 598 187832 626
rect 190656 598 191052 626
rect 184020 536 184072 542
rect 190656 513 190684 598
rect 184020 478 184072 484
rect 190642 504 190698 513
rect 184032 338 184060 478
rect 184020 332 184072 338
rect 184020 274 184072 280
rect 183928 196 183980 202
rect 183928 138 183980 144
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190642 439 190698 448
rect 190798 -960 190910 480
rect 191024 252 191052 598
rect 191116 388 191144 700
rect 191300 700 191604 728
rect 191668 700 193628 728
rect 191300 513 191328 700
rect 191668 626 191696 700
rect 191392 598 191696 626
rect 191852 598 193444 626
rect 191286 504 191342 513
rect 191286 439 191342 448
rect 191392 388 191420 598
rect 191116 360 191420 388
rect 191852 252 191880 598
rect 191024 224 191880 252
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 193416 456 193444 598
rect 193496 468 193548 474
rect 193416 428 193496 456
rect 193496 410 193548 416
rect 193600 406 193628 700
rect 194612 660 194640 734
rect 194612 632 195836 660
rect 193588 400 193640 406
rect 193588 342 193640 348
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 195808 388 195836 632
rect 196624 400 196676 406
rect 195808 360 196624 388
rect 196624 342 196676 348
rect 196778 -960 196890 480
rect 197004 406 197032 870
rect 198186 912 198242 921
rect 197782 870 198186 898
rect 197726 847 197782 856
rect 198186 847 198242 856
rect 197542 776 197598 785
rect 198646 776 198702 785
rect 197598 734 197676 762
rect 197542 711 197598 720
rect 197358 640 197414 649
rect 197358 575 197414 584
rect 196992 400 197044 406
rect 197372 388 197400 575
rect 197648 513 197676 734
rect 198646 711 198702 720
rect 198462 640 198518 649
rect 197740 598 198462 626
rect 197634 504 197690 513
rect 197634 439 197690 448
rect 197740 388 197768 598
rect 198462 575 198518 584
rect 198186 504 198242 513
rect 197372 360 197768 388
rect 196992 342 197044 348
rect 197974 -960 198086 480
rect 198186 439 198242 448
rect 198370 504 198426 513
rect 198370 439 198372 448
rect 198200 406 198228 439
rect 198424 439 198426 448
rect 198464 468 198516 474
rect 198372 410 198424 416
rect 198464 410 198516 416
rect 198188 400 198240 406
rect 198188 342 198240 348
rect 198280 400 198332 406
rect 198280 342 198332 348
rect 198476 354 198504 410
rect 198660 354 198688 711
rect 198752 474 198780 1006
rect 198844 598 202920 626
rect 198740 468 198792 474
rect 198740 410 198792 416
rect 198292 82 198320 342
rect 198476 326 198688 354
rect 198370 232 198426 241
rect 198554 232 198610 241
rect 198426 190 198554 218
rect 198370 167 198426 176
rect 198554 167 198610 176
rect 198844 82 198872 598
rect 198292 54 198872 82
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 202892 354 202920 598
rect 203168 474 203196 1414
rect 204640 1306 204668 1498
rect 204824 1494 204852 1527
rect 204812 1488 204864 1494
rect 204812 1430 204864 1436
rect 204272 1278 204668 1306
rect 204272 649 204300 1278
rect 204364 1006 205206 1034
rect 204364 678 204392 1006
rect 205284 898 205312 1550
rect 205454 1527 205510 1536
rect 207294 1592 207350 1601
rect 207294 1527 207350 1536
rect 207478 1592 207534 1601
rect 207534 1550 207888 1578
rect 207478 1527 207534 1536
rect 207308 1442 207336 1527
rect 207754 1456 207810 1465
rect 207308 1414 207754 1442
rect 207754 1391 207810 1400
rect 204548 870 205312 898
rect 204352 672 204404 678
rect 204258 640 204314 649
rect 203260 598 204116 626
rect 203156 468 203208 474
rect 203156 410 203208 416
rect 203260 354 203288 598
rect 204088 490 204116 598
rect 204548 649 204576 870
rect 207860 796 207888 1550
rect 208030 1320 208086 1329
rect 208030 1255 208086 1264
rect 204640 768 207888 796
rect 208044 796 208072 1255
rect 208964 1068 208992 1652
rect 211342 1592 211398 1601
rect 211342 1527 211398 1536
rect 211356 1494 211384 1527
rect 211344 1488 211396 1494
rect 209884 1414 211292 1442
rect 211344 1430 211396 1436
rect 211448 1442 211476 1652
rect 220176 1692 220450 1698
rect 216772 1634 216824 1640
rect 216876 1652 218652 1680
rect 214196 1624 214248 1630
rect 212552 1584 214196 1612
rect 212170 1456 212226 1465
rect 211448 1414 212170 1442
rect 209884 1329 209912 1414
rect 211160 1352 211212 1358
rect 209870 1320 209926 1329
rect 209056 1278 209360 1306
rect 209056 1193 209084 1278
rect 209042 1184 209098 1193
rect 209042 1119 209098 1128
rect 209226 1184 209282 1193
rect 209332 1170 209360 1278
rect 211160 1294 211212 1300
rect 211264 1306 211292 1414
rect 212170 1391 212226 1400
rect 212552 1306 212580 1584
rect 214196 1566 214248 1572
rect 214472 1624 214524 1630
rect 214932 1624 214984 1630
rect 214472 1566 214524 1572
rect 214852 1584 214932 1612
rect 214378 1456 214434 1465
rect 214484 1442 214512 1566
rect 214434 1414 214512 1442
rect 214378 1391 214434 1400
rect 209870 1255 209926 1264
rect 209502 1184 209558 1193
rect 209332 1142 209502 1170
rect 209226 1119 209282 1128
rect 209502 1119 209558 1128
rect 209240 1068 209268 1119
rect 208964 1040 209268 1068
rect 211172 1034 211200 1294
rect 211264 1278 212580 1306
rect 214380 1352 214432 1358
rect 214748 1352 214800 1358
rect 214432 1300 214682 1306
rect 214380 1294 214682 1300
rect 214852 1329 214880 1584
rect 214932 1566 214984 1572
rect 216588 1624 216640 1630
rect 216876 1578 216904 1652
rect 216640 1572 216904 1578
rect 216588 1566 216904 1572
rect 216600 1550 216904 1566
rect 217704 1584 218560 1612
rect 216770 1456 216826 1465
rect 216954 1456 217010 1465
rect 216826 1414 216954 1442
rect 216770 1391 216826 1400
rect 217704 1426 217732 1584
rect 218072 1516 218468 1544
rect 218072 1426 218100 1516
rect 218150 1456 218206 1465
rect 216954 1391 217010 1400
rect 217692 1420 217744 1426
rect 217692 1362 217744 1368
rect 218060 1420 218112 1426
rect 218206 1414 218376 1442
rect 218440 1426 218468 1516
rect 218150 1391 218206 1400
rect 218060 1362 218112 1368
rect 214748 1294 214800 1300
rect 214838 1320 214894 1329
rect 214392 1278 214682 1294
rect 211894 1184 211950 1193
rect 214760 1170 214788 1294
rect 215022 1320 215078 1329
rect 214838 1255 214894 1264
rect 214944 1278 215022 1306
rect 214944 1170 214972 1278
rect 215022 1255 215078 1264
rect 217414 1320 217470 1329
rect 217414 1255 217470 1264
rect 217966 1320 218022 1329
rect 218348 1306 218376 1414
rect 218428 1420 218480 1426
rect 218532 1408 218560 1584
rect 218624 1544 218652 1652
rect 220228 1686 220450 1692
rect 232134 1728 232190 1737
rect 220450 1663 220506 1672
rect 220176 1634 220228 1640
rect 224788 1652 225828 1680
rect 236552 1760 236604 1766
rect 234066 1728 234122 1737
rect 233568 1708 233726 1714
rect 233516 1702 233726 1708
rect 233528 1686 233726 1702
rect 232134 1663 232190 1672
rect 240140 1760 240192 1766
rect 236604 1720 238248 1748
rect 236552 1702 236604 1708
rect 234066 1663 234122 1672
rect 218624 1516 221688 1544
rect 218796 1420 218848 1426
rect 218532 1380 218796 1408
rect 218428 1362 218480 1368
rect 218796 1362 218848 1368
rect 221660 1329 221688 1516
rect 223946 1456 224002 1465
rect 223946 1391 224002 1400
rect 224498 1456 224554 1465
rect 224554 1414 224632 1442
rect 224498 1391 224554 1400
rect 221646 1320 221702 1329
rect 218348 1278 221596 1306
rect 217966 1255 218022 1264
rect 214760 1142 214972 1170
rect 217428 1170 217456 1255
rect 217874 1184 217930 1193
rect 217428 1142 217874 1170
rect 211950 1128 213960 1136
rect 211894 1119 213960 1128
rect 217980 1154 218008 1255
rect 217874 1119 217930 1128
rect 217968 1148 218020 1154
rect 211908 1108 213960 1119
rect 211172 1006 213868 1034
rect 208320 870 209452 898
rect 208216 808 208268 814
rect 208044 768 208216 796
rect 204352 614 204404 620
rect 204534 640 204590 649
rect 204258 575 204314 584
rect 204534 575 204590 584
rect 204640 490 204668 768
rect 208216 750 208268 756
rect 207756 672 207808 678
rect 205086 640 205142 649
rect 205142 598 207704 626
rect 207848 672 207900 678
rect 207756 614 207808 620
rect 207846 640 207848 649
rect 207900 640 207902 649
rect 205086 575 205142 584
rect 202892 326 203288 354
rect 203862 -960 203974 480
rect 204088 462 204668 490
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 207676 354 207704 598
rect 207768 490 207796 614
rect 207846 575 207902 584
rect 208320 490 208348 870
rect 209424 796 209452 870
rect 212092 870 213776 898
rect 209424 768 211568 796
rect 208596 734 209360 762
rect 208596 626 208624 734
rect 207768 462 208348 490
rect 208504 598 208624 626
rect 209332 626 209360 734
rect 211434 640 211490 649
rect 209332 598 211434 626
rect 208504 354 208532 598
rect 211434 575 211490 584
rect 207676 326 208532 354
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 211540 354 211568 768
rect 212092 728 212120 870
rect 212000 700 212120 728
rect 212000 474 212028 700
rect 213748 660 213776 870
rect 213840 814 213868 1006
rect 213932 898 213960 1108
rect 217968 1090 218020 1096
rect 214852 1006 220860 1034
rect 214852 898 214880 1006
rect 220832 898 220860 1006
rect 213932 870 214880 898
rect 217612 870 219664 898
rect 220832 870 221504 898
rect 213828 808 213880 814
rect 213828 750 213880 756
rect 217612 678 217640 870
rect 219348 808 219400 814
rect 219348 750 219400 756
rect 219440 808 219492 814
rect 219440 750 219492 756
rect 217704 700 217916 728
rect 214104 672 214156 678
rect 213748 632 214104 660
rect 212092 598 213684 626
rect 215024 672 215076 678
rect 215022 640 215024 649
rect 217600 672 217652 678
rect 215076 640 215078 649
rect 214104 614 214156 620
rect 211988 468 212040 474
rect 211988 410 212040 416
rect 212092 354 212120 598
rect 213656 524 213684 598
rect 214208 598 214880 626
rect 214208 524 214236 598
rect 213656 496 214236 524
rect 214852 524 214880 598
rect 215206 640 215262 649
rect 215022 575 215078 584
rect 215128 598 215206 626
rect 215128 524 215156 598
rect 217600 614 217652 620
rect 215206 575 215262 584
rect 217704 542 217732 700
rect 217782 640 217838 649
rect 217888 626 217916 700
rect 219360 649 219388 750
rect 219452 678 219480 750
rect 219636 678 219664 870
rect 221094 776 221150 785
rect 221094 711 221150 720
rect 221372 740 221424 746
rect 221108 678 221136 711
rect 221372 682 221424 688
rect 219440 672 219492 678
rect 217966 640 218022 649
rect 217888 598 217966 626
rect 217782 575 217838 584
rect 217966 575 218022 584
rect 219346 640 219402 649
rect 219440 614 219492 620
rect 219624 672 219676 678
rect 219624 614 219676 620
rect 221096 672 221148 678
rect 221384 649 221412 682
rect 221476 660 221504 870
rect 221568 796 221596 1278
rect 221646 1255 221702 1264
rect 223764 1148 223816 1154
rect 223764 1090 223816 1096
rect 223856 1148 223908 1154
rect 223960 1136 223988 1391
rect 224040 1148 224092 1154
rect 223960 1108 224040 1136
rect 223856 1090 223908 1096
rect 224040 1090 224092 1096
rect 223776 898 223804 1090
rect 223868 1034 223896 1090
rect 223868 1006 224250 1034
rect 223776 870 224540 898
rect 221568 768 224356 796
rect 224224 672 224276 678
rect 221096 614 221148 620
rect 221370 640 221426 649
rect 219346 575 219402 584
rect 221476 632 224224 660
rect 224224 614 224276 620
rect 221370 575 221426 584
rect 217796 542 217824 575
rect 214852 496 215156 524
rect 217508 536 217560 542
rect 211540 326 212120 354
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 217508 478 217560 484
rect 217692 536 217744 542
rect 217692 478 217744 484
rect 217784 536 217836 542
rect 217968 536 218020 542
rect 217784 478 217836 484
rect 217888 496 217968 524
rect 217520 354 217548 478
rect 217888 354 217916 496
rect 224328 524 224356 768
rect 224406 776 224462 785
rect 224406 711 224462 720
rect 224420 678 224448 711
rect 224408 672 224460 678
rect 224512 660 224540 870
rect 224604 785 224632 1414
rect 224788 1306 224816 1652
rect 225694 1592 225750 1601
rect 225064 1550 225644 1578
rect 225064 1329 225092 1550
rect 225418 1456 225474 1465
rect 225418 1391 225474 1400
rect 224696 1278 224816 1306
rect 225050 1320 225106 1329
rect 224590 776 224646 785
rect 224590 711 224646 720
rect 224592 672 224644 678
rect 224512 632 224592 660
rect 224408 614 224460 620
rect 224592 614 224644 620
rect 224696 524 224724 1278
rect 225050 1255 225106 1264
rect 225234 1320 225290 1329
rect 225234 1255 225290 1264
rect 224776 1216 224828 1222
rect 224776 1158 224828 1164
rect 224958 1184 225014 1193
rect 224788 898 224816 1158
rect 225142 1184 225198 1193
rect 225064 1154 225142 1170
rect 224958 1119 225014 1128
rect 225052 1148 225142 1154
rect 224972 1034 225000 1119
rect 225104 1142 225142 1148
rect 225248 1154 225276 1255
rect 225326 1184 225382 1193
rect 225142 1119 225198 1128
rect 225236 1148 225288 1154
rect 225052 1090 225104 1096
rect 225326 1119 225382 1128
rect 225236 1090 225288 1096
rect 225340 1034 225368 1119
rect 224972 1006 225368 1034
rect 225432 1034 225460 1391
rect 225512 1352 225564 1358
rect 225512 1294 225564 1300
rect 225524 1154 225552 1294
rect 225616 1170 225644 1550
rect 225800 1578 225828 1652
rect 232044 1624 232096 1630
rect 225878 1592 225934 1601
rect 225800 1550 225878 1578
rect 225694 1527 225750 1536
rect 225878 1527 225934 1536
rect 231766 1592 231822 1601
rect 231766 1527 231822 1536
rect 231964 1584 232044 1612
rect 225708 1306 225736 1527
rect 231780 1476 231808 1527
rect 231964 1476 231992 1584
rect 232044 1566 232096 1572
rect 231780 1448 231992 1476
rect 230492 1414 231716 1442
rect 225984 1329 227484 1340
rect 225786 1320 225842 1329
rect 225708 1278 225786 1306
rect 225786 1255 225842 1264
rect 225984 1320 227498 1329
rect 225984 1312 227442 1320
rect 225984 1170 226012 1312
rect 227442 1255 227498 1264
rect 225512 1148 225564 1154
rect 225616 1142 226012 1170
rect 226614 1184 226670 1193
rect 230492 1170 230520 1414
rect 226670 1142 230520 1170
rect 226614 1119 226670 1128
rect 225512 1090 225564 1096
rect 231688 1068 231716 1414
rect 232148 1329 232176 1663
rect 234080 1630 234108 1663
rect 232504 1624 232556 1630
rect 234068 1624 234120 1630
rect 232556 1584 232636 1612
rect 232504 1566 232556 1572
rect 232608 1494 232636 1584
rect 234068 1566 234120 1572
rect 237932 1624 237984 1630
rect 237932 1566 237984 1572
rect 238116 1624 238168 1630
rect 238116 1566 238168 1572
rect 232596 1488 232648 1494
rect 232596 1430 232648 1436
rect 233148 1488 233200 1494
rect 233200 1448 233280 1476
rect 233148 1430 233200 1436
rect 232134 1320 232190 1329
rect 232502 1320 232558 1329
rect 232134 1255 232190 1264
rect 232412 1284 232464 1290
rect 232502 1255 232558 1264
rect 233056 1284 233108 1290
rect 232412 1226 232464 1232
rect 232424 1068 232452 1226
rect 231688 1040 232084 1068
rect 232056 1034 232084 1040
rect 232148 1040 232452 1068
rect 232148 1034 232176 1040
rect 225432 1006 231624 1034
rect 232056 1006 232176 1034
rect 231490 912 231546 921
rect 224788 870 231490 898
rect 231596 898 231624 1006
rect 231596 870 231808 898
rect 231490 847 231546 856
rect 231780 796 231808 870
rect 232516 796 232544 1255
rect 233056 1226 233108 1232
rect 233148 1284 233200 1290
rect 233148 1226 233200 1232
rect 231306 776 231362 785
rect 225340 734 231306 762
rect 225340 678 225368 734
rect 231780 768 232544 796
rect 232964 808 233016 814
rect 233068 796 233096 1226
rect 233160 921 233188 1226
rect 233146 912 233202 921
rect 233252 898 233280 1448
rect 237944 1068 237972 1566
rect 238022 1320 238078 1329
rect 238128 1290 238156 1566
rect 238220 1442 238248 1720
rect 238390 1728 238446 1737
rect 238446 1708 240140 1714
rect 238446 1702 240192 1708
rect 241520 1760 241572 1766
rect 250168 1760 250220 1766
rect 247788 1737 250116 1748
rect 245474 1728 245530 1737
rect 241572 1708 242480 1714
rect 241520 1702 242480 1708
rect 238446 1686 240180 1702
rect 241532 1686 242480 1702
rect 238390 1663 238446 1672
rect 238668 1624 238720 1630
rect 238760 1624 238812 1630
rect 238720 1584 238760 1612
rect 238668 1566 238720 1572
rect 238760 1566 238812 1572
rect 238942 1592 238998 1601
rect 242070 1592 242126 1601
rect 238998 1550 239904 1578
rect 238942 1527 238998 1536
rect 238944 1488 238996 1494
rect 238666 1456 238722 1465
rect 238220 1414 238666 1442
rect 238944 1430 238996 1436
rect 238666 1391 238722 1400
rect 238206 1320 238262 1329
rect 238022 1255 238078 1264
rect 238116 1284 238168 1290
rect 238036 1222 238064 1255
rect 238206 1255 238262 1264
rect 238312 1278 238616 1306
rect 238116 1226 238168 1232
rect 238024 1216 238076 1222
rect 238024 1158 238076 1164
rect 238220 1068 238248 1255
rect 237944 1040 238248 1068
rect 233804 1006 234016 1034
rect 233330 912 233386 921
rect 233252 870 233330 898
rect 233146 847 233202 856
rect 233330 847 233386 856
rect 233804 796 233832 1006
rect 233068 768 233832 796
rect 232964 750 233016 756
rect 231306 711 231362 720
rect 225328 672 225380 678
rect 225328 614 225380 620
rect 231492 672 231544 678
rect 231676 672 231728 678
rect 231544 632 231676 660
rect 231492 614 231544 620
rect 232976 649 233004 750
rect 233148 672 233200 678
rect 231676 614 231728 620
rect 232962 640 233018 649
rect 232962 575 233018 584
rect 233146 640 233148 649
rect 233988 660 234016 1006
rect 238206 776 238262 785
rect 238312 762 238340 1278
rect 238588 1222 238616 1278
rect 238956 1222 238984 1430
rect 239140 1414 239444 1442
rect 239140 1290 239168 1414
rect 239128 1284 239180 1290
rect 239128 1226 239180 1232
rect 239312 1284 239364 1290
rect 239312 1226 239364 1232
rect 238392 1216 238444 1222
rect 238392 1158 238444 1164
rect 238576 1216 238628 1222
rect 238576 1158 238628 1164
rect 238944 1216 238996 1222
rect 238944 1158 238996 1164
rect 238404 785 238432 1158
rect 239220 1080 239272 1086
rect 239220 1022 239272 1028
rect 239232 814 239260 1022
rect 238484 808 238536 814
rect 238262 734 238340 762
rect 238390 776 238446 785
rect 238206 711 238262 720
rect 239220 808 239272 814
rect 238484 750 238536 756
rect 239126 776 239182 785
rect 238390 711 238446 720
rect 238496 660 238524 750
rect 239324 785 239352 1226
rect 239220 750 239272 756
rect 239310 776 239366 785
rect 239126 711 239182 720
rect 239416 762 239444 1414
rect 239876 1290 239904 1550
rect 240152 1550 241928 1578
rect 239772 1284 239824 1290
rect 239772 1226 239824 1232
rect 239864 1284 239916 1290
rect 239864 1226 239916 1232
rect 239784 1034 239812 1226
rect 240152 1034 240180 1550
rect 241336 1488 241388 1494
rect 241336 1430 241388 1436
rect 241348 1290 241376 1430
rect 241244 1284 241296 1290
rect 241244 1226 241296 1232
rect 241336 1284 241388 1290
rect 241336 1226 241388 1232
rect 241256 1170 241284 1226
rect 241256 1142 241836 1170
rect 239784 1006 240180 1034
rect 239416 734 241560 762
rect 239310 711 239366 720
rect 241532 728 241560 734
rect 233200 640 233202 649
rect 233988 632 238524 660
rect 239140 626 239168 711
rect 241532 700 241744 728
rect 239140 598 241560 626
rect 233146 575 233202 584
rect 224328 496 224724 524
rect 217968 478 218020 484
rect 217520 326 217916 354
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 224314 368 224370 377
rect 224682 368 224738 377
rect 224314 303 224370 312
rect 224604 326 224682 354
rect 224328 218 224356 303
rect 224604 218 224632 326
rect 224682 303 224738 312
rect 224328 190 224632 218
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241532 354 241560 598
rect 241716 474 241744 700
rect 241808 660 241836 1142
rect 241900 898 241928 1550
rect 242070 1527 242126 1536
rect 242084 1136 242112 1527
rect 241992 1108 242112 1136
rect 241992 1018 242020 1108
rect 241980 1012 242032 1018
rect 241980 954 242032 960
rect 242452 932 242480 1686
rect 245396 1686 245474 1714
rect 242898 1456 242954 1465
rect 245290 1456 245346 1465
rect 242954 1414 243202 1442
rect 243280 1414 245290 1442
rect 242898 1391 242954 1400
rect 243280 932 243308 1414
rect 245290 1391 245346 1400
rect 245396 1068 245424 1686
rect 247682 1728 247738 1737
rect 245474 1663 245530 1672
rect 245672 1686 247682 1714
rect 245568 1080 245620 1086
rect 242452 904 243308 932
rect 243464 1040 245424 1068
rect 245488 1040 245568 1068
rect 241900 870 242020 898
rect 241992 796 242020 870
rect 241992 768 242112 796
rect 242084 762 242112 768
rect 243464 762 243492 1040
rect 245488 796 245516 1040
rect 245568 1022 245620 1028
rect 245028 785 245516 796
rect 242084 734 243492 762
rect 245014 776 245516 785
rect 245070 768 245516 776
rect 245014 711 245070 720
rect 245672 660 245700 1686
rect 247682 1663 247738 1672
rect 247788 1728 250130 1737
rect 247788 1720 250074 1728
rect 247788 1578 247816 1720
rect 250168 1702 250220 1708
rect 253664 1760 253716 1766
rect 253664 1702 253716 1708
rect 257068 1760 257120 1766
rect 262312 1760 262364 1766
rect 257068 1702 257120 1708
rect 258078 1728 258134 1737
rect 250074 1663 250130 1672
rect 250180 1578 250208 1702
rect 247144 1550 247816 1578
rect 249076 1550 250208 1578
rect 250272 1550 250852 1578
rect 247144 1086 247172 1550
rect 248970 1456 249026 1465
rect 247236 1414 248970 1442
rect 247132 1080 247184 1086
rect 241808 632 245700 660
rect 246592 1006 246896 1034
rect 247132 1022 247184 1028
rect 246592 542 246620 1006
rect 246762 912 246818 921
rect 246868 898 246896 1006
rect 246946 912 247002 921
rect 246868 870 246946 898
rect 246762 847 246818 856
rect 246946 847 247002 856
rect 246776 796 246804 847
rect 246776 768 247080 796
rect 247052 542 247080 768
rect 241796 536 241848 542
rect 241796 478 241848 484
rect 246580 536 246632 542
rect 241704 468 241756 474
rect 241704 410 241756 416
rect 241808 354 241836 478
rect 241532 326 241836 354
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246580 478 246632 484
rect 247040 536 247092 542
rect 246734 -960 246846 480
rect 247040 478 247092 484
rect 247236 474 247264 1414
rect 248970 1391 249026 1400
rect 247314 1320 247370 1329
rect 247314 1255 247370 1264
rect 247328 898 247356 1255
rect 249076 1170 249104 1550
rect 249892 1488 249944 1494
rect 247880 1142 249104 1170
rect 249168 1436 249892 1442
rect 249168 1430 249944 1436
rect 249982 1456 250038 1465
rect 249168 1414 249932 1430
rect 247500 1080 247552 1086
rect 247406 1048 247462 1057
rect 247462 1028 247500 1034
rect 247462 1022 247552 1028
rect 247774 1048 247830 1057
rect 247462 1006 247540 1022
rect 247406 983 247462 992
rect 247880 1034 247908 1142
rect 247830 1006 247908 1034
rect 248236 1080 248288 1086
rect 249168 1068 249196 1414
rect 250272 1442 250300 1550
rect 250038 1414 250300 1442
rect 250720 1488 250772 1494
rect 250720 1430 250772 1436
rect 250824 1442 250852 1550
rect 251546 1456 251602 1465
rect 249982 1391 250038 1400
rect 250626 1320 250682 1329
rect 248288 1040 249196 1068
rect 250180 1278 250626 1306
rect 248236 1022 248288 1028
rect 247774 983 247830 992
rect 250180 921 250208 1278
rect 250626 1255 250682 1264
rect 250732 1057 250760 1430
rect 250824 1414 251546 1442
rect 251546 1391 251602 1400
rect 252756 1414 253336 1442
rect 252756 1329 252784 1414
rect 252742 1320 252798 1329
rect 250824 1278 251404 1306
rect 250534 1048 250590 1057
rect 250534 983 250590 992
rect 250718 1048 250774 1057
rect 250718 983 250774 992
rect 250166 912 250222 921
rect 247328 870 248000 898
rect 247866 776 247922 785
rect 247512 734 247866 762
rect 247512 542 247540 734
rect 247972 762 248000 870
rect 250548 898 250576 983
rect 250824 898 250852 1278
rect 251376 1222 251404 1278
rect 253308 1290 253336 1414
rect 252742 1255 252798 1264
rect 253112 1284 253164 1290
rect 253112 1226 253164 1232
rect 253296 1284 253348 1290
rect 253296 1226 253348 1232
rect 251364 1216 251416 1222
rect 251364 1158 251416 1164
rect 252742 1184 252798 1193
rect 253018 1184 253074 1193
rect 252798 1142 253018 1170
rect 252742 1119 252798 1128
rect 253018 1119 253074 1128
rect 251638 1048 251694 1057
rect 251638 983 251694 992
rect 252112 1006 252678 1034
rect 250548 870 250852 898
rect 251652 898 251680 983
rect 251652 870 252048 898
rect 250166 847 250222 856
rect 247972 734 251220 762
rect 247866 711 247922 720
rect 251192 660 251220 734
rect 252020 678 252048 870
rect 251916 672 251968 678
rect 247604 649 248460 660
rect 247590 640 248474 649
rect 247646 632 248418 640
rect 247590 575 247646 584
rect 251192 632 251772 660
rect 248418 575 248474 584
rect 247500 536 247552 542
rect 247500 478 247552 484
rect 247224 468 247276 474
rect 247224 410 247276 416
rect 247930 -960 248042 480
rect 248326 368 248382 377
rect 248786 368 248842 377
rect 248382 326 248786 354
rect 248326 303 248382 312
rect 248786 303 248842 312
rect 248418 232 248474 241
rect 248694 232 248750 241
rect 248474 190 248694 218
rect 248418 167 248474 176
rect 248694 167 248750 176
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 251744 474 251772 632
rect 251916 614 251968 620
rect 252008 672 252060 678
rect 252008 614 252060 620
rect 251928 524 251956 614
rect 252112 524 252140 1006
rect 252466 912 252522 921
rect 252926 912 252982 921
rect 252466 847 252522 856
rect 252756 870 252926 898
rect 252480 762 252508 847
rect 252756 762 252784 870
rect 252926 847 252982 856
rect 252480 734 252784 762
rect 252836 672 252888 678
rect 252836 614 252888 620
rect 251928 496 252140 524
rect 251732 468 251784 474
rect 251732 410 251784 416
rect 252622 -960 252734 480
rect 252848 474 252876 614
rect 253124 474 253152 1226
rect 253294 1048 253350 1057
rect 253294 983 253350 992
rect 253308 660 253336 983
rect 253676 921 253704 1702
rect 256606 1592 256662 1601
rect 256606 1527 256662 1536
rect 254030 1456 254086 1465
rect 254214 1456 254270 1465
rect 254086 1414 254164 1442
rect 254030 1391 254086 1400
rect 253846 1320 253902 1329
rect 253846 1255 253902 1264
rect 254030 1320 254086 1329
rect 254136 1290 254164 1414
rect 254214 1391 254270 1400
rect 254030 1255 254032 1264
rect 253860 1170 253888 1255
rect 254084 1255 254086 1264
rect 254124 1284 254176 1290
rect 254032 1226 254084 1232
rect 254124 1226 254176 1232
rect 254228 1170 254256 1391
rect 256514 1320 256570 1329
rect 256620 1290 256648 1527
rect 257080 1465 257108 1702
rect 262034 1728 262090 1737
rect 258736 1698 260788 1714
rect 258448 1692 258500 1698
rect 258134 1672 258448 1680
rect 258078 1663 258448 1672
rect 258092 1652 258448 1663
rect 258448 1634 258500 1640
rect 258736 1692 260800 1698
rect 258736 1686 260748 1692
rect 258736 1578 258764 1686
rect 260748 1634 260800 1640
rect 261300 1692 261352 1698
rect 261300 1634 261352 1640
rect 261760 1692 261812 1698
rect 261812 1672 262034 1680
rect 280068 1760 280120 1766
rect 262364 1720 262536 1748
rect 262312 1702 262364 1708
rect 261812 1663 262090 1672
rect 261812 1652 262076 1663
rect 261760 1634 261812 1640
rect 261312 1578 261340 1634
rect 262312 1624 262364 1630
rect 262034 1592 262090 1601
rect 258092 1550 258764 1578
rect 260392 1550 260604 1578
rect 261312 1550 262034 1578
rect 258092 1465 258120 1550
rect 257066 1456 257122 1465
rect 257066 1391 257122 1400
rect 258078 1456 258134 1465
rect 258078 1391 258134 1400
rect 259090 1456 259146 1465
rect 259090 1391 259092 1400
rect 259144 1391 259146 1400
rect 259184 1420 259236 1426
rect 259092 1362 259144 1368
rect 259184 1362 259236 1368
rect 256514 1255 256516 1264
rect 256568 1255 256570 1264
rect 256608 1284 256660 1290
rect 256516 1226 256568 1232
rect 256608 1226 256660 1232
rect 253860 1142 254256 1170
rect 255870 1048 255926 1057
rect 255870 983 255926 992
rect 253662 912 253718 921
rect 253662 847 253718 856
rect 255884 762 255912 983
rect 255962 776 256018 785
rect 255884 734 255962 762
rect 258354 776 258410 785
rect 255962 711 256018 720
rect 256068 734 258354 762
rect 256068 660 256096 734
rect 258354 711 258410 720
rect 253308 632 256096 660
rect 252836 468 252888 474
rect 252836 410 252888 416
rect 253112 468 253164 474
rect 253112 410 253164 416
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259196 474 259224 1362
rect 260392 1290 260420 1550
rect 260470 1456 260526 1465
rect 260576 1442 260604 1550
rect 262312 1566 262364 1572
rect 262034 1527 262090 1536
rect 260654 1456 260710 1465
rect 260576 1414 260654 1442
rect 260470 1391 260526 1400
rect 260654 1391 260710 1400
rect 260852 1414 261432 1442
rect 260484 1290 260512 1391
rect 260380 1284 260432 1290
rect 260380 1226 260432 1232
rect 260472 1284 260524 1290
rect 260472 1226 260524 1232
rect 260564 1216 260616 1222
rect 260564 1158 260616 1164
rect 260576 898 260604 1158
rect 260852 898 260880 1414
rect 261404 1329 261432 1414
rect 261206 1320 261262 1329
rect 261206 1255 261262 1264
rect 261390 1320 261446 1329
rect 261390 1255 261446 1264
rect 261220 1204 261248 1255
rect 261220 1176 261892 1204
rect 260576 870 260880 898
rect 261864 785 261892 1176
rect 262324 1057 262352 1566
rect 262508 1057 262536 1720
rect 268474 1728 268530 1737
rect 265544 1686 268474 1714
rect 262600 1550 265112 1578
rect 261942 1048 261998 1057
rect 262310 1048 262366 1057
rect 261998 1006 262246 1034
rect 261942 983 261998 992
rect 262310 983 262366 992
rect 262494 1048 262550 1057
rect 262494 983 262550 992
rect 260838 776 260894 785
rect 261850 776 261906 785
rect 260894 734 261800 762
rect 260838 711 260894 720
rect 259276 672 259328 678
rect 261576 672 261628 678
rect 261574 640 261576 649
rect 261628 640 261630 649
rect 259328 620 260052 626
rect 259276 614 260052 620
rect 259288 598 260052 614
rect 259184 468 259236 474
rect 259184 410 259236 416
rect 259798 -960 259910 480
rect 260024 474 260052 598
rect 260576 598 261248 626
rect 260576 474 260604 598
rect 260012 468 260064 474
rect 260012 410 260064 416
rect 260564 468 260616 474
rect 260564 410 260616 416
rect 260994 -960 261106 480
rect 261220 474 261248 598
rect 261574 575 261630 584
rect 261772 542 261800 734
rect 261850 711 261906 720
rect 262600 649 262628 1550
rect 263048 1488 263100 1494
rect 265084 1476 265112 1550
rect 265164 1488 265216 1494
rect 265084 1448 265164 1476
rect 263100 1436 265020 1442
rect 263048 1430 265020 1436
rect 265164 1430 265216 1436
rect 265440 1488 265492 1494
rect 265440 1430 265492 1436
rect 263060 1414 265020 1430
rect 262678 1320 262734 1329
rect 264992 1306 265020 1414
rect 265346 1320 265402 1329
rect 262734 1278 262812 1306
rect 264992 1278 265346 1306
rect 262678 1255 262734 1264
rect 262784 1170 262812 1278
rect 265346 1255 265402 1264
rect 265452 1170 265480 1430
rect 262784 1142 265112 1170
rect 265084 1034 265112 1142
rect 265360 1142 265480 1170
rect 265360 1034 265388 1142
rect 265084 1006 265388 1034
rect 262678 776 262734 785
rect 262678 711 262734 720
rect 262862 776 262918 785
rect 262862 711 262918 720
rect 262586 640 262642 649
rect 262586 575 262642 584
rect 261760 536 261812 542
rect 261760 478 261812 484
rect 261208 468 261260 474
rect 261208 410 261260 416
rect 262190 -960 262302 480
rect 262692 354 262720 711
rect 262876 474 262904 711
rect 265544 626 265572 1686
rect 268842 1728 268898 1737
rect 268474 1663 268530 1672
rect 268672 1686 268842 1714
rect 268382 1592 268438 1601
rect 268672 1578 268700 1686
rect 279330 1728 279386 1737
rect 268842 1663 268898 1672
rect 272260 1686 273484 1714
rect 272156 1624 272208 1630
rect 270958 1592 271014 1601
rect 268438 1550 268700 1578
rect 268764 1550 270724 1578
rect 268382 1527 268438 1536
rect 265624 1488 265676 1494
rect 268660 1488 268712 1494
rect 265624 1430 265676 1436
rect 268014 1456 268070 1465
rect 265452 598 265572 626
rect 265452 542 265480 598
rect 265440 536 265492 542
rect 262864 468 262916 474
rect 262864 410 262916 416
rect 262956 468 263008 474
rect 262956 410 263008 416
rect 262968 354 262996 410
rect 262692 326 262996 354
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265440 478 265492 484
rect 264888 468 264940 474
rect 264888 410 264940 416
rect 264900 354 264928 410
rect 265636 388 265664 1430
rect 268764 1476 268792 1550
rect 268712 1448 268792 1476
rect 268844 1488 268896 1494
rect 268842 1456 268844 1465
rect 269488 1488 269540 1494
rect 268896 1456 268898 1465
rect 268660 1430 268712 1436
rect 269026 1456 269082 1465
rect 268014 1391 268070 1400
rect 268842 1391 268898 1400
rect 268948 1414 269026 1442
rect 268028 1170 268056 1391
rect 268948 1170 268976 1414
rect 270696 1476 270724 1550
rect 270958 1527 271014 1536
rect 271878 1592 271934 1601
rect 272156 1566 272208 1572
rect 271878 1527 271934 1536
rect 270696 1448 270816 1476
rect 269488 1430 269540 1436
rect 269026 1391 269082 1400
rect 269210 1184 269266 1193
rect 268028 1142 268976 1170
rect 269040 1142 269210 1170
rect 265990 776 266046 785
rect 266266 776 266322 785
rect 266046 734 266266 762
rect 265990 711 266046 720
rect 269040 762 269068 1142
rect 269210 1119 269266 1128
rect 266266 711 266322 720
rect 266832 734 269068 762
rect 266832 649 266860 734
rect 267004 672 267056 678
rect 266818 640 266874 649
rect 266818 575 266874 584
rect 267002 640 267004 649
rect 267188 672 267240 678
rect 267056 640 267058 649
rect 267188 614 267240 620
rect 267002 575 267058 584
rect 267200 490 267228 614
rect 267384 598 269068 626
rect 267384 490 267412 598
rect 265084 360 265664 388
rect 265084 354 265112 360
rect 264900 326 265112 354
rect 265070 232 265126 241
rect 265070 167 265126 176
rect 265622 232 265678 241
rect 265622 167 265678 176
rect 265084 82 265112 167
rect 265636 82 265664 167
rect 265084 54 265664 82
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 267200 462 267412 490
rect 268078 -960 268190 480
rect 269040 474 269068 598
rect 269028 468 269080 474
rect 269028 410 269080 416
rect 269274 -960 269386 480
rect 269500 474 269528 1430
rect 270788 1222 270816 1448
rect 270972 1442 271000 1527
rect 271328 1488 271380 1494
rect 271234 1456 271290 1465
rect 270972 1414 271234 1442
rect 271328 1430 271380 1436
rect 271234 1391 271290 1400
rect 271340 1290 271368 1430
rect 271418 1320 271474 1329
rect 271328 1284 271380 1290
rect 271474 1278 271722 1306
rect 271418 1255 271474 1264
rect 271328 1226 271380 1232
rect 270592 1216 270644 1222
rect 270776 1216 270828 1222
rect 270644 1164 270724 1170
rect 270592 1158 270724 1164
rect 270776 1158 270828 1164
rect 270604 1142 270724 1158
rect 269488 468 269540 474
rect 269488 410 269540 416
rect 270470 -960 270582 480
rect 270696 474 270724 1142
rect 271050 776 271106 785
rect 271234 776 271290 785
rect 271106 746 271184 762
rect 271106 740 271196 746
rect 271106 734 271144 740
rect 271050 711 271106 720
rect 271234 711 271290 720
rect 271144 682 271196 688
rect 270960 672 271012 678
rect 271248 626 271276 711
rect 271012 620 271276 626
rect 270960 614 271276 620
rect 270972 598 271276 614
rect 271892 542 271920 1527
rect 272168 1290 272196 1566
rect 272260 1494 272288 1686
rect 272248 1488 272300 1494
rect 272248 1430 272300 1436
rect 272340 1488 272392 1494
rect 272340 1430 272392 1436
rect 272352 1290 272380 1430
rect 272156 1284 272208 1290
rect 272156 1226 272208 1232
rect 272340 1284 272392 1290
rect 272340 1226 272392 1232
rect 273456 1193 273484 1686
rect 279330 1663 279386 1672
rect 279436 1708 280068 1714
rect 280252 1760 280304 1766
rect 279436 1702 280120 1708
rect 280172 1720 280252 1748
rect 279436 1686 280108 1702
rect 273904 1624 273956 1630
rect 273904 1566 273956 1572
rect 273996 1624 274048 1630
rect 273996 1566 274048 1572
rect 273812 1488 273864 1494
rect 273534 1456 273590 1465
rect 273812 1430 273864 1436
rect 273534 1391 273590 1400
rect 273258 1184 273314 1193
rect 273442 1184 273498 1193
rect 273314 1142 273392 1170
rect 273258 1119 273314 1128
rect 273364 746 273392 1142
rect 273548 1170 273576 1391
rect 273824 1290 273852 1430
rect 273916 1290 273944 1566
rect 273812 1284 273864 1290
rect 273812 1226 273864 1232
rect 273904 1284 273956 1290
rect 273904 1226 273956 1232
rect 274008 1170 274036 1566
rect 273548 1142 274036 1170
rect 273442 1119 273498 1128
rect 273352 740 273404 746
rect 273352 682 273404 688
rect 279344 542 279372 1663
rect 279436 1193 279464 1686
rect 280172 1601 280200 1720
rect 290280 1760 290332 1766
rect 285770 1728 285826 1737
rect 280252 1702 280304 1708
rect 280356 1686 281120 1714
rect 280252 1624 280304 1630
rect 279790 1592 279846 1601
rect 279974 1592 280030 1601
rect 279846 1550 279974 1578
rect 279790 1527 279846 1536
rect 279974 1527 280030 1536
rect 280158 1592 280214 1601
rect 280356 1612 280384 1686
rect 280304 1584 280384 1612
rect 280528 1624 280580 1630
rect 280526 1592 280528 1601
rect 280580 1592 280582 1601
rect 280252 1566 280304 1572
rect 280158 1527 280214 1536
rect 280526 1527 280582 1536
rect 279516 1488 279568 1494
rect 279516 1430 279568 1436
rect 280252 1488 280304 1494
rect 280252 1430 280304 1436
rect 279528 1290 279556 1430
rect 279516 1284 279568 1290
rect 279516 1226 279568 1232
rect 279884 1216 279936 1222
rect 279422 1184 279478 1193
rect 280264 1204 280292 1430
rect 280540 1414 280936 1442
rect 280540 1329 280568 1414
rect 280526 1320 280582 1329
rect 280526 1255 280582 1264
rect 280264 1176 280384 1204
rect 279936 1164 280016 1170
rect 279884 1158 280016 1164
rect 279896 1142 280016 1158
rect 279422 1119 279478 1128
rect 279882 776 279938 785
rect 279988 762 280016 1142
rect 280250 776 280306 785
rect 279988 734 280200 762
rect 279882 711 279938 720
rect 279896 626 279924 711
rect 280068 672 280120 678
rect 279896 620 280068 626
rect 280172 660 280200 734
rect 280356 762 280384 1176
rect 280908 1170 280936 1414
rect 280986 1320 281042 1329
rect 281092 1306 281120 1686
rect 281552 1686 285770 1714
rect 281552 1465 281580 1686
rect 337844 1760 337896 1766
rect 294602 1728 294658 1737
rect 290280 1702 290332 1708
rect 285770 1663 285826 1672
rect 281644 1550 282224 1578
rect 285784 1562 289768 1578
rect 281538 1456 281594 1465
rect 281538 1391 281594 1400
rect 281042 1278 281120 1306
rect 280986 1255 281042 1264
rect 280908 1142 281198 1170
rect 280306 734 280384 762
rect 280250 711 280306 720
rect 281540 672 281592 678
rect 280172 632 280384 660
rect 279896 614 280120 620
rect 279896 598 280108 614
rect 270776 536 270828 542
rect 270776 478 270828 484
rect 271880 536 271932 542
rect 270684 468 270736 474
rect 270684 410 270736 416
rect 270788 406 270816 478
rect 270776 400 270828 406
rect 270776 342 270828 348
rect 271666 -960 271778 480
rect 271880 478 271932 484
rect 279332 536 279384 542
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 279332 478 279384 484
rect 280038 -960 280150 480
rect 280356 474 280384 632
rect 281644 660 281672 1550
rect 282196 1494 282224 1550
rect 285772 1556 289780 1562
rect 285824 1550 289728 1556
rect 285772 1498 285824 1504
rect 289728 1498 289780 1504
rect 281724 1488 281776 1494
rect 281722 1456 281724 1465
rect 282092 1488 282144 1494
rect 281776 1456 281778 1465
rect 282092 1430 282144 1436
rect 282184 1488 282236 1494
rect 289360 1488 289412 1494
rect 282184 1430 282236 1436
rect 285310 1456 285366 1465
rect 281722 1391 281778 1400
rect 282104 1306 282132 1430
rect 285954 1456 286010 1465
rect 285366 1414 285954 1442
rect 285310 1391 285366 1400
rect 285954 1391 286010 1400
rect 288912 1436 289360 1442
rect 288912 1430 289412 1436
rect 288912 1414 289400 1430
rect 282104 1278 285444 1306
rect 281908 1216 281960 1222
rect 281908 1158 281960 1164
rect 281920 785 281948 1158
rect 281906 776 281962 785
rect 281906 711 281962 720
rect 282090 776 282146 785
rect 282090 711 282146 720
rect 285310 776 285366 785
rect 285416 762 285444 1278
rect 287518 1184 287574 1193
rect 287794 1184 287850 1193
rect 287518 1119 287574 1128
rect 287624 1142 287794 1170
rect 285678 1048 285734 1057
rect 285734 1006 286364 1034
rect 285678 983 285734 992
rect 286232 876 286284 882
rect 285876 836 286232 864
rect 285770 776 285826 785
rect 285416 734 285770 762
rect 285310 711 285366 720
rect 285770 711 285826 720
rect 281592 632 281672 660
rect 281540 614 281592 620
rect 282104 490 282132 711
rect 285324 626 285352 711
rect 285876 626 285904 836
rect 286232 818 286284 824
rect 286336 762 286364 1006
rect 287532 882 287560 1119
rect 287520 876 287572 882
rect 287520 818 287572 824
rect 287624 762 287652 1142
rect 287794 1119 287850 1128
rect 286336 734 287652 762
rect 285324 598 285628 626
rect 280344 468 280396 474
rect 280344 410 280396 416
rect 281234 -960 281346 480
rect 281552 474 282132 490
rect 281540 468 282132 474
rect 281592 462 282132 468
rect 281540 410 281592 416
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285600 474 285628 598
rect 285692 598 285904 626
rect 286048 672 286100 678
rect 286100 620 288572 626
rect 286048 614 288572 620
rect 286060 598 288572 614
rect 285692 474 285720 598
rect 285588 468 285640 474
rect 285588 410 285640 416
rect 285680 468 285732 474
rect 285680 410 285732 416
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 288544 218 288572 598
rect 288912 338 288940 1414
rect 289634 1320 289690 1329
rect 289372 1278 289634 1306
rect 288900 332 288952 338
rect 288900 274 288952 280
rect 289372 218 289400 1278
rect 289634 1255 289690 1264
rect 290188 1216 290240 1222
rect 289542 1184 289598 1193
rect 290188 1158 290240 1164
rect 289542 1119 289598 1128
rect 289556 762 289584 1119
rect 289648 882 289860 898
rect 289636 876 289860 882
rect 289688 870 289860 876
rect 289832 864 289860 870
rect 289832 836 290136 864
rect 289636 818 289688 824
rect 289556 734 289768 762
rect 289740 678 289768 734
rect 289728 672 289780 678
rect 289728 614 289780 620
rect 290108 542 290136 836
rect 290096 536 290148 542
rect 288544 190 289400 218
rect 289514 -960 289626 480
rect 290096 478 290148 484
rect 290200 474 290228 1158
rect 290292 746 290320 1702
rect 290936 1686 291148 1714
rect 290936 1630 290964 1686
rect 290372 1624 290424 1630
rect 290924 1624 290976 1630
rect 290424 1572 290766 1578
rect 290372 1566 290766 1572
rect 290924 1566 290976 1572
rect 290384 1550 290766 1566
rect 290372 1488 290424 1494
rect 290372 1430 290424 1436
rect 290384 1193 290412 1430
rect 290556 1216 290608 1222
rect 290370 1184 290426 1193
rect 290556 1158 290608 1164
rect 291016 1216 291068 1222
rect 291016 1158 291068 1164
rect 290370 1119 290426 1128
rect 290568 898 290596 1158
rect 291028 898 291056 1158
rect 291120 1034 291148 1686
rect 294970 1728 295026 1737
rect 294602 1663 294658 1672
rect 294708 1686 294970 1714
rect 293684 1624 293736 1630
rect 293736 1584 294000 1612
rect 293684 1566 293736 1572
rect 293972 1494 294000 1584
rect 293960 1488 294012 1494
rect 293960 1430 294012 1436
rect 294616 1204 294644 1663
rect 294708 1329 294736 1686
rect 309966 1728 310022 1737
rect 296824 1698 298692 1714
rect 299952 1698 300164 1714
rect 296812 1692 298692 1698
rect 294970 1663 295026 1672
rect 295076 1652 295748 1680
rect 295076 1578 295104 1652
rect 294800 1550 295104 1578
rect 295614 1592 295670 1601
rect 294800 1494 294828 1550
rect 295720 1578 295748 1652
rect 296864 1686 298692 1692
rect 296812 1634 296864 1640
rect 295798 1592 295854 1601
rect 295720 1550 295798 1578
rect 295614 1527 295670 1536
rect 296258 1592 296314 1601
rect 295798 1527 295854 1536
rect 296180 1550 296258 1578
rect 294788 1488 294840 1494
rect 295340 1488 295392 1494
rect 294788 1430 294840 1436
rect 294984 1448 295340 1476
rect 294984 1329 295012 1448
rect 295340 1430 295392 1436
rect 295628 1442 295656 1527
rect 296180 1442 296208 1550
rect 296258 1527 296314 1536
rect 296732 1562 298600 1578
rect 296732 1556 298612 1562
rect 296732 1550 298560 1556
rect 295628 1414 296208 1442
rect 294694 1320 294750 1329
rect 294694 1255 294750 1264
rect 294970 1320 295026 1329
rect 294970 1255 295026 1264
rect 295154 1320 295210 1329
rect 296732 1290 296760 1550
rect 298560 1498 298612 1504
rect 296812 1488 296864 1494
rect 296812 1430 296864 1436
rect 295154 1255 295210 1264
rect 296720 1284 296772 1290
rect 294616 1176 294828 1204
rect 293866 1048 293922 1057
rect 291120 1006 293866 1034
rect 293866 983 293922 992
rect 290568 870 291056 898
rect 293788 882 294736 898
rect 293776 876 294736 882
rect 293828 870 294736 876
rect 293776 818 293828 824
rect 290370 776 290426 785
rect 290280 740 290332 746
rect 290370 711 290372 720
rect 290280 682 290332 688
rect 290424 711 290426 720
rect 290372 682 290424 688
rect 294708 626 294736 870
rect 294800 785 294828 1176
rect 294786 776 294842 785
rect 295168 746 295196 1255
rect 296720 1226 296772 1232
rect 296718 1184 296774 1193
rect 296824 1170 296852 1430
rect 296774 1142 296852 1170
rect 296718 1119 296774 1128
rect 296902 1048 296958 1057
rect 296902 983 296904 992
rect 296956 983 296958 992
rect 296904 954 296956 960
rect 298664 898 298692 1686
rect 299940 1692 300164 1698
rect 299992 1686 300164 1692
rect 300136 1680 300164 1686
rect 300228 1680 300256 1700
rect 300136 1652 300256 1680
rect 321742 1728 321798 1737
rect 309966 1663 310022 1672
rect 314752 1692 314804 1698
rect 299940 1634 299992 1640
rect 305642 1592 305698 1601
rect 305552 1556 305604 1562
rect 305826 1592 305882 1601
rect 305642 1527 305644 1536
rect 305552 1498 305604 1504
rect 305696 1527 305698 1536
rect 305748 1550 305826 1578
rect 305644 1498 305696 1504
rect 299940 1488 299992 1494
rect 299940 1430 299992 1436
rect 305564 1442 305592 1498
rect 305748 1442 305776 1550
rect 305826 1527 305882 1536
rect 307022 1592 307078 1601
rect 307022 1527 307078 1536
rect 307206 1592 307262 1601
rect 307206 1527 307262 1536
rect 309230 1592 309286 1601
rect 309230 1527 309286 1536
rect 299952 1057 299980 1430
rect 305564 1414 305776 1442
rect 300676 1216 300728 1222
rect 300676 1158 300728 1164
rect 299938 1048 299994 1057
rect 300688 1034 300716 1158
rect 303434 1048 303490 1057
rect 300688 1006 303434 1034
rect 299938 983 299994 992
rect 303434 983 303490 992
rect 306930 1048 306986 1057
rect 307036 1034 307064 1527
rect 307114 1048 307170 1057
rect 307036 1006 307114 1034
rect 306930 983 306932 992
rect 306984 983 306986 992
rect 307114 983 307170 992
rect 306932 954 306984 960
rect 298664 870 300532 898
rect 295246 776 295302 785
rect 294786 711 294842 720
rect 295156 740 295208 746
rect 295246 711 295302 720
rect 295352 734 297036 762
rect 295156 682 295208 688
rect 295260 626 295288 711
rect 293880 598 294552 626
rect 294708 598 295288 626
rect 293880 542 293908 598
rect 293868 536 293920 542
rect 290188 468 290240 474
rect 290188 410 290240 416
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 293868 478 293920 484
rect 294524 490 294552 598
rect 295352 490 295380 734
rect 297008 678 297036 734
rect 296996 672 297048 678
rect 296996 614 297048 620
rect 294298 -960 294410 480
rect 294524 462 295380 490
rect 300504 490 300532 870
rect 306748 876 306800 882
rect 307220 864 307248 1527
rect 309244 1494 309272 1527
rect 309980 1494 310008 1663
rect 314752 1634 314804 1640
rect 319720 1692 319772 1698
rect 321742 1663 321798 1672
rect 321926 1728 321982 1737
rect 352932 1760 352984 1766
rect 347410 1728 347466 1737
rect 337896 1708 338238 1714
rect 337844 1702 338238 1708
rect 337856 1686 338238 1702
rect 321926 1663 321982 1672
rect 348330 1728 348386 1737
rect 347466 1686 347714 1714
rect 347410 1663 347466 1672
rect 352932 1702 352984 1708
rect 366364 1760 366416 1766
rect 375932 1760 375984 1766
rect 373722 1728 373778 1737
rect 366416 1708 366758 1714
rect 366364 1702 366758 1708
rect 348330 1663 348386 1672
rect 348700 1692 348752 1698
rect 319720 1634 319772 1640
rect 309232 1488 309284 1494
rect 309968 1488 310020 1494
rect 309232 1430 309284 1436
rect 309336 1426 309718 1442
rect 309968 1430 310020 1436
rect 309324 1420 309718 1426
rect 309376 1414 309718 1420
rect 309784 1420 309836 1426
rect 309324 1362 309376 1368
rect 309784 1362 309836 1368
rect 308954 1184 309010 1193
rect 306800 836 307248 864
rect 307312 1142 308954 1170
rect 306748 818 306800 824
rect 307312 762 307340 1142
rect 308954 1119 309010 1128
rect 309322 1048 309378 1057
rect 309322 983 309378 992
rect 300688 734 307340 762
rect 309336 762 309364 983
rect 309796 921 309824 1362
rect 309966 1184 310022 1193
rect 309966 1119 310022 1128
rect 309782 912 309838 921
rect 309980 882 310008 1119
rect 314764 921 314792 1634
rect 319732 1601 319760 1634
rect 319534 1592 319590 1601
rect 318904 1562 319194 1578
rect 318892 1556 319194 1562
rect 318944 1550 319194 1556
rect 319534 1527 319590 1536
rect 319718 1592 319774 1601
rect 319718 1527 319774 1536
rect 318892 1498 318944 1504
rect 318432 1488 318484 1494
rect 318432 1430 318484 1436
rect 317694 1320 317750 1329
rect 317694 1255 317750 1264
rect 318338 1320 318394 1329
rect 318338 1255 318394 1264
rect 317708 950 317736 1255
rect 317696 944 317748 950
rect 314750 912 314806 921
rect 309782 847 309838 856
rect 309968 876 310020 882
rect 309968 818 310020 824
rect 310060 876 310112 882
rect 317696 886 317748 892
rect 314750 847 314806 856
rect 310060 818 310112 824
rect 310072 762 310100 818
rect 309336 734 310100 762
rect 300688 678 300716 734
rect 300676 672 300728 678
rect 300676 614 300728 620
rect 300768 672 300820 678
rect 300768 614 300820 620
rect 300780 490 300808 614
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 300504 462 300808 490
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 318352 354 318380 1255
rect 318444 1222 318472 1430
rect 318614 1320 318670 1329
rect 318614 1255 318670 1264
rect 318432 1216 318484 1222
rect 318432 1158 318484 1164
rect 318628 1018 318656 1255
rect 319548 1018 319576 1527
rect 320272 1488 320324 1494
rect 319824 1448 320272 1476
rect 318616 1012 318668 1018
rect 318616 954 318668 960
rect 319444 1012 319496 1018
rect 319444 954 319496 960
rect 319536 1012 319588 1018
rect 319536 954 319588 960
rect 319456 898 319484 954
rect 319456 870 319760 898
rect 319732 814 319760 870
rect 319720 808 319772 814
rect 319720 750 319772 756
rect 319824 626 319852 1448
rect 320272 1430 320324 1436
rect 321756 1034 321784 1663
rect 321940 1193 321968 1663
rect 329748 1488 329800 1494
rect 322952 1414 324912 1442
rect 322952 1329 322980 1414
rect 322938 1320 322994 1329
rect 323122 1320 323178 1329
rect 322938 1255 322994 1264
rect 323044 1278 323122 1306
rect 321926 1184 321982 1193
rect 322110 1184 322166 1193
rect 321926 1119 321982 1128
rect 322032 1142 322110 1170
rect 322032 1034 322060 1142
rect 322110 1119 322166 1128
rect 321756 1006 322060 1034
rect 318904 598 319852 626
rect 318904 474 318932 598
rect 318892 468 318944 474
rect 318892 410 318944 416
rect 318984 468 319036 474
rect 318984 410 319036 416
rect 318996 354 319024 410
rect 318352 326 319024 354
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 323044 474 323072 1278
rect 324884 1306 324912 1414
rect 329576 1436 329748 1442
rect 329576 1430 329800 1436
rect 329576 1414 329788 1430
rect 324962 1320 325018 1329
rect 324884 1278 324962 1306
rect 323122 1255 323178 1264
rect 324962 1255 325018 1264
rect 327538 1320 327594 1329
rect 327538 1255 327540 1264
rect 327592 1255 327594 1264
rect 327722 1320 327778 1329
rect 327722 1255 327778 1264
rect 327906 1320 327962 1329
rect 327906 1255 327962 1264
rect 327540 1226 327592 1232
rect 326908 1142 327212 1170
rect 326908 1057 326936 1142
rect 326894 1048 326950 1057
rect 326894 983 326950 992
rect 327078 1048 327134 1057
rect 327184 1034 327212 1142
rect 327262 1048 327318 1057
rect 327184 1006 327262 1034
rect 327078 983 327134 992
rect 327736 1018 327764 1255
rect 327262 983 327318 992
rect 327724 1012 327776 1018
rect 327092 898 327120 983
rect 327724 954 327776 960
rect 327816 1012 327868 1018
rect 327816 954 327868 960
rect 327828 898 327856 954
rect 327092 870 327856 898
rect 327920 542 327948 1255
rect 328826 1184 328882 1193
rect 328826 1119 328882 1128
rect 328748 950 328776 1020
rect 328840 950 328868 1119
rect 329576 1018 329604 1414
rect 329656 1284 329708 1290
rect 329656 1226 329708 1232
rect 329668 1170 329696 1226
rect 338304 1216 338356 1222
rect 329746 1184 329802 1193
rect 329668 1142 329746 1170
rect 329746 1119 329802 1128
rect 331770 1184 331826 1193
rect 331954 1184 332010 1193
rect 331770 1119 331826 1128
rect 331876 1142 331954 1170
rect 331784 1018 331812 1119
rect 329564 1012 329616 1018
rect 329564 954 329616 960
rect 331680 1012 331732 1018
rect 331680 954 331732 960
rect 331772 1012 331824 1018
rect 331772 954 331824 960
rect 328736 944 328788 950
rect 328550 912 328606 921
rect 328736 886 328788 892
rect 328828 944 328880 950
rect 329748 944 329800 950
rect 328828 886 328880 892
rect 329654 912 329710 921
rect 328550 847 328606 856
rect 329710 892 329748 898
rect 329710 886 329800 892
rect 329838 912 329894 921
rect 329710 870 329788 886
rect 329654 847 329710 856
rect 331692 898 331720 954
rect 331876 898 331904 1142
rect 331954 1119 332010 1128
rect 335818 1184 335874 1193
rect 335818 1119 335874 1128
rect 336002 1184 336058 1193
rect 336002 1119 336058 1128
rect 337856 1142 338160 1170
rect 348344 1193 348372 1663
rect 348700 1634 348752 1640
rect 338304 1158 338356 1164
rect 348330 1184 348386 1193
rect 335832 1018 335860 1119
rect 335728 1012 335780 1018
rect 335728 954 335780 960
rect 335820 1012 335872 1018
rect 335820 954 335872 960
rect 331692 870 331904 898
rect 329838 847 329894 856
rect 328564 762 328592 847
rect 329852 762 329880 847
rect 335740 762 335768 954
rect 336016 921 336044 1119
rect 336002 912 336058 921
rect 336002 847 336058 856
rect 336186 912 336242 921
rect 336186 847 336242 856
rect 328564 734 329880 762
rect 335372 734 335584 762
rect 335740 734 336136 762
rect 335372 678 335400 734
rect 335556 678 335584 734
rect 335360 672 335412 678
rect 335360 614 335412 620
rect 335544 672 335596 678
rect 335544 614 335596 620
rect 327908 536 327960 542
rect 336108 524 336136 734
rect 336200 649 336228 847
rect 336186 640 336242 649
rect 336370 640 336426 649
rect 336186 575 336242 584
rect 336292 598 336370 626
rect 336292 524 336320 598
rect 336370 575 336426 584
rect 336108 496 336320 524
rect 323032 468 323084 474
rect 323032 410 323084 416
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 327908 478 327960 484
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 337856 474 337884 1142
rect 338132 932 338160 1142
rect 338316 932 338344 1158
rect 348330 1119 348386 1128
rect 338132 904 338344 932
rect 343088 944 343140 950
rect 343088 886 343140 892
rect 343100 649 343128 886
rect 348712 785 348740 1634
rect 352944 1601 352972 1702
rect 358176 1692 358228 1698
rect 366376 1686 366758 1702
rect 373722 1663 373778 1672
rect 373906 1728 373962 1737
rect 404452 1760 404504 1766
rect 380162 1728 380218 1737
rect 375984 1708 376234 1714
rect 375932 1702 376234 1708
rect 375944 1686 376234 1702
rect 373906 1663 373962 1672
rect 380162 1663 380218 1672
rect 380346 1728 380402 1737
rect 380346 1663 380402 1672
rect 389086 1728 389142 1737
rect 389086 1663 389142 1672
rect 395434 1728 395490 1737
rect 395434 1663 395490 1672
rect 398654 1728 398710 1737
rect 398654 1663 398710 1672
rect 399574 1728 399630 1737
rect 399574 1663 399630 1672
rect 403714 1728 403770 1737
rect 474924 1760 474976 1766
rect 415674 1728 415730 1737
rect 404504 1708 404754 1714
rect 404452 1702 404754 1708
rect 404464 1686 404754 1702
rect 413848 1698 414230 1714
rect 413836 1692 414230 1698
rect 403714 1663 403770 1672
rect 358176 1634 358228 1640
rect 352930 1592 352986 1601
rect 352930 1527 352986 1536
rect 356336 1488 356388 1494
rect 356336 1430 356388 1436
rect 354036 1216 354088 1222
rect 354036 1158 354088 1164
rect 352196 1080 352248 1086
rect 352196 1022 352248 1028
rect 349528 944 349580 950
rect 349526 912 349528 921
rect 352208 921 352236 1022
rect 349580 912 349582 921
rect 349526 847 349582 856
rect 352194 912 352250 921
rect 352194 847 352250 856
rect 354048 785 354076 1158
rect 356244 944 356296 950
rect 356242 912 356244 921
rect 356296 912 356298 921
rect 356348 898 356376 1430
rect 356808 1426 357190 1442
rect 356796 1420 357190 1426
rect 356848 1414 357190 1420
rect 356796 1362 356848 1368
rect 357992 1284 358044 1290
rect 357992 1226 358044 1232
rect 356980 1216 357032 1222
rect 356980 1158 357032 1164
rect 356426 912 356482 921
rect 356348 870 356426 898
rect 356242 847 356298 856
rect 356426 847 356482 856
rect 356520 808 356572 814
rect 348698 776 348754 785
rect 348698 711 348754 720
rect 354034 776 354090 785
rect 356520 750 356572 756
rect 354034 711 354090 720
rect 356532 649 356560 750
rect 356992 649 357020 1158
rect 358004 898 358032 1226
rect 357636 870 358032 898
rect 357636 785 357664 870
rect 357622 776 357678 785
rect 357622 711 357678 720
rect 343086 640 343142 649
rect 343086 575 343142 584
rect 356518 640 356574 649
rect 356518 575 356574 584
rect 356978 640 357034 649
rect 356978 575 357034 584
rect 337844 468 337896 474
rect 337844 410 337896 416
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358188 377 358216 1634
rect 365994 1592 366050 1601
rect 365994 1527 366050 1536
rect 366178 1592 366234 1601
rect 366178 1527 366234 1536
rect 366008 1329 366036 1527
rect 364706 1320 364762 1329
rect 365994 1320 366050 1329
rect 364706 1255 364762 1264
rect 365260 1284 365312 1290
rect 364720 785 364748 1255
rect 365994 1255 366050 1264
rect 365260 1226 365312 1232
rect 364706 776 364762 785
rect 364706 711 364762 720
rect 365272 649 365300 1226
rect 366192 1193 366220 1527
rect 373354 1320 373410 1329
rect 373354 1255 373410 1264
rect 366178 1184 366234 1193
rect 366178 1119 366234 1128
rect 372526 1184 372582 1193
rect 372526 1119 372582 1128
rect 372540 814 372568 1119
rect 372804 1080 372856 1086
rect 372856 1028 373120 1034
rect 372804 1022 373120 1028
rect 372816 1006 373120 1022
rect 373092 882 373120 1006
rect 373080 876 373132 882
rect 373080 818 373132 824
rect 372528 808 372580 814
rect 373368 785 373396 1255
rect 373736 1193 373764 1663
rect 373722 1184 373778 1193
rect 373722 1119 373778 1128
rect 373920 950 373948 1663
rect 380176 950 380204 1663
rect 373908 944 373960 950
rect 373908 886 373960 892
rect 380164 944 380216 950
rect 380164 886 380216 892
rect 372528 750 372580 756
rect 373354 776 373410 785
rect 373354 711 373410 720
rect 376758 776 376814 785
rect 376758 711 376814 720
rect 365074 640 365130 649
rect 365074 575 365130 584
rect 365258 640 365314 649
rect 365258 575 365314 584
rect 358174 368 358230 377
rect 358174 303 358230 312
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365088 377 365116 575
rect 376668 536 376720 542
rect 376772 490 376800 711
rect 380360 649 380388 1663
rect 385316 1488 385368 1494
rect 385368 1436 385710 1442
rect 385316 1430 385710 1436
rect 385328 1414 385710 1430
rect 389100 1193 389128 1663
rect 395448 1630 395476 1663
rect 398668 1630 398696 1663
rect 399588 1630 399616 1663
rect 403728 1630 403756 1663
rect 413888 1686 414230 1692
rect 415674 1663 415676 1672
rect 413836 1634 413888 1640
rect 415728 1663 415730 1672
rect 418802 1728 418858 1737
rect 418802 1663 418804 1672
rect 415676 1634 415728 1640
rect 418856 1663 418858 1672
rect 432326 1728 432382 1737
rect 432326 1663 432328 1672
rect 418804 1634 418856 1640
rect 432380 1663 432382 1672
rect 436006 1728 436062 1737
rect 436006 1663 436062 1672
rect 443458 1728 443514 1737
rect 443458 1663 443514 1672
rect 443642 1728 443698 1737
rect 443642 1663 443644 1672
rect 432328 1634 432380 1640
rect 394884 1624 394936 1630
rect 395436 1624 395488 1630
rect 394936 1572 395186 1578
rect 394884 1566 395186 1572
rect 395436 1566 395488 1572
rect 398656 1624 398708 1630
rect 398656 1566 398708 1572
rect 399576 1624 399628 1630
rect 399576 1566 399628 1572
rect 403716 1624 403768 1630
rect 432972 1624 433024 1630
rect 403716 1566 403768 1572
rect 406842 1592 406898 1601
rect 394896 1550 395186 1566
rect 406842 1527 406898 1536
rect 407026 1592 407082 1601
rect 407026 1527 407082 1536
rect 415122 1592 415178 1601
rect 415122 1527 415178 1536
rect 418802 1592 418858 1601
rect 423416 1562 423706 1578
rect 433024 1572 433274 1578
rect 432972 1566 433274 1572
rect 418802 1527 418858 1536
rect 423404 1556 423706 1562
rect 406856 1329 406884 1527
rect 406658 1320 406714 1329
rect 406658 1255 406714 1264
rect 406842 1320 406898 1329
rect 406842 1255 406898 1264
rect 389086 1184 389142 1193
rect 389086 1119 389142 1128
rect 389362 1184 389418 1193
rect 389362 1119 389418 1128
rect 389376 950 389404 1119
rect 389364 944 389416 950
rect 389364 886 389416 892
rect 406108 808 406160 814
rect 381542 776 381598 785
rect 381542 711 381598 720
rect 406106 776 406108 785
rect 406160 776 406162 785
rect 406106 711 406162 720
rect 406382 776 406438 785
rect 406382 711 406438 720
rect 380346 640 380402 649
rect 380346 575 380402 584
rect 381556 542 381584 711
rect 386050 640 386106 649
rect 386050 575 386106 584
rect 393410 640 393466 649
rect 393410 575 393466 584
rect 376720 484 376800 490
rect 365074 368 365130 377
rect 365074 303 365130 312
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 376668 478 376800 484
rect 381544 536 381596 542
rect 376680 462 376800 478
rect 376668 400 376720 406
rect 377036 400 377088 406
rect 376720 348 377036 354
rect 376668 342 377088 348
rect 376680 326 377076 342
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 381544 478 381596 484
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 386064 377 386092 575
rect 393424 542 393452 575
rect 393412 536 393464 542
rect 386050 368 386106 377
rect 386050 303 386106 312
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 393412 478 393464 484
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 406396 377 406424 711
rect 406672 377 406700 1255
rect 407040 814 407068 1527
rect 413652 1080 413704 1086
rect 413652 1022 413704 1028
rect 407028 808 407080 814
rect 407028 750 407080 756
rect 411260 808 411312 814
rect 411260 750 411312 756
rect 411272 649 411300 750
rect 411258 640 411314 649
rect 411258 575 411314 584
rect 406382 368 406438 377
rect 406382 303 406438 312
rect 406658 368 406714 377
rect 406658 303 406714 312
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 413664 377 413692 1022
rect 415136 649 415164 1527
rect 418816 1329 418844 1527
rect 423456 1550 423706 1556
rect 425060 1556 425112 1562
rect 423404 1498 423456 1504
rect 432984 1550 433274 1566
rect 425060 1498 425112 1504
rect 418802 1320 418858 1329
rect 425072 1306 425100 1498
rect 436020 1329 436048 1663
rect 443472 1630 443500 1663
rect 443696 1663 443698 1672
rect 453302 1728 453358 1737
rect 453302 1663 453304 1672
rect 443644 1634 443696 1640
rect 453356 1663 453358 1672
rect 462870 1728 462926 1737
rect 462870 1663 462872 1672
rect 453304 1634 453356 1640
rect 462924 1663 462926 1672
rect 474922 1728 474924 1737
rect 481272 1760 481324 1766
rect 474976 1728 474978 1737
rect 474922 1663 474978 1672
rect 481270 1728 481272 1737
rect 489000 1760 489052 1766
rect 481324 1728 481326 1737
rect 481270 1663 481326 1672
rect 488998 1728 489000 1737
rect 501788 1760 501840 1766
rect 489052 1728 489054 1737
rect 488998 1663 489054 1672
rect 501786 1728 501788 1737
rect 512368 1760 512420 1766
rect 501840 1728 501842 1737
rect 512366 1728 512368 1737
rect 529388 1760 529440 1766
rect 512420 1728 512422 1737
rect 501786 1663 501842 1672
rect 509056 1692 509108 1698
rect 462872 1634 462924 1640
rect 512366 1663 512422 1672
rect 522578 1728 522634 1737
rect 522578 1663 522634 1672
rect 529386 1728 529388 1737
rect 559104 1760 559156 1766
rect 529440 1728 529442 1737
rect 567292 1760 567344 1766
rect 559104 1702 559156 1708
rect 567290 1728 567292 1737
rect 567344 1728 567346 1737
rect 529386 1663 529442 1672
rect 558000 1692 558052 1698
rect 509056 1634 509108 1640
rect 443460 1624 443512 1630
rect 440698 1592 440754 1601
rect 453212 1624 453264 1630
rect 443460 1566 443512 1572
rect 453210 1592 453212 1601
rect 453264 1592 453266 1601
rect 440698 1527 440754 1536
rect 453210 1527 453266 1536
rect 462594 1592 462650 1601
rect 471518 1592 471574 1601
rect 471270 1550 471518 1578
rect 462594 1527 462650 1536
rect 471518 1527 471574 1536
rect 424980 1290 425100 1306
rect 418802 1255 418858 1264
rect 424968 1284 425100 1290
rect 425020 1278 425100 1284
rect 436006 1320 436062 1329
rect 436006 1255 436062 1264
rect 424968 1226 425020 1232
rect 440712 1193 440740 1527
rect 451924 1488 451976 1494
rect 451976 1436 452226 1442
rect 451924 1430 452226 1436
rect 451936 1414 452226 1430
rect 462608 1329 462636 1527
rect 443182 1320 443238 1329
rect 443182 1255 443238 1264
rect 453302 1320 453358 1329
rect 453302 1255 453358 1264
rect 460570 1320 460626 1329
rect 460570 1255 460626 1264
rect 462594 1320 462650 1329
rect 462594 1255 462650 1264
rect 476394 1320 476450 1329
rect 476394 1255 476450 1264
rect 476578 1320 476634 1329
rect 482190 1320 482246 1329
rect 476578 1255 476634 1264
rect 480168 1284 480220 1290
rect 440698 1184 440754 1193
rect 440698 1119 440754 1128
rect 425704 808 425756 814
rect 425704 750 425756 756
rect 434994 776 435050 785
rect 415122 640 415178 649
rect 415122 575 415178 584
rect 413650 368 413706 377
rect 413650 303 413706 312
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 425716 377 425744 750
rect 434994 711 434996 720
rect 435048 711 435050 720
rect 434996 682 435048 688
rect 427818 640 427874 649
rect 427818 575 427874 584
rect 425702 368 425758 377
rect 425702 303 425758 312
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 427832 377 427860 575
rect 442736 513 442764 1020
rect 442816 740 442868 746
rect 442816 682 442868 688
rect 442828 649 442856 682
rect 442814 640 442870 649
rect 442814 575 442870 584
rect 442722 504 442778 513
rect 427818 368 427874 377
rect 427818 303 427874 312
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442722 439 442778 448
rect 442970 -960 443082 480
rect 443196 377 443224 1255
rect 453316 1086 453344 1255
rect 453304 1080 453356 1086
rect 453304 1022 453356 1028
rect 460584 785 460612 1255
rect 460570 776 460626 785
rect 460570 711 460626 720
rect 443182 368 443238 377
rect 443182 303 443238 312
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 461688 241 461716 1020
rect 476408 746 476436 1255
rect 476592 785 476620 1255
rect 501326 1320 501382 1329
rect 482190 1255 482246 1264
rect 492496 1284 492548 1290
rect 480168 1226 480220 1232
rect 480180 1086 480208 1226
rect 480168 1080 480220 1086
rect 480168 1022 480220 1028
rect 476764 808 476816 814
rect 476578 776 476634 785
rect 476396 740 476448 746
rect 476764 750 476816 756
rect 476578 711 476634 720
rect 476396 682 476448 688
rect 476776 649 476804 750
rect 476762 640 476818 649
rect 480732 610 480760 1020
rect 482204 785 482232 1255
rect 492496 1226 492548 1232
rect 492680 1284 492732 1290
rect 501326 1255 501382 1264
rect 504178 1320 504234 1329
rect 504178 1255 504234 1264
rect 492680 1226 492732 1232
rect 492508 1068 492536 1226
rect 492692 1068 492720 1226
rect 493968 1216 494020 1222
rect 494244 1216 494296 1222
rect 494020 1164 494244 1170
rect 493968 1158 494296 1164
rect 493980 1142 494284 1158
rect 501340 1086 501368 1255
rect 492508 1040 492720 1068
rect 501328 1080 501380 1086
rect 489840 1006 490222 1034
rect 501328 1022 501380 1028
rect 486148 808 486200 814
rect 482190 776 482246 785
rect 486148 750 486200 756
rect 482190 711 482246 720
rect 476762 575 476818 584
rect 480720 604 480772 610
rect 480720 546 480772 552
rect 461674 232 461730 241
rect 461674 167 461730 176
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473358 232 473414 241
rect 473358 167 473414 176
rect 473726 232 473782 241
rect 473726 167 473782 176
rect 473372 66 473400 167
rect 473740 66 473768 167
rect 473360 60 473412 66
rect 473360 2 473412 8
rect 473728 60 473780 66
rect 473728 2 473780 8
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486160 241 486188 750
rect 486146 232 486202 241
rect 486146 167 486202 176
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 489840 474 489868 1006
rect 490196 740 490248 746
rect 490196 682 490248 688
rect 490208 649 490236 682
rect 490194 640 490250 649
rect 490194 575 490250 584
rect 489828 468 489880 474
rect 489828 410 489880 416
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 499684 338 499712 1020
rect 504192 785 504220 1255
rect 504178 776 504234 785
rect 504178 711 504234 720
rect 509068 649 509096 1634
rect 515588 1624 515640 1630
rect 515588 1566 515640 1572
rect 512000 1284 512052 1290
rect 512000 1226 512052 1232
rect 509054 640 509110 649
rect 509054 575 509110 584
rect 499672 332 499724 338
rect 499672 274 499724 280
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509252 270 509280 1020
rect 512012 950 512040 1226
rect 512644 1080 512696 1086
rect 512644 1022 512696 1028
rect 512000 944 512052 950
rect 512000 886 512052 892
rect 512656 785 512684 1022
rect 515600 785 515628 1566
rect 516690 1320 516746 1329
rect 516690 1255 516746 1264
rect 516874 1320 516930 1329
rect 516874 1255 516930 1264
rect 516704 785 516732 1255
rect 512642 776 512698 785
rect 512642 711 512698 720
rect 515586 776 515642 785
rect 515586 711 515642 720
rect 516690 776 516746 785
rect 516690 711 516746 720
rect 516888 610 516916 1255
rect 518728 814 518756 1020
rect 518716 808 518768 814
rect 518716 750 518768 756
rect 522592 649 522620 1663
rect 558000 1634 558052 1640
rect 528836 1624 528888 1630
rect 528836 1566 528888 1572
rect 549260 1624 549312 1630
rect 549260 1566 549312 1572
rect 522578 640 522634 649
rect 509884 604 509936 610
rect 509884 546 509936 552
rect 516876 604 516928 610
rect 522578 575 522634 584
rect 516876 546 516928 552
rect 509896 513 509924 546
rect 509882 504 509938 513
rect 509240 264 509292 270
rect 509240 206 509292 212
rect 509578 -960 509690 480
rect 509882 439 509938 448
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528204 406 528232 1020
rect 528192 400 528244 406
rect 528192 342 528244 348
rect 528622 -960 528734 480
rect 528848 377 528876 1566
rect 537312 1414 537694 1442
rect 537312 1329 537340 1414
rect 537298 1320 537354 1329
rect 535368 1284 535420 1290
rect 537298 1255 537354 1264
rect 538770 1320 538826 1329
rect 549272 1306 549300 1566
rect 556434 1456 556490 1465
rect 556490 1414 556738 1442
rect 556434 1391 556490 1400
rect 549180 1290 549300 1306
rect 538770 1255 538826 1264
rect 549168 1284 549300 1290
rect 535368 1226 535420 1232
rect 531778 1184 531834 1193
rect 531778 1119 531834 1128
rect 531792 785 531820 1119
rect 535380 1086 535408 1226
rect 535368 1080 535420 1086
rect 535368 1022 535420 1028
rect 531778 776 531834 785
rect 536930 776 536986 785
rect 531778 711 531834 720
rect 536760 734 536930 762
rect 536760 649 536788 734
rect 536930 711 536986 720
rect 536746 640 536802 649
rect 536746 575 536802 584
rect 528834 368 528890 377
rect 528834 303 528890 312
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 538784 377 538812 1255
rect 549220 1278 549300 1284
rect 552478 1320 552534 1329
rect 552478 1255 552534 1264
rect 549168 1226 549220 1232
rect 552492 1170 552520 1255
rect 558012 1193 558040 1634
rect 559116 1601 559144 1702
rect 567290 1663 567346 1672
rect 559102 1592 559158 1601
rect 559102 1527 559158 1536
rect 559378 1592 559434 1601
rect 559378 1527 559434 1536
rect 565818 1592 565874 1601
rect 565874 1550 566214 1578
rect 565818 1527 565874 1536
rect 552754 1184 552810 1193
rect 552492 1142 552754 1170
rect 552754 1119 552810 1128
rect 557998 1184 558054 1193
rect 557998 1119 558054 1128
rect 538956 944 539008 950
rect 538956 886 539008 892
rect 538968 377 538996 886
rect 547248 678 547276 1020
rect 547236 672 547288 678
rect 547236 614 547288 620
rect 545670 504 545726 513
rect 538770 368 538826 377
rect 538770 303 538826 312
rect 538954 368 539010 377
rect 538954 303 539010 312
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 545670 439 545726 448
rect 545684 241 545712 439
rect 545670 232 545726 241
rect 545670 167 545726 176
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559392 377 559420 1527
rect 565818 1456 565874 1465
rect 565818 1391 565820 1400
rect 565872 1391 565874 1400
rect 565820 1362 565872 1368
rect 559562 1320 559618 1329
rect 559562 1255 559618 1264
rect 564438 1320 564494 1329
rect 564438 1255 564440 1264
rect 559576 785 559604 1255
rect 564492 1255 564494 1264
rect 564440 1226 564492 1232
rect 568224 1018 568252 40004
rect 568408 38570 568436 49014
rect 568592 40202 568620 49694
rect 568776 40440 568804 63022
rect 569420 61588 569448 64654
rect 569972 61742 570000 64790
rect 569960 61736 570012 61742
rect 570156 61690 570184 66098
rect 569960 61678 570012 61684
rect 570064 61662 570184 61690
rect 569960 61600 570012 61606
rect 569420 61560 569960 61588
rect 569960 61542 570012 61548
rect 570064 61418 570092 61662
rect 570144 61600 570196 61606
rect 570144 61542 570196 61548
rect 568868 61390 570092 61418
rect 568868 41018 568896 61390
rect 570052 61328 570104 61334
rect 570052 61270 570104 61276
rect 569960 60784 570012 60790
rect 568960 60732 569960 60738
rect 568960 60726 570012 60732
rect 568960 60710 570000 60726
rect 568960 41120 568988 60710
rect 570064 60636 570092 61270
rect 569052 60608 570092 60636
rect 569052 41290 569080 60608
rect 570156 60228 570184 61542
rect 569144 60200 570184 60228
rect 569144 41426 569172 60200
rect 570248 60092 570276 68342
rect 580170 64560 580226 64569
rect 580170 64495 580226 64504
rect 580184 63578 580212 64495
rect 574744 63572 574796 63578
rect 574744 63514 574796 63520
rect 580172 63572 580224 63578
rect 580172 63514 580224 63520
rect 569236 60064 570276 60092
rect 569236 41562 569264 60064
rect 569960 59968 570012 59974
rect 569328 59916 569960 59922
rect 569328 59910 570012 59916
rect 569328 59894 570000 59910
rect 569328 41698 569356 59894
rect 569960 58880 570012 58886
rect 569420 58828 569960 58834
rect 569420 58822 570012 58828
rect 569420 58806 570000 58822
rect 569420 41800 569448 58806
rect 569960 58744 570012 58750
rect 569512 58692 569960 58698
rect 569512 58686 570012 58692
rect 569512 58670 570000 58686
rect 569512 42786 569540 58670
rect 569960 56976 570012 56982
rect 569604 56924 569960 56930
rect 569604 56918 570012 56924
rect 569604 56902 570000 56918
rect 569604 43058 569632 56902
rect 569696 56766 570000 56794
rect 569696 43194 569724 56766
rect 569972 56710 570000 56766
rect 569960 56704 570012 56710
rect 569960 56646 570012 56652
rect 569960 56568 570012 56574
rect 569960 56510 570012 56516
rect 569972 53938 570000 56510
rect 569788 53910 570000 53938
rect 569788 45370 569816 53910
rect 569880 53786 570000 53802
rect 569880 53780 570012 53786
rect 569880 53774 569960 53780
rect 569880 45540 569908 53774
rect 569960 53722 570012 53728
rect 569960 45552 570012 45558
rect 569880 45512 569960 45540
rect 569960 45494 570012 45500
rect 570328 45552 570380 45558
rect 570328 45494 570380 45500
rect 569788 45342 570000 45370
rect 569972 43314 570000 45342
rect 569960 43308 570012 43314
rect 569960 43250 570012 43256
rect 569696 43166 570000 43194
rect 569604 43030 569908 43058
rect 569512 42758 569724 42786
rect 569696 42106 569724 42758
rect 569880 42208 569908 43030
rect 569972 42362 570000 43166
rect 569960 42356 570012 42362
rect 569960 42298 570012 42304
rect 569960 42220 570012 42226
rect 569880 42180 569960 42208
rect 569960 42162 570012 42168
rect 569696 42078 570276 42106
rect 569960 41812 570012 41818
rect 569420 41772 569960 41800
rect 569960 41754 570012 41760
rect 569328 41682 570000 41698
rect 569328 41676 570012 41682
rect 569328 41670 569960 41676
rect 569960 41618 570012 41624
rect 569236 41534 570000 41562
rect 569144 41398 569540 41426
rect 569052 41262 569448 41290
rect 568960 41092 569172 41120
rect 568868 40990 568988 41018
rect 568960 40712 568988 40990
rect 569144 40712 569172 41092
rect 569420 40882 569448 41262
rect 569512 40984 569540 41398
rect 569972 41138 570000 41534
rect 569960 41132 570012 41138
rect 569960 41074 570012 41080
rect 569960 40996 570012 41002
rect 569512 40956 569960 40984
rect 569960 40938 570012 40944
rect 569420 40854 570184 40882
rect 569960 40724 570012 40730
rect 568960 40684 569080 40712
rect 569144 40684 569960 40712
rect 569052 40610 569080 40684
rect 569960 40666 570012 40672
rect 569052 40582 570092 40610
rect 569960 40452 570012 40458
rect 568776 40412 569960 40440
rect 569960 40394 570012 40400
rect 569960 40316 570012 40322
rect 568868 40276 569960 40304
rect 568868 40202 568896 40276
rect 569960 40258 570012 40264
rect 568592 40174 568896 40202
rect 569960 40180 570012 40186
rect 569236 40140 569960 40168
rect 569236 39658 569264 40140
rect 569960 40122 570012 40128
rect 569960 40044 570012 40050
rect 568868 39630 569264 39658
rect 569420 40004 569960 40032
rect 568868 39420 568896 39630
rect 568868 39392 569080 39420
rect 568408 38542 568528 38570
rect 568500 6610 568528 38542
rect 569052 31362 569080 39392
rect 569420 39250 569448 40004
rect 569960 39986 570012 39992
rect 569960 39908 570012 39914
rect 568868 31334 569080 31362
rect 569144 39222 569448 39250
rect 569512 39868 569960 39896
rect 568868 31226 568896 31334
rect 568776 31198 568896 31226
rect 568776 30818 568804 31198
rect 568776 30790 569080 30818
rect 569052 30138 569080 30790
rect 568592 30110 569080 30138
rect 568592 24698 568620 30110
rect 569144 30002 569172 39222
rect 569512 35442 569540 39868
rect 569960 39850 570012 39856
rect 570064 39794 570092 40582
rect 569696 39766 570092 39794
rect 569696 39658 569724 39766
rect 569960 39704 570012 39710
rect 569880 39664 569960 39692
rect 569880 39658 569908 39664
rect 568684 29974 569172 30002
rect 569328 35414 569540 35442
rect 569604 39630 569724 39658
rect 569788 39630 569908 39658
rect 569960 39646 570012 39652
rect 568684 24868 568712 29974
rect 569328 29730 569356 35414
rect 569604 35306 569632 39630
rect 568776 29702 569356 29730
rect 569420 35278 569632 35306
rect 568776 25140 568804 29702
rect 569420 25650 569448 35278
rect 569788 35170 569816 39630
rect 570156 39522 570184 40854
rect 569512 35142 569816 35170
rect 569880 39494 570184 39522
rect 569512 26330 569540 35142
rect 569880 26500 569908 39494
rect 569960 39432 570012 39438
rect 570248 39386 570276 42078
rect 569960 39374 570012 39380
rect 569972 28370 570000 39374
rect 570156 39358 570276 39386
rect 570156 31074 570184 39358
rect 570236 39092 570288 39098
rect 570236 39034 570288 39040
rect 570144 31068 570196 31074
rect 570144 31010 570196 31016
rect 570248 28370 570276 39034
rect 570340 34921 570368 45494
rect 574756 41857 574784 63514
rect 574742 41848 574798 41857
rect 574742 41783 574798 41792
rect 570326 34912 570382 34921
rect 570326 34847 570382 34856
rect 570328 34808 570380 34814
rect 570328 34750 570380 34756
rect 569972 28342 570092 28370
rect 569960 26512 570012 26518
rect 569880 26472 569960 26500
rect 569960 26454 570012 26460
rect 569512 26302 570000 26330
rect 569972 25770 570000 26302
rect 569960 25764 570012 25770
rect 569960 25706 570012 25712
rect 569420 25622 570000 25650
rect 569972 25566 570000 25622
rect 569960 25560 570012 25566
rect 569960 25502 570012 25508
rect 569960 25152 570012 25158
rect 568776 25112 569960 25140
rect 569960 25094 570012 25100
rect 568684 24840 568988 24868
rect 568592 24670 568896 24698
rect 568868 18714 568896 24670
rect 568316 6582 568528 6610
rect 568684 18686 568896 18714
rect 568316 1766 568344 6582
rect 568684 4978 568712 18686
rect 568960 18442 568988 24840
rect 569960 24336 570012 24342
rect 568408 4950 568712 4978
rect 568776 18414 568988 18442
rect 569052 24296 569960 24324
rect 568304 1760 568356 1766
rect 568304 1702 568356 1708
rect 568304 1624 568356 1630
rect 568304 1566 568356 1572
rect 568316 1358 568344 1566
rect 568304 1352 568356 1358
rect 568304 1294 568356 1300
rect 568408 1193 568436 4950
rect 568776 4842 568804 18414
rect 569052 16130 569080 24296
rect 569960 24278 570012 24284
rect 569960 24200 570012 24206
rect 568592 4814 568804 4842
rect 568868 16102 569080 16130
rect 569144 24148 569960 24154
rect 569144 24142 570012 24148
rect 569144 24126 570000 24142
rect 568592 2258 568620 4814
rect 568500 2230 568620 2258
rect 568500 1562 568528 2230
rect 568868 1986 568896 16102
rect 569144 15994 569172 24126
rect 569960 23792 570012 23798
rect 568684 1958 568896 1986
rect 568960 15966 569172 15994
rect 569236 23740 569960 23746
rect 569236 23734 570012 23740
rect 569236 23718 570000 23734
rect 568684 1630 568712 1958
rect 568960 1714 568988 15966
rect 569236 15858 569264 23718
rect 569052 15830 569264 15858
rect 569420 23594 570000 23610
rect 569420 23588 570012 23594
rect 569420 23582 569960 23588
rect 569052 1834 569080 15830
rect 569420 15722 569448 23582
rect 569960 23530 570012 23536
rect 570064 23338 570092 28342
rect 569788 23310 570092 23338
rect 570156 28342 570276 28370
rect 569788 18034 569816 23310
rect 569960 23248 570012 23254
rect 569960 23190 570012 23196
rect 569604 18006 569816 18034
rect 569604 17932 569632 18006
rect 569236 15694 569448 15722
rect 569512 17904 569632 17932
rect 569236 15586 569264 15694
rect 569144 15558 569264 15586
rect 569040 1828 569092 1834
rect 569040 1770 569092 1776
rect 568960 1686 569080 1714
rect 568672 1624 568724 1630
rect 568672 1566 568724 1572
rect 568488 1556 568540 1562
rect 568488 1498 568540 1504
rect 568764 1556 568816 1562
rect 568764 1498 568816 1504
rect 568776 1306 568804 1498
rect 568684 1278 568804 1306
rect 568394 1184 568450 1193
rect 568394 1119 568450 1128
rect 568684 1057 568712 1278
rect 568670 1048 568726 1057
rect 568212 1012 568264 1018
rect 568670 983 568726 992
rect 568212 954 568264 960
rect 559562 776 559618 785
rect 559562 711 559618 720
rect 569052 626 569080 1686
rect 569144 785 569172 15558
rect 569512 15450 569540 17904
rect 569972 17762 570000 23190
rect 570156 21434 570184 28342
rect 570236 25152 570288 25158
rect 570236 25094 570288 25100
rect 570248 23594 570276 25094
rect 570340 24342 570368 34750
rect 570328 24336 570380 24342
rect 570328 24278 570380 24284
rect 570236 23588 570288 23594
rect 570236 23530 570288 23536
rect 569236 15422 569540 15450
rect 569604 17734 570000 17762
rect 570064 21406 570184 21434
rect 569236 6882 569264 15422
rect 569604 15178 569632 17734
rect 569960 17672 570012 17678
rect 569512 15150 569632 15178
rect 569696 17632 569960 17660
rect 569512 8514 569540 15150
rect 569696 12322 569724 17632
rect 569960 17614 570012 17620
rect 569604 12294 569724 12322
rect 569604 9602 569632 12294
rect 569604 9574 569724 9602
rect 569696 8650 569724 9574
rect 569696 8634 570000 8650
rect 569696 8628 570012 8634
rect 569696 8622 569960 8628
rect 569960 8570 570012 8576
rect 569512 8486 569632 8514
rect 569604 8242 569632 8486
rect 569512 8214 569632 8242
rect 569236 6854 569448 6882
rect 569224 1828 569276 1834
rect 569224 1770 569276 1776
rect 569130 776 569186 785
rect 569130 711 569186 720
rect 568868 598 569080 626
rect 559378 368 559434 377
rect 559378 303 559434 312
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 568868 134 568896 598
rect 568856 128 568908 134
rect 568856 70 568908 76
rect 569010 -960 569122 480
rect 569236 202 569264 1770
rect 569420 950 569448 6854
rect 569512 1222 569540 8214
rect 569960 8152 570012 8158
rect 569604 8100 569960 8106
rect 569604 8094 570012 8100
rect 569604 8078 570000 8094
rect 569604 1737 569632 8078
rect 570064 7970 570092 21406
rect 580170 17640 580226 17649
rect 580170 17575 580226 17584
rect 580184 15162 580212 17575
rect 571616 15156 571668 15162
rect 571616 15098 571668 15104
rect 580172 15156 580224 15162
rect 580172 15098 580224 15104
rect 570328 14748 570380 14754
rect 570328 14690 570380 14696
rect 570340 12345 570368 14690
rect 571628 14657 571656 15098
rect 571614 14648 571670 14657
rect 571614 14583 571670 14592
rect 570326 12336 570382 12345
rect 570326 12271 570382 12280
rect 570328 8628 570380 8634
rect 570328 8570 570380 8576
rect 569696 7942 570092 7970
rect 569590 1728 569646 1737
rect 569590 1663 569646 1672
rect 569500 1216 569552 1222
rect 569500 1158 569552 1164
rect 569408 944 569460 950
rect 569408 886 569460 892
rect 569224 196 569276 202
rect 569224 138 569276 144
rect 569696 105 569724 7942
rect 569960 7880 570012 7886
rect 569788 7840 569960 7868
rect 569788 1698 569816 7840
rect 569960 7822 570012 7828
rect 570340 4457 570368 8570
rect 570326 4448 570382 4457
rect 570326 4383 570382 4392
rect 569776 1692 569828 1698
rect 569776 1634 569828 1640
rect 569682 96 569738 105
rect 569682 31 569738 40
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 1398 682216 1454 682272
rect 325606 680448 325662 680504
rect 296718 680332 296774 680368
rect 345018 680584 345074 680640
rect 296718 680312 296720 680332
rect 296720 680312 296772 680332
rect 296772 680312 296774 680332
rect 364798 680332 364854 680368
rect 364798 680312 364800 680332
rect 364800 680312 364852 680332
rect 364852 680312 364854 680332
rect 370226 680332 370282 680368
rect 379426 680604 379482 680640
rect 379426 680584 379428 680604
rect 379428 680584 379480 680604
rect 379480 680584 379482 680604
rect 380070 680348 380072 680368
rect 380072 680348 380124 680368
rect 380124 680348 380126 680368
rect 370226 680312 370228 680332
rect 370228 680312 370280 680332
rect 370280 680312 370282 680332
rect 380070 680312 380126 680348
rect 381634 680312 381690 680368
rect 394698 680348 394700 680368
rect 394700 680348 394752 680368
rect 394752 680348 394754 680368
rect 394698 680312 394754 680348
rect 403162 680348 403164 680368
rect 403164 680348 403216 680368
rect 403216 680348 403218 680368
rect 403162 680312 403218 680348
rect 439502 680856 439558 680912
rect 412730 680348 412732 680368
rect 412732 680348 412784 680368
rect 412784 680348 412786 680368
rect 412730 680312 412786 680348
rect 418618 680348 418620 680368
rect 418620 680348 418672 680368
rect 418672 680348 418674 680368
rect 418618 680312 418674 680348
rect 428186 680348 428188 680368
rect 428188 680348 428240 680368
rect 428240 680348 428242 680368
rect 428186 680312 428242 680348
rect 466642 680468 466698 680504
rect 466642 680448 466644 680468
rect 466644 680448 466696 680468
rect 466696 680448 466698 680468
rect 437754 680348 437756 680368
rect 437756 680348 437808 680368
rect 437808 680348 437810 680368
rect 437754 680312 437810 680348
rect 439502 680312 439558 680368
rect 451370 680348 451372 680368
rect 451372 680348 451424 680368
rect 451424 680348 451426 680368
rect 451370 680312 451426 680348
rect 457166 680348 457168 680368
rect 457168 680348 457220 680368
rect 457220 680348 457222 680368
rect 457166 680312 457222 680348
rect 463698 680312 463754 680368
rect 564714 680992 564770 681048
rect 543830 680584 543886 680640
rect 557446 680604 557502 680640
rect 557446 680584 557448 680604
rect 557448 680584 557500 680604
rect 557500 680584 557502 680604
rect 466550 680348 466552 680368
rect 466552 680348 466604 680368
rect 466604 680348 466606 680368
rect 466550 680312 466606 680348
rect 481178 680332 481234 680368
rect 481178 680312 481180 680332
rect 481180 680312 481232 680332
rect 481232 680312 481234 680332
rect 485778 680332 485834 680368
rect 495438 680348 495440 680368
rect 495440 680348 495492 680368
rect 495492 680348 495494 680368
rect 485778 680312 485780 680332
rect 485780 680312 485832 680332
rect 485832 680312 485834 680332
rect 495438 680312 495494 680348
rect 505926 680348 505928 680368
rect 505928 680348 505980 680368
rect 505980 680348 505982 680368
rect 505926 680312 505982 680348
rect 515402 680348 515404 680368
rect 515404 680348 515456 680368
rect 515456 680348 515458 680368
rect 515402 680312 515458 680348
rect 524418 680348 524420 680368
rect 524420 680348 524472 680368
rect 524472 680348 524474 680368
rect 524418 680312 524474 680348
rect 534354 680348 534356 680368
rect 534356 680348 534408 680368
rect 534408 680348 534410 680368
rect 534354 680312 534410 680348
rect 559378 680584 559434 680640
rect 554778 680448 554834 680504
rect 559194 680448 559250 680504
rect 543830 680312 543886 680368
rect 544014 680348 544016 680368
rect 544016 680348 544068 680368
rect 544068 680348 544070 680368
rect 544014 680312 544070 680348
rect 554870 680332 554926 680368
rect 554870 680312 554872 680332
rect 554872 680312 554924 680332
rect 554924 680312 554926 680332
rect 558550 680332 558606 680368
rect 561586 680448 561642 680504
rect 561770 680448 561826 680504
rect 563242 680448 563298 680504
rect 564714 680448 564770 680504
rect 558550 680312 558552 680332
rect 558552 680312 558604 680332
rect 558604 680312 558606 680332
rect 560758 680332 560814 680368
rect 560758 680312 560760 680332
rect 560760 680312 560812 680332
rect 560812 680312 560814 680332
rect 561218 680312 561274 680368
rect 561862 680332 561918 680368
rect 561862 680312 561864 680332
rect 561864 680312 561916 680332
rect 561916 680312 561918 680332
rect 562506 680332 562562 680368
rect 562506 680312 562508 680332
rect 562508 680312 562560 680332
rect 562560 680312 562562 680332
rect 566370 680332 566426 680368
rect 566370 680312 566372 680332
rect 566372 680312 566424 680332
rect 566424 680312 566426 680332
rect 18 624552 74 624608
rect 110 352144 166 352200
rect 18 215736 74 215792
rect 1122 669432 1178 669488
rect 754 442312 810 442368
rect 570 374312 626 374368
rect 662 329024 718 329080
rect 570 208120 626 208176
rect 18 36080 74 36136
rect 202 584 258 640
rect 938 397296 994 397352
rect 478 103400 534 103456
rect 570 78920 626 78976
rect 478 17992 534 18048
rect 1214 646720 1270 646776
rect 662 32272 718 32328
rect 754 19896 810 19952
rect 570 7792 626 7848
rect 386 448 442 504
rect 580170 674600 580226 674656
rect 572718 667392 572774 667448
rect 1582 623736 1638 623792
rect 1582 601024 1638 601080
rect 572718 640192 572774 640248
rect 579710 627680 579766 627736
rect 1582 578312 1638 578368
rect 1306 567296 1362 567352
rect 1582 556180 1584 556200
rect 1584 556180 1636 556200
rect 1636 556180 1638 556200
rect 1582 556144 1638 556180
rect 1582 533024 1638 533080
rect 1490 510584 1546 510640
rect 1398 465024 1454 465080
rect 1398 452376 1454 452432
rect 1398 419736 1454 419792
rect 1398 394984 1454 395040
rect 1306 337456 1362 337512
rect 1398 306312 1454 306368
rect 1398 294344 1454 294400
rect 1398 283736 1454 283792
rect 1398 261024 1454 261080
rect 1398 251232 1454 251288
rect 1306 238312 1362 238368
rect 1398 221484 1400 221504
rect 1400 221484 1452 221504
rect 1452 221484 1454 221504
rect 1398 221448 1454 221484
rect 1306 214512 1362 214568
rect 1398 198228 1400 198248
rect 1400 198228 1452 198248
rect 1452 198228 1454 198248
rect 1398 198192 1454 198228
rect 1306 193024 1362 193080
rect 1582 509904 1638 509960
rect 1582 487736 1638 487792
rect 1490 173032 1546 173088
rect 1490 170312 1546 170368
rect 1398 167592 1454 167648
rect 1398 165008 1454 165064
rect 570326 612448 570382 612504
rect 572718 585792 572774 585848
rect 1582 148688 1638 148744
rect 1582 146920 1638 146976
rect 1490 138644 1546 138680
rect 1490 138624 1492 138644
rect 1492 138624 1544 138644
rect 1544 138624 1546 138644
rect 580262 580760 580318 580816
rect 572718 558592 572774 558648
rect 3146 339632 3202 339688
rect 3146 321000 3202 321056
rect 580170 533840 580226 533896
rect 570326 530848 570382 530904
rect 570326 503648 570382 503704
rect 579802 486784 579858 486840
rect 570326 476448 570382 476504
rect 570326 449248 570382 449304
rect 580170 439864 580226 439920
rect 572718 422592 572774 422648
rect 570326 394848 570382 394904
rect 570326 367648 570382 367704
rect 572718 340992 572774 341048
rect 572718 313792 572774 313848
rect 570418 286048 570474 286104
rect 568394 248376 568450 248432
rect 570510 284588 570512 284608
rect 570512 284588 570564 284608
rect 570564 284588 570566 284608
rect 570510 284552 570566 284588
rect 569222 260072 569278 260128
rect 580170 392944 580226 393000
rect 574742 259392 574798 259448
rect 2870 185272 2926 185328
rect 568854 222264 568910 222320
rect 568578 193568 568634 193624
rect 568302 193432 568358 193488
rect 570326 193568 570382 193624
rect 1306 122032 1362 122088
rect 1214 108160 1270 108216
rect 1214 107072 1270 107128
rect 1306 99592 1362 99648
rect 1214 80824 1270 80880
rect 1306 57976 1362 58032
rect 1306 45872 1362 45928
rect 1214 33224 1270 33280
rect 1214 26988 1270 27024
rect 1214 26968 1216 26988
rect 1216 26968 1268 26988
rect 1268 26968 1270 26988
rect 1214 26832 1270 26888
rect 1122 12844 1178 12880
rect 1122 12824 1124 12844
rect 1124 12824 1176 12844
rect 1176 12824 1178 12844
rect 1122 12144 1178 12200
rect 1582 126384 1638 126440
rect 1398 35400 1454 35456
rect 1490 30232 1546 30288
rect 1398 29688 1454 29744
rect 1490 25744 1546 25800
rect 1398 20032 1454 20088
rect 1398 19760 1454 19816
rect 754 1264 810 1320
rect 662 720 718 776
rect 294 312 350 368
rect 1214 4392 1270 4448
rect 1214 992 1270 1048
rect 1582 8764 1638 8800
rect 1582 8744 1584 8764
rect 1584 8744 1636 8764
rect 1636 8744 1638 8764
rect 568486 174528 568542 174584
rect 569222 178472 569278 178528
rect 3514 96056 3570 96112
rect 3790 40296 3846 40352
rect 1490 1400 1546 1456
rect 1858 1536 1914 1592
rect 1766 856 1822 912
rect 1950 312 2006 368
rect 580170 346024 580226 346080
rect 574834 232192 574890 232248
rect 580170 299104 580226 299160
rect 574926 204992 574982 205048
rect 574742 150592 574798 150648
rect 580170 252184 580226 252240
rect 580170 205264 580226 205320
rect 575018 177792 575074 177848
rect 580170 158344 580226 158400
rect 572718 123392 572774 123448
rect 570326 99320 570382 99376
rect 572718 96192 572774 96248
rect 570326 90072 570382 90128
rect 580170 111424 580226 111480
rect 574742 68992 574798 69048
rect 20074 13232 20130 13288
rect 19982 7928 20038 7984
rect 225694 6432 225750 6488
rect 225786 5072 225842 5128
rect 124310 3712 124366 3768
rect 177946 3712 178002 3768
rect 268382 3712 268438 3768
rect 6090 1672 6146 1728
rect 6826 1672 6882 1728
rect 3698 1400 3754 1456
rect 5906 1420 5962 1456
rect 5906 1400 5908 1420
rect 5908 1400 5960 1420
rect 5960 1400 5962 1420
rect 6090 1400 6146 1456
rect 4986 584 5042 640
rect 3422 176 3478 232
rect 5630 584 5686 640
rect 7378 448 7434 504
rect 11242 1672 11298 1728
rect 14462 1672 14518 1728
rect 10414 1128 10470 1184
rect 10230 720 10286 776
rect 9862 76 9864 96
rect 9864 76 9916 96
rect 9916 76 9918 96
rect 9862 40 9918 76
rect 14462 1400 14518 1456
rect 14646 1400 14702 1456
rect 13634 856 13690 912
rect 14462 856 14518 912
rect 10690 312 10746 368
rect 10230 40 10286 96
rect 13266 584 13322 640
rect 13450 604 13506 640
rect 13450 584 13452 604
rect 13452 584 13504 604
rect 13504 584 13506 604
rect 12622 312 12678 368
rect 13082 176 13138 232
rect 14646 312 14702 368
rect 14554 176 14610 232
rect 15842 312 15898 368
rect 15014 176 15070 232
rect 22098 856 22154 912
rect 19338 176 19394 232
rect 20718 584 20774 640
rect 21914 584 21970 640
rect 37370 1672 37426 1728
rect 37738 1692 37794 1728
rect 37738 1672 37740 1692
rect 37740 1672 37792 1692
rect 37792 1672 37794 1692
rect 26422 1536 26478 1592
rect 26606 1536 26662 1592
rect 29734 1536 29790 1592
rect 32678 1536 32734 1592
rect 28262 1400 28318 1456
rect 26882 992 26938 1048
rect 27894 992 27950 1048
rect 23110 720 23166 776
rect 24306 720 24362 776
rect 19798 312 19854 368
rect 19706 176 19762 232
rect 27894 856 27950 912
rect 31482 1400 31538 1456
rect 28354 312 28410 368
rect 34978 856 35034 912
rect 30470 312 30526 368
rect 33690 448 33746 504
rect 35162 448 35218 504
rect 39394 1536 39450 1592
rect 40958 1672 41014 1728
rect 41142 1672 41198 1728
rect 48686 1708 48688 1728
rect 48688 1708 48740 1728
rect 48740 1708 48742 1728
rect 39302 1400 39358 1456
rect 39762 1536 39818 1592
rect 39302 1128 39358 1184
rect 38566 856 38622 912
rect 38198 756 38200 776
rect 38200 756 38252 776
rect 38252 756 38254 776
rect 38198 720 38254 756
rect 38382 720 38438 776
rect 48686 1672 48742 1708
rect 42522 1572 42524 1592
rect 42524 1572 42576 1592
rect 42576 1572 42578 1592
rect 42522 1536 42578 1572
rect 42706 1536 42762 1592
rect 42246 1400 42302 1456
rect 44086 1400 44142 1456
rect 45466 1400 45522 1456
rect 48042 1536 48098 1592
rect 48686 1536 48742 1592
rect 49330 1536 49386 1592
rect 45650 1400 45706 1456
rect 42062 1128 42118 1184
rect 42246 1128 42302 1184
rect 46570 992 46626 1048
rect 46754 992 46810 1048
rect 47030 992 47086 1048
rect 46294 720 46350 776
rect 46570 720 46626 776
rect 45558 448 45614 504
rect 47950 856 48006 912
rect 55034 1672 55090 1728
rect 55218 1672 55274 1728
rect 50802 1536 50858 1592
rect 50986 1536 51042 1592
rect 48134 856 48190 912
rect 46662 448 46718 504
rect 55034 1400 55090 1456
rect 48962 720 49018 776
rect 49514 720 49570 776
rect 49882 448 49938 504
rect 49514 176 49570 232
rect 50710 448 50766 504
rect 51814 176 51870 232
rect 55954 856 56010 912
rect 55678 720 55734 776
rect 56598 1400 56654 1456
rect 59082 1672 59138 1728
rect 59266 1672 59322 1728
rect 57886 1536 57942 1592
rect 58438 1536 58494 1592
rect 58530 1400 58586 1456
rect 64878 1672 64934 1728
rect 61014 1536 61070 1592
rect 61198 1536 61254 1592
rect 58162 1128 58218 1184
rect 58346 1128 58402 1184
rect 55954 176 56010 232
rect 56138 176 56194 232
rect 60278 1264 60334 1320
rect 60830 1264 60886 1320
rect 60738 1128 60794 1184
rect 57426 176 57482 232
rect 57794 176 57850 232
rect 62394 1400 62450 1456
rect 62946 1400 63002 1456
rect 63038 1264 63094 1320
rect 63314 1128 63370 1184
rect 63774 1264 63830 1320
rect 63498 992 63554 1048
rect 63866 1128 63922 1184
rect 61382 176 61438 232
rect 64510 1536 64566 1592
rect 65338 1536 65394 1592
rect 68834 1672 68890 1728
rect 72422 1672 72478 1728
rect 73710 1672 73766 1728
rect 66902 1556 66958 1592
rect 66902 1536 66904 1556
rect 66904 1536 66956 1556
rect 66956 1536 66958 1556
rect 66902 1400 66958 1456
rect 64786 1128 64842 1184
rect 66718 1128 66774 1184
rect 67086 1400 67142 1456
rect 64418 176 64474 232
rect 65338 448 65394 504
rect 65062 312 65118 368
rect 65338 312 65394 368
rect 66718 176 66774 232
rect 66902 212 66904 232
rect 66904 212 66956 232
rect 66956 212 66958 232
rect 66902 176 66958 212
rect 68098 448 68154 504
rect 68466 448 68522 504
rect 74078 1536 74134 1592
rect 73986 1400 74042 1456
rect 75366 1536 75422 1592
rect 76194 1536 76250 1592
rect 73342 992 73398 1048
rect 74262 992 74318 1048
rect 74446 992 74502 1048
rect 72606 448 72662 504
rect 72790 448 72846 504
rect 73342 312 73398 368
rect 73802 312 73858 368
rect 73526 212 73528 232
rect 73528 212 73580 232
rect 73580 212 73582 232
rect 73526 176 73582 212
rect 74078 448 74134 504
rect 74078 176 74134 232
rect 73894 40 73950 96
rect 74538 40 74594 96
rect 75734 448 75790 504
rect 75918 448 75974 504
rect 76194 448 76250 504
rect 77114 1536 77170 1592
rect 78402 1536 78458 1592
rect 78586 1536 78642 1592
rect 82266 1536 82322 1592
rect 77666 176 77722 232
rect 78494 448 78550 504
rect 78218 176 78274 232
rect 82174 1128 82230 1184
rect 82634 1672 82690 1728
rect 83738 1672 83794 1728
rect 85670 1672 85726 1728
rect 83186 1400 83242 1456
rect 83370 1400 83426 1456
rect 83646 1400 83702 1456
rect 78862 40 78918 96
rect 79230 448 79286 504
rect 80426 448 80482 504
rect 82450 856 82506 912
rect 82174 176 82230 232
rect 81622 40 81678 96
rect 82910 40 82966 96
rect 84198 176 84254 232
rect 84382 176 84438 232
rect 92570 1536 92626 1592
rect 92754 1536 92810 1592
rect 91926 1400 91982 1456
rect 85854 1264 85910 1320
rect 86038 1264 86094 1320
rect 92202 1264 92258 1320
rect 96434 1536 96490 1592
rect 96618 1536 96674 1592
rect 96986 1536 97042 1592
rect 100482 1672 100538 1728
rect 101678 1556 101734 1592
rect 101678 1536 101680 1556
rect 101680 1536 101732 1556
rect 101732 1536 101734 1556
rect 100942 1400 100998 1456
rect 101126 1400 101182 1456
rect 101310 1400 101366 1456
rect 96618 1264 96674 1320
rect 84198 40 84254 96
rect 87510 176 87566 232
rect 90730 1128 90786 1184
rect 92202 1164 92204 1184
rect 92204 1164 92256 1184
rect 92256 1164 92258 1184
rect 92202 1128 92258 1164
rect 91466 856 91522 912
rect 92110 856 92166 912
rect 91742 720 91798 776
rect 92018 720 92074 776
rect 92478 312 92534 368
rect 92662 312 92718 368
rect 93582 176 93638 232
rect 93766 176 93822 232
rect 97078 992 97134 1048
rect 97262 992 97318 1048
rect 93858 40 93914 96
rect 94134 40 94190 96
rect 97906 1264 97962 1320
rect 100206 1264 100262 1320
rect 101402 1264 101458 1320
rect 102782 1400 102838 1456
rect 103058 1400 103114 1456
rect 102322 1264 102378 1320
rect 101402 1128 101458 1184
rect 102598 1264 102654 1320
rect 97814 176 97870 232
rect 98274 176 98330 232
rect 103058 1264 103114 1320
rect 101034 40 101090 96
rect 102230 720 102286 776
rect 102690 740 102746 776
rect 102690 720 102692 740
rect 102692 720 102744 740
rect 102744 720 102746 740
rect 103426 1536 103482 1592
rect 103518 1264 103574 1320
rect 106738 1264 106794 1320
rect 104622 1164 104624 1184
rect 104624 1164 104676 1184
rect 104676 1164 104678 1184
rect 104622 1128 104678 1164
rect 104806 1148 104862 1184
rect 104806 1128 104808 1148
rect 104808 1128 104860 1148
rect 104860 1128 104862 1148
rect 103794 720 103850 776
rect 103978 720 104034 776
rect 101770 40 101826 96
rect 101954 40 102010 96
rect 106830 1128 106886 1184
rect 107106 992 107162 1048
rect 107382 1128 107438 1184
rect 109038 992 109094 1048
rect 111430 1672 111486 1728
rect 110786 1400 110842 1456
rect 111246 1536 111302 1592
rect 112166 1572 112168 1592
rect 112168 1572 112220 1592
rect 112220 1572 112222 1592
rect 112166 1536 112222 1572
rect 111246 1436 111248 1456
rect 111248 1436 111300 1456
rect 111300 1436 111302 1456
rect 111246 1400 111302 1436
rect 111430 1420 111486 1456
rect 111430 1400 111432 1420
rect 111432 1400 111484 1420
rect 111484 1400 111486 1420
rect 111982 1400 112038 1456
rect 110326 1128 110382 1184
rect 109222 992 109278 1048
rect 110510 1164 110512 1184
rect 110512 1164 110564 1184
rect 110564 1164 110566 1184
rect 110510 1128 110566 1164
rect 111614 1128 111670 1184
rect 112626 1128 112682 1184
rect 107382 720 107438 776
rect 107842 740 107898 776
rect 107842 720 107844 740
rect 107844 720 107896 740
rect 107896 720 107898 740
rect 108578 40 108634 96
rect 111614 584 111670 640
rect 111798 584 111854 640
rect 108946 176 109002 232
rect 111890 448 111946 504
rect 111706 176 111762 232
rect 112074 584 112130 640
rect 112350 584 112406 640
rect 112074 448 112130 504
rect 113730 756 113732 776
rect 113732 756 113784 776
rect 113784 756 113786 776
rect 113730 720 113786 756
rect 114098 584 114154 640
rect 120630 1672 120686 1728
rect 116858 1264 116914 1320
rect 117042 1264 117098 1320
rect 120170 1536 120226 1592
rect 120630 1400 120686 1456
rect 120906 1400 120962 1456
rect 120354 1128 120410 1184
rect 116398 720 116454 776
rect 116582 720 116638 776
rect 115754 584 115810 640
rect 115938 584 115994 640
rect 112626 40 112682 96
rect 116582 176 116638 232
rect 116858 176 116914 232
rect 122286 1672 122342 1728
rect 124310 1672 124366 1728
rect 121918 1536 121974 1592
rect 121826 1264 121882 1320
rect 122010 1264 122066 1320
rect 125782 1672 125838 1728
rect 128266 1708 128268 1728
rect 128268 1708 128320 1728
rect 128320 1708 128322 1728
rect 128266 1672 128322 1708
rect 127806 1536 127862 1592
rect 127714 1400 127770 1456
rect 127990 1536 128046 1592
rect 127898 1400 127954 1456
rect 129002 1672 129058 1728
rect 135166 1692 135222 1728
rect 135166 1672 135168 1692
rect 135168 1672 135220 1692
rect 135220 1672 135222 1692
rect 134890 1536 134946 1592
rect 135350 1672 135406 1728
rect 135626 1672 135682 1728
rect 136270 1672 136326 1728
rect 135074 1536 135130 1592
rect 129002 1400 129058 1456
rect 120906 584 120962 640
rect 121182 584 121238 640
rect 122746 720 122802 776
rect 119618 40 119674 96
rect 122654 312 122710 368
rect 123298 312 123354 368
rect 125506 1128 125562 1184
rect 126702 1128 126758 1184
rect 128450 1128 128506 1184
rect 123574 992 123630 1048
rect 123758 992 123814 1048
rect 128818 992 128874 1048
rect 123758 584 123814 640
rect 123942 584 123998 640
rect 129094 720 129150 776
rect 134798 1420 134854 1456
rect 134798 1400 134800 1420
rect 134800 1400 134852 1420
rect 134852 1400 134854 1420
rect 131302 1264 131358 1320
rect 124218 584 124274 640
rect 129646 720 129702 776
rect 131486 1264 131542 1320
rect 131486 992 131542 1048
rect 131670 1264 131726 1320
rect 134706 1264 134762 1320
rect 135534 1400 135590 1456
rect 135074 1264 135130 1320
rect 135902 1264 135958 1320
rect 136362 1264 136418 1320
rect 136546 1536 136602 1592
rect 136914 1400 136970 1456
rect 136914 1264 136970 1320
rect 138386 1692 138442 1728
rect 138386 1672 138388 1692
rect 138388 1672 138440 1692
rect 138440 1672 138442 1692
rect 137190 1264 137246 1320
rect 135534 1128 135590 1184
rect 131670 1012 131726 1048
rect 131670 992 131672 1012
rect 131672 992 131724 1012
rect 131724 992 131726 1012
rect 135810 992 135866 1048
rect 138386 856 138442 912
rect 129278 448 129334 504
rect 129922 448 129978 504
rect 136086 720 136142 776
rect 139214 1420 139270 1456
rect 139214 1400 139216 1420
rect 139216 1400 139268 1420
rect 139268 1400 139270 1420
rect 139582 1400 139638 1456
rect 139766 1128 139822 1184
rect 140042 1400 140098 1456
rect 140226 1400 140282 1456
rect 139030 992 139086 1048
rect 139398 856 139454 912
rect 139582 856 139638 912
rect 139398 720 139454 776
rect 139582 720 139638 776
rect 135350 584 135406 640
rect 141146 1672 141202 1728
rect 144366 1672 144422 1728
rect 145102 1672 145158 1728
rect 140778 1536 140834 1592
rect 140962 1536 141018 1592
rect 141238 1400 141294 1456
rect 141514 1400 141570 1456
rect 141330 1128 141386 1184
rect 140042 584 140098 640
rect 142250 720 142306 776
rect 142434 720 142490 776
rect 145010 1536 145066 1592
rect 145654 1672 145710 1728
rect 145838 1708 145840 1728
rect 145840 1708 145892 1728
rect 145892 1708 145894 1728
rect 145838 1672 145894 1708
rect 146206 1708 146208 1728
rect 146208 1708 146260 1728
rect 146260 1708 146262 1728
rect 146206 1672 146262 1708
rect 145838 1536 145894 1592
rect 147402 1536 147458 1592
rect 145286 1128 145342 1184
rect 145470 1128 145526 1184
rect 144182 720 144238 776
rect 148046 1672 148102 1728
rect 147862 1264 147918 1320
rect 148966 1672 149022 1728
rect 148690 1536 148746 1592
rect 148690 1264 148746 1320
rect 148874 1264 148930 1320
rect 148598 1128 148654 1184
rect 149150 1672 149206 1728
rect 149058 1264 149114 1320
rect 149242 1128 149298 1184
rect 145746 720 145802 776
rect 146942 720 146998 776
rect 154302 1672 154358 1728
rect 151542 1400 151598 1456
rect 151818 1400 151874 1456
rect 153934 1536 153990 1592
rect 152002 1264 152058 1320
rect 150898 1128 150954 1184
rect 150254 620 150256 640
rect 150256 620 150308 640
rect 150308 620 150310 640
rect 150254 584 150310 620
rect 151174 856 151230 912
rect 152370 1264 152426 1320
rect 152554 1264 152610 1320
rect 158810 1672 158866 1728
rect 158994 1672 159050 1728
rect 154118 1264 154174 1320
rect 151082 584 151138 640
rect 150806 448 150862 504
rect 151450 584 151506 640
rect 153382 992 153438 1048
rect 153566 992 153622 1048
rect 157522 1264 157578 1320
rect 157982 1400 158038 1456
rect 158166 1400 158222 1456
rect 157062 992 157118 1048
rect 157246 992 157302 1048
rect 157890 1128 157946 1184
rect 158074 1128 158130 1184
rect 158442 1148 158498 1184
rect 158442 1128 158444 1148
rect 158444 1128 158496 1148
rect 158496 1128 158498 1148
rect 158626 1128 158682 1184
rect 150990 176 151046 232
rect 151818 176 151874 232
rect 153106 312 153162 368
rect 153290 312 153346 368
rect 157154 584 157210 640
rect 157614 620 157616 640
rect 157616 620 157668 640
rect 157668 620 157670 640
rect 156878 448 156934 504
rect 157154 448 157210 504
rect 156878 312 156934 368
rect 157614 584 157670 620
rect 158994 1400 159050 1456
rect 160282 1556 160338 1592
rect 160282 1536 160284 1556
rect 160284 1536 160336 1556
rect 160336 1536 160338 1556
rect 161202 1536 161258 1592
rect 159638 1400 159694 1456
rect 159362 1264 159418 1320
rect 159546 1264 159602 1320
rect 159270 1128 159326 1184
rect 159454 1128 159510 1184
rect 161846 1264 161902 1320
rect 164238 1400 164294 1456
rect 163778 1264 163834 1320
rect 166814 1672 166870 1728
rect 169114 1692 169170 1728
rect 169114 1672 169116 1692
rect 169116 1672 169168 1692
rect 169168 1672 169170 1692
rect 157890 584 157946 640
rect 157338 312 157394 368
rect 158074 584 158130 640
rect 157798 312 157854 368
rect 166354 1128 166410 1184
rect 163686 992 163742 1048
rect 166630 992 166686 1048
rect 166814 992 166870 1048
rect 161478 720 161534 776
rect 161754 720 161810 776
rect 163134 720 163190 776
rect 161386 312 161442 368
rect 161754 584 161810 640
rect 163686 720 163742 776
rect 163870 740 163926 776
rect 163870 720 163872 740
rect 163872 720 163924 740
rect 163924 720 163926 740
rect 163502 584 163558 640
rect 169022 1400 169078 1456
rect 169206 1420 169262 1456
rect 169206 1400 169208 1420
rect 169208 1400 169260 1420
rect 169260 1400 169262 1420
rect 168930 1264 168986 1320
rect 168654 1128 168710 1184
rect 169114 1264 169170 1320
rect 169390 1128 169446 1184
rect 169574 1128 169630 1184
rect 170770 1264 170826 1320
rect 170494 1128 170550 1184
rect 171046 1536 171102 1592
rect 171598 1536 171654 1592
rect 173346 1400 173402 1456
rect 173806 1264 173862 1320
rect 173254 1128 173310 1184
rect 176290 1128 176346 1184
rect 177118 1128 177174 1184
rect 169666 584 169722 640
rect 169850 584 169906 640
rect 170034 584 170090 640
rect 163134 312 163190 368
rect 163318 312 163374 368
rect 176014 740 176070 776
rect 176014 720 176016 740
rect 176016 720 176068 740
rect 176068 720 176070 740
rect 176198 720 176254 776
rect 178774 1672 178830 1728
rect 179050 1692 179106 1728
rect 179050 1672 179052 1692
rect 179052 1672 179104 1692
rect 179104 1672 179106 1692
rect 177670 1536 177726 1592
rect 177762 1264 177818 1320
rect 178038 1284 178094 1320
rect 178314 1400 178370 1456
rect 178038 1264 178040 1284
rect 178040 1264 178092 1284
rect 178092 1264 178094 1284
rect 177670 1128 177726 1184
rect 178682 1400 178738 1456
rect 179142 1128 179198 1184
rect 179326 1128 179382 1184
rect 179878 1536 179934 1592
rect 179694 1264 179750 1320
rect 181718 1536 181774 1592
rect 184662 1536 184718 1592
rect 183742 1400 183798 1456
rect 184386 1400 184442 1456
rect 180246 1264 180302 1320
rect 180798 1128 180854 1184
rect 177394 584 177450 640
rect 177946 620 177948 640
rect 177948 620 178000 640
rect 178000 620 178002 640
rect 177946 584 178002 620
rect 182638 1264 182694 1320
rect 182914 1128 182970 1184
rect 184202 1128 184258 1184
rect 183926 992 183982 1048
rect 184294 992 184350 1048
rect 184202 720 184258 776
rect 184386 720 184442 776
rect 190642 1672 190698 1728
rect 190642 1536 190698 1592
rect 189630 1264 189686 1320
rect 185858 1128 185914 1184
rect 186502 1128 186558 1184
rect 190366 1128 190422 1184
rect 189906 992 189962 1048
rect 190918 1672 190974 1728
rect 192206 1672 192262 1728
rect 196438 1672 196494 1728
rect 196714 1672 196770 1728
rect 190918 1400 190974 1456
rect 190826 1128 190882 1184
rect 191102 1264 191158 1320
rect 191562 1128 191618 1184
rect 191378 992 191434 1048
rect 190458 720 190514 776
rect 195978 1536 196034 1592
rect 196714 1128 196770 1184
rect 197174 992 197230 1048
rect 198094 1128 198150 1184
rect 198738 1672 198794 1728
rect 200026 1672 200082 1728
rect 207294 1672 207350 1728
rect 208122 1672 208178 1728
rect 199106 1556 199162 1592
rect 199106 1536 199108 1556
rect 199108 1536 199160 1556
rect 199160 1536 199162 1556
rect 199750 1536 199806 1592
rect 204442 1536 204498 1592
rect 216678 1672 216734 1728
rect 204810 1536 204866 1592
rect 200302 1400 200358 1456
rect 198370 992 198426 1048
rect 190642 448 190698 504
rect 191286 448 191342 504
rect 197726 856 197782 912
rect 198186 856 198242 912
rect 197542 720 197598 776
rect 197358 584 197414 640
rect 198646 720 198702 776
rect 197634 448 197690 504
rect 198462 584 198518 640
rect 198186 448 198242 504
rect 198370 468 198426 504
rect 198370 448 198372 468
rect 198372 448 198424 468
rect 198424 448 198426 468
rect 198370 176 198426 232
rect 198554 176 198610 232
rect 205454 1536 205510 1592
rect 207294 1536 207350 1592
rect 207478 1536 207534 1592
rect 207754 1400 207810 1456
rect 204258 584 204314 640
rect 208030 1264 208086 1320
rect 211342 1536 211398 1592
rect 209042 1128 209098 1184
rect 209226 1128 209282 1184
rect 209870 1264 209926 1320
rect 212170 1400 212226 1456
rect 214378 1400 214434 1456
rect 209502 1128 209558 1184
rect 216770 1400 216826 1456
rect 216954 1400 217010 1456
rect 218150 1400 218206 1456
rect 211894 1128 211950 1184
rect 214838 1264 214894 1320
rect 215022 1264 215078 1320
rect 217414 1264 217470 1320
rect 217966 1264 218022 1320
rect 220450 1672 220506 1728
rect 232134 1672 232190 1728
rect 234066 1672 234122 1728
rect 223946 1400 224002 1456
rect 224498 1400 224554 1456
rect 217874 1128 217930 1184
rect 204534 584 204590 640
rect 205086 584 205142 640
rect 207846 620 207848 640
rect 207848 620 207900 640
rect 207900 620 207902 640
rect 207846 584 207902 620
rect 211434 584 211490 640
rect 215022 620 215024 640
rect 215024 620 215076 640
rect 215076 620 215078 640
rect 215022 584 215078 620
rect 215206 584 215262 640
rect 217782 584 217838 640
rect 221094 720 221150 776
rect 217966 584 218022 640
rect 219346 584 219402 640
rect 221646 1264 221702 1320
rect 221370 584 221426 640
rect 224406 720 224462 776
rect 225418 1400 225474 1456
rect 224590 720 224646 776
rect 225050 1264 225106 1320
rect 225234 1264 225290 1320
rect 224958 1128 225014 1184
rect 225142 1128 225198 1184
rect 225326 1128 225382 1184
rect 225694 1536 225750 1592
rect 225878 1536 225934 1592
rect 231766 1536 231822 1592
rect 225786 1264 225842 1320
rect 227442 1264 227498 1320
rect 226614 1128 226670 1184
rect 232134 1264 232190 1320
rect 232502 1264 232558 1320
rect 231490 856 231546 912
rect 231306 720 231362 776
rect 233146 856 233202 912
rect 238022 1264 238078 1320
rect 238390 1672 238446 1728
rect 238942 1536 238998 1592
rect 238666 1400 238722 1456
rect 238206 1264 238262 1320
rect 233330 856 233386 912
rect 232962 584 233018 640
rect 238206 720 238262 776
rect 238390 720 238446 776
rect 239126 720 239182 776
rect 239310 720 239366 776
rect 233146 620 233148 640
rect 233148 620 233200 640
rect 233200 620 233202 640
rect 233146 584 233202 620
rect 224314 312 224370 368
rect 224682 312 224738 368
rect 242070 1536 242126 1592
rect 242898 1400 242954 1456
rect 245290 1400 245346 1456
rect 245474 1672 245530 1728
rect 245014 720 245070 776
rect 247682 1672 247738 1728
rect 250074 1672 250130 1728
rect 246762 856 246818 912
rect 246946 856 247002 912
rect 248970 1400 249026 1456
rect 247314 1264 247370 1320
rect 247406 992 247462 1048
rect 247774 992 247830 1048
rect 249982 1400 250038 1456
rect 250626 1264 250682 1320
rect 251546 1400 251602 1456
rect 250534 992 250590 1048
rect 250718 992 250774 1048
rect 247866 720 247922 776
rect 250166 856 250222 912
rect 252742 1264 252798 1320
rect 252742 1128 252798 1184
rect 253018 1128 253074 1184
rect 251638 992 251694 1048
rect 247590 584 247646 640
rect 248418 584 248474 640
rect 248326 312 248382 368
rect 248786 312 248842 368
rect 248418 176 248474 232
rect 248694 176 248750 232
rect 252466 856 252522 912
rect 252926 856 252982 912
rect 253294 992 253350 1048
rect 256606 1536 256662 1592
rect 254030 1400 254086 1456
rect 253846 1264 253902 1320
rect 254030 1284 254086 1320
rect 254214 1400 254270 1456
rect 254030 1264 254032 1284
rect 254032 1264 254084 1284
rect 254084 1264 254086 1284
rect 256514 1284 256570 1320
rect 258078 1672 258134 1728
rect 262034 1672 262090 1728
rect 257066 1400 257122 1456
rect 258078 1400 258134 1456
rect 259090 1420 259146 1456
rect 259090 1400 259092 1420
rect 259092 1400 259144 1420
rect 259144 1400 259146 1420
rect 256514 1264 256516 1284
rect 256516 1264 256568 1284
rect 256568 1264 256570 1284
rect 255870 992 255926 1048
rect 253662 856 253718 912
rect 255962 720 256018 776
rect 258354 720 258410 776
rect 260470 1400 260526 1456
rect 262034 1536 262090 1592
rect 260654 1400 260710 1456
rect 261206 1264 261262 1320
rect 261390 1264 261446 1320
rect 261942 992 261998 1048
rect 262310 992 262366 1048
rect 262494 992 262550 1048
rect 260838 720 260894 776
rect 261574 620 261576 640
rect 261576 620 261628 640
rect 261628 620 261630 640
rect 261574 584 261630 620
rect 261850 720 261906 776
rect 262678 1264 262734 1320
rect 265346 1264 265402 1320
rect 262678 720 262734 776
rect 262862 720 262918 776
rect 262586 584 262642 640
rect 268474 1672 268530 1728
rect 268382 1536 268438 1592
rect 268842 1672 268898 1728
rect 268014 1400 268070 1456
rect 268842 1436 268844 1456
rect 268844 1436 268896 1456
rect 268896 1436 268898 1456
rect 268842 1400 268898 1436
rect 269026 1400 269082 1456
rect 270958 1536 271014 1592
rect 271878 1536 271934 1592
rect 265990 720 266046 776
rect 266266 720 266322 776
rect 269210 1128 269266 1184
rect 266818 584 266874 640
rect 267002 620 267004 640
rect 267004 620 267056 640
rect 267056 620 267058 640
rect 267002 584 267058 620
rect 265070 176 265126 232
rect 265622 176 265678 232
rect 271234 1400 271290 1456
rect 271418 1264 271474 1320
rect 271050 720 271106 776
rect 271234 720 271290 776
rect 279330 1672 279386 1728
rect 273534 1400 273590 1456
rect 273258 1128 273314 1184
rect 273442 1128 273498 1184
rect 279790 1536 279846 1592
rect 279974 1536 280030 1592
rect 280158 1536 280214 1592
rect 280526 1572 280528 1592
rect 280528 1572 280580 1592
rect 280580 1572 280582 1592
rect 280526 1536 280582 1572
rect 279422 1128 279478 1184
rect 280526 1264 280582 1320
rect 279882 720 279938 776
rect 280250 720 280306 776
rect 280986 1264 281042 1320
rect 285770 1672 285826 1728
rect 281538 1400 281594 1456
rect 281722 1436 281724 1456
rect 281724 1436 281776 1456
rect 281776 1436 281778 1456
rect 281722 1400 281778 1436
rect 285310 1400 285366 1456
rect 285954 1400 286010 1456
rect 281906 720 281962 776
rect 282090 720 282146 776
rect 285310 720 285366 776
rect 287518 1128 287574 1184
rect 285678 992 285734 1048
rect 285770 720 285826 776
rect 287794 1128 287850 1184
rect 289634 1264 289690 1320
rect 289542 1128 289598 1184
rect 290370 1128 290426 1184
rect 294602 1672 294658 1728
rect 294970 1672 295026 1728
rect 295614 1536 295670 1592
rect 295798 1536 295854 1592
rect 296258 1536 296314 1592
rect 294694 1264 294750 1320
rect 294970 1264 295026 1320
rect 295154 1264 295210 1320
rect 293866 992 293922 1048
rect 290370 740 290426 776
rect 290370 720 290372 740
rect 290372 720 290424 740
rect 290424 720 290426 740
rect 294786 720 294842 776
rect 296718 1128 296774 1184
rect 296902 1012 296958 1048
rect 296902 992 296904 1012
rect 296904 992 296956 1012
rect 296956 992 296958 1012
rect 309966 1672 310022 1728
rect 305642 1556 305698 1592
rect 305642 1536 305644 1556
rect 305644 1536 305696 1556
rect 305696 1536 305698 1556
rect 305826 1536 305882 1592
rect 307022 1536 307078 1592
rect 307206 1536 307262 1592
rect 309230 1536 309286 1592
rect 299938 992 299994 1048
rect 303434 992 303490 1048
rect 306930 1012 306986 1048
rect 306930 992 306932 1012
rect 306932 992 306984 1012
rect 306984 992 306986 1012
rect 307114 992 307170 1048
rect 295246 720 295302 776
rect 321742 1672 321798 1728
rect 321926 1672 321982 1728
rect 347410 1672 347466 1728
rect 348330 1672 348386 1728
rect 308954 1128 309010 1184
rect 309322 992 309378 1048
rect 309966 1128 310022 1184
rect 309782 856 309838 912
rect 319534 1536 319590 1592
rect 319718 1536 319774 1592
rect 317694 1264 317750 1320
rect 318338 1264 318394 1320
rect 314750 856 314806 912
rect 318614 1264 318670 1320
rect 322938 1264 322994 1320
rect 321926 1128 321982 1184
rect 322110 1128 322166 1184
rect 323122 1264 323178 1320
rect 324962 1264 325018 1320
rect 327538 1284 327594 1320
rect 327538 1264 327540 1284
rect 327540 1264 327592 1284
rect 327592 1264 327594 1284
rect 327722 1264 327778 1320
rect 327906 1264 327962 1320
rect 326894 992 326950 1048
rect 327078 992 327134 1048
rect 327262 992 327318 1048
rect 328826 1128 328882 1184
rect 329746 1128 329802 1184
rect 331770 1128 331826 1184
rect 328550 856 328606 912
rect 329654 856 329710 912
rect 329838 856 329894 912
rect 331954 1128 332010 1184
rect 335818 1128 335874 1184
rect 336002 1128 336058 1184
rect 336002 856 336058 912
rect 336186 856 336242 912
rect 336186 584 336242 640
rect 336370 584 336426 640
rect 348330 1128 348386 1184
rect 373722 1672 373778 1728
rect 373906 1672 373962 1728
rect 380162 1672 380218 1728
rect 380346 1672 380402 1728
rect 389086 1672 389142 1728
rect 395434 1672 395490 1728
rect 398654 1672 398710 1728
rect 399574 1672 399630 1728
rect 403714 1672 403770 1728
rect 352930 1536 352986 1592
rect 349526 892 349528 912
rect 349528 892 349580 912
rect 349580 892 349582 912
rect 349526 856 349582 892
rect 352194 856 352250 912
rect 356242 892 356244 912
rect 356244 892 356296 912
rect 356296 892 356298 912
rect 356242 856 356298 892
rect 356426 856 356482 912
rect 348698 720 348754 776
rect 354034 720 354090 776
rect 357622 720 357678 776
rect 343086 584 343142 640
rect 356518 584 356574 640
rect 356978 584 357034 640
rect 365994 1536 366050 1592
rect 366178 1536 366234 1592
rect 364706 1264 364762 1320
rect 365994 1264 366050 1320
rect 364706 720 364762 776
rect 373354 1264 373410 1320
rect 366178 1128 366234 1184
rect 372526 1128 372582 1184
rect 373722 1128 373778 1184
rect 373354 720 373410 776
rect 376758 720 376814 776
rect 365074 584 365130 640
rect 365258 584 365314 640
rect 358174 312 358230 368
rect 415674 1692 415730 1728
rect 415674 1672 415676 1692
rect 415676 1672 415728 1692
rect 415728 1672 415730 1692
rect 418802 1692 418858 1728
rect 418802 1672 418804 1692
rect 418804 1672 418856 1692
rect 418856 1672 418858 1692
rect 432326 1692 432382 1728
rect 432326 1672 432328 1692
rect 432328 1672 432380 1692
rect 432380 1672 432382 1692
rect 436006 1672 436062 1728
rect 443458 1672 443514 1728
rect 443642 1692 443698 1728
rect 443642 1672 443644 1692
rect 443644 1672 443696 1692
rect 443696 1672 443698 1692
rect 406842 1536 406898 1592
rect 407026 1536 407082 1592
rect 415122 1536 415178 1592
rect 418802 1536 418858 1592
rect 406658 1264 406714 1320
rect 406842 1264 406898 1320
rect 389086 1128 389142 1184
rect 389362 1128 389418 1184
rect 381542 720 381598 776
rect 406106 756 406108 776
rect 406108 756 406160 776
rect 406160 756 406162 776
rect 406106 720 406162 756
rect 406382 720 406438 776
rect 380346 584 380402 640
rect 386050 584 386106 640
rect 393410 584 393466 640
rect 365074 312 365130 368
rect 386050 312 386106 368
rect 411258 584 411314 640
rect 406382 312 406438 368
rect 406658 312 406714 368
rect 418802 1264 418858 1320
rect 453302 1692 453358 1728
rect 453302 1672 453304 1692
rect 453304 1672 453356 1692
rect 453356 1672 453358 1692
rect 462870 1692 462926 1728
rect 462870 1672 462872 1692
rect 462872 1672 462924 1692
rect 462924 1672 462926 1692
rect 474922 1708 474924 1728
rect 474924 1708 474976 1728
rect 474976 1708 474978 1728
rect 474922 1672 474978 1708
rect 481270 1708 481272 1728
rect 481272 1708 481324 1728
rect 481324 1708 481326 1728
rect 481270 1672 481326 1708
rect 488998 1708 489000 1728
rect 489000 1708 489052 1728
rect 489052 1708 489054 1728
rect 488998 1672 489054 1708
rect 501786 1708 501788 1728
rect 501788 1708 501840 1728
rect 501840 1708 501842 1728
rect 501786 1672 501842 1708
rect 512366 1708 512368 1728
rect 512368 1708 512420 1728
rect 512420 1708 512422 1728
rect 512366 1672 512422 1708
rect 522578 1672 522634 1728
rect 529386 1708 529388 1728
rect 529388 1708 529440 1728
rect 529440 1708 529442 1728
rect 529386 1672 529442 1708
rect 567290 1708 567292 1728
rect 567292 1708 567344 1728
rect 567344 1708 567346 1728
rect 440698 1536 440754 1592
rect 453210 1572 453212 1592
rect 453212 1572 453264 1592
rect 453264 1572 453266 1592
rect 453210 1536 453266 1572
rect 462594 1536 462650 1592
rect 471518 1536 471574 1592
rect 436006 1264 436062 1320
rect 443182 1264 443238 1320
rect 453302 1264 453358 1320
rect 460570 1264 460626 1320
rect 462594 1264 462650 1320
rect 476394 1264 476450 1320
rect 476578 1264 476634 1320
rect 440698 1128 440754 1184
rect 415122 584 415178 640
rect 413650 312 413706 368
rect 434994 740 435050 776
rect 434994 720 434996 740
rect 434996 720 435048 740
rect 435048 720 435050 740
rect 427818 584 427874 640
rect 425702 312 425758 368
rect 442814 584 442870 640
rect 427818 312 427874 368
rect 442722 448 442778 504
rect 460570 720 460626 776
rect 443182 312 443238 368
rect 482190 1264 482246 1320
rect 476578 720 476634 776
rect 476762 584 476818 640
rect 501326 1264 501382 1320
rect 504178 1264 504234 1320
rect 482190 720 482246 776
rect 461674 176 461730 232
rect 473358 176 473414 232
rect 473726 176 473782 232
rect 486146 176 486202 232
rect 490194 584 490250 640
rect 504178 720 504234 776
rect 509054 584 509110 640
rect 516690 1264 516746 1320
rect 516874 1264 516930 1320
rect 512642 720 512698 776
rect 515586 720 515642 776
rect 516690 720 516746 776
rect 522578 584 522634 640
rect 509882 448 509938 504
rect 537298 1264 537354 1320
rect 538770 1264 538826 1320
rect 556434 1400 556490 1456
rect 531778 1128 531834 1184
rect 531778 720 531834 776
rect 536930 720 536986 776
rect 536746 584 536802 640
rect 528834 312 528890 368
rect 552478 1264 552534 1320
rect 567290 1672 567346 1708
rect 559102 1536 559158 1592
rect 559378 1536 559434 1592
rect 565818 1536 565874 1592
rect 552754 1128 552810 1184
rect 557998 1128 558054 1184
rect 538770 312 538826 368
rect 538954 312 539010 368
rect 545670 448 545726 504
rect 545670 176 545726 232
rect 565818 1420 565874 1456
rect 565818 1400 565820 1420
rect 565820 1400 565872 1420
rect 565872 1400 565874 1420
rect 559562 1264 559618 1320
rect 564438 1284 564494 1320
rect 564438 1264 564440 1284
rect 564440 1264 564492 1284
rect 564492 1264 564494 1284
rect 580170 64504 580226 64560
rect 574742 41792 574798 41848
rect 570326 34856 570382 34912
rect 568394 1128 568450 1184
rect 568670 992 568726 1048
rect 559562 720 559618 776
rect 569130 720 569186 776
rect 559378 312 559434 368
rect 580170 17584 580226 17640
rect 571614 14592 571670 14648
rect 570326 12280 570382 12336
rect 569590 1672 569646 1728
rect 570326 4392 570382 4448
rect 569682 40 569738 96
<< metal3 >>
rect 583520 697900 584960 698140
rect -960 696540 480 696780
rect 583520 686204 584960 686444
rect -960 682274 480 682364
rect 1393 682274 1459 682277
rect -960 682272 1459 682274
rect -960 682216 1398 682272
rect 1454 682216 1459 682272
rect -960 682214 1459 682216
rect -960 682124 480 682214
rect 1393 682211 1459 682214
rect 550582 680988 550588 681052
rect 550652 681050 550658 681052
rect 564709 681050 564775 681053
rect 550652 681048 564775 681050
rect 550652 680992 564714 681048
rect 564770 680992 564775 681048
rect 550652 680990 564775 680992
rect 550652 680988 550658 680990
rect 564709 680987 564775 680990
rect 434662 680852 434668 680916
rect 434732 680914 434738 680916
rect 439497 680914 439563 680917
rect 434732 680912 439563 680914
rect 434732 680856 439502 680912
rect 439558 680856 439563 680912
rect 434732 680854 439563 680856
rect 434732 680852 434738 680854
rect 439497 680851 439563 680854
rect 559782 680778 559788 680780
rect 364382 680718 366098 680778
rect 344870 680580 344876 680644
rect 344940 680642 344946 680644
rect 345013 680642 345079 680645
rect 344940 680640 345079 680642
rect 344940 680584 345018 680640
rect 345074 680584 345079 680640
rect 344940 680582 345079 680584
rect 344940 680580 344946 680582
rect 345013 680579 345079 680582
rect 325601 680506 325667 680509
rect 364382 680506 364442 680718
rect 325601 680504 364442 680506
rect 325601 680448 325606 680504
rect 325662 680448 364442 680504
rect 325601 680446 364442 680448
rect 325601 680443 325667 680446
rect 296713 680370 296779 680373
rect 364793 680370 364859 680373
rect 296713 680368 364859 680370
rect 296713 680312 296718 680368
rect 296774 680312 364798 680368
rect 364854 680312 364859 680368
rect 296713 680310 364859 680312
rect 366038 680370 366098 680718
rect 418110 680718 419642 680778
rect 379421 680642 379487 680645
rect 369902 680640 379487 680642
rect 369902 680584 379426 680640
rect 379482 680584 379487 680640
rect 369902 680582 379487 680584
rect 369902 680370 369962 680582
rect 379421 680579 379487 680582
rect 418110 680506 418170 680718
rect 393454 680446 403450 680506
rect 366038 680310 369962 680370
rect 370221 680370 370287 680373
rect 380065 680370 380131 680373
rect 370221 680368 380131 680370
rect 370221 680312 370226 680368
rect 370282 680312 380070 680368
rect 380126 680312 380131 680368
rect 370221 680310 380131 680312
rect 296713 680307 296779 680310
rect 364793 680307 364859 680310
rect 370221 680307 370287 680310
rect 380065 680307 380131 680310
rect 381629 680370 381695 680373
rect 393454 680370 393514 680446
rect 381629 680368 393514 680370
rect 381629 680312 381634 680368
rect 381690 680312 393514 680368
rect 381629 680310 393514 680312
rect 394693 680370 394759 680373
rect 403157 680370 403223 680373
rect 394693 680368 403223 680370
rect 394693 680312 394698 680368
rect 394754 680312 403162 680368
rect 403218 680312 403223 680368
rect 394693 680310 403223 680312
rect 403390 680370 403450 680446
rect 412590 680446 418170 680506
rect 412590 680370 412650 680446
rect 403390 680310 412650 680370
rect 412725 680370 412791 680373
rect 418613 680370 418679 680373
rect 412725 680368 418679 680370
rect 412725 680312 412730 680368
rect 412786 680312 418618 680368
rect 418674 680312 418679 680368
rect 412725 680310 418679 680312
rect 419582 680370 419642 680718
rect 456750 680718 458282 680778
rect 434662 680642 434668 680644
rect 427862 680582 434668 680642
rect 427862 680370 427922 680582
rect 434662 680580 434668 680582
rect 434732 680580 434738 680644
rect 456750 680506 456810 680718
rect 451230 680446 456810 680506
rect 419582 680310 427922 680370
rect 428181 680370 428247 680373
rect 437749 680370 437815 680373
rect 428181 680368 437815 680370
rect 428181 680312 428186 680368
rect 428242 680312 437754 680368
rect 437810 680312 437815 680368
rect 428181 680310 437815 680312
rect 381629 680307 381695 680310
rect 394693 680307 394759 680310
rect 403157 680307 403223 680310
rect 412725 680307 412791 680310
rect 418613 680307 418679 680310
rect 428181 680307 428247 680310
rect 437749 680307 437815 680310
rect 439497 680370 439563 680373
rect 451230 680370 451290 680446
rect 439497 680368 451290 680370
rect 439497 680312 439502 680368
rect 439558 680312 451290 680368
rect 439497 680310 451290 680312
rect 451365 680370 451431 680373
rect 457161 680370 457227 680373
rect 451365 680368 457227 680370
rect 451365 680312 451370 680368
rect 451426 680312 457166 680368
rect 457222 680312 457227 680368
rect 451365 680310 457227 680312
rect 458222 680370 458282 680718
rect 534030 680718 535562 680778
rect 466637 680506 466703 680509
rect 534030 680506 534090 680718
rect 466637 680504 495818 680506
rect 466637 680448 466642 680504
rect 466698 680448 495818 680504
rect 466637 680446 495818 680448
rect 466637 680443 466703 680446
rect 463693 680370 463759 680373
rect 458222 680368 463759 680370
rect 458222 680312 463698 680368
rect 463754 680312 463759 680368
rect 458222 680310 463759 680312
rect 439497 680307 439563 680310
rect 451365 680307 451431 680310
rect 457161 680307 457227 680310
rect 463693 680307 463759 680310
rect 466545 680370 466611 680373
rect 481173 680370 481239 680373
rect 466545 680368 481239 680370
rect 466545 680312 466550 680368
rect 466606 680312 481178 680368
rect 481234 680312 481239 680368
rect 466545 680310 481239 680312
rect 466545 680307 466611 680310
rect 481173 680307 481239 680310
rect 485773 680370 485839 680373
rect 495433 680370 495499 680373
rect 485773 680368 495499 680370
rect 485773 680312 485778 680368
rect 485834 680312 495438 680368
rect 495494 680312 495499 680368
rect 485773 680310 495499 680312
rect 495758 680370 495818 680446
rect 505142 680446 534090 680506
rect 505142 680370 505202 680446
rect 495758 680310 505202 680370
rect 505921 680370 505987 680373
rect 515397 680370 515463 680373
rect 505921 680368 515463 680370
rect 505921 680312 505926 680368
rect 505982 680312 515402 680368
rect 515458 680312 515463 680368
rect 505921 680310 515463 680312
rect 485773 680307 485839 680310
rect 495433 680307 495499 680310
rect 505921 680307 505987 680310
rect 515397 680307 515463 680310
rect 524413 680370 524479 680373
rect 534349 680370 534415 680373
rect 524413 680368 534415 680370
rect 524413 680312 524418 680368
rect 524474 680312 534354 680368
rect 534410 680312 534415 680368
rect 524413 680310 534415 680312
rect 535502 680370 535562 680718
rect 557582 680718 559788 680778
rect 543825 680642 543891 680645
rect 550582 680642 550588 680644
rect 543825 680640 550588 680642
rect 543825 680584 543830 680640
rect 543886 680584 550588 680640
rect 543825 680582 550588 680584
rect 543825 680579 543891 680582
rect 550582 680580 550588 680582
rect 550652 680580 550658 680644
rect 557441 680642 557507 680645
rect 553902 680640 557507 680642
rect 553902 680584 557446 680640
rect 557502 680584 557507 680640
rect 553902 680582 557507 680584
rect 543825 680370 543891 680373
rect 535502 680368 543891 680370
rect 535502 680312 543830 680368
rect 543886 680312 543891 680368
rect 535502 680310 543891 680312
rect 524413 680307 524479 680310
rect 534349 680307 534415 680310
rect 543825 680307 543891 680310
rect 544009 680370 544075 680373
rect 553902 680370 553962 680582
rect 557441 680579 557507 680582
rect 554773 680506 554839 680509
rect 557582 680506 557642 680718
rect 559782 680716 559788 680718
rect 559852 680716 559858 680780
rect 559373 680642 559439 680645
rect 561990 680642 561996 680644
rect 559373 680640 561996 680642
rect 559373 680584 559378 680640
rect 559434 680584 561996 680640
rect 559373 680582 561996 680584
rect 559373 680579 559439 680582
rect 561990 680580 561996 680582
rect 562060 680580 562066 680644
rect 559046 680506 559052 680508
rect 554773 680504 557642 680506
rect 554773 680448 554778 680504
rect 554834 680448 557642 680504
rect 554773 680446 557642 680448
rect 558318 680446 559052 680506
rect 554773 680443 554839 680446
rect 544009 680368 553962 680370
rect 544009 680312 544014 680368
rect 544070 680312 553962 680368
rect 544009 680310 553962 680312
rect 554865 680370 554931 680373
rect 558318 680370 558378 680446
rect 559046 680444 559052 680446
rect 559116 680444 559122 680508
rect 559189 680506 559255 680509
rect 561581 680508 561647 680509
rect 561254 680506 561260 680508
rect 559189 680504 561260 680506
rect 559189 680448 559194 680504
rect 559250 680448 561260 680504
rect 559189 680446 561260 680448
rect 559189 680443 559255 680446
rect 561254 680444 561260 680446
rect 561324 680444 561330 680508
rect 561581 680506 561628 680508
rect 561536 680504 561628 680506
rect 561536 680448 561586 680504
rect 561536 680446 561628 680448
rect 561581 680444 561628 680446
rect 561692 680444 561698 680508
rect 561765 680506 561831 680509
rect 563094 680506 563100 680508
rect 561765 680504 563100 680506
rect 561765 680448 561770 680504
rect 561826 680448 563100 680504
rect 561765 680446 563100 680448
rect 561581 680443 561647 680444
rect 561765 680443 561831 680446
rect 563094 680444 563100 680446
rect 563164 680444 563170 680508
rect 563237 680506 563303 680509
rect 564566 680506 564572 680508
rect 563237 680504 564572 680506
rect 563237 680448 563242 680504
rect 563298 680448 564572 680504
rect 563237 680446 564572 680448
rect 563237 680443 563303 680446
rect 564566 680444 564572 680446
rect 564636 680444 564642 680508
rect 564709 680506 564775 680509
rect 567142 680506 567148 680508
rect 564709 680504 567148 680506
rect 564709 680448 564714 680504
rect 564770 680448 567148 680504
rect 564709 680446 567148 680448
rect 564709 680443 564775 680446
rect 567142 680444 567148 680446
rect 567212 680444 567218 680508
rect 554865 680368 558378 680370
rect 554865 680312 554870 680368
rect 554926 680312 558378 680368
rect 554865 680310 558378 680312
rect 558545 680370 558611 680373
rect 560753 680372 560819 680373
rect 559414 680370 559420 680372
rect 558545 680368 559420 680370
rect 558545 680312 558550 680368
rect 558606 680312 559420 680368
rect 558545 680310 559420 680312
rect 544009 680307 544075 680310
rect 554865 680307 554931 680310
rect 558545 680307 558611 680310
rect 559414 680308 559420 680310
rect 559484 680308 559490 680372
rect 560702 680370 560708 680372
rect 560662 680310 560708 680370
rect 560772 680368 560819 680372
rect 560814 680312 560819 680368
rect 560702 680308 560708 680310
rect 560772 680308 560819 680312
rect 561070 680308 561076 680372
rect 561140 680370 561146 680372
rect 561213 680370 561279 680373
rect 561140 680368 561279 680370
rect 561140 680312 561218 680368
rect 561274 680312 561279 680368
rect 561140 680310 561279 680312
rect 561140 680308 561146 680310
rect 560753 680307 560819 680308
rect 561213 680307 561279 680310
rect 561857 680370 561923 680373
rect 562358 680370 562364 680372
rect 561857 680368 562364 680370
rect 561857 680312 561862 680368
rect 561918 680312 562364 680368
rect 561857 680310 562364 680312
rect 561857 680307 561923 680310
rect 562358 680308 562364 680310
rect 562428 680308 562434 680372
rect 562501 680370 562567 680373
rect 566365 680372 566431 680373
rect 563646 680370 563652 680372
rect 562501 680368 563652 680370
rect 562501 680312 562506 680368
rect 562562 680312 563652 680368
rect 562501 680310 563652 680312
rect 562501 680307 562567 680310
rect 563646 680308 563652 680310
rect 563716 680308 563722 680372
rect 566365 680370 566412 680372
rect 566320 680368 566412 680370
rect 566320 680312 566370 680368
rect 566320 680310 566412 680312
rect 566365 680308 566412 680310
rect 566476 680308 566482 680372
rect 566365 680307 566431 680308
rect 580165 674658 580231 674661
rect 583520 674658 584960 674748
rect 580165 674656 584960 674658
rect 580165 674600 580170 674656
rect 580226 674600 584960 674656
rect 580165 674598 584960 674600
rect 580165 674595 580231 674598
rect 583520 674508 584960 674598
rect 1166 669493 1226 669596
rect 1117 669488 1226 669493
rect 1117 669432 1122 669488
rect 1178 669432 1226 669488
rect 1117 669430 1226 669432
rect 1117 669427 1183 669430
rect -960 667844 480 668084
rect 572713 667450 572779 667453
rect 570860 667448 572779 667450
rect 570860 667392 572718 667448
rect 572774 667392 572779 667448
rect 570860 667390 572779 667392
rect 572713 667387 572779 667390
rect 583520 662676 584960 662916
rect -960 653428 480 653668
rect 583520 650980 584960 651220
rect 1166 646781 1226 646884
rect 1166 646776 1275 646781
rect 1166 646720 1214 646776
rect 1270 646720 1275 646776
rect 1166 646718 1275 646720
rect 1209 646715 1275 646718
rect 572713 640250 572779 640253
rect 570860 640248 572779 640250
rect 570860 640192 572718 640248
rect 572774 640192 572779 640248
rect 570860 640190 572779 640192
rect 572713 640187 572779 640190
rect 583520 639284 584960 639524
rect -960 639012 480 639252
rect 579705 627738 579771 627741
rect 583520 627738 584960 627828
rect 579705 627736 584960 627738
rect 579705 627680 579710 627736
rect 579766 627680 584960 627736
rect 579705 627678 584960 627680
rect 579705 627675 579771 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect -960 624822 674 624882
rect -960 624732 480 624822
rect 13 624610 79 624613
rect 614 624610 674 624822
rect 13 624608 674 624610
rect 13 624552 18 624608
rect 74 624552 674 624608
rect 13 624550 674 624552
rect 13 624547 79 624550
rect 1534 623797 1594 624308
rect 1534 623792 1643 623797
rect 1534 623736 1582 623792
rect 1638 623736 1643 623792
rect 1534 623734 1643 623736
rect 1577 623731 1643 623734
rect 583520 615756 584960 615996
rect 570278 612509 570338 613020
rect 570278 612504 570387 612509
rect 570278 612448 570326 612504
rect 570382 612448 570387 612504
rect 570278 612446 570387 612448
rect 570321 612443 570387 612446
rect -960 610316 480 610556
rect 583520 604060 584960 604300
rect 1534 601085 1594 601596
rect 1534 601080 1643 601085
rect 1534 601024 1582 601080
rect 1638 601024 1643 601080
rect 1534 601022 1643 601024
rect 1577 601019 1643 601022
rect -960 595900 480 596140
rect 583520 592364 584960 592604
rect 572713 585850 572779 585853
rect 570860 585848 572779 585850
rect 570860 585792 572718 585848
rect 572774 585792 572779 585848
rect 570860 585790 572779 585792
rect 572713 585787 572779 585790
rect -960 581620 480 581860
rect 580257 580818 580323 580821
rect 583520 580818 584960 580908
rect 580257 580816 584960 580818
rect 580257 580760 580262 580816
rect 580318 580760 584960 580816
rect 580257 580758 584960 580760
rect 580257 580755 580323 580758
rect 583520 580668 584960 580758
rect 1534 578373 1594 578884
rect 1534 578368 1643 578373
rect 1534 578312 1582 578368
rect 1638 578312 1643 578368
rect 1534 578310 1643 578312
rect 1577 578307 1643 578310
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 1301 567354 1367 567357
rect -960 567352 1367 567354
rect -960 567296 1306 567352
rect 1362 567296 1367 567352
rect -960 567294 1367 567296
rect -960 567204 480 567294
rect 1301 567291 1367 567294
rect 572713 558650 572779 558653
rect 570860 558648 572779 558650
rect 570860 558592 572718 558648
rect 572774 558592 572779 558648
rect 570860 558590 572779 558592
rect 572713 558587 572779 558590
rect 583520 557140 584960 557380
rect 1534 556205 1594 556308
rect 1534 556200 1643 556205
rect 1534 556144 1582 556200
rect 1638 556144 1643 556200
rect 1534 556142 1643 556144
rect 1577 556139 1643 556142
rect -960 552924 480 553164
rect 583520 545444 584960 545684
rect -960 538508 480 538748
rect 580165 533898 580231 533901
rect 583520 533898 584960 533988
rect 580165 533896 584960 533898
rect 580165 533840 580170 533896
rect 580226 533840 584960 533896
rect 580165 533838 584960 533840
rect 580165 533835 580231 533838
rect 583520 533748 584960 533838
rect 1534 533085 1594 533596
rect 1534 533080 1643 533085
rect 1534 533024 1582 533080
rect 1638 533024 1643 533080
rect 1534 533022 1643 533024
rect 1577 533019 1643 533022
rect 570278 530909 570338 531420
rect 570278 530904 570387 530909
rect 570278 530848 570326 530904
rect 570382 530848 570387 530904
rect 570278 530846 570387 530848
rect 570321 530843 570387 530846
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 1534 510645 1594 510884
rect 1485 510640 1594 510645
rect 1485 510584 1490 510640
rect 1546 510584 1594 510640
rect 1485 510582 1594 510584
rect 1485 510579 1551 510582
rect 583520 510220 584960 510460
rect -960 509962 480 510052
rect 1577 509962 1643 509965
rect -960 509960 1643 509962
rect -960 509904 1582 509960
rect 1638 509904 1643 509960
rect -960 509902 1643 509904
rect -960 509812 480 509902
rect 1577 509899 1643 509902
rect 570278 503709 570338 504220
rect 570278 503704 570387 503709
rect 570278 503648 570326 503704
rect 570382 503648 570387 503704
rect 570278 503646 570387 503648
rect 570321 503643 570387 503646
rect 583520 498524 584960 498764
rect -960 495396 480 495636
rect 1534 487797 1594 488308
rect 1534 487792 1643 487797
rect 1534 487736 1582 487792
rect 1638 487736 1643 487792
rect 1534 487734 1643 487736
rect 1577 487731 1643 487734
rect 579797 486842 579863 486845
rect 583520 486842 584960 486932
rect 579797 486840 584960 486842
rect 579797 486784 579802 486840
rect 579858 486784 584960 486840
rect 579797 486782 584960 486784
rect 579797 486779 579863 486782
rect 583520 486692 584960 486782
rect -960 480980 480 481220
rect 570278 476509 570338 477020
rect 570278 476504 570387 476509
rect 570278 476448 570326 476504
rect 570382 476448 570387 476504
rect 570278 476446 570387 476448
rect 570321 476443 570387 476446
rect 583520 474996 584960 475236
rect -960 466700 480 466940
rect 1350 465085 1410 465596
rect 1350 465080 1459 465085
rect 1350 465024 1398 465080
rect 1454 465024 1459 465080
rect 1350 465022 1459 465024
rect 1393 465019 1459 465022
rect 583520 463300 584960 463540
rect -960 452434 480 452524
rect 1393 452434 1459 452437
rect -960 452432 1459 452434
rect -960 452376 1398 452432
rect 1454 452376 1459 452432
rect -960 452374 1459 452376
rect -960 452284 480 452374
rect 1393 452371 1459 452374
rect 583520 451604 584960 451844
rect 570278 449309 570338 449820
rect 570278 449304 570387 449309
rect 570278 449248 570326 449304
rect 570382 449248 570387 449304
rect 570278 449246 570387 449248
rect 570321 449243 570387 449246
rect 749 442370 815 442373
rect 1166 442370 1226 442884
rect 749 442368 1226 442370
rect 749 442312 754 442368
rect 810 442312 1226 442368
rect 749 442310 1226 442312
rect 749 442307 815 442310
rect 580165 439922 580231 439925
rect 583520 439922 584960 440012
rect 580165 439920 584960 439922
rect 580165 439864 580170 439920
rect 580226 439864 584960 439920
rect 580165 439862 584960 439864
rect 580165 439859 580231 439862
rect 583520 439772 584960 439862
rect -960 437868 480 438108
rect 583520 428076 584960 428316
rect -960 423588 480 423828
rect 572713 422650 572779 422653
rect 570860 422648 572779 422650
rect 570860 422592 572718 422648
rect 572774 422592 572779 422648
rect 570860 422590 572779 422592
rect 572713 422587 572779 422590
rect 1350 419797 1410 420308
rect 1350 419792 1459 419797
rect 1350 419736 1398 419792
rect 1454 419736 1459 419792
rect 1350 419734 1459 419736
rect 1393 419731 1459 419734
rect 583520 416380 584960 416620
rect -960 409172 480 409412
rect 583520 404684 584960 404924
rect 933 397354 999 397357
rect 1166 397354 1226 397596
rect 933 397352 1226 397354
rect 933 397296 938 397352
rect 994 397296 1226 397352
rect 933 397294 1226 397296
rect 933 397291 999 397294
rect -960 395042 480 395132
rect 1393 395042 1459 395045
rect -960 395040 1459 395042
rect -960 394984 1398 395040
rect 1454 394984 1459 395040
rect -960 394982 1459 394984
rect -960 394892 480 394982
rect 1393 394979 1459 394982
rect 570278 394909 570338 395420
rect 570278 394904 570387 394909
rect 570278 394848 570326 394904
rect 570382 394848 570387 394904
rect 570278 394846 570387 394848
rect 570321 394843 570387 394846
rect 580165 393002 580231 393005
rect 583520 393002 584960 393092
rect 580165 393000 584960 393002
rect 580165 392944 580170 393000
rect 580226 392944 584960 393000
rect 580165 392942 584960 392944
rect 580165 392939 580231 392942
rect 583520 392852 584960 392942
rect 583520 381156 584960 381396
rect -960 380476 480 380716
rect 565 374370 631 374373
rect 1166 374370 1226 374884
rect 565 374368 1226 374370
rect 565 374312 570 374368
rect 626 374312 1226 374368
rect 565 374310 1226 374312
rect 565 374307 631 374310
rect 583520 369460 584960 369700
rect 570278 367709 570338 368220
rect 570278 367704 570387 367709
rect 570278 367648 570326 367704
rect 570382 367648 570387 367704
rect 570278 367646 570387 367648
rect 570321 367643 570387 367646
rect -960 366060 480 366300
rect 583520 357764 584960 358004
rect 105 352202 171 352205
rect 1166 352202 1226 352308
rect 105 352200 1226 352202
rect 105 352144 110 352200
rect 166 352144 1226 352200
rect 105 352142 1226 352144
rect 105 352139 171 352142
rect -960 351780 480 352020
rect 580165 346082 580231 346085
rect 583520 346082 584960 346172
rect 580165 346080 584960 346082
rect 580165 346024 580170 346080
rect 580226 346024 584960 346080
rect 580165 346022 584960 346024
rect 580165 346019 580231 346022
rect 583520 345932 584960 346022
rect 572713 341050 572779 341053
rect 570860 341048 572779 341050
rect 570860 340992 572718 341048
rect 572774 340992 572779 341048
rect 570860 340990 572779 340992
rect 572713 340987 572779 340990
rect 3141 339692 3207 339693
rect 3136 339690 3142 339692
rect 3050 339630 3142 339690
rect 3136 339628 3142 339630
rect 3206 339628 3212 339692
rect 3141 339627 3207 339628
rect -960 337514 480 337604
rect 1301 337514 1367 337517
rect -960 337512 1367 337514
rect -960 337456 1306 337512
rect 1362 337456 1367 337512
rect -960 337454 1367 337456
rect -960 337364 480 337454
rect 1301 337451 1367 337454
rect 583520 334236 584960 334476
rect 657 329082 723 329085
rect 1166 329082 1226 329596
rect 657 329080 1226 329082
rect 657 329024 662 329080
rect 718 329024 1226 329080
rect 657 329022 1226 329024
rect 657 329019 723 329022
rect -960 322948 480 323188
rect 583520 322540 584960 322780
rect 3141 321060 3207 321061
rect 3136 321058 3142 321060
rect 3050 320998 3142 321058
rect 3136 320996 3142 320998
rect 3206 320996 3212 321060
rect 3141 320995 3207 320996
rect 572713 313850 572779 313853
rect 570860 313848 572779 313850
rect 570860 313792 572718 313848
rect 572774 313792 572779 313848
rect 570860 313790 572779 313792
rect 572713 313787 572779 313790
rect 583520 310708 584960 310948
rect -960 308668 480 308908
rect 1350 306373 1410 306884
rect 1350 306368 1459 306373
rect 1350 306312 1398 306368
rect 1454 306312 1459 306368
rect 1350 306310 1459 306312
rect 1393 306307 1459 306310
rect 580165 299162 580231 299165
rect 583520 299162 584960 299252
rect 580165 299160 584960 299162
rect 580165 299104 580170 299160
rect 580226 299104 584960 299160
rect 580165 299102 584960 299104
rect 580165 299099 580231 299102
rect 583520 299012 584960 299102
rect -960 294402 480 294492
rect 1393 294402 1459 294405
rect -960 294400 1459 294402
rect -960 294344 1398 294400
rect 1454 294344 1459 294400
rect -960 294342 1459 294344
rect -960 294252 480 294342
rect 1393 294339 1459 294342
rect 583520 287316 584960 287556
rect 570462 286109 570522 286620
rect 570413 286104 570522 286109
rect 570413 286048 570418 286104
rect 570474 286048 570522 286104
rect 570413 286046 570522 286048
rect 570413 286043 570479 286046
rect 570505 284612 570571 284613
rect 570454 284548 570460 284612
rect 570524 284610 570571 284612
rect 570524 284608 570616 284610
rect 570566 284552 570616 284608
rect 570524 284550 570616 284552
rect 570524 284548 570571 284550
rect 570505 284547 570571 284548
rect 1350 283797 1410 284308
rect 1350 283792 1459 283797
rect 1350 283736 1398 283792
rect 1454 283736 1459 283792
rect 1350 283734 1459 283736
rect 1393 283731 1459 283734
rect -960 279972 480 280212
rect 583520 275620 584960 275860
rect -960 265556 480 265796
rect 583520 263788 584960 264028
rect 1350 261085 1410 261596
rect 1350 261080 1459 261085
rect 1350 261024 1398 261080
rect 1454 261024 1459 261080
rect 1350 261022 1459 261024
rect 1393 261019 1459 261022
rect 569217 260132 569283 260133
rect 569212 260068 569218 260132
rect 569282 260130 569288 260132
rect 569282 260070 569374 260130
rect 569282 260068 569288 260070
rect 569217 260067 569283 260068
rect 574737 259450 574803 259453
rect 570860 259448 574803 259450
rect 570860 259392 574742 259448
rect 574798 259392 574803 259448
rect 570860 259390 574803 259392
rect 574737 259387 574803 259390
rect 580165 252242 580231 252245
rect 583520 252242 584960 252332
rect 580165 252240 584960 252242
rect 580165 252184 580170 252240
rect 580226 252184 584960 252240
rect 580165 252182 584960 252184
rect 580165 252179 580231 252182
rect 583520 252092 584960 252182
rect -960 251290 480 251380
rect 1393 251290 1459 251293
rect -960 251288 1459 251290
rect -960 251232 1398 251288
rect 1454 251232 1459 251288
rect -960 251230 1459 251232
rect -960 251140 480 251230
rect 1393 251227 1459 251230
rect 568389 248436 568455 248437
rect 568384 248434 568390 248436
rect 568298 248374 568390 248434
rect 568384 248372 568390 248374
rect 568454 248372 568460 248436
rect 568389 248371 568455 248372
rect 583520 240396 584960 240636
rect 1350 238373 1410 238884
rect 1301 238368 1410 238373
rect 1301 238312 1306 238368
rect 1362 238312 1410 238368
rect 1301 238310 1410 238312
rect 1301 238307 1367 238310
rect -960 236860 480 237100
rect 574829 232250 574895 232253
rect 570860 232248 574895 232250
rect 570860 232192 574834 232248
rect 574890 232192 574895 232248
rect 570860 232190 574895 232192
rect 574829 232187 574895 232190
rect 583520 228700 584960 228940
rect -960 222444 480 222684
rect 568849 222324 568915 222325
rect 568844 222260 568850 222324
rect 568914 222322 568920 222324
rect 568914 222262 569006 222322
rect 568914 222260 568920 222262
rect 568849 222259 568915 222260
rect 1393 221508 1459 221509
rect 1342 221506 1348 221508
rect 1302 221446 1348 221506
rect 1412 221504 1459 221508
rect 1454 221448 1459 221504
rect 1342 221444 1348 221446
rect 1412 221444 1459 221448
rect 1393 221443 1459 221444
rect 583520 216868 584960 217108
rect 13 215794 79 215797
rect 1166 215794 1226 216308
rect 13 215792 1226 215794
rect 13 215736 18 215792
rect 74 215736 1226 215792
rect 13 215734 1226 215736
rect 13 215731 79 215734
rect 1301 214572 1367 214573
rect 1301 214570 1348 214572
rect 1256 214568 1348 214570
rect 1256 214512 1306 214568
rect 1256 214510 1348 214512
rect 1301 214508 1348 214510
rect 1412 214508 1418 214572
rect 1301 214507 1367 214508
rect -960 208178 480 208268
rect 565 208178 631 208181
rect -960 208176 631 208178
rect -960 208120 570 208176
rect 626 208120 631 208176
rect -960 208118 631 208120
rect -960 208028 480 208118
rect 565 208115 631 208118
rect 580165 205322 580231 205325
rect 583520 205322 584960 205412
rect 580165 205320 584960 205322
rect 580165 205264 580170 205320
rect 580226 205264 584960 205320
rect 580165 205262 584960 205264
rect 580165 205259 580231 205262
rect 583520 205172 584960 205262
rect 574921 205050 574987 205053
rect 570860 205048 574987 205050
rect 570860 204992 574926 205048
rect 574982 204992 574987 205048
rect 570860 204990 574987 204992
rect 574921 204987 574987 204990
rect 1393 198250 1459 198253
rect 1526 198250 1532 198252
rect 1393 198248 1532 198250
rect 1393 198192 1398 198248
rect 1454 198192 1532 198248
rect 1393 198190 1532 198192
rect 1393 198187 1459 198190
rect 1526 198188 1532 198190
rect 1596 198188 1602 198252
rect -960 193748 480 193988
rect 568573 193628 568639 193629
rect 570321 193628 570387 193629
rect 1350 193085 1410 193596
rect 568568 193564 568574 193628
rect 568638 193626 568644 193628
rect 568638 193566 568730 193626
rect 568638 193564 568644 193566
rect 570270 193564 570276 193628
rect 570340 193626 570387 193628
rect 570340 193624 570432 193626
rect 570382 193568 570432 193624
rect 570340 193566 570432 193568
rect 570340 193564 570387 193566
rect 568573 193563 568639 193564
rect 570321 193563 570387 193564
rect 568297 193492 568363 193493
rect 568292 193428 568298 193492
rect 568362 193490 568368 193492
rect 568362 193430 568454 193490
rect 568362 193428 568368 193430
rect 570454 193428 570460 193492
rect 570524 193490 570530 193492
rect 570638 193490 570644 193492
rect 570524 193430 570644 193490
rect 570524 193428 570530 193430
rect 570638 193428 570644 193430
rect 570708 193428 570714 193492
rect 583520 193476 584960 193716
rect 568297 193427 568363 193428
rect 1301 193080 1410 193085
rect 1301 193024 1306 193080
rect 1362 193024 1410 193080
rect 1301 193022 1410 193024
rect 1301 193019 1367 193022
rect 2865 185332 2931 185333
rect 2860 185268 2866 185332
rect 2930 185330 2936 185332
rect 2930 185270 3022 185330
rect 2930 185268 2936 185270
rect 2865 185267 2931 185268
rect 583520 181780 584960 182020
rect -960 179332 480 179572
rect 569217 178532 569283 178533
rect 569166 178530 569172 178532
rect 569126 178470 569172 178530
rect 569236 178528 569283 178532
rect 569278 178472 569283 178528
rect 569166 178468 569172 178470
rect 569236 178468 569283 178472
rect 569217 178467 569283 178468
rect 575013 177850 575079 177853
rect 570860 177848 575079 177850
rect 570860 177792 575018 177848
rect 575074 177792 575079 177848
rect 570860 177790 575079 177792
rect 575013 177787 575079 177790
rect 568481 174588 568547 174589
rect 568476 174524 568482 174588
rect 568546 174586 568552 174588
rect 568546 174526 568638 174586
rect 568546 174524 568552 174526
rect 568481 174523 568547 174524
rect 1485 173092 1551 173093
rect 1485 173090 1532 173092
rect 1440 173088 1532 173090
rect 1440 173032 1490 173088
rect 1440 173030 1532 173032
rect 1485 173028 1532 173030
rect 1596 173028 1602 173092
rect 1485 173027 1551 173028
rect 1534 170373 1594 170884
rect 1485 170368 1594 170373
rect 1485 170312 1490 170368
rect 1546 170312 1594 170368
rect 1485 170310 1594 170312
rect 1485 170307 1551 170310
rect 583520 169948 584960 170188
rect 1393 167650 1459 167653
rect 1526 167650 1532 167652
rect 1393 167648 1532 167650
rect 1393 167592 1398 167648
rect 1454 167592 1532 167648
rect 1393 167590 1532 167592
rect 1393 167587 1459 167590
rect 1526 167588 1532 167590
rect 1596 167588 1602 167652
rect -960 165066 480 165156
rect 1393 165066 1459 165069
rect -960 165064 1459 165066
rect -960 165008 1398 165064
rect 1454 165008 1459 165064
rect -960 165006 1459 165008
rect -960 164916 480 165006
rect 1393 165003 1459 165006
rect 580165 158402 580231 158405
rect 583520 158402 584960 158492
rect 580165 158400 584960 158402
rect 580165 158344 580170 158400
rect 580226 158344 584960 158400
rect 580165 158342 584960 158344
rect 580165 158339 580231 158342
rect 583520 158252 584960 158342
rect -960 150636 480 150876
rect 574737 150650 574803 150653
rect 570860 150648 574803 150650
rect 570860 150592 574742 150648
rect 574798 150592 574803 150648
rect 570860 150590 574803 150592
rect 574737 150587 574803 150590
rect 1577 148746 1643 148749
rect 1534 148744 1643 148746
rect 1534 148688 1582 148744
rect 1638 148688 1643 148744
rect 1534 148683 1643 148688
rect 1534 148308 1594 148683
rect 1577 146980 1643 146981
rect 1526 146978 1532 146980
rect 1486 146918 1532 146978
rect 1596 146976 1643 146980
rect 1638 146920 1643 146976
rect 1526 146916 1532 146918
rect 1596 146916 1643 146920
rect 1577 146915 1643 146916
rect 583520 146556 584960 146796
rect 1485 138684 1551 138685
rect 1485 138680 1532 138684
rect 1596 138682 1602 138684
rect 1485 138624 1490 138680
rect 1485 138620 1532 138624
rect 1596 138622 1642 138682
rect 1596 138620 1602 138622
rect 1485 138619 1551 138620
rect -960 136220 480 136460
rect 583520 134724 584960 134964
rect 1577 126442 1643 126445
rect 1534 126440 1643 126442
rect 1534 126384 1582 126440
rect 1638 126384 1643 126440
rect 1534 126379 1643 126384
rect 1534 125596 1594 126379
rect 572713 123450 572779 123453
rect 570860 123448 572779 123450
rect 570860 123392 572718 123448
rect 572774 123392 572779 123448
rect 570860 123390 572779 123392
rect 572713 123387 572779 123390
rect 583520 123028 584960 123268
rect -960 122090 480 122180
rect 1301 122090 1367 122093
rect -960 122088 1367 122090
rect -960 122032 1306 122088
rect 1362 122032 1367 122088
rect -960 122030 1367 122032
rect -960 121940 480 122030
rect 1301 122027 1367 122030
rect 580165 111482 580231 111485
rect 583520 111482 584960 111572
rect 580165 111480 584960 111482
rect 580165 111424 580170 111480
rect 580226 111424 584960 111480
rect 580165 111422 584960 111424
rect 580165 111419 580231 111422
rect 583520 111332 584960 111422
rect 1209 108218 1275 108221
rect 1342 108218 1348 108220
rect 1209 108216 1348 108218
rect 1209 108160 1214 108216
rect 1270 108160 1348 108216
rect 1209 108158 1348 108160
rect 1209 108155 1275 108158
rect 1342 108156 1348 108158
rect 1412 108156 1418 108220
rect -960 107524 480 107764
rect 1209 107130 1275 107133
rect 1526 107130 1532 107132
rect 1209 107128 1532 107130
rect 1209 107072 1214 107128
rect 1270 107072 1532 107128
rect 1209 107070 1532 107072
rect 1209 107067 1275 107070
rect 1526 107068 1532 107070
rect 1596 107068 1602 107132
rect 473 103458 539 103461
rect 473 103456 1042 103458
rect 473 103400 478 103456
rect 534 103400 1042 103456
rect 473 103398 1042 103400
rect 473 103395 539 103398
rect 982 102884 1042 103398
rect 1301 99650 1367 99653
rect 1526 99650 1532 99652
rect 1301 99648 1532 99650
rect 1301 99592 1306 99648
rect 1362 99592 1532 99648
rect 1301 99590 1532 99592
rect 1301 99587 1367 99590
rect 1526 99588 1532 99590
rect 1596 99588 1602 99652
rect 583520 99636 584960 99876
rect 570321 99380 570387 99381
rect 570270 99316 570276 99380
rect 570340 99378 570387 99380
rect 570340 99376 570432 99378
rect 570382 99320 570432 99376
rect 570340 99318 570432 99320
rect 570340 99316 570387 99318
rect 570321 99315 570387 99316
rect 572713 96250 572779 96253
rect 570860 96248 572779 96250
rect 570860 96192 572718 96248
rect 572774 96192 572779 96248
rect 570860 96190 572779 96192
rect 572713 96187 572779 96190
rect 3509 96116 3575 96117
rect 3504 96114 3510 96116
rect 3418 96054 3510 96114
rect 3504 96052 3510 96054
rect 3574 96052 3580 96116
rect 3509 96051 3575 96052
rect -960 93108 480 93348
rect 570321 90130 570387 90133
rect 570454 90130 570460 90132
rect 570321 90128 570460 90130
rect 570321 90072 570326 90128
rect 570382 90072 570460 90128
rect 570321 90070 570460 90072
rect 570321 90067 570387 90070
rect 570454 90068 570460 90070
rect 570524 90068 570530 90132
rect 583520 87804 584960 88044
rect 1209 80882 1275 80885
rect 1166 80880 1275 80882
rect 1166 80824 1214 80880
rect 1270 80824 1275 80880
rect 1166 80819 1275 80824
rect 1166 80308 1226 80819
rect -960 78978 480 79068
rect 565 78978 631 78981
rect -960 78976 631 78978
rect -960 78920 570 78976
rect 626 78920 631 78976
rect -960 78918 631 78920
rect -960 78828 480 78918
rect 565 78915 631 78918
rect 583520 76108 584960 76348
rect 574737 69050 574803 69053
rect 570860 69048 574803 69050
rect 570860 68992 574742 69048
rect 574798 68992 574803 69048
rect 570860 68990 574803 68992
rect 574737 68987 574803 68990
rect -960 64412 480 64652
rect 580165 64562 580231 64565
rect 583520 64562 584960 64652
rect 580165 64560 584960 64562
rect 580165 64504 580170 64560
rect 580226 64504 584960 64560
rect 580165 64502 584960 64504
rect 580165 64499 580231 64502
rect 583520 64412 584960 64502
rect 1301 58034 1367 58037
rect 1301 58032 1410 58034
rect 1301 57976 1306 58032
rect 1362 57976 1410 58032
rect 1301 57971 1410 57976
rect 1350 57596 1410 57971
rect 583520 52716 584960 52956
rect -960 49996 480 50236
rect 1301 45930 1367 45933
rect 1526 45930 1532 45932
rect 1301 45928 1532 45930
rect 1301 45872 1306 45928
rect 1362 45872 1532 45928
rect 1301 45870 1532 45872
rect 1301 45867 1367 45870
rect 1526 45868 1532 45870
rect 1596 45868 1602 45932
rect 574737 41850 574803 41853
rect 570860 41848 574803 41850
rect 570860 41792 574742 41848
rect 574798 41792 574803 41848
rect 570860 41790 574803 41792
rect 574737 41787 574803 41790
rect 583520 40884 584960 41124
rect 3785 40356 3851 40357
rect 3734 40292 3740 40356
rect 3804 40354 3851 40356
rect 3804 40352 3896 40354
rect 3846 40296 3896 40352
rect 3804 40294 3896 40296
rect 3804 40292 3851 40294
rect 3785 40291 3851 40292
rect 13 36138 79 36141
rect 13 36136 674 36138
rect 13 36080 18 36136
rect 74 36080 674 36136
rect 13 36078 674 36080
rect 13 36075 79 36078
rect -960 35866 480 35956
rect 614 35866 674 36078
rect -960 35806 674 35866
rect -960 35716 480 35806
rect 1393 35458 1459 35461
rect 1350 35456 1459 35458
rect 1350 35400 1398 35456
rect 1454 35400 1459 35456
rect 1350 35395 1459 35400
rect 1350 34884 1410 35395
rect 570321 34916 570387 34917
rect 570270 34852 570276 34916
rect 570340 34914 570387 34916
rect 570340 34912 570432 34914
rect 570382 34856 570432 34912
rect 570340 34854 570432 34856
rect 570340 34852 570387 34854
rect 570321 34851 570387 34852
rect 1209 33282 1275 33285
rect 1526 33282 1532 33284
rect 1209 33280 1532 33282
rect 1209 33224 1214 33280
rect 1270 33224 1532 33280
rect 1209 33222 1532 33224
rect 1209 33219 1275 33222
rect 1526 33220 1532 33222
rect 1596 33220 1602 33284
rect 657 32332 723 32333
rect 606 32268 612 32332
rect 676 32330 723 32332
rect 676 32328 768 32330
rect 718 32272 768 32328
rect 676 32270 768 32272
rect 676 32268 723 32270
rect 657 32267 723 32268
rect 1485 30292 1551 30293
rect 1485 30288 1532 30292
rect 1596 30290 1602 30292
rect 1485 30232 1490 30288
rect 1485 30228 1532 30232
rect 1596 30230 1642 30290
rect 1596 30228 1602 30230
rect 1485 30227 1551 30228
rect 1393 29748 1459 29749
rect 1342 29746 1348 29748
rect 1302 29686 1348 29746
rect 1412 29744 1459 29748
rect 1454 29688 1459 29744
rect 1342 29684 1348 29686
rect 1412 29684 1459 29688
rect 1393 29683 1459 29684
rect 583520 29188 584960 29428
rect 1209 27026 1275 27029
rect 1526 27026 1532 27028
rect 1209 27024 1532 27026
rect 1209 26968 1214 27024
rect 1270 26968 1532 27024
rect 1209 26966 1532 26968
rect 1209 26963 1275 26966
rect 1526 26964 1532 26966
rect 1596 26964 1602 27028
rect 1209 26890 1275 26893
rect 1342 26890 1348 26892
rect 1209 26888 1348 26890
rect 1209 26832 1214 26888
rect 1270 26832 1348 26888
rect 1209 26830 1348 26832
rect 1209 26827 1275 26830
rect 1342 26828 1348 26830
rect 1412 26828 1418 26892
rect 974 25740 980 25804
rect 1044 25802 1050 25804
rect 1485 25802 1551 25805
rect 1044 25800 1551 25802
rect 1044 25744 1490 25800
rect 1546 25744 1551 25800
rect 1044 25742 1551 25744
rect 1044 25740 1050 25742
rect 1485 25739 1551 25742
rect -960 21300 480 21540
rect 1393 20090 1459 20093
rect 1526 20090 1532 20092
rect 1393 20088 1532 20090
rect 1393 20032 1398 20088
rect 1454 20032 1532 20088
rect 1393 20030 1532 20032
rect 1393 20027 1459 20030
rect 1526 20028 1532 20030
rect 1596 20028 1602 20092
rect 749 19954 815 19957
rect 1342 19954 1348 19956
rect 749 19952 1348 19954
rect 749 19896 754 19952
rect 810 19896 1348 19952
rect 749 19894 1348 19896
rect 749 19891 815 19894
rect 1342 19892 1348 19894
rect 1412 19892 1418 19956
rect 1158 19756 1164 19820
rect 1228 19818 1234 19820
rect 1393 19818 1459 19821
rect 1228 19816 1459 19818
rect 1228 19760 1398 19816
rect 1454 19760 1459 19816
rect 1228 19758 1459 19760
rect 1228 19756 1234 19758
rect 1393 19755 1459 19758
rect 473 18050 539 18053
rect 1526 18050 1532 18052
rect 473 18048 1532 18050
rect 473 17992 478 18048
rect 534 17992 1532 18048
rect 473 17990 1532 17992
rect 473 17987 539 17990
rect 1526 17988 1532 17990
rect 1596 17988 1602 18052
rect 580165 17642 580231 17645
rect 583520 17642 584960 17732
rect 580165 17640 584960 17642
rect 580165 17584 580170 17640
rect 580226 17584 584960 17640
rect 580165 17582 584960 17584
rect 580165 17579 580231 17582
rect 583520 17492 584960 17582
rect 571609 14650 571675 14653
rect 570860 14648 571675 14650
rect 570860 14592 571614 14648
rect 571670 14592 571675 14648
rect 570860 14590 571675 14592
rect 571609 14587 571675 14590
rect 20069 13292 20135 13293
rect 20069 13288 20116 13292
rect 20180 13290 20186 13292
rect 20069 13232 20074 13288
rect 20069 13228 20116 13232
rect 20180 13230 20226 13290
rect 20180 13228 20186 13230
rect 20069 13227 20135 13228
rect 974 12820 980 12884
rect 1044 12882 1050 12884
rect 1117 12882 1183 12885
rect 1044 12880 1183 12882
rect 1044 12824 1122 12880
rect 1178 12824 1183 12880
rect 1044 12822 1183 12824
rect 1044 12820 1050 12822
rect 1117 12819 1183 12822
rect 570321 12340 570387 12341
rect 1166 12205 1226 12308
rect 570270 12276 570276 12340
rect 570340 12338 570387 12340
rect 570340 12336 570432 12338
rect 570382 12280 570432 12336
rect 570340 12278 570432 12280
rect 570340 12276 570387 12278
rect 570321 12275 570387 12276
rect 1117 12200 1226 12205
rect 1117 12144 1122 12200
rect 1178 12144 1226 12200
rect 1117 12142 1226 12144
rect 1117 12139 1183 12142
rect 1577 8804 1643 8805
rect 1526 8740 1532 8804
rect 1596 8802 1643 8804
rect 1596 8800 1688 8802
rect 1638 8744 1688 8800
rect 1596 8742 1688 8744
rect 1596 8740 1643 8742
rect 1577 8739 1643 8740
rect 19977 7988 20043 7989
rect 19926 7924 19932 7988
rect 19996 7986 20043 7988
rect 19996 7984 20088 7986
rect 20038 7928 20088 7984
rect 19996 7926 20088 7928
rect 19996 7924 20043 7926
rect 19977 7923 20043 7924
rect 565 7852 631 7853
rect 565 7850 612 7852
rect 520 7848 612 7850
rect 520 7792 570 7848
rect 520 7790 612 7792
rect 565 7788 612 7790
rect 676 7788 682 7852
rect 565 7787 631 7788
rect -960 7020 480 7260
rect 225689 6490 225755 6493
rect 225822 6490 225828 6492
rect 225689 6488 225828 6490
rect 225689 6432 225694 6488
rect 225750 6432 225828 6488
rect 225689 6430 225828 6432
rect 225689 6427 225755 6430
rect 225822 6428 225828 6430
rect 225892 6428 225898 6492
rect 583520 5796 584960 6036
rect 225781 5132 225847 5133
rect 225781 5130 225828 5132
rect 225736 5128 225828 5130
rect 225736 5072 225786 5128
rect 225736 5070 225828 5072
rect 225781 5068 225828 5070
rect 225892 5068 225898 5132
rect 225781 5067 225847 5068
rect 1209 4450 1275 4453
rect 1342 4450 1348 4452
rect 1209 4448 1348 4450
rect 1209 4392 1214 4448
rect 1270 4392 1348 4448
rect 1209 4390 1348 4392
rect 1209 4387 1275 4390
rect 1342 4388 1348 4390
rect 1412 4388 1418 4452
rect 570321 4450 570387 4453
rect 570454 4450 570460 4452
rect 570321 4448 570460 4450
rect 570321 4392 570326 4448
rect 570382 4392 570460 4448
rect 570321 4390 570460 4392
rect 570321 4387 570387 4390
rect 570454 4388 570460 4390
rect 570524 4388 570530 4452
rect 124305 3772 124371 3773
rect 177941 3772 178007 3773
rect 268377 3772 268443 3773
rect 124300 3708 124306 3772
rect 124370 3770 124376 3772
rect 177936 3770 177942 3772
rect 124370 3710 124462 3770
rect 177850 3710 177942 3770
rect 124370 3708 124376 3710
rect 177936 3708 177942 3710
rect 178006 3708 178012 3772
rect 268372 3708 268378 3772
rect 268442 3770 268448 3772
rect 268442 3710 268534 3770
rect 268442 3708 268448 3710
rect 124305 3707 124371 3708
rect 177941 3707 178007 3708
rect 268377 3707 268443 3708
rect 91732 1804 91738 1868
rect 91802 1866 91808 1868
rect 91802 1806 91984 1866
rect 91802 1804 91808 1806
rect 2998 1668 3004 1732
rect 3068 1730 3074 1732
rect 6085 1730 6151 1733
rect 3068 1728 6151 1730
rect 3068 1672 6090 1728
rect 6146 1672 6151 1728
rect 3068 1670 6151 1672
rect 3068 1668 3074 1670
rect 6085 1667 6151 1670
rect 6821 1730 6887 1733
rect 11237 1730 11303 1733
rect 6821 1728 11303 1730
rect 6821 1672 6826 1728
rect 6882 1672 11242 1728
rect 11298 1672 11303 1728
rect 6821 1670 11303 1672
rect 6821 1667 6887 1670
rect 11237 1667 11303 1670
rect 14457 1730 14523 1733
rect 37365 1730 37431 1733
rect 14457 1728 37431 1730
rect 14457 1672 14462 1728
rect 14518 1672 37370 1728
rect 37426 1672 37431 1728
rect 14457 1670 37431 1672
rect 14457 1667 14523 1670
rect 37365 1667 37431 1670
rect 37733 1730 37799 1733
rect 40953 1730 41019 1733
rect 37733 1728 41019 1730
rect 37733 1672 37738 1728
rect 37794 1672 40958 1728
rect 41014 1672 41019 1728
rect 37733 1670 41019 1672
rect 37733 1667 37799 1670
rect 40953 1667 41019 1670
rect 41137 1730 41203 1733
rect 48681 1730 48747 1733
rect 55029 1730 55095 1733
rect 41137 1728 48747 1730
rect 41137 1672 41142 1728
rect 41198 1672 48686 1728
rect 48742 1672 48747 1728
rect 41137 1670 48747 1672
rect 41137 1667 41203 1670
rect 48681 1667 48747 1670
rect 49190 1728 55095 1730
rect 49190 1672 55034 1728
rect 55090 1672 55095 1728
rect 49190 1670 55095 1672
rect 1853 1594 1919 1597
rect 26417 1594 26483 1597
rect 1853 1592 26483 1594
rect 1853 1536 1858 1592
rect 1914 1536 26422 1592
rect 26478 1536 26483 1592
rect 1853 1534 26483 1536
rect 1853 1531 1919 1534
rect 26417 1531 26483 1534
rect 26601 1594 26667 1597
rect 29729 1594 29795 1597
rect 26601 1592 29795 1594
rect 26601 1536 26606 1592
rect 26662 1536 29734 1592
rect 29790 1536 29795 1592
rect 26601 1534 29795 1536
rect 26601 1531 26667 1534
rect 29729 1531 29795 1534
rect 32673 1594 32739 1597
rect 39389 1594 39455 1597
rect 32673 1592 39455 1594
rect 32673 1536 32678 1592
rect 32734 1536 39394 1592
rect 39450 1536 39455 1592
rect 32673 1534 39455 1536
rect 32673 1531 32739 1534
rect 39389 1531 39455 1534
rect 39757 1594 39823 1597
rect 42517 1594 42583 1597
rect 39757 1592 42583 1594
rect 39757 1536 39762 1592
rect 39818 1536 42522 1592
rect 42578 1536 42583 1592
rect 39757 1534 42583 1536
rect 39757 1531 39823 1534
rect 42517 1531 42583 1534
rect 42701 1594 42767 1597
rect 48037 1594 48103 1597
rect 42701 1592 48103 1594
rect 42701 1536 42706 1592
rect 42762 1536 48042 1592
rect 48098 1536 48103 1592
rect 42701 1534 48103 1536
rect 42701 1531 42767 1534
rect 48037 1531 48103 1534
rect 48681 1594 48747 1597
rect 49190 1594 49250 1670
rect 55029 1667 55095 1670
rect 55213 1730 55279 1733
rect 59077 1730 59143 1733
rect 55213 1728 59143 1730
rect 55213 1672 55218 1728
rect 55274 1672 59082 1728
rect 59138 1672 59143 1728
rect 55213 1670 59143 1672
rect 55213 1667 55279 1670
rect 59077 1667 59143 1670
rect 59261 1730 59327 1733
rect 64873 1730 64939 1733
rect 59261 1728 64939 1730
rect 59261 1672 59266 1728
rect 59322 1672 64878 1728
rect 64934 1672 64939 1728
rect 59261 1670 64939 1672
rect 59261 1667 59327 1670
rect 64873 1667 64939 1670
rect 65006 1668 65012 1732
rect 65076 1730 65082 1732
rect 68686 1730 68692 1732
rect 65076 1670 68692 1730
rect 65076 1668 65082 1670
rect 68686 1668 68692 1670
rect 68756 1668 68762 1732
rect 68829 1730 68895 1733
rect 72417 1730 72483 1733
rect 68829 1728 72483 1730
rect 68829 1672 68834 1728
rect 68890 1672 72422 1728
rect 72478 1672 72483 1728
rect 68829 1670 72483 1672
rect 68829 1667 68895 1670
rect 72417 1667 72483 1670
rect 72550 1668 72556 1732
rect 72620 1730 72626 1732
rect 73705 1730 73771 1733
rect 75310 1730 75316 1732
rect 72620 1728 73771 1730
rect 72620 1672 73710 1728
rect 73766 1672 73771 1728
rect 72620 1670 73771 1672
rect 72620 1668 72626 1670
rect 73705 1667 73771 1670
rect 73846 1670 75316 1730
rect 48681 1592 49250 1594
rect 48681 1536 48686 1592
rect 48742 1536 49250 1592
rect 48681 1534 49250 1536
rect 49325 1594 49391 1597
rect 50797 1594 50863 1597
rect 49325 1592 50863 1594
rect 49325 1536 49330 1592
rect 49386 1536 50802 1592
rect 50858 1536 50863 1592
rect 49325 1534 50863 1536
rect 48681 1531 48747 1534
rect 49325 1531 49391 1534
rect 50797 1531 50863 1534
rect 50981 1594 51047 1597
rect 52310 1594 52316 1596
rect 50981 1592 52316 1594
rect 50981 1536 50986 1592
rect 51042 1536 52316 1592
rect 50981 1534 52316 1536
rect 50981 1531 51047 1534
rect 52310 1532 52316 1534
rect 52380 1532 52386 1596
rect 57881 1594 57947 1597
rect 58433 1594 58499 1597
rect 54894 1592 57947 1594
rect 54894 1536 57886 1592
rect 57942 1536 57947 1592
rect 54894 1534 57947 1536
rect 1485 1458 1551 1461
rect 2998 1458 3004 1460
rect 1485 1456 3004 1458
rect 1485 1400 1490 1456
rect 1546 1400 3004 1456
rect 1485 1398 3004 1400
rect 1485 1395 1551 1398
rect 2998 1396 3004 1398
rect 3068 1396 3074 1460
rect 3693 1458 3759 1461
rect 5901 1458 5967 1461
rect 3693 1456 5967 1458
rect 3693 1400 3698 1456
rect 3754 1400 5906 1456
rect 5962 1400 5967 1456
rect 3693 1398 5967 1400
rect 3693 1395 3759 1398
rect 5901 1395 5967 1398
rect 6085 1458 6151 1461
rect 14457 1458 14523 1461
rect 6085 1456 14523 1458
rect 6085 1400 6090 1456
rect 6146 1400 14462 1456
rect 14518 1400 14523 1456
rect 6085 1398 14523 1400
rect 6085 1395 6151 1398
rect 14457 1395 14523 1398
rect 14641 1458 14707 1461
rect 28257 1458 28323 1461
rect 14641 1456 28323 1458
rect 14641 1400 14646 1456
rect 14702 1400 28262 1456
rect 28318 1400 28323 1456
rect 14641 1398 28323 1400
rect 14641 1395 14707 1398
rect 28257 1395 28323 1398
rect 31477 1458 31543 1461
rect 39062 1458 39068 1460
rect 31477 1456 39068 1458
rect 31477 1400 31482 1456
rect 31538 1400 39068 1456
rect 31477 1398 39068 1400
rect 31477 1395 31543 1398
rect 39062 1396 39068 1398
rect 39132 1396 39138 1460
rect 39297 1458 39363 1461
rect 42241 1458 42307 1461
rect 39297 1456 42307 1458
rect 39297 1400 39302 1456
rect 39358 1400 42246 1456
rect 42302 1400 42307 1456
rect 39297 1398 42307 1400
rect 39297 1395 39363 1398
rect 42241 1395 42307 1398
rect 44081 1458 44147 1461
rect 45461 1458 45527 1461
rect 44081 1456 45527 1458
rect 44081 1400 44086 1456
rect 44142 1400 45466 1456
rect 45522 1400 45527 1456
rect 44081 1398 45527 1400
rect 44081 1395 44147 1398
rect 45461 1395 45527 1398
rect 45645 1458 45711 1461
rect 54894 1458 54954 1534
rect 57881 1531 57947 1534
rect 58022 1592 58499 1594
rect 58022 1536 58438 1592
rect 58494 1536 58499 1592
rect 58022 1534 58499 1536
rect 45645 1456 54954 1458
rect 45645 1400 45650 1456
rect 45706 1400 54954 1456
rect 45645 1398 54954 1400
rect 55029 1458 55095 1461
rect 56358 1458 56364 1460
rect 55029 1456 56364 1458
rect 55029 1400 55034 1456
rect 55090 1400 56364 1456
rect 55029 1398 56364 1400
rect 45645 1395 45711 1398
rect 55029 1395 55095 1398
rect 56358 1396 56364 1398
rect 56428 1396 56434 1460
rect 56593 1458 56659 1461
rect 58022 1458 58082 1534
rect 58433 1531 58499 1534
rect 58566 1532 58572 1596
rect 58636 1594 58642 1596
rect 61009 1594 61075 1597
rect 58636 1592 61075 1594
rect 58636 1536 61014 1592
rect 61070 1536 61075 1592
rect 58636 1534 61075 1536
rect 58636 1532 58642 1534
rect 61009 1531 61075 1534
rect 61193 1594 61259 1597
rect 64505 1594 64571 1597
rect 61193 1592 64571 1594
rect 61193 1536 61198 1592
rect 61254 1536 64510 1592
rect 64566 1536 64571 1592
rect 61193 1534 64571 1536
rect 61193 1531 61259 1534
rect 64505 1531 64571 1534
rect 65333 1594 65399 1597
rect 66662 1594 66668 1596
rect 65333 1592 66668 1594
rect 65333 1536 65338 1592
rect 65394 1536 66668 1592
rect 65333 1534 66668 1536
rect 65333 1531 65399 1534
rect 66662 1532 66668 1534
rect 66732 1532 66738 1596
rect 66897 1594 66963 1597
rect 73102 1594 73108 1596
rect 66897 1592 73108 1594
rect 66897 1536 66902 1592
rect 66958 1536 73108 1592
rect 66897 1534 73108 1536
rect 66897 1531 66963 1534
rect 73102 1532 73108 1534
rect 73172 1532 73178 1596
rect 73286 1532 73292 1596
rect 73356 1594 73362 1596
rect 73846 1594 73906 1670
rect 75310 1668 75316 1670
rect 75380 1668 75386 1732
rect 76046 1668 76052 1732
rect 76116 1730 76122 1732
rect 76782 1730 76788 1732
rect 76116 1670 76788 1730
rect 76116 1668 76122 1670
rect 76782 1668 76788 1670
rect 76852 1668 76858 1732
rect 82486 1730 82492 1732
rect 76974 1670 82492 1730
rect 73356 1534 73906 1594
rect 74073 1594 74139 1597
rect 75361 1594 75427 1597
rect 74073 1592 75427 1594
rect 74073 1536 74078 1592
rect 74134 1536 75366 1592
rect 75422 1536 75427 1592
rect 74073 1534 75427 1536
rect 73356 1532 73362 1534
rect 74073 1531 74139 1534
rect 75361 1531 75427 1534
rect 75494 1532 75500 1596
rect 75564 1594 75570 1596
rect 76189 1594 76255 1597
rect 75564 1592 76255 1594
rect 75564 1536 76194 1592
rect 76250 1536 76255 1592
rect 75564 1534 76255 1536
rect 75564 1532 75570 1534
rect 76189 1531 76255 1534
rect 76414 1532 76420 1596
rect 76484 1594 76490 1596
rect 76974 1594 77034 1670
rect 82486 1668 82492 1670
rect 82556 1668 82562 1732
rect 82629 1730 82695 1733
rect 83590 1730 83596 1732
rect 82629 1728 83596 1730
rect 82629 1672 82634 1728
rect 82690 1672 83596 1728
rect 82629 1670 83596 1672
rect 82629 1667 82695 1670
rect 83590 1668 83596 1670
rect 83660 1668 83666 1732
rect 83733 1730 83799 1733
rect 85665 1730 85731 1733
rect 83733 1728 85731 1730
rect 83733 1672 83738 1728
rect 83794 1672 85670 1728
rect 85726 1672 85731 1728
rect 83733 1670 85731 1672
rect 83733 1667 83799 1670
rect 85665 1667 85731 1670
rect 85798 1668 85804 1732
rect 85868 1730 85874 1732
rect 88006 1730 88012 1732
rect 85868 1670 88012 1730
rect 85868 1668 85874 1670
rect 88006 1668 88012 1670
rect 88076 1668 88082 1732
rect 88190 1668 88196 1732
rect 88260 1730 88266 1732
rect 91924 1730 91984 1806
rect 92790 1730 92796 1732
rect 88260 1670 91524 1730
rect 91924 1670 92796 1730
rect 88260 1668 88266 1670
rect 76484 1534 77034 1594
rect 77109 1594 77175 1597
rect 78397 1594 78463 1597
rect 77109 1592 78463 1594
rect 77109 1536 77114 1592
rect 77170 1536 78402 1592
rect 78458 1536 78463 1592
rect 77109 1534 78463 1536
rect 76484 1532 76490 1534
rect 77109 1531 77175 1534
rect 78397 1531 78463 1534
rect 78581 1594 78647 1597
rect 82261 1594 82327 1597
rect 78581 1592 82327 1594
rect 78581 1536 78586 1592
rect 78642 1536 82266 1592
rect 82322 1536 82327 1592
rect 78581 1534 82327 1536
rect 78581 1531 78647 1534
rect 82261 1531 82327 1534
rect 83038 1532 83044 1596
rect 83108 1594 83114 1596
rect 91464 1594 91524 1670
rect 92790 1668 92796 1670
rect 92860 1668 92866 1732
rect 92974 1668 92980 1732
rect 93044 1730 93050 1732
rect 94446 1730 94452 1732
rect 93044 1670 94452 1730
rect 93044 1668 93050 1670
rect 94446 1668 94452 1670
rect 94516 1668 94522 1732
rect 95366 1730 95372 1732
rect 94638 1670 95372 1730
rect 92565 1594 92631 1597
rect 83108 1534 91386 1594
rect 91464 1592 92631 1594
rect 91464 1536 92570 1592
rect 92626 1536 92631 1592
rect 91464 1534 92631 1536
rect 83108 1532 83114 1534
rect 56593 1456 58082 1458
rect 56593 1400 56598 1456
rect 56654 1400 58082 1456
rect 56593 1398 58082 1400
rect 58525 1458 58591 1461
rect 62389 1458 62455 1461
rect 58525 1456 62455 1458
rect 58525 1400 58530 1456
rect 58586 1400 62394 1456
rect 62450 1400 62455 1456
rect 58525 1398 62455 1400
rect 56593 1395 56659 1398
rect 58525 1395 58591 1398
rect 62389 1395 62455 1398
rect 62941 1458 63007 1461
rect 66897 1458 66963 1461
rect 62941 1456 66963 1458
rect 62941 1400 62946 1456
rect 63002 1400 66902 1456
rect 66958 1400 66963 1456
rect 62941 1398 66963 1400
rect 62941 1395 63007 1398
rect 66897 1395 66963 1398
rect 67081 1458 67147 1461
rect 73470 1458 73476 1460
rect 67081 1456 73476 1458
rect 67081 1400 67086 1456
rect 67142 1400 73476 1456
rect 67081 1398 73476 1400
rect 67081 1395 67147 1398
rect 73470 1396 73476 1398
rect 73540 1396 73546 1460
rect 73981 1458 74047 1461
rect 83181 1458 83247 1461
rect 83365 1460 83431 1461
rect 83365 1458 83412 1460
rect 73981 1456 83247 1458
rect 73981 1400 73986 1456
rect 74042 1400 83186 1456
rect 83242 1400 83247 1456
rect 73981 1398 83247 1400
rect 83320 1456 83412 1458
rect 83320 1400 83370 1456
rect 83320 1398 83412 1400
rect 73981 1395 74047 1398
rect 83181 1395 83247 1398
rect 83365 1396 83412 1398
rect 83476 1396 83482 1460
rect 83641 1458 83707 1461
rect 91326 1458 91386 1534
rect 92565 1531 92631 1534
rect 92749 1594 92815 1597
rect 94638 1594 94698 1670
rect 95366 1668 95372 1670
rect 95436 1668 95442 1732
rect 95550 1668 95556 1732
rect 95620 1730 95626 1732
rect 100334 1730 100340 1732
rect 95620 1670 100340 1730
rect 95620 1668 95626 1670
rect 100334 1668 100340 1670
rect 100404 1668 100410 1732
rect 100477 1730 100543 1733
rect 102734 1730 103116 1764
rect 111425 1730 111491 1733
rect 100477 1728 111491 1730
rect 100477 1672 100482 1728
rect 100538 1704 111430 1728
rect 100538 1672 102794 1704
rect 100477 1670 102794 1672
rect 103056 1672 111430 1704
rect 111486 1672 111491 1728
rect 103056 1670 111491 1672
rect 100477 1667 100543 1670
rect 111425 1667 111491 1670
rect 111558 1668 111564 1732
rect 111628 1730 111634 1732
rect 120625 1730 120691 1733
rect 111628 1728 120691 1730
rect 111628 1672 120630 1728
rect 120686 1672 120691 1728
rect 111628 1670 120691 1672
rect 111628 1668 111634 1670
rect 120625 1667 120691 1670
rect 120758 1668 120764 1732
rect 120828 1730 120834 1732
rect 122281 1730 122347 1733
rect 124305 1730 124371 1733
rect 120828 1670 122160 1730
rect 120828 1668 120834 1670
rect 92749 1592 94698 1594
rect 92749 1536 92754 1592
rect 92810 1536 94698 1592
rect 92749 1534 94698 1536
rect 92749 1531 92815 1534
rect 94814 1532 94820 1596
rect 94884 1594 94890 1596
rect 95734 1594 95740 1596
rect 94884 1534 95740 1594
rect 94884 1532 94890 1534
rect 95734 1532 95740 1534
rect 95804 1532 95810 1596
rect 96429 1594 96495 1597
rect 96613 1594 96679 1597
rect 96429 1592 96679 1594
rect 96429 1536 96434 1592
rect 96490 1536 96618 1592
rect 96674 1536 96679 1592
rect 96429 1534 96679 1536
rect 96429 1531 96495 1534
rect 96613 1531 96679 1534
rect 96981 1594 97047 1597
rect 101673 1594 101739 1597
rect 96981 1592 101739 1594
rect 96981 1536 96986 1592
rect 97042 1536 101678 1592
rect 101734 1536 101739 1592
rect 96981 1534 101739 1536
rect 96981 1531 97047 1534
rect 101673 1531 101739 1534
rect 101806 1532 101812 1596
rect 101876 1594 101882 1596
rect 103278 1594 103284 1596
rect 101876 1534 103284 1594
rect 101876 1532 101882 1534
rect 103278 1532 103284 1534
rect 103348 1532 103354 1596
rect 103421 1594 103487 1597
rect 111241 1596 111307 1597
rect 103421 1592 111120 1594
rect 103421 1536 103426 1592
rect 103482 1536 111120 1592
rect 103421 1534 111120 1536
rect 103421 1531 103487 1534
rect 91921 1458 91987 1461
rect 100937 1458 101003 1461
rect 101121 1460 101187 1461
rect 83641 1456 91202 1458
rect 83641 1400 83646 1456
rect 83702 1400 91202 1456
rect 83641 1398 91202 1400
rect 91326 1456 91987 1458
rect 91326 1400 91926 1456
rect 91982 1400 91987 1456
rect 91326 1398 91987 1400
rect 83365 1395 83431 1396
rect 83641 1395 83707 1398
rect 749 1322 815 1325
rect 60273 1322 60339 1325
rect 749 1320 60339 1322
rect 749 1264 754 1320
rect 810 1264 60278 1320
rect 60334 1264 60339 1320
rect 749 1262 60339 1264
rect 749 1259 815 1262
rect 60273 1259 60339 1262
rect 60825 1322 60891 1325
rect 63033 1322 63099 1325
rect 60825 1320 63099 1322
rect 60825 1264 60830 1320
rect 60886 1264 63038 1320
rect 63094 1264 63099 1320
rect 60825 1262 63099 1264
rect 60825 1259 60891 1262
rect 63033 1259 63099 1262
rect 63769 1322 63835 1325
rect 83038 1322 83044 1324
rect 63769 1320 83044 1322
rect 63769 1264 63774 1320
rect 63830 1264 83044 1320
rect 63769 1262 83044 1264
rect 63769 1259 63835 1262
rect 83038 1260 83044 1262
rect 83108 1260 83114 1324
rect 83222 1260 83228 1324
rect 83292 1322 83298 1324
rect 85849 1322 85915 1325
rect 83292 1320 85915 1322
rect 83292 1264 85854 1320
rect 85910 1264 85915 1320
rect 83292 1262 85915 1264
rect 83292 1260 83298 1262
rect 85849 1259 85915 1262
rect 86033 1322 86099 1325
rect 90950 1322 90956 1324
rect 86033 1320 90956 1322
rect 86033 1264 86038 1320
rect 86094 1264 90956 1320
rect 86033 1262 90956 1264
rect 86033 1259 86099 1262
rect 90950 1260 90956 1262
rect 91020 1260 91026 1324
rect 91142 1322 91202 1398
rect 91921 1395 91987 1398
rect 92062 1456 101003 1458
rect 92062 1400 100942 1456
rect 100998 1400 101003 1456
rect 92062 1398 101003 1400
rect 92062 1322 92122 1398
rect 100937 1395 101003 1398
rect 101070 1396 101076 1460
rect 101140 1458 101187 1460
rect 101305 1458 101371 1461
rect 102777 1458 102843 1461
rect 101140 1456 101232 1458
rect 101182 1400 101232 1456
rect 101140 1398 101232 1400
rect 101305 1456 102843 1458
rect 101305 1400 101310 1456
rect 101366 1400 102782 1456
rect 102838 1400 102843 1456
rect 101305 1398 102843 1400
rect 101140 1396 101187 1398
rect 101121 1395 101187 1396
rect 101305 1395 101371 1398
rect 102777 1395 102843 1398
rect 102910 1396 102916 1460
rect 102980 1396 102986 1460
rect 103053 1458 103119 1461
rect 110781 1458 110847 1461
rect 103053 1456 110847 1458
rect 103053 1400 103058 1456
rect 103114 1400 110786 1456
rect 110842 1400 110847 1456
rect 103053 1398 110847 1400
rect 111060 1458 111120 1534
rect 111190 1532 111196 1596
rect 111260 1594 111307 1596
rect 112161 1594 112227 1597
rect 120165 1594 120231 1597
rect 121913 1594 121979 1597
rect 111260 1592 111352 1594
rect 111302 1536 111352 1592
rect 111260 1534 111352 1536
rect 112161 1592 120231 1594
rect 112161 1536 112166 1592
rect 112222 1536 120170 1592
rect 120226 1536 120231 1592
rect 112161 1534 120231 1536
rect 111260 1532 111307 1534
rect 111241 1531 111307 1532
rect 112161 1531 112227 1534
rect 120165 1531 120231 1534
rect 120766 1592 121979 1594
rect 120766 1536 121918 1592
rect 121974 1536 121979 1592
rect 120766 1534 121979 1536
rect 122100 1594 122160 1670
rect 122281 1728 124371 1730
rect 122281 1672 122286 1728
rect 122342 1672 124310 1728
rect 124366 1672 124371 1728
rect 122281 1670 124371 1672
rect 122281 1667 122347 1670
rect 124305 1667 124371 1670
rect 124438 1668 124444 1732
rect 124508 1730 124514 1732
rect 125777 1730 125843 1733
rect 124508 1728 125843 1730
rect 124508 1672 125782 1728
rect 125838 1672 125843 1728
rect 124508 1670 125843 1672
rect 124508 1668 124514 1670
rect 125777 1667 125843 1670
rect 125910 1668 125916 1732
rect 125980 1730 125986 1732
rect 127934 1730 127940 1732
rect 125980 1670 127940 1730
rect 125980 1668 125986 1670
rect 127934 1668 127940 1670
rect 128004 1668 128010 1732
rect 128261 1730 128327 1733
rect 128854 1730 128860 1732
rect 128261 1728 128860 1730
rect 128261 1672 128266 1728
rect 128322 1672 128860 1728
rect 128261 1670 128860 1672
rect 128261 1667 128327 1670
rect 128854 1668 128860 1670
rect 128924 1668 128930 1732
rect 128997 1730 129063 1733
rect 135161 1730 135227 1733
rect 135345 1732 135411 1733
rect 128997 1728 135227 1730
rect 128997 1672 129002 1728
rect 129058 1672 135166 1728
rect 135222 1672 135227 1728
rect 128997 1670 135227 1672
rect 128997 1667 129063 1670
rect 135161 1667 135227 1670
rect 135294 1668 135300 1732
rect 135364 1730 135411 1732
rect 135621 1732 135687 1733
rect 135364 1728 135456 1730
rect 135406 1672 135456 1728
rect 135364 1670 135456 1672
rect 135621 1728 135668 1732
rect 135732 1730 135738 1732
rect 135621 1672 135626 1728
rect 135364 1668 135411 1670
rect 135345 1667 135411 1668
rect 135621 1668 135668 1672
rect 135732 1670 135778 1730
rect 135732 1668 135738 1670
rect 136076 1668 136082 1732
rect 136146 1730 136152 1732
rect 136265 1730 136331 1733
rect 136146 1728 136331 1730
rect 136146 1672 136270 1728
rect 136326 1672 136331 1728
rect 136146 1670 136331 1672
rect 136146 1668 136152 1670
rect 135621 1667 135687 1668
rect 136265 1667 136331 1670
rect 136398 1668 136404 1732
rect 136468 1730 136474 1732
rect 138381 1730 138447 1733
rect 136468 1728 138447 1730
rect 136468 1672 138386 1728
rect 138442 1672 138447 1728
rect 136468 1670 138447 1672
rect 136468 1668 136474 1670
rect 138381 1667 138447 1670
rect 139342 1668 139348 1732
rect 139412 1730 139418 1732
rect 140998 1730 141004 1732
rect 139412 1670 141004 1730
rect 139412 1668 139418 1670
rect 140998 1668 141004 1670
rect 141068 1668 141074 1732
rect 141141 1730 141207 1733
rect 141141 1728 141572 1730
rect 141141 1672 141146 1728
rect 141202 1672 141572 1728
rect 141141 1670 141572 1672
rect 141141 1667 141207 1670
rect 127801 1594 127867 1597
rect 122100 1592 127867 1594
rect 122100 1536 127806 1592
rect 127862 1536 127867 1592
rect 122100 1534 127867 1536
rect 111241 1458 111307 1461
rect 111060 1456 111307 1458
rect 111060 1400 111246 1456
rect 111302 1400 111307 1456
rect 111060 1398 111307 1400
rect 91142 1262 92122 1322
rect 92197 1322 92263 1325
rect 96470 1322 96476 1324
rect 92197 1320 96476 1322
rect 92197 1264 92202 1320
rect 92258 1264 96476 1320
rect 92197 1262 96476 1264
rect 92197 1259 92263 1262
rect 96470 1260 96476 1262
rect 96540 1260 96546 1324
rect 96613 1322 96679 1325
rect 97758 1322 97764 1324
rect 96613 1320 97764 1322
rect 96613 1264 96618 1320
rect 96674 1264 97764 1320
rect 96613 1262 97764 1264
rect 96613 1259 96679 1262
rect 97758 1260 97764 1262
rect 97828 1260 97834 1324
rect 97901 1322 97967 1325
rect 100201 1322 100267 1325
rect 97901 1320 100267 1322
rect 97901 1264 97906 1320
rect 97962 1264 100206 1320
rect 100262 1264 100267 1320
rect 97901 1262 100267 1264
rect 97901 1259 97967 1262
rect 100201 1259 100267 1262
rect 100334 1260 100340 1324
rect 100404 1322 100410 1324
rect 101254 1322 101260 1324
rect 100404 1262 101260 1322
rect 100404 1260 100410 1262
rect 101254 1260 101260 1262
rect 101324 1260 101330 1324
rect 101397 1322 101463 1325
rect 102317 1324 102383 1325
rect 102174 1322 102180 1324
rect 101397 1320 102180 1322
rect 101397 1264 101402 1320
rect 101458 1264 102180 1320
rect 101397 1262 102180 1264
rect 101397 1259 101463 1262
rect 102174 1260 102180 1262
rect 102244 1260 102250 1324
rect 102317 1320 102364 1324
rect 102428 1322 102434 1324
rect 102593 1322 102659 1325
rect 102918 1322 102978 1396
rect 103053 1395 103119 1398
rect 110781 1395 110847 1398
rect 111241 1395 111307 1398
rect 111425 1458 111491 1461
rect 111742 1458 111748 1460
rect 111425 1456 111748 1458
rect 111425 1400 111430 1456
rect 111486 1400 111748 1456
rect 111425 1398 111748 1400
rect 111425 1395 111491 1398
rect 111742 1396 111748 1398
rect 111812 1396 111818 1460
rect 111977 1458 112043 1461
rect 120625 1458 120691 1461
rect 120766 1460 120826 1534
rect 121913 1531 121979 1534
rect 127801 1531 127867 1534
rect 127985 1594 128051 1597
rect 128486 1594 128492 1596
rect 127985 1592 128492 1594
rect 127985 1536 127990 1592
rect 128046 1536 128492 1592
rect 127985 1534 128492 1536
rect 127985 1531 128051 1534
rect 128486 1532 128492 1534
rect 128556 1532 128562 1596
rect 134885 1594 134951 1597
rect 128816 1592 134951 1594
rect 128816 1536 134890 1592
rect 134946 1536 134951 1592
rect 128816 1534 134951 1536
rect 128816 1492 128876 1534
rect 134885 1531 134951 1534
rect 135069 1594 135135 1597
rect 136541 1594 136607 1597
rect 140773 1594 140839 1597
rect 135069 1592 136607 1594
rect 135069 1536 135074 1592
rect 135130 1536 136546 1592
rect 136602 1536 136607 1592
rect 135069 1534 136607 1536
rect 135069 1531 135135 1534
rect 136541 1531 136607 1534
rect 136728 1592 140839 1594
rect 136728 1536 140778 1592
rect 140834 1536 140839 1592
rect 136728 1534 140839 1536
rect 111977 1456 120691 1458
rect 111977 1400 111982 1456
rect 112038 1400 120630 1456
rect 120686 1400 120691 1456
rect 111977 1398 120691 1400
rect 111977 1395 112043 1398
rect 120625 1395 120691 1398
rect 120758 1396 120764 1460
rect 120828 1396 120834 1460
rect 120901 1458 120967 1461
rect 127709 1458 127775 1461
rect 120901 1456 127775 1458
rect 120901 1400 120906 1456
rect 120962 1400 127714 1456
rect 127770 1400 127775 1456
rect 120901 1398 127775 1400
rect 120901 1395 120967 1398
rect 127709 1395 127775 1398
rect 127893 1458 127959 1461
rect 128678 1458 128876 1492
rect 127893 1456 128876 1458
rect 127893 1400 127898 1456
rect 127954 1432 128876 1456
rect 128997 1458 129063 1461
rect 134793 1458 134859 1461
rect 135110 1458 135116 1460
rect 128997 1456 134859 1458
rect 127954 1400 128738 1432
rect 127893 1398 128738 1400
rect 128997 1400 129002 1456
rect 129058 1400 134798 1456
rect 134854 1400 134859 1456
rect 128997 1398 134859 1400
rect 127893 1395 127959 1398
rect 128997 1395 129063 1398
rect 134793 1395 134859 1398
rect 134934 1398 135116 1458
rect 102317 1264 102322 1320
rect 102317 1260 102364 1264
rect 102428 1262 102474 1322
rect 102593 1320 102978 1322
rect 102593 1264 102598 1320
rect 102654 1264 102978 1320
rect 102593 1262 102978 1264
rect 103053 1322 103119 1325
rect 103278 1322 103284 1324
rect 103053 1320 103284 1322
rect 103053 1264 103058 1320
rect 103114 1264 103284 1320
rect 103053 1262 103284 1264
rect 102428 1260 102434 1262
rect 102317 1259 102383 1260
rect 102593 1259 102659 1262
rect 103053 1259 103119 1262
rect 103278 1260 103284 1262
rect 103348 1260 103354 1324
rect 103513 1322 103579 1325
rect 106733 1322 106799 1325
rect 116853 1322 116919 1325
rect 103513 1320 106799 1322
rect 103513 1264 103518 1320
rect 103574 1264 106738 1320
rect 106794 1264 106799 1320
rect 103513 1262 106799 1264
rect 103513 1259 103579 1262
rect 106733 1259 106799 1262
rect 106966 1320 116919 1322
rect 106966 1264 116858 1320
rect 116914 1264 116919 1320
rect 106966 1262 116919 1264
rect 2814 1124 2820 1188
rect 2884 1186 2890 1188
rect 10409 1186 10475 1189
rect 2884 1184 10475 1186
rect 2884 1128 10414 1184
rect 10470 1128 10475 1184
rect 2884 1126 10475 1128
rect 2884 1124 2890 1126
rect 10409 1123 10475 1126
rect 10910 1124 10916 1188
rect 10980 1186 10986 1188
rect 39297 1186 39363 1189
rect 10980 1184 39363 1186
rect 10980 1128 39302 1184
rect 39358 1128 39363 1184
rect 10980 1126 39363 1128
rect 10980 1124 10986 1126
rect 39297 1123 39363 1126
rect 39430 1124 39436 1188
rect 39500 1186 39506 1188
rect 42057 1186 42123 1189
rect 39500 1184 42123 1186
rect 39500 1128 42062 1184
rect 42118 1128 42123 1184
rect 39500 1126 42123 1128
rect 39500 1124 39506 1126
rect 42057 1123 42123 1126
rect 42241 1186 42307 1189
rect 58157 1186 58223 1189
rect 42241 1184 58223 1186
rect 42241 1128 42246 1184
rect 42302 1128 58162 1184
rect 58218 1128 58223 1184
rect 42241 1126 58223 1128
rect 42241 1123 42307 1126
rect 58157 1123 58223 1126
rect 58341 1186 58407 1189
rect 60590 1186 60596 1188
rect 58341 1184 60596 1186
rect 58341 1128 58346 1184
rect 58402 1128 60596 1184
rect 58341 1126 60596 1128
rect 58341 1123 58407 1126
rect 60590 1124 60596 1126
rect 60660 1124 60666 1188
rect 60733 1186 60799 1189
rect 63309 1186 63375 1189
rect 60733 1184 63375 1186
rect 60733 1128 60738 1184
rect 60794 1128 63314 1184
rect 63370 1128 63375 1184
rect 60733 1126 63375 1128
rect 60733 1123 60799 1126
rect 63309 1123 63375 1126
rect 63861 1186 63927 1189
rect 64638 1186 64644 1188
rect 63861 1184 64644 1186
rect 63861 1128 63866 1184
rect 63922 1128 64644 1184
rect 63861 1126 64644 1128
rect 63861 1123 63927 1126
rect 64638 1124 64644 1126
rect 64708 1124 64714 1188
rect 64781 1186 64847 1189
rect 66713 1186 66779 1189
rect 64781 1184 66779 1186
rect 64781 1128 64786 1184
rect 64842 1128 66718 1184
rect 66774 1128 66779 1184
rect 64781 1126 66779 1128
rect 64781 1123 64847 1126
rect 66713 1123 66779 1126
rect 66846 1124 66852 1188
rect 66916 1186 66922 1188
rect 82169 1186 82235 1189
rect 66916 1184 82235 1186
rect 66916 1128 82174 1184
rect 82230 1128 82235 1184
rect 66916 1126 82235 1128
rect 66916 1124 66922 1126
rect 82169 1123 82235 1126
rect 82302 1124 82308 1188
rect 82372 1124 82378 1188
rect 82670 1124 82676 1188
rect 82740 1186 82746 1188
rect 90582 1186 90588 1188
rect 82740 1126 90588 1186
rect 82740 1124 82746 1126
rect 90582 1124 90588 1126
rect 90652 1124 90658 1188
rect 90725 1186 90791 1189
rect 92197 1186 92263 1189
rect 90725 1184 92263 1186
rect 90725 1128 90730 1184
rect 90786 1128 92202 1184
rect 92258 1128 92263 1184
rect 90725 1126 92263 1128
rect 1209 1050 1275 1053
rect 26877 1050 26943 1053
rect 1209 1048 26943 1050
rect 1209 992 1214 1048
rect 1270 992 26882 1048
rect 26938 992 26943 1048
rect 1209 990 26943 992
rect 1209 987 1275 990
rect 26877 987 26943 990
rect 27889 1050 27955 1053
rect 46565 1050 46631 1053
rect 46749 1052 46815 1053
rect 46749 1050 46796 1052
rect 27889 1048 46631 1050
rect 27889 992 27894 1048
rect 27950 992 46570 1048
rect 46626 992 46631 1048
rect 27889 990 46631 992
rect 46704 1048 46796 1050
rect 46704 992 46754 1048
rect 46704 990 46796 992
rect 27889 987 27955 990
rect 46565 987 46631 990
rect 46749 988 46796 990
rect 46860 988 46866 1052
rect 47025 1050 47091 1053
rect 63493 1050 63559 1053
rect 47025 1048 63559 1050
rect 47025 992 47030 1048
rect 47086 992 63498 1048
rect 63554 992 63559 1048
rect 47025 990 63559 992
rect 46749 987 46815 988
rect 47025 987 47091 990
rect 63493 987 63559 990
rect 63718 988 63724 1052
rect 63788 1050 63794 1052
rect 72918 1050 72924 1052
rect 63788 990 72924 1050
rect 63788 988 63794 990
rect 72918 988 72924 990
rect 72988 988 72994 1052
rect 73102 988 73108 1052
rect 73172 1050 73178 1052
rect 73337 1050 73403 1053
rect 73172 1048 73403 1050
rect 73172 992 73342 1048
rect 73398 992 73403 1048
rect 73172 990 73403 992
rect 73172 988 73178 990
rect 73337 987 73403 990
rect 73470 988 73476 1052
rect 73540 1050 73546 1052
rect 74257 1050 74323 1053
rect 73540 1048 74323 1050
rect 73540 992 74262 1048
rect 74318 992 74323 1048
rect 73540 990 74323 992
rect 73540 988 73546 990
rect 74257 987 74323 990
rect 74441 1050 74507 1053
rect 82310 1050 82370 1124
rect 90725 1123 90791 1126
rect 92197 1123 92263 1126
rect 92422 1124 92428 1188
rect 92492 1186 92498 1188
rect 101254 1186 101260 1188
rect 92492 1126 101260 1186
rect 92492 1124 92498 1126
rect 101254 1124 101260 1126
rect 101324 1124 101330 1188
rect 101397 1186 101463 1189
rect 104617 1186 104683 1189
rect 101397 1184 104683 1186
rect 101397 1128 101402 1184
rect 101458 1128 104622 1184
rect 104678 1128 104683 1184
rect 101397 1126 104683 1128
rect 101397 1123 101463 1126
rect 104617 1123 104683 1126
rect 104801 1186 104867 1189
rect 106825 1186 106891 1189
rect 104801 1184 106891 1186
rect 104801 1128 104806 1184
rect 104862 1128 106830 1184
rect 106886 1128 106891 1184
rect 104801 1126 106891 1128
rect 104801 1123 104867 1126
rect 106825 1123 106891 1126
rect 83222 1050 83228 1052
rect 74441 1048 82370 1050
rect 74441 992 74446 1048
rect 74502 992 82370 1048
rect 74441 990 82370 992
rect 82494 990 83228 1050
rect 74441 987 74507 990
rect 82494 917 82554 990
rect 83222 988 83228 990
rect 83292 988 83298 1052
rect 83406 988 83412 1052
rect 83476 1050 83482 1052
rect 97073 1050 97139 1053
rect 83476 1048 97139 1050
rect 83476 992 97078 1048
rect 97134 992 97139 1048
rect 83476 990 97139 992
rect 83476 988 83482 990
rect 97073 987 97139 990
rect 97257 1050 97323 1053
rect 106966 1050 107026 1262
rect 116853 1259 116919 1262
rect 117037 1322 117103 1325
rect 121821 1322 121887 1325
rect 117037 1320 121887 1322
rect 117037 1264 117042 1320
rect 117098 1264 121826 1320
rect 121882 1264 121887 1320
rect 117037 1262 121887 1264
rect 117037 1259 117103 1262
rect 121821 1259 121887 1262
rect 122005 1322 122071 1325
rect 131297 1322 131363 1325
rect 131481 1324 131547 1325
rect 122005 1320 131363 1322
rect 122005 1264 122010 1320
rect 122066 1264 131302 1320
rect 131358 1264 131363 1320
rect 122005 1262 131363 1264
rect 122005 1259 122071 1262
rect 131297 1259 131363 1262
rect 131430 1260 131436 1324
rect 131500 1322 131547 1324
rect 131665 1322 131731 1325
rect 134374 1322 134380 1324
rect 131500 1320 131592 1322
rect 131542 1264 131592 1320
rect 131500 1262 131592 1264
rect 131665 1320 134380 1322
rect 131665 1264 131670 1320
rect 131726 1264 134380 1320
rect 131665 1262 134380 1264
rect 131500 1260 131547 1262
rect 131481 1259 131547 1260
rect 131665 1259 131731 1262
rect 134374 1260 134380 1262
rect 134444 1260 134450 1324
rect 134701 1322 134767 1325
rect 134934 1322 134994 1398
rect 135110 1396 135116 1398
rect 135180 1396 135186 1460
rect 135529 1458 135595 1461
rect 136582 1458 136588 1460
rect 135529 1456 136588 1458
rect 135529 1400 135534 1456
rect 135590 1400 136588 1456
rect 135529 1398 136588 1400
rect 135529 1395 135595 1398
rect 136582 1396 136588 1398
rect 136652 1396 136658 1460
rect 134701 1320 134994 1322
rect 134701 1264 134706 1320
rect 134762 1264 134994 1320
rect 134701 1262 134994 1264
rect 135069 1322 135135 1325
rect 135897 1322 135963 1325
rect 135069 1320 135963 1322
rect 135069 1264 135074 1320
rect 135130 1264 135902 1320
rect 135958 1264 135963 1320
rect 135069 1262 135963 1264
rect 134701 1259 134767 1262
rect 135069 1259 135135 1262
rect 135897 1259 135963 1262
rect 136357 1322 136423 1325
rect 136728 1322 136788 1534
rect 140773 1531 140839 1534
rect 140957 1594 141023 1597
rect 141512 1594 141572 1670
rect 141734 1668 141740 1732
rect 141804 1730 141810 1732
rect 144361 1730 144427 1733
rect 141804 1728 144427 1730
rect 141804 1672 144366 1728
rect 144422 1672 144427 1728
rect 141804 1670 144427 1672
rect 141804 1668 141810 1670
rect 144361 1667 144427 1670
rect 145097 1730 145163 1733
rect 145649 1730 145715 1733
rect 145833 1732 145899 1733
rect 146201 1732 146267 1733
rect 145097 1728 145715 1730
rect 145097 1672 145102 1728
rect 145158 1672 145654 1728
rect 145710 1672 145715 1728
rect 145097 1670 145715 1672
rect 145097 1667 145163 1670
rect 145649 1667 145715 1670
rect 145782 1668 145788 1732
rect 145852 1730 145899 1732
rect 146150 1730 146156 1732
rect 145852 1728 145944 1730
rect 145894 1672 145944 1728
rect 145852 1670 145944 1672
rect 146110 1670 146156 1730
rect 146220 1728 146267 1732
rect 146262 1672 146267 1728
rect 145852 1668 145899 1670
rect 146150 1668 146156 1670
rect 146220 1668 146267 1672
rect 146334 1668 146340 1732
rect 146404 1730 146410 1732
rect 148041 1730 148107 1733
rect 146404 1728 148107 1730
rect 146404 1672 148046 1728
rect 148102 1672 148107 1728
rect 146404 1670 148107 1672
rect 146404 1668 146410 1670
rect 145833 1667 145899 1668
rect 146201 1667 146267 1668
rect 148041 1667 148107 1670
rect 148174 1668 148180 1732
rect 148244 1730 148250 1732
rect 148961 1730 149027 1733
rect 148244 1728 149027 1730
rect 148244 1672 148966 1728
rect 149022 1672 149027 1728
rect 148244 1670 149027 1672
rect 148244 1668 148250 1670
rect 148961 1667 149027 1670
rect 149145 1730 149211 1733
rect 152222 1730 152228 1732
rect 149145 1728 152228 1730
rect 149145 1672 149150 1728
rect 149206 1672 152228 1728
rect 149145 1670 152228 1672
rect 149145 1667 149211 1670
rect 152222 1668 152228 1670
rect 152292 1668 152298 1732
rect 154297 1730 154363 1733
rect 152782 1728 154363 1730
rect 152782 1672 154302 1728
rect 154358 1672 154363 1728
rect 152782 1670 154363 1672
rect 144862 1594 144868 1596
rect 140957 1592 141434 1594
rect 140957 1536 140962 1592
rect 141018 1536 141434 1592
rect 140957 1534 141434 1536
rect 141512 1534 144868 1594
rect 140957 1531 141023 1534
rect 136909 1458 136975 1461
rect 138606 1458 138612 1460
rect 136909 1456 138612 1458
rect 136909 1400 136914 1456
rect 136970 1400 138612 1456
rect 136909 1398 138612 1400
rect 136909 1395 136975 1398
rect 138606 1396 138612 1398
rect 138676 1396 138682 1460
rect 138790 1396 138796 1460
rect 138860 1458 138866 1460
rect 139209 1458 139275 1461
rect 138860 1456 139275 1458
rect 138860 1400 139214 1456
rect 139270 1400 139275 1456
rect 138860 1398 139275 1400
rect 138860 1396 138866 1398
rect 139209 1395 139275 1398
rect 139577 1458 139643 1461
rect 140037 1458 140103 1461
rect 139577 1456 140103 1458
rect 139577 1400 139582 1456
rect 139638 1400 140042 1456
rect 140098 1400 140103 1456
rect 139577 1398 140103 1400
rect 139577 1395 139643 1398
rect 140037 1395 140103 1398
rect 140221 1458 140287 1461
rect 141233 1458 141299 1461
rect 140221 1456 141299 1458
rect 140221 1400 140226 1456
rect 140282 1400 141238 1456
rect 141294 1400 141299 1456
rect 140221 1398 141299 1400
rect 140221 1395 140287 1398
rect 141233 1395 141299 1398
rect 136909 1324 136975 1325
rect 136909 1322 136956 1324
rect 136357 1320 136788 1322
rect 136357 1264 136362 1320
rect 136418 1264 136788 1320
rect 136357 1262 136788 1264
rect 136864 1320 136956 1322
rect 136864 1264 136914 1320
rect 136864 1262 136956 1264
rect 136357 1259 136423 1262
rect 136909 1260 136956 1262
rect 137020 1260 137026 1324
rect 137185 1322 137251 1325
rect 141182 1322 141188 1324
rect 137185 1320 141188 1322
rect 137185 1264 137190 1320
rect 137246 1264 141188 1320
rect 137185 1262 141188 1264
rect 136909 1259 136975 1260
rect 137185 1259 137251 1262
rect 141182 1260 141188 1262
rect 141252 1260 141258 1324
rect 141374 1322 141434 1534
rect 144862 1532 144868 1534
rect 144932 1532 144938 1596
rect 145005 1594 145071 1597
rect 145833 1594 145899 1597
rect 145005 1592 145899 1594
rect 145005 1536 145010 1592
rect 145066 1536 145838 1592
rect 145894 1536 145899 1592
rect 145005 1534 145899 1536
rect 145005 1531 145071 1534
rect 145833 1531 145899 1534
rect 145966 1532 145972 1596
rect 146036 1594 146042 1596
rect 147254 1594 147260 1596
rect 146036 1534 147260 1594
rect 146036 1532 146042 1534
rect 147254 1532 147260 1534
rect 147324 1532 147330 1596
rect 147397 1594 147463 1597
rect 147806 1594 147812 1596
rect 147397 1592 147812 1594
rect 147397 1536 147402 1592
rect 147458 1536 147812 1592
rect 147397 1534 147812 1536
rect 147397 1531 147463 1534
rect 147806 1532 147812 1534
rect 147876 1532 147882 1596
rect 148685 1594 148751 1597
rect 152782 1594 152842 1670
rect 154297 1667 154363 1670
rect 154430 1668 154436 1732
rect 154500 1730 154506 1732
rect 156086 1730 156092 1732
rect 154500 1670 156092 1730
rect 154500 1668 154506 1670
rect 156086 1668 156092 1670
rect 156156 1668 156162 1732
rect 158478 1668 158484 1732
rect 158548 1730 158554 1732
rect 158805 1730 158871 1733
rect 158548 1728 158871 1730
rect 158548 1672 158810 1728
rect 158866 1672 158871 1728
rect 158548 1670 158871 1672
rect 158548 1668 158554 1670
rect 158805 1667 158871 1670
rect 158989 1730 159055 1733
rect 166809 1730 166875 1733
rect 158989 1728 166875 1730
rect 158989 1672 158994 1728
rect 159050 1672 166814 1728
rect 166870 1672 166875 1728
rect 158989 1670 166875 1672
rect 158989 1667 159055 1670
rect 166809 1667 166875 1670
rect 166942 1668 166948 1732
rect 167012 1730 167018 1732
rect 168966 1730 168972 1732
rect 167012 1670 168972 1730
rect 167012 1668 167018 1670
rect 168966 1668 168972 1670
rect 169036 1668 169042 1732
rect 169109 1730 169175 1733
rect 169109 1728 169586 1730
rect 169109 1672 169114 1728
rect 169170 1672 169586 1728
rect 169109 1670 169586 1672
rect 169109 1667 169175 1670
rect 148685 1592 152842 1594
rect 148685 1536 148690 1592
rect 148746 1536 152842 1592
rect 148685 1534 152842 1536
rect 153929 1594 153995 1597
rect 153929 1592 157810 1594
rect 153929 1536 153934 1592
rect 153990 1536 157810 1592
rect 153929 1534 157810 1536
rect 148685 1531 148751 1534
rect 153929 1531 153995 1534
rect 141509 1458 141575 1461
rect 151537 1458 151603 1461
rect 141509 1456 151603 1458
rect 141509 1400 141514 1456
rect 141570 1400 151542 1456
rect 151598 1400 151603 1456
rect 141509 1398 151603 1400
rect 141509 1395 141575 1398
rect 151537 1395 151603 1398
rect 151813 1458 151879 1461
rect 157558 1458 157564 1460
rect 151813 1456 157564 1458
rect 151813 1400 151818 1456
rect 151874 1400 157564 1456
rect 151813 1398 157564 1400
rect 151813 1395 151879 1398
rect 157558 1396 157564 1398
rect 157628 1396 157634 1460
rect 147857 1322 147923 1325
rect 147990 1322 147996 1324
rect 141374 1262 147690 1322
rect 107142 1124 107148 1188
rect 107212 1186 107218 1188
rect 107377 1186 107443 1189
rect 107212 1184 107443 1186
rect 107212 1128 107382 1184
rect 107438 1128 107443 1184
rect 107212 1126 107443 1128
rect 107212 1124 107218 1126
rect 107377 1123 107443 1126
rect 107510 1124 107516 1188
rect 107580 1186 107586 1188
rect 110321 1186 110387 1189
rect 107580 1184 110387 1186
rect 107580 1128 110326 1184
rect 110382 1128 110387 1184
rect 107580 1126 110387 1128
rect 107580 1124 107586 1126
rect 110321 1123 110387 1126
rect 110505 1186 110571 1189
rect 111609 1188 111675 1189
rect 111374 1186 111380 1188
rect 110505 1184 111380 1186
rect 110505 1128 110510 1184
rect 110566 1128 111380 1184
rect 110505 1126 111380 1128
rect 110505 1123 110571 1126
rect 111374 1124 111380 1126
rect 111444 1124 111450 1188
rect 111558 1124 111564 1188
rect 111628 1186 111675 1188
rect 111628 1184 111720 1186
rect 111670 1128 111720 1184
rect 111628 1126 111720 1128
rect 111628 1124 111675 1126
rect 111788 1124 111794 1188
rect 111858 1186 111864 1188
rect 112478 1186 112484 1188
rect 111858 1126 112484 1186
rect 111858 1124 111864 1126
rect 112478 1124 112484 1126
rect 112548 1124 112554 1188
rect 112621 1186 112687 1189
rect 120206 1186 120212 1188
rect 112621 1184 120212 1186
rect 112621 1128 112626 1184
rect 112682 1128 120212 1184
rect 112621 1126 120212 1128
rect 111609 1123 111675 1124
rect 112621 1123 112687 1126
rect 120206 1124 120212 1126
rect 120276 1124 120282 1188
rect 120349 1186 120415 1189
rect 125358 1186 125364 1188
rect 120349 1184 125364 1186
rect 120349 1128 120354 1184
rect 120410 1128 125364 1184
rect 120349 1126 125364 1128
rect 120349 1123 120415 1126
rect 125358 1124 125364 1126
rect 125428 1124 125434 1188
rect 125501 1186 125567 1189
rect 126697 1186 126763 1189
rect 125501 1184 126763 1186
rect 125501 1128 125506 1184
rect 125562 1128 126702 1184
rect 126758 1128 126763 1184
rect 125501 1126 126763 1128
rect 125501 1123 125567 1126
rect 126697 1123 126763 1126
rect 126830 1124 126836 1188
rect 126900 1186 126906 1188
rect 128302 1186 128308 1188
rect 126900 1126 128308 1186
rect 126900 1124 126906 1126
rect 128302 1124 128308 1126
rect 128372 1124 128378 1188
rect 128445 1186 128511 1189
rect 135529 1186 135595 1189
rect 128445 1184 135595 1186
rect 128445 1128 128450 1184
rect 128506 1128 135534 1184
rect 135590 1128 135595 1184
rect 128445 1126 135595 1128
rect 128445 1123 128511 1126
rect 135529 1123 135595 1126
rect 135670 1126 139226 1186
rect 97257 1048 107026 1050
rect 97257 992 97262 1048
rect 97318 992 107026 1048
rect 97257 990 107026 992
rect 107101 1050 107167 1053
rect 109033 1050 109099 1053
rect 107101 1048 109099 1050
rect 107101 992 107106 1048
rect 107162 992 109038 1048
rect 109094 992 109099 1048
rect 107101 990 109099 992
rect 97257 987 97323 990
rect 107101 987 107167 990
rect 109033 987 109099 990
rect 109217 1050 109283 1053
rect 123569 1050 123635 1053
rect 123753 1052 123819 1053
rect 109217 1048 123635 1050
rect 109217 992 109222 1048
rect 109278 992 123574 1048
rect 123630 992 123635 1048
rect 109217 990 123635 992
rect 109217 987 109283 990
rect 123569 987 123635 990
rect 123702 988 123708 1052
rect 123772 1050 123819 1052
rect 123772 1048 123864 1050
rect 123814 992 123864 1048
rect 123772 990 123864 992
rect 123772 988 123819 990
rect 124070 988 124076 1052
rect 124140 1050 124146 1052
rect 128670 1050 128676 1052
rect 124140 990 128676 1050
rect 124140 988 124146 990
rect 128670 988 128676 990
rect 128740 988 128746 1052
rect 128813 1050 128879 1053
rect 128813 1048 129842 1050
rect 128813 992 128818 1048
rect 128874 992 129842 1048
rect 128813 990 129842 992
rect 123753 987 123819 988
rect 128813 987 128879 990
rect 1761 914 1827 917
rect 1761 912 10426 914
rect 1761 856 1766 912
rect 1822 856 10426 912
rect 1761 854 10426 856
rect 1761 851 1827 854
rect 657 778 723 781
rect 10225 778 10291 781
rect 657 776 10291 778
rect 657 720 662 776
rect 718 720 10230 776
rect 10286 720 10291 776
rect 657 718 10291 720
rect 10366 778 10426 854
rect 10542 852 10548 916
rect 10612 914 10618 916
rect 13629 914 13695 917
rect 10612 912 13695 914
rect 10612 856 13634 912
rect 13690 856 13695 912
rect 10612 854 13695 856
rect 10612 852 10618 854
rect 13629 851 13695 854
rect 14457 914 14523 917
rect 19190 914 19196 916
rect 14457 912 19196 914
rect 14457 856 14462 912
rect 14518 856 19196 912
rect 14457 854 19196 856
rect 14457 851 14523 854
rect 19190 852 19196 854
rect 19260 852 19266 916
rect 22093 914 22159 917
rect 27889 914 27955 917
rect 22093 912 27955 914
rect 22093 856 22098 912
rect 22154 856 27894 912
rect 27950 856 27955 912
rect 22093 854 27955 856
rect 22093 851 22159 854
rect 27889 851 27955 854
rect 28206 852 28212 916
rect 28276 914 28282 916
rect 34973 914 35039 917
rect 28276 912 35039 914
rect 28276 856 34978 912
rect 35034 856 35039 912
rect 28276 854 35039 856
rect 28276 852 28282 854
rect 34973 851 35039 854
rect 38561 914 38627 917
rect 47945 914 48011 917
rect 38561 912 48011 914
rect 38561 856 38566 912
rect 38622 856 47950 912
rect 48006 856 48011 912
rect 38561 854 48011 856
rect 38561 851 38627 854
rect 47945 851 48011 854
rect 48129 914 48195 917
rect 55949 914 56015 917
rect 82302 914 82308 916
rect 48129 912 55874 914
rect 48129 856 48134 912
rect 48190 856 55874 912
rect 48129 854 55874 856
rect 48129 851 48195 854
rect 23105 778 23171 781
rect 10366 776 23171 778
rect 10366 720 23110 776
rect 23166 720 23171 776
rect 10366 718 23171 720
rect 657 715 723 718
rect 10225 715 10291 718
rect 23105 715 23171 718
rect 24301 778 24367 781
rect 38193 778 38259 781
rect 24301 776 38259 778
rect 24301 720 24306 776
rect 24362 720 38198 776
rect 38254 720 38259 776
rect 24301 718 38259 720
rect 24301 715 24367 718
rect 38193 715 38259 718
rect 38377 778 38443 781
rect 46289 778 46355 781
rect 38377 776 46355 778
rect 38377 720 38382 776
rect 38438 720 46294 776
rect 46350 720 46355 776
rect 38377 718 46355 720
rect 38377 715 38443 718
rect 46289 715 46355 718
rect 46565 778 46631 781
rect 48957 778 49023 781
rect 46565 776 49023 778
rect 46565 720 46570 776
rect 46626 720 48962 776
rect 49018 720 49023 776
rect 46565 718 49023 720
rect 46565 715 46631 718
rect 48957 715 49023 718
rect 49509 778 49575 781
rect 55673 778 55739 781
rect 49509 776 55739 778
rect 49509 720 49514 776
rect 49570 720 55678 776
rect 55734 720 55739 776
rect 49509 718 55739 720
rect 55814 778 55874 854
rect 55949 912 82308 914
rect 55949 856 55954 912
rect 56010 856 82308 912
rect 55949 854 82308 856
rect 55949 851 56015 854
rect 82302 852 82308 854
rect 82372 852 82378 916
rect 82445 912 82554 917
rect 82445 856 82450 912
rect 82506 856 82554 912
rect 82445 854 82554 856
rect 82445 851 82511 854
rect 82670 852 82676 916
rect 82740 914 82746 916
rect 91318 914 91324 916
rect 82740 854 91324 914
rect 82740 852 82746 854
rect 91318 852 91324 854
rect 91388 852 91394 916
rect 91461 914 91527 917
rect 91686 914 91692 916
rect 91461 912 91692 914
rect 91461 856 91466 912
rect 91522 856 91692 912
rect 91461 854 91692 856
rect 91461 851 91527 854
rect 91686 852 91692 854
rect 91756 852 91762 916
rect 92105 914 92171 917
rect 91878 912 92171 914
rect 91878 856 92110 912
rect 92166 856 92171 912
rect 91878 854 92171 856
rect 91737 778 91803 781
rect 91878 780 91938 854
rect 92105 851 92171 854
rect 92238 852 92244 916
rect 92308 914 92314 916
rect 129590 914 129596 916
rect 92308 854 129596 914
rect 92308 852 92314 854
rect 129590 852 129596 854
rect 129660 852 129666 916
rect 55814 776 91803 778
rect 55814 720 91742 776
rect 91798 720 91803 776
rect 55814 718 91803 720
rect 49509 715 49575 718
rect 55673 715 55739 718
rect 91737 715 91803 718
rect 91870 716 91876 780
rect 91940 716 91946 780
rect 92013 778 92079 781
rect 102225 778 102291 781
rect 92013 776 102291 778
rect 92013 720 92018 776
rect 92074 720 102230 776
rect 102286 720 102291 776
rect 92013 718 102291 720
rect 92013 715 92079 718
rect 102225 715 102291 718
rect 102358 716 102364 780
rect 102428 778 102434 780
rect 102685 778 102751 781
rect 102428 776 102751 778
rect 102428 720 102690 776
rect 102746 720 102751 776
rect 102428 718 102751 720
rect 102428 716 102434 718
rect 102685 715 102751 718
rect 102910 716 102916 780
rect 102980 778 102986 780
rect 103789 778 103855 781
rect 102980 776 103855 778
rect 102980 720 103794 776
rect 103850 720 103855 776
rect 102980 718 103855 720
rect 102980 716 102986 718
rect 103789 715 103855 718
rect 103973 778 104039 781
rect 106958 778 106964 780
rect 103973 776 106964 778
rect 103973 720 103978 776
rect 104034 720 106964 776
rect 103973 718 106964 720
rect 103973 715 104039 718
rect 106958 716 106964 718
rect 107028 716 107034 780
rect 107377 778 107443 781
rect 107694 778 107700 780
rect 107377 776 107700 778
rect 107377 720 107382 776
rect 107438 720 107700 776
rect 107377 718 107700 720
rect 107377 715 107443 718
rect 107694 716 107700 718
rect 107764 716 107770 780
rect 107837 778 107903 781
rect 111558 778 111564 780
rect 107837 776 111564 778
rect 107837 720 107842 776
rect 107898 720 111564 776
rect 107837 718 111564 720
rect 107837 715 107903 718
rect 111558 716 111564 718
rect 111628 716 111634 780
rect 111742 716 111748 780
rect 111812 778 111818 780
rect 113725 778 113791 781
rect 116393 778 116459 781
rect 111812 776 113791 778
rect 111812 720 113730 776
rect 113786 720 113791 776
rect 111812 718 113791 720
rect 111812 716 111818 718
rect 113725 715 113791 718
rect 113958 776 116459 778
rect 113958 720 116398 776
rect 116454 720 116459 776
rect 113958 718 116459 720
rect 197 642 263 645
rect 4981 642 5047 645
rect 197 640 5047 642
rect 197 584 202 640
rect 258 584 4986 640
rect 5042 584 5047 640
rect 197 582 5047 584
rect 197 579 263 582
rect 4981 579 5047 582
rect 5625 642 5691 645
rect 13261 642 13327 645
rect 5625 640 13327 642
rect 5625 584 5630 640
rect 5686 584 13266 640
rect 13322 584 13327 640
rect 5625 582 13327 584
rect 5625 579 5691 582
rect 13261 579 13327 582
rect 13445 642 13511 645
rect 20713 642 20779 645
rect 13445 640 20779 642
rect 13445 584 13450 640
rect 13506 584 20718 640
rect 20774 584 20779 640
rect 13445 582 20779 584
rect 13445 579 13511 582
rect 20713 579 20779 582
rect 21909 642 21975 645
rect 111609 642 111675 645
rect 21909 640 102794 642
rect 21909 584 21914 640
rect 21970 584 102794 640
rect 21909 582 102794 584
rect 21909 579 21975 582
rect 381 506 447 509
rect 7373 506 7439 509
rect 33685 506 33751 509
rect 381 504 7439 506
rect 381 448 386 504
rect 442 448 7378 504
rect 7434 448 7439 504
rect 381 446 7439 448
rect 381 443 447 446
rect 7373 443 7439 446
rect 10918 504 33751 506
rect 10918 448 33690 504
rect 33746 448 33751 504
rect 10918 446 33751 448
rect 289 370 355 373
rect 422 370 428 372
rect 289 368 428 370
rect 289 312 294 368
rect 350 312 428 368
rect 289 310 428 312
rect 289 307 355 310
rect 422 308 428 310
rect 492 308 498 372
rect 1945 370 2011 373
rect 10685 370 10751 373
rect 1945 368 10751 370
rect 1945 312 1950 368
rect 2006 312 10690 368
rect 10746 312 10751 368
rect 1945 310 10751 312
rect 1945 307 2011 310
rect 10685 307 10751 310
rect 3417 234 3483 237
rect 10918 234 10978 446
rect 33685 443 33751 446
rect 35157 506 35223 509
rect 45553 506 45619 509
rect 35157 504 45619 506
rect 35157 448 35162 504
rect 35218 448 45558 504
rect 45614 448 45619 504
rect 35157 446 45619 448
rect 35157 443 35223 446
rect 45553 443 45619 446
rect 46657 506 46723 509
rect 49877 506 49943 509
rect 46657 504 49943 506
rect 46657 448 46662 504
rect 46718 448 49882 504
rect 49938 448 49943 504
rect 46657 446 49943 448
rect 46657 443 46723 446
rect 49877 443 49943 446
rect 50705 506 50771 509
rect 65333 506 65399 509
rect 68093 506 68159 509
rect 50705 504 65258 506
rect 50705 448 50710 504
rect 50766 448 65258 504
rect 50705 446 65258 448
rect 50705 443 50771 446
rect 12617 370 12683 373
rect 14641 370 14707 373
rect 12617 368 14707 370
rect 12617 312 12622 368
rect 12678 312 14646 368
rect 14702 312 14707 368
rect 12617 310 14707 312
rect 12617 307 12683 310
rect 14641 307 14707 310
rect 14958 308 14964 372
rect 15028 370 15034 372
rect 15837 370 15903 373
rect 15028 368 15903 370
rect 15028 312 15842 368
rect 15898 312 15903 368
rect 15028 310 15903 312
rect 15028 308 15034 310
rect 15837 307 15903 310
rect 19793 370 19859 373
rect 28349 370 28415 373
rect 19793 368 28415 370
rect 19793 312 19798 368
rect 19854 312 28354 368
rect 28410 312 28415 368
rect 19793 310 28415 312
rect 19793 307 19859 310
rect 28349 307 28415 310
rect 30465 370 30531 373
rect 65057 370 65123 373
rect 30465 368 65123 370
rect 30465 312 30470 368
rect 30526 312 65062 368
rect 65118 312 65123 368
rect 30465 310 65123 312
rect 30465 307 30531 310
rect 65057 307 65123 310
rect 3417 232 10978 234
rect 3417 176 3422 232
rect 3478 176 10978 232
rect 3417 174 10978 176
rect 13077 234 13143 237
rect 14549 234 14615 237
rect 13077 232 14615 234
rect 13077 176 13082 232
rect 13138 176 14554 232
rect 14610 176 14615 232
rect 13077 174 14615 176
rect 3417 171 3483 174
rect 13077 171 13143 174
rect 14549 171 14615 174
rect 15009 234 15075 237
rect 19333 234 19399 237
rect 15009 232 19399 234
rect 15009 176 15014 232
rect 15070 176 19338 232
rect 19394 176 19399 232
rect 15009 174 19399 176
rect 15009 171 15075 174
rect 19333 171 19399 174
rect 19701 234 19767 237
rect 49509 234 49575 237
rect 19701 232 49575 234
rect 19701 176 19706 232
rect 19762 176 49514 232
rect 49570 176 49575 232
rect 19701 174 49575 176
rect 19701 171 19767 174
rect 49509 171 49575 174
rect 51809 234 51875 237
rect 55949 234 56015 237
rect 51809 232 56015 234
rect 51809 176 51814 232
rect 51870 176 55954 232
rect 56010 176 56015 232
rect 51809 174 56015 176
rect 51809 171 51875 174
rect 55949 171 56015 174
rect 56133 234 56199 237
rect 57421 234 57487 237
rect 56133 232 57487 234
rect 56133 176 56138 232
rect 56194 176 57426 232
rect 57482 176 57487 232
rect 56133 174 57487 176
rect 56133 171 56199 174
rect 57421 171 57487 174
rect 57789 234 57855 237
rect 61142 234 61148 236
rect 57789 232 61148 234
rect 57789 176 57794 232
rect 57850 176 61148 232
rect 57789 174 61148 176
rect 57789 171 57855 174
rect 61142 172 61148 174
rect 61212 172 61218 236
rect 61377 234 61443 237
rect 64413 234 64479 237
rect 61377 232 64479 234
rect 61377 176 61382 232
rect 61438 176 64418 232
rect 64474 176 64479 232
rect 61377 174 64479 176
rect 65198 234 65258 446
rect 65333 504 68159 506
rect 65333 448 65338 504
rect 65394 448 68098 504
rect 68154 448 68159 504
rect 65333 446 68159 448
rect 65333 443 65399 446
rect 68093 443 68159 446
rect 68461 506 68527 509
rect 72601 506 72667 509
rect 68461 504 72667 506
rect 68461 448 68466 504
rect 68522 448 72606 504
rect 72662 448 72667 504
rect 68461 446 72667 448
rect 68461 443 68527 446
rect 72601 443 72667 446
rect 72785 506 72851 509
rect 74073 506 74139 509
rect 72785 504 74139 506
rect 72785 448 72790 504
rect 72846 448 74078 504
rect 74134 448 74139 504
rect 72785 446 74139 448
rect 72785 443 72851 446
rect 74073 443 74139 446
rect 74206 444 74212 508
rect 74276 506 74282 508
rect 75729 506 75795 509
rect 74276 504 75795 506
rect 74276 448 75734 504
rect 75790 448 75795 504
rect 74276 446 75795 448
rect 74276 444 74282 446
rect 75729 443 75795 446
rect 75913 506 75979 509
rect 76046 506 76052 508
rect 75913 504 76052 506
rect 75913 448 75918 504
rect 75974 448 76052 504
rect 75913 446 76052 448
rect 75913 443 75979 446
rect 76046 444 76052 446
rect 76116 444 76122 508
rect 76189 506 76255 509
rect 78489 506 78555 509
rect 76189 504 78555 506
rect 76189 448 76194 504
rect 76250 448 78494 504
rect 78550 448 78555 504
rect 76189 446 78555 448
rect 76189 443 76255 446
rect 78489 443 78555 446
rect 78622 444 78628 508
rect 78692 506 78698 508
rect 79225 506 79291 509
rect 78692 504 79291 506
rect 78692 448 79230 504
rect 79286 448 79291 504
rect 78692 446 79291 448
rect 78692 444 78698 446
rect 79225 443 79291 446
rect 79358 444 79364 508
rect 79428 506 79434 508
rect 80278 506 80284 508
rect 79428 446 80284 506
rect 79428 444 79434 446
rect 80278 444 80284 446
rect 80348 444 80354 508
rect 80421 506 80487 509
rect 102542 506 102548 508
rect 80421 504 102548 506
rect 80421 448 80426 504
rect 80482 448 102548 504
rect 80421 446 102548 448
rect 80421 443 80487 446
rect 102542 444 102548 446
rect 102612 444 102618 508
rect 102734 506 102794 582
rect 103102 640 111675 642
rect 103102 584 111614 640
rect 111670 584 111675 640
rect 103102 582 111675 584
rect 103102 506 103162 582
rect 111609 579 111675 582
rect 111793 642 111859 645
rect 112069 642 112135 645
rect 111793 640 112135 642
rect 111793 584 111798 640
rect 111854 584 112074 640
rect 112130 584 112135 640
rect 111793 582 112135 584
rect 111793 579 111859 582
rect 112069 579 112135 582
rect 112345 642 112411 645
rect 113958 642 114018 718
rect 116393 715 116459 718
rect 116577 778 116643 781
rect 122741 778 122807 781
rect 116577 776 122807 778
rect 116577 720 116582 776
rect 116638 720 122746 776
rect 122802 720 122807 776
rect 116577 718 122807 720
rect 116577 715 116643 718
rect 122741 715 122807 718
rect 122966 716 122972 780
rect 123036 778 123042 780
rect 129089 778 129155 781
rect 123036 776 129155 778
rect 123036 720 129094 776
rect 129150 720 129155 776
rect 123036 718 129155 720
rect 123036 716 123042 718
rect 129089 715 129155 718
rect 129222 716 129228 780
rect 129292 778 129298 780
rect 129641 778 129707 781
rect 129292 776 129707 778
rect 129292 720 129646 776
rect 129702 720 129707 776
rect 129292 718 129707 720
rect 129782 778 129842 990
rect 129958 988 129964 1052
rect 130028 1050 130034 1052
rect 131481 1050 131547 1053
rect 130028 1048 131547 1050
rect 130028 992 131486 1048
rect 131542 992 131547 1048
rect 130028 990 131547 992
rect 130028 988 130034 990
rect 131481 987 131547 990
rect 131665 1050 131731 1053
rect 135478 1050 135484 1052
rect 131665 1048 135484 1050
rect 131665 992 131670 1048
rect 131726 992 135484 1048
rect 131665 990 135484 992
rect 131665 987 131731 990
rect 135478 988 135484 990
rect 135548 988 135554 1052
rect 129958 852 129964 916
rect 130028 914 130034 916
rect 135670 914 135730 1126
rect 135805 1050 135871 1053
rect 139025 1050 139091 1053
rect 135805 1048 139091 1050
rect 135805 992 135810 1048
rect 135866 992 139030 1048
rect 139086 992 139091 1048
rect 135805 990 139091 992
rect 139166 1050 139226 1126
rect 139572 1124 139578 1188
rect 139642 1186 139648 1188
rect 139761 1186 139827 1189
rect 139642 1184 139827 1186
rect 139642 1128 139766 1184
rect 139822 1128 139827 1184
rect 139642 1126 139827 1128
rect 139642 1124 139648 1126
rect 139761 1123 139827 1126
rect 139894 1124 139900 1188
rect 139964 1186 139970 1188
rect 141182 1186 141188 1188
rect 139964 1126 141188 1186
rect 139964 1124 139970 1126
rect 141182 1124 141188 1126
rect 141252 1124 141258 1188
rect 141325 1186 141391 1189
rect 145281 1186 145347 1189
rect 141325 1184 145347 1186
rect 141325 1128 141330 1184
rect 141386 1128 145286 1184
rect 145342 1128 145347 1184
rect 141325 1126 145347 1128
rect 141325 1123 141391 1126
rect 145281 1123 145347 1126
rect 145465 1186 145531 1189
rect 147438 1186 147444 1188
rect 145465 1184 147444 1186
rect 145465 1128 145470 1184
rect 145526 1128 147444 1184
rect 145465 1126 147444 1128
rect 145465 1123 145531 1126
rect 147438 1124 147444 1126
rect 147508 1124 147514 1188
rect 147630 1186 147690 1262
rect 147857 1320 147996 1322
rect 147857 1264 147862 1320
rect 147918 1264 147996 1320
rect 147857 1262 147996 1264
rect 147857 1259 147923 1262
rect 147990 1260 147996 1262
rect 148060 1260 148066 1324
rect 148174 1260 148180 1324
rect 148244 1322 148250 1324
rect 148685 1322 148751 1325
rect 148244 1320 148751 1322
rect 148244 1264 148690 1320
rect 148746 1264 148751 1320
rect 148244 1262 148751 1264
rect 148244 1260 148250 1262
rect 148685 1259 148751 1262
rect 148869 1320 148935 1325
rect 148869 1264 148874 1320
rect 148930 1264 148935 1320
rect 148869 1259 148935 1264
rect 149053 1322 149119 1325
rect 151997 1322 152063 1325
rect 152365 1322 152431 1325
rect 149053 1320 151508 1322
rect 149053 1264 149058 1320
rect 149114 1264 151508 1320
rect 149053 1262 151508 1264
rect 149053 1259 149119 1262
rect 148593 1186 148659 1189
rect 147630 1184 148659 1186
rect 147630 1128 148598 1184
rect 148654 1128 148659 1184
rect 147630 1126 148659 1128
rect 148593 1123 148659 1126
rect 148726 1124 148732 1188
rect 148796 1186 148802 1188
rect 148872 1186 148932 1259
rect 148796 1126 148932 1186
rect 149237 1186 149303 1189
rect 150750 1186 150756 1188
rect 149237 1184 150756 1186
rect 149237 1128 149242 1184
rect 149298 1128 150756 1184
rect 149237 1126 150756 1128
rect 148796 1124 148802 1126
rect 149237 1123 149303 1126
rect 150750 1124 150756 1126
rect 150820 1124 150826 1188
rect 150893 1186 150959 1189
rect 151302 1186 151308 1188
rect 150893 1184 151308 1186
rect 150893 1128 150898 1184
rect 150954 1128 151308 1184
rect 150893 1126 151308 1128
rect 150893 1123 150959 1126
rect 151302 1124 151308 1126
rect 151372 1124 151378 1188
rect 151448 1186 151508 1262
rect 151997 1320 152431 1322
rect 151997 1264 152002 1320
rect 152058 1264 152370 1320
rect 152426 1264 152431 1320
rect 151997 1262 152431 1264
rect 151997 1259 152063 1262
rect 152365 1259 152431 1262
rect 152549 1322 152615 1325
rect 153878 1322 153884 1324
rect 152549 1320 153884 1322
rect 152549 1264 152554 1320
rect 152610 1264 153884 1320
rect 152549 1262 153884 1264
rect 152549 1259 152615 1262
rect 153878 1260 153884 1262
rect 153948 1260 153954 1324
rect 154113 1322 154179 1325
rect 157517 1322 157583 1325
rect 154113 1320 157583 1322
rect 154113 1264 154118 1320
rect 154174 1264 157522 1320
rect 157578 1264 157583 1320
rect 154113 1262 157583 1264
rect 157750 1322 157810 1534
rect 157926 1532 157932 1596
rect 157996 1594 158002 1596
rect 160134 1594 160140 1596
rect 157996 1534 160140 1594
rect 157996 1532 158002 1534
rect 160134 1532 160140 1534
rect 160204 1532 160210 1596
rect 160277 1594 160343 1597
rect 161054 1594 161060 1596
rect 160277 1592 161060 1594
rect 160277 1536 160282 1592
rect 160338 1536 161060 1592
rect 160277 1534 161060 1536
rect 160277 1531 160343 1534
rect 161054 1532 161060 1534
rect 161124 1532 161130 1596
rect 161197 1594 161263 1597
rect 169334 1594 169340 1596
rect 161197 1592 169340 1594
rect 161197 1536 161202 1592
rect 161258 1536 169340 1592
rect 161197 1534 169340 1536
rect 161197 1531 161263 1534
rect 169334 1532 169340 1534
rect 169404 1532 169410 1596
rect 169526 1594 169586 1670
rect 169886 1668 169892 1732
rect 169956 1730 169962 1732
rect 175774 1730 175780 1732
rect 169956 1670 175780 1730
rect 169956 1668 169962 1670
rect 175774 1668 175780 1670
rect 175844 1668 175850 1732
rect 175958 1668 175964 1732
rect 176028 1730 176034 1732
rect 178166 1730 178172 1732
rect 176028 1670 178172 1730
rect 176028 1668 176034 1670
rect 178166 1668 178172 1670
rect 178236 1668 178242 1732
rect 178769 1730 178835 1733
rect 178902 1730 178908 1732
rect 178769 1728 178908 1730
rect 178769 1672 178774 1728
rect 178830 1672 178908 1728
rect 178769 1670 178908 1672
rect 178769 1667 178835 1670
rect 178902 1668 178908 1670
rect 178972 1668 178978 1732
rect 179045 1730 179111 1733
rect 179045 1728 184858 1730
rect 179045 1672 179050 1728
rect 179106 1672 184858 1728
rect 179045 1670 184858 1672
rect 179045 1667 179111 1670
rect 171041 1594 171107 1597
rect 169526 1592 171107 1594
rect 169526 1536 171046 1592
rect 171102 1536 171107 1592
rect 169526 1534 171107 1536
rect 171041 1531 171107 1534
rect 171174 1532 171180 1596
rect 171244 1594 171250 1596
rect 171593 1594 171659 1597
rect 171244 1592 171659 1594
rect 171244 1536 171598 1592
rect 171654 1536 171659 1592
rect 171244 1534 171659 1536
rect 171244 1532 171250 1534
rect 171593 1531 171659 1534
rect 171726 1532 171732 1596
rect 171796 1594 171802 1596
rect 173014 1594 173020 1596
rect 171796 1534 173020 1594
rect 171796 1532 171802 1534
rect 173014 1532 173020 1534
rect 173084 1532 173090 1596
rect 177665 1594 177731 1597
rect 178166 1594 178172 1596
rect 173206 1592 177731 1594
rect 173206 1536 177670 1592
rect 177726 1536 177731 1592
rect 173206 1534 177731 1536
rect 157977 1460 158043 1461
rect 157926 1458 157932 1460
rect 157886 1398 157932 1458
rect 157996 1456 158043 1460
rect 158038 1400 158043 1456
rect 157926 1396 157932 1398
rect 157996 1396 158043 1400
rect 157977 1395 158043 1396
rect 158161 1458 158227 1461
rect 158989 1458 159055 1461
rect 158161 1456 159055 1458
rect 158161 1400 158166 1456
rect 158222 1400 158994 1456
rect 159050 1400 159055 1456
rect 158161 1398 159055 1400
rect 158161 1395 158227 1398
rect 158989 1395 159055 1398
rect 159398 1396 159404 1460
rect 159468 1458 159474 1460
rect 159633 1458 159699 1461
rect 159468 1456 159699 1458
rect 159468 1400 159638 1456
rect 159694 1400 159699 1456
rect 159468 1398 159699 1400
rect 159468 1396 159474 1398
rect 159633 1395 159699 1398
rect 159766 1396 159772 1460
rect 159836 1458 159842 1460
rect 161238 1458 161244 1460
rect 159836 1398 161244 1458
rect 159836 1396 159842 1398
rect 161238 1396 161244 1398
rect 161308 1396 161314 1460
rect 161606 1396 161612 1460
rect 161676 1458 161682 1460
rect 163998 1458 164004 1460
rect 161676 1398 164004 1458
rect 161676 1396 161682 1398
rect 163998 1396 164004 1398
rect 164068 1396 164074 1460
rect 164233 1458 164299 1461
rect 169017 1458 169083 1461
rect 164233 1456 169083 1458
rect 164233 1400 164238 1456
rect 164294 1400 169022 1456
rect 169078 1400 169083 1456
rect 164233 1398 169083 1400
rect 164233 1395 164299 1398
rect 169017 1395 169083 1398
rect 169201 1458 169267 1461
rect 173206 1458 173266 1534
rect 177665 1531 177731 1534
rect 177806 1534 178172 1594
rect 169201 1456 173266 1458
rect 169201 1400 169206 1456
rect 169262 1400 173266 1456
rect 169201 1398 173266 1400
rect 173341 1458 173407 1461
rect 176878 1458 176884 1460
rect 173341 1456 176884 1458
rect 173341 1400 173346 1456
rect 173402 1400 176884 1456
rect 173341 1398 176884 1400
rect 169201 1395 169267 1398
rect 173341 1395 173407 1398
rect 176878 1396 176884 1398
rect 176948 1396 176954 1460
rect 177062 1396 177068 1460
rect 177132 1458 177138 1460
rect 177806 1458 177866 1534
rect 178166 1532 178172 1534
rect 178236 1532 178242 1596
rect 178350 1532 178356 1596
rect 178420 1594 178426 1596
rect 179638 1594 179644 1596
rect 178420 1534 179644 1594
rect 178420 1532 178426 1534
rect 179638 1532 179644 1534
rect 179708 1532 179714 1596
rect 179873 1594 179939 1597
rect 181713 1594 181779 1597
rect 179873 1592 181779 1594
rect 179873 1536 179878 1592
rect 179934 1536 181718 1592
rect 181774 1536 181779 1592
rect 179873 1534 181779 1536
rect 179873 1531 179939 1534
rect 181713 1531 181779 1534
rect 181846 1532 181852 1596
rect 181916 1594 181922 1596
rect 181916 1534 183984 1594
rect 181916 1532 181922 1534
rect 177132 1398 177866 1458
rect 177132 1396 177138 1398
rect 177982 1396 177988 1460
rect 178052 1458 178058 1460
rect 178309 1458 178375 1461
rect 178052 1456 178375 1458
rect 178052 1400 178314 1456
rect 178370 1400 178375 1456
rect 178052 1398 178375 1400
rect 178052 1396 178058 1398
rect 178309 1395 178375 1398
rect 178677 1458 178743 1461
rect 183737 1458 183803 1461
rect 178677 1456 183803 1458
rect 178677 1400 178682 1456
rect 178738 1400 183742 1456
rect 183798 1400 183803 1456
rect 178677 1398 183803 1400
rect 178677 1395 178743 1398
rect 183737 1395 183803 1398
rect 159357 1322 159423 1325
rect 157750 1320 159423 1322
rect 157750 1264 159362 1320
rect 159418 1264 159423 1320
rect 157750 1262 159423 1264
rect 154113 1259 154179 1262
rect 157517 1259 157583 1262
rect 159357 1259 159423 1262
rect 159541 1322 159607 1325
rect 161841 1322 161907 1325
rect 159541 1320 161907 1322
rect 159541 1264 159546 1320
rect 159602 1264 161846 1320
rect 161902 1264 161907 1320
rect 159541 1262 161907 1264
rect 159541 1259 159607 1262
rect 161841 1259 161907 1262
rect 161974 1260 161980 1324
rect 162044 1322 162050 1324
rect 163446 1322 163452 1324
rect 162044 1262 163452 1322
rect 162044 1260 162050 1262
rect 163446 1260 163452 1262
rect 163516 1260 163522 1324
rect 163773 1322 163839 1325
rect 168925 1322 168991 1325
rect 163773 1320 168991 1322
rect 163773 1264 163778 1320
rect 163834 1264 168930 1320
rect 168986 1264 168991 1320
rect 163773 1262 168991 1264
rect 163773 1259 163839 1262
rect 168925 1259 168991 1262
rect 169109 1322 169175 1325
rect 169886 1322 169892 1324
rect 169109 1320 169892 1322
rect 169109 1264 169114 1320
rect 169170 1264 169892 1320
rect 169109 1262 169892 1264
rect 169109 1259 169175 1262
rect 169886 1260 169892 1262
rect 169956 1260 169962 1324
rect 170070 1260 170076 1324
rect 170140 1322 170146 1324
rect 170765 1322 170831 1325
rect 173801 1322 173867 1325
rect 170140 1262 170690 1322
rect 170140 1260 170146 1262
rect 157885 1186 157951 1189
rect 151448 1184 157951 1186
rect 151448 1128 157890 1184
rect 157946 1128 157951 1184
rect 151448 1126 157951 1128
rect 157885 1123 157951 1126
rect 158069 1186 158135 1189
rect 158437 1186 158503 1189
rect 158069 1184 158503 1186
rect 158069 1128 158074 1184
rect 158130 1128 158442 1184
rect 158498 1128 158503 1184
rect 158069 1126 158503 1128
rect 158069 1123 158135 1126
rect 158437 1123 158503 1126
rect 158621 1186 158687 1189
rect 159265 1186 159331 1189
rect 158621 1184 159331 1186
rect 158621 1128 158626 1184
rect 158682 1128 159270 1184
rect 159326 1128 159331 1184
rect 158621 1126 159331 1128
rect 158621 1123 158687 1126
rect 159265 1123 159331 1126
rect 159449 1186 159515 1189
rect 166206 1186 166212 1188
rect 159449 1184 166212 1186
rect 159449 1128 159454 1184
rect 159510 1128 166212 1184
rect 159449 1126 166212 1128
rect 159449 1123 159515 1126
rect 166206 1124 166212 1126
rect 166276 1124 166282 1188
rect 166349 1186 166415 1189
rect 168649 1186 168715 1189
rect 166349 1184 168715 1186
rect 166349 1128 166354 1184
rect 166410 1128 168654 1184
rect 168710 1128 168715 1184
rect 166349 1126 168715 1128
rect 166349 1123 166415 1126
rect 168649 1123 168715 1126
rect 168782 1124 168788 1188
rect 168852 1186 168858 1188
rect 169385 1186 169451 1189
rect 168852 1184 169451 1186
rect 168852 1128 169390 1184
rect 169446 1128 169451 1184
rect 168852 1126 169451 1128
rect 168852 1124 168858 1126
rect 169385 1123 169451 1126
rect 169569 1186 169635 1189
rect 170489 1186 170555 1189
rect 169569 1184 170555 1186
rect 169569 1128 169574 1184
rect 169630 1128 170494 1184
rect 170550 1128 170555 1184
rect 169569 1126 170555 1128
rect 170630 1186 170690 1262
rect 170765 1320 173867 1322
rect 170765 1264 170770 1320
rect 170826 1264 173806 1320
rect 173862 1264 173867 1320
rect 170765 1262 173867 1264
rect 170765 1259 170831 1262
rect 173801 1259 173867 1262
rect 173934 1260 173940 1324
rect 174004 1322 174010 1324
rect 175958 1322 175964 1324
rect 174004 1262 175964 1322
rect 174004 1260 174010 1262
rect 175958 1260 175964 1262
rect 176028 1260 176034 1324
rect 176326 1260 176332 1324
rect 176396 1322 176402 1324
rect 177757 1322 177823 1325
rect 176396 1320 177823 1322
rect 176396 1264 177762 1320
rect 177818 1264 177823 1320
rect 176396 1262 177823 1264
rect 176396 1260 176402 1262
rect 177757 1259 177823 1262
rect 178033 1322 178099 1325
rect 179454 1322 179460 1324
rect 178033 1320 179460 1322
rect 178033 1264 178038 1320
rect 178094 1264 179460 1320
rect 178033 1262 179460 1264
rect 178033 1259 178099 1262
rect 179454 1260 179460 1262
rect 179524 1260 179530 1324
rect 179689 1322 179755 1325
rect 180241 1322 180307 1325
rect 179689 1320 180307 1322
rect 179689 1264 179694 1320
rect 179750 1264 180246 1320
rect 180302 1264 180307 1320
rect 179689 1262 180307 1264
rect 179689 1259 179755 1262
rect 180241 1259 180307 1262
rect 180374 1260 180380 1324
rect 180444 1322 180450 1324
rect 182633 1322 182699 1325
rect 183686 1322 183692 1324
rect 180444 1320 182699 1322
rect 180444 1264 182638 1320
rect 182694 1264 182699 1320
rect 180444 1262 182699 1264
rect 180444 1260 180450 1262
rect 182633 1259 182699 1262
rect 182774 1262 183692 1322
rect 173249 1186 173315 1189
rect 170630 1184 173315 1186
rect 170630 1128 173254 1184
rect 173310 1128 173315 1184
rect 170630 1126 173315 1128
rect 169569 1123 169635 1126
rect 170489 1123 170555 1126
rect 173249 1123 173315 1126
rect 173382 1124 173388 1188
rect 173452 1186 173458 1188
rect 176142 1186 176148 1188
rect 173452 1126 176148 1186
rect 173452 1124 173458 1126
rect 176142 1124 176148 1126
rect 176212 1124 176218 1188
rect 176285 1186 176351 1189
rect 177113 1186 177179 1189
rect 176285 1184 177179 1186
rect 176285 1128 176290 1184
rect 176346 1128 177118 1184
rect 177174 1128 177179 1184
rect 176285 1126 177179 1128
rect 176285 1123 176351 1126
rect 177113 1123 177179 1126
rect 177665 1186 177731 1189
rect 179137 1186 179203 1189
rect 177665 1184 179203 1186
rect 177665 1128 177670 1184
rect 177726 1128 179142 1184
rect 179198 1128 179203 1184
rect 177665 1126 179203 1128
rect 177665 1123 177731 1126
rect 179137 1123 179203 1126
rect 179321 1186 179387 1189
rect 180793 1186 180859 1189
rect 179321 1184 180859 1186
rect 179321 1128 179326 1184
rect 179382 1128 180798 1184
rect 180854 1128 180859 1184
rect 179321 1126 180859 1128
rect 179321 1123 179387 1126
rect 180793 1123 180859 1126
rect 180926 1124 180932 1188
rect 180996 1186 181002 1188
rect 182774 1186 182834 1262
rect 183686 1260 183692 1262
rect 183756 1260 183762 1324
rect 183924 1322 183984 1534
rect 184054 1532 184060 1596
rect 184124 1594 184130 1596
rect 184657 1594 184723 1597
rect 184124 1592 184723 1594
rect 184124 1536 184662 1592
rect 184718 1536 184723 1592
rect 184124 1534 184723 1536
rect 184798 1594 184858 1670
rect 184974 1668 184980 1732
rect 185044 1730 185050 1732
rect 190637 1730 190703 1733
rect 185044 1728 190703 1730
rect 185044 1672 190642 1728
rect 190698 1672 190703 1728
rect 185044 1670 190703 1672
rect 185044 1668 185050 1670
rect 190637 1667 190703 1670
rect 190913 1730 190979 1733
rect 192201 1730 192267 1733
rect 190913 1728 192267 1730
rect 190913 1672 190918 1728
rect 190974 1672 192206 1728
rect 192262 1672 192267 1728
rect 190913 1670 192267 1672
rect 190913 1667 190979 1670
rect 192201 1667 192267 1670
rect 192334 1668 192340 1732
rect 192404 1730 192410 1732
rect 194726 1730 194732 1732
rect 192404 1670 194732 1730
rect 192404 1668 192410 1670
rect 194726 1668 194732 1670
rect 194796 1668 194802 1732
rect 194910 1668 194916 1732
rect 194980 1730 194986 1732
rect 196433 1730 196499 1733
rect 194980 1728 196499 1730
rect 194980 1672 196438 1728
rect 196494 1672 196499 1728
rect 194980 1670 196499 1672
rect 194980 1668 194986 1670
rect 196433 1667 196499 1670
rect 196709 1730 196775 1733
rect 198733 1730 198799 1733
rect 200021 1730 200087 1733
rect 207289 1730 207355 1733
rect 207974 1730 207980 1732
rect 196709 1728 198612 1730
rect 196709 1672 196714 1728
rect 196770 1672 198612 1728
rect 196709 1670 198612 1672
rect 196709 1667 196775 1670
rect 190494 1594 190500 1596
rect 184798 1534 190500 1594
rect 184124 1532 184130 1534
rect 184657 1531 184723 1534
rect 190494 1532 190500 1534
rect 190564 1532 190570 1596
rect 190637 1594 190703 1597
rect 195830 1594 195836 1596
rect 190637 1592 195836 1594
rect 190637 1536 190642 1592
rect 190698 1536 195836 1592
rect 190637 1534 195836 1536
rect 190637 1531 190703 1534
rect 195830 1532 195836 1534
rect 195900 1532 195906 1596
rect 195973 1594 196039 1597
rect 197118 1594 197124 1596
rect 195973 1592 197124 1594
rect 195973 1536 195978 1592
rect 196034 1536 197124 1592
rect 195973 1534 197124 1536
rect 195973 1531 196039 1534
rect 197118 1532 197124 1534
rect 197188 1532 197194 1596
rect 198406 1594 198412 1596
rect 197310 1534 198412 1594
rect 184381 1458 184447 1461
rect 190913 1458 190979 1461
rect 184381 1456 190979 1458
rect 184381 1400 184386 1456
rect 184442 1400 190918 1456
rect 190974 1400 190979 1456
rect 184381 1398 190979 1400
rect 184381 1395 184447 1398
rect 190913 1395 190979 1398
rect 191046 1396 191052 1460
rect 191116 1458 191122 1460
rect 197310 1458 197370 1534
rect 198406 1532 198412 1534
rect 198476 1532 198482 1596
rect 198552 1594 198612 1670
rect 198733 1728 199946 1730
rect 198733 1672 198738 1728
rect 198794 1672 199946 1728
rect 198733 1670 199946 1672
rect 198733 1667 198799 1670
rect 199101 1594 199167 1597
rect 199745 1594 199811 1597
rect 198552 1534 199026 1594
rect 191116 1398 197370 1458
rect 191116 1396 191122 1398
rect 197486 1396 197492 1460
rect 197556 1458 197562 1460
rect 198774 1458 198780 1460
rect 197556 1398 198780 1458
rect 197556 1396 197562 1398
rect 198774 1396 198780 1398
rect 198844 1396 198850 1460
rect 198966 1458 199026 1534
rect 199101 1592 199811 1594
rect 199101 1536 199106 1592
rect 199162 1536 199750 1592
rect 199806 1536 199811 1592
rect 199101 1534 199811 1536
rect 199886 1594 199946 1670
rect 200021 1728 207355 1730
rect 200021 1672 200026 1728
rect 200082 1672 207294 1728
rect 207350 1672 207355 1728
rect 200021 1670 207355 1672
rect 200021 1667 200087 1670
rect 207289 1667 207355 1670
rect 207476 1670 207980 1730
rect 207476 1597 207536 1670
rect 207974 1668 207980 1670
rect 208044 1668 208050 1732
rect 208117 1730 208183 1733
rect 216673 1730 216739 1733
rect 208117 1728 216739 1730
rect 208117 1672 208122 1728
rect 208178 1672 216678 1728
rect 216734 1672 216739 1728
rect 208117 1670 216739 1672
rect 208117 1667 208183 1670
rect 216673 1667 216739 1670
rect 216806 1668 216812 1732
rect 216876 1730 216882 1732
rect 220302 1730 220308 1732
rect 216876 1670 220308 1730
rect 216876 1668 216882 1670
rect 220302 1668 220308 1670
rect 220372 1668 220378 1732
rect 220445 1730 220511 1733
rect 232129 1730 232195 1733
rect 234061 1730 234127 1733
rect 220445 1728 231962 1730
rect 220445 1672 220450 1728
rect 220506 1672 231962 1728
rect 220445 1670 231962 1672
rect 220445 1667 220511 1670
rect 200982 1594 200988 1596
rect 199886 1534 200988 1594
rect 199101 1531 199167 1534
rect 199745 1531 199811 1534
rect 200982 1532 200988 1534
rect 201052 1532 201058 1596
rect 203190 1532 203196 1596
rect 203260 1594 203266 1596
rect 204294 1594 204300 1596
rect 203260 1534 204300 1594
rect 203260 1532 203266 1534
rect 204294 1532 204300 1534
rect 204364 1532 204370 1596
rect 204437 1594 204503 1597
rect 204805 1596 204871 1597
rect 204662 1594 204668 1596
rect 204437 1592 204668 1594
rect 204437 1536 204442 1592
rect 204498 1536 204668 1592
rect 204437 1534 204668 1536
rect 204437 1531 204503 1534
rect 204662 1532 204668 1534
rect 204732 1532 204738 1596
rect 204805 1592 204852 1596
rect 204916 1594 204922 1596
rect 205449 1594 205515 1597
rect 207289 1594 207355 1597
rect 204805 1536 204810 1592
rect 204805 1532 204852 1536
rect 204916 1534 204962 1594
rect 205449 1592 207355 1594
rect 205449 1536 205454 1592
rect 205510 1536 207294 1592
rect 207350 1536 207355 1592
rect 205449 1534 207355 1536
rect 204916 1532 204922 1534
rect 204805 1531 204871 1532
rect 205449 1531 205515 1534
rect 207289 1531 207355 1534
rect 207473 1592 207539 1597
rect 207473 1536 207478 1592
rect 207534 1536 207539 1592
rect 207473 1531 207539 1536
rect 207614 1534 210066 1594
rect 200297 1458 200363 1461
rect 198966 1456 200363 1458
rect 198966 1400 200302 1456
rect 200358 1400 200363 1456
rect 198966 1398 200363 1400
rect 200297 1395 200363 1398
rect 200430 1396 200436 1460
rect 200500 1458 200506 1460
rect 207614 1458 207674 1534
rect 200500 1398 207674 1458
rect 207749 1458 207815 1461
rect 207749 1456 208226 1458
rect 207749 1400 207754 1456
rect 207810 1400 208226 1456
rect 207749 1398 208226 1400
rect 200500 1396 200506 1398
rect 207749 1395 207815 1398
rect 189625 1322 189691 1325
rect 183924 1320 189691 1322
rect 183924 1264 189630 1320
rect 189686 1264 189691 1320
rect 183924 1262 189691 1264
rect 189625 1259 189691 1262
rect 189758 1260 189764 1324
rect 189828 1322 189834 1324
rect 191097 1322 191163 1325
rect 189828 1320 191163 1322
rect 189828 1264 191102 1320
rect 191158 1264 191163 1320
rect 189828 1262 191163 1264
rect 189828 1260 189834 1262
rect 191097 1259 191163 1262
rect 191230 1260 191236 1324
rect 191300 1322 191306 1324
rect 208025 1322 208091 1325
rect 191300 1320 208091 1322
rect 191300 1264 208030 1320
rect 208086 1264 208091 1320
rect 191300 1262 208091 1264
rect 208166 1322 208226 1398
rect 208342 1396 208348 1460
rect 208412 1458 208418 1460
rect 209814 1458 209820 1460
rect 208412 1398 209820 1458
rect 208412 1396 208418 1398
rect 209814 1396 209820 1398
rect 209884 1396 209890 1460
rect 210006 1458 210066 1534
rect 210182 1532 210188 1596
rect 210252 1594 210258 1596
rect 211337 1594 211403 1597
rect 210252 1534 211170 1594
rect 210252 1532 210258 1534
rect 210918 1458 210924 1460
rect 210006 1398 210924 1458
rect 210918 1396 210924 1398
rect 210988 1396 210994 1460
rect 211110 1458 211170 1534
rect 211337 1592 224740 1594
rect 211337 1536 211342 1592
rect 211398 1536 224740 1592
rect 211337 1534 224740 1536
rect 211337 1531 211403 1534
rect 212022 1458 212028 1460
rect 211110 1398 212028 1458
rect 212022 1396 212028 1398
rect 212092 1396 212098 1460
rect 212165 1458 212231 1461
rect 214373 1458 214439 1461
rect 216765 1458 216831 1461
rect 212165 1456 214439 1458
rect 212165 1400 212170 1456
rect 212226 1400 214378 1456
rect 214434 1400 214439 1456
rect 212165 1398 214439 1400
rect 212165 1395 212231 1398
rect 214373 1395 214439 1398
rect 214606 1456 216831 1458
rect 214606 1400 216770 1456
rect 216826 1400 216831 1456
rect 214606 1398 216831 1400
rect 209865 1322 209931 1325
rect 208166 1320 209931 1322
rect 208166 1264 209870 1320
rect 209926 1264 209931 1320
rect 208166 1262 209931 1264
rect 191300 1260 191306 1262
rect 208025 1259 208091 1262
rect 209865 1259 209931 1262
rect 209998 1260 210004 1324
rect 210068 1322 210074 1324
rect 214606 1322 214666 1398
rect 216765 1395 216831 1398
rect 216949 1458 217015 1461
rect 218145 1458 218211 1461
rect 216949 1456 218211 1458
rect 216949 1400 216954 1456
rect 217010 1400 218150 1456
rect 218206 1400 218211 1456
rect 216949 1398 218211 1400
rect 216949 1395 217015 1398
rect 218145 1395 218211 1398
rect 218278 1396 218284 1460
rect 218348 1458 218354 1460
rect 223941 1458 224007 1461
rect 224493 1460 224559 1461
rect 224493 1458 224540 1460
rect 218348 1456 224007 1458
rect 218348 1400 223946 1456
rect 224002 1400 224007 1456
rect 218348 1398 224007 1400
rect 224448 1456 224540 1458
rect 224448 1400 224498 1456
rect 224448 1398 224540 1400
rect 218348 1396 218354 1398
rect 223941 1395 224007 1398
rect 224493 1396 224540 1398
rect 224604 1396 224610 1460
rect 224680 1458 224740 1534
rect 224902 1532 224908 1596
rect 224972 1594 224978 1596
rect 225689 1594 225755 1597
rect 224972 1592 225755 1594
rect 224972 1536 225694 1592
rect 225750 1536 225755 1592
rect 224972 1534 225755 1536
rect 224972 1532 224978 1534
rect 225689 1531 225755 1534
rect 225873 1594 225939 1597
rect 231761 1594 231827 1597
rect 225873 1592 231827 1594
rect 225873 1536 225878 1592
rect 225934 1536 231766 1592
rect 231822 1536 231827 1592
rect 225873 1534 231827 1536
rect 231902 1594 231962 1670
rect 232129 1728 234127 1730
rect 232129 1672 232134 1728
rect 232190 1672 234066 1728
rect 234122 1672 234127 1728
rect 232129 1670 234127 1672
rect 232129 1667 232195 1670
rect 234061 1667 234127 1670
rect 234286 1668 234292 1732
rect 234356 1730 234362 1732
rect 237966 1730 237972 1732
rect 234356 1670 237972 1730
rect 234356 1668 234362 1670
rect 237966 1668 237972 1670
rect 238036 1668 238042 1732
rect 238385 1730 238451 1733
rect 245326 1730 245332 1732
rect 238158 1728 238451 1730
rect 238158 1672 238390 1728
rect 238446 1672 238451 1728
rect 238158 1670 238451 1672
rect 238158 1594 238218 1670
rect 238385 1667 238451 1670
rect 238526 1670 245332 1730
rect 231902 1534 238218 1594
rect 225873 1531 225939 1534
rect 231761 1531 231827 1534
rect 225413 1458 225479 1461
rect 238526 1458 238586 1670
rect 245326 1668 245332 1670
rect 245396 1668 245402 1732
rect 245469 1730 245535 1733
rect 247534 1730 247540 1732
rect 245469 1728 247540 1730
rect 245469 1672 245474 1728
rect 245530 1672 247540 1728
rect 245469 1670 247540 1672
rect 245469 1667 245535 1670
rect 247534 1668 247540 1670
rect 247604 1668 247610 1732
rect 247677 1730 247743 1733
rect 250069 1730 250135 1733
rect 258073 1730 258139 1733
rect 261702 1730 261708 1732
rect 247677 1728 249994 1730
rect 247677 1672 247682 1728
rect 247738 1672 249994 1728
rect 247677 1670 249994 1672
rect 247677 1667 247743 1670
rect 238702 1532 238708 1596
rect 238772 1594 238778 1596
rect 238937 1594 239003 1597
rect 238772 1592 239003 1594
rect 238772 1536 238942 1592
rect 238998 1536 239003 1592
rect 238772 1534 239003 1536
rect 238772 1532 238778 1534
rect 238937 1531 239003 1534
rect 239070 1532 239076 1596
rect 239140 1594 239146 1596
rect 241830 1594 241836 1596
rect 239140 1534 241836 1594
rect 239140 1532 239146 1534
rect 241830 1532 241836 1534
rect 241900 1532 241906 1596
rect 242065 1594 242131 1597
rect 249742 1594 249748 1596
rect 242065 1592 249748 1594
rect 242065 1536 242070 1592
rect 242126 1536 249748 1592
rect 242065 1534 249748 1536
rect 242065 1531 242131 1534
rect 249742 1532 249748 1534
rect 249812 1532 249818 1596
rect 249934 1594 249994 1670
rect 250069 1728 258139 1730
rect 250069 1672 250074 1728
rect 250130 1672 258078 1728
rect 258134 1672 258139 1728
rect 250069 1670 258139 1672
rect 250069 1667 250135 1670
rect 258073 1667 258139 1670
rect 258214 1670 261708 1730
rect 249934 1534 253122 1594
rect 224680 1456 225479 1458
rect 224680 1400 225418 1456
rect 225474 1400 225479 1456
rect 224680 1398 225479 1400
rect 224493 1395 224559 1396
rect 225413 1395 225479 1398
rect 225646 1398 238586 1458
rect 238661 1458 238727 1461
rect 242893 1458 242959 1461
rect 238661 1456 242959 1458
rect 238661 1400 238666 1456
rect 238722 1400 242898 1456
rect 242954 1400 242959 1456
rect 238661 1398 242959 1400
rect 214833 1324 214899 1325
rect 214782 1322 214788 1324
rect 210068 1262 214666 1322
rect 214742 1262 214788 1322
rect 214852 1320 214899 1324
rect 214894 1264 214899 1320
rect 210068 1260 210074 1262
rect 214782 1260 214788 1262
rect 214852 1260 214899 1264
rect 214833 1259 214899 1260
rect 215017 1322 215083 1325
rect 217409 1322 217475 1325
rect 215017 1320 217475 1322
rect 215017 1264 215022 1320
rect 215078 1264 217414 1320
rect 217470 1264 217475 1320
rect 215017 1262 217475 1264
rect 215017 1259 215083 1262
rect 217409 1259 217475 1262
rect 217542 1260 217548 1324
rect 217612 1322 217618 1324
rect 217961 1322 218027 1325
rect 217612 1320 218027 1322
rect 217612 1264 217966 1320
rect 218022 1264 218027 1320
rect 217612 1262 218027 1264
rect 217612 1260 217618 1262
rect 217961 1259 218027 1262
rect 221641 1322 221707 1325
rect 225045 1322 225111 1325
rect 221641 1320 225111 1322
rect 221641 1264 221646 1320
rect 221702 1264 225050 1320
rect 225106 1264 225111 1320
rect 221641 1262 225111 1264
rect 221641 1259 221707 1262
rect 225045 1259 225111 1262
rect 225229 1322 225295 1325
rect 225646 1322 225706 1398
rect 238661 1395 238727 1398
rect 242893 1395 242959 1398
rect 243118 1396 243124 1460
rect 243188 1458 243194 1460
rect 245142 1458 245148 1460
rect 243188 1398 245148 1458
rect 243188 1396 243194 1398
rect 245142 1396 245148 1398
rect 245212 1396 245218 1460
rect 245285 1458 245351 1461
rect 246614 1458 246620 1460
rect 245285 1456 246620 1458
rect 245285 1400 245290 1456
rect 245346 1400 246620 1456
rect 245285 1398 246620 1400
rect 245285 1395 245351 1398
rect 246614 1396 246620 1398
rect 246684 1396 246690 1460
rect 246798 1396 246804 1460
rect 246868 1458 246874 1460
rect 248822 1458 248828 1460
rect 246868 1398 248828 1458
rect 246868 1396 246874 1398
rect 248822 1396 248828 1398
rect 248892 1396 248898 1460
rect 248965 1458 249031 1461
rect 249977 1458 250043 1461
rect 248965 1456 250043 1458
rect 248965 1400 248970 1456
rect 249026 1400 249982 1456
rect 250038 1400 250043 1456
rect 248965 1398 250043 1400
rect 248965 1395 249031 1398
rect 249977 1395 250043 1398
rect 250110 1396 250116 1460
rect 250180 1458 250186 1460
rect 251541 1458 251607 1461
rect 253062 1458 253122 1534
rect 253238 1532 253244 1596
rect 253308 1594 253314 1596
rect 253308 1534 253674 1594
rect 253308 1532 253314 1534
rect 253422 1458 253428 1460
rect 250180 1398 251466 1458
rect 250180 1396 250186 1398
rect 225229 1320 225706 1322
rect 225229 1264 225234 1320
rect 225290 1264 225706 1320
rect 225229 1262 225706 1264
rect 225781 1322 225847 1325
rect 227437 1324 227503 1325
rect 227110 1322 227116 1324
rect 225781 1320 227116 1322
rect 225781 1264 225786 1320
rect 225842 1264 227116 1320
rect 225781 1262 227116 1264
rect 225229 1259 225295 1262
rect 225781 1259 225847 1262
rect 227110 1260 227116 1262
rect 227180 1260 227186 1324
rect 227437 1322 227484 1324
rect 227392 1320 227484 1322
rect 227392 1264 227442 1320
rect 227392 1262 227484 1264
rect 227437 1260 227484 1262
rect 227548 1260 227554 1324
rect 227662 1260 227668 1324
rect 227732 1322 227738 1324
rect 229134 1322 229140 1324
rect 227732 1262 229140 1322
rect 227732 1260 227738 1262
rect 229134 1260 229140 1262
rect 229204 1260 229210 1324
rect 229318 1260 229324 1324
rect 229388 1322 229394 1324
rect 232129 1322 232195 1325
rect 229388 1320 232195 1322
rect 229388 1264 232134 1320
rect 232190 1264 232195 1320
rect 229388 1262 232195 1264
rect 229388 1260 229394 1262
rect 227437 1259 227503 1260
rect 232129 1259 232195 1262
rect 232497 1322 232563 1325
rect 238017 1322 238083 1325
rect 232497 1320 238083 1322
rect 232497 1264 232502 1320
rect 232558 1264 238022 1320
rect 238078 1264 238083 1320
rect 232497 1262 238083 1264
rect 232497 1259 232563 1262
rect 238017 1259 238083 1262
rect 238201 1322 238267 1325
rect 245510 1322 245516 1324
rect 238201 1320 245516 1322
rect 238201 1264 238206 1320
rect 238262 1264 245516 1320
rect 238201 1262 245516 1264
rect 238201 1259 238267 1262
rect 245510 1260 245516 1262
rect 245580 1260 245586 1324
rect 245694 1260 245700 1324
rect 245764 1322 245770 1324
rect 247309 1322 247375 1325
rect 245764 1320 247375 1322
rect 245764 1264 247314 1320
rect 247370 1264 247375 1320
rect 245764 1262 247375 1264
rect 245764 1260 245770 1262
rect 247309 1259 247375 1262
rect 247902 1260 247908 1324
rect 247972 1322 247978 1324
rect 250478 1322 250484 1324
rect 247972 1262 250484 1322
rect 247972 1260 247978 1262
rect 250478 1260 250484 1262
rect 250548 1260 250554 1324
rect 250621 1322 250687 1325
rect 251214 1322 251220 1324
rect 250621 1320 251220 1322
rect 250621 1264 250626 1320
rect 250682 1264 251220 1320
rect 250621 1262 251220 1264
rect 250621 1259 250687 1262
rect 251214 1260 251220 1262
rect 251284 1260 251290 1324
rect 251406 1322 251466 1398
rect 251541 1456 252938 1458
rect 251541 1400 251546 1456
rect 251602 1400 252938 1456
rect 251541 1398 252938 1400
rect 253062 1398 253428 1458
rect 251541 1395 251607 1398
rect 252737 1322 252803 1325
rect 251406 1320 252803 1322
rect 251406 1264 252742 1320
rect 252798 1264 252803 1320
rect 251406 1262 252803 1264
rect 252737 1259 252803 1262
rect 180996 1126 182834 1186
rect 182909 1186 182975 1189
rect 184197 1186 184263 1189
rect 185853 1186 185919 1189
rect 182909 1184 184122 1186
rect 182909 1128 182914 1184
rect 182970 1128 184122 1184
rect 182909 1126 184122 1128
rect 180996 1124 181002 1126
rect 182909 1123 182975 1126
rect 153377 1050 153443 1053
rect 139166 1048 153443 1050
rect 139166 992 153382 1048
rect 153438 992 153443 1048
rect 139166 990 153443 992
rect 135805 987 135871 990
rect 139025 987 139091 990
rect 153377 987 153443 990
rect 153561 1050 153627 1053
rect 157057 1050 157123 1053
rect 153561 1048 157123 1050
rect 153561 992 153566 1048
rect 153622 992 157062 1048
rect 157118 992 157123 1048
rect 153561 990 157123 992
rect 153561 987 153627 990
rect 157057 987 157123 990
rect 157241 1050 157307 1053
rect 163681 1050 163747 1053
rect 157241 1048 163747 1050
rect 157241 992 157246 1048
rect 157302 992 163686 1048
rect 163742 992 163747 1048
rect 157241 990 163747 992
rect 157241 987 157307 990
rect 163681 987 163747 990
rect 163814 988 163820 1052
rect 163884 1050 163890 1052
rect 166625 1050 166691 1053
rect 163884 1048 166691 1050
rect 163884 992 166630 1048
rect 166686 992 166691 1048
rect 163884 990 166691 992
rect 163884 988 163890 990
rect 166625 987 166691 990
rect 166809 1050 166875 1053
rect 183921 1050 183987 1053
rect 166809 1048 183987 1050
rect 166809 992 166814 1048
rect 166870 992 183926 1048
rect 183982 992 183987 1048
rect 166809 990 183987 992
rect 184062 1050 184122 1126
rect 184197 1184 185919 1186
rect 184197 1128 184202 1184
rect 184258 1128 185858 1184
rect 185914 1128 185919 1184
rect 184197 1126 185919 1128
rect 184197 1123 184263 1126
rect 185853 1123 185919 1126
rect 186497 1186 186563 1189
rect 190361 1186 190427 1189
rect 186497 1184 190427 1186
rect 186497 1128 186502 1184
rect 186558 1128 190366 1184
rect 190422 1128 190427 1184
rect 186497 1126 190427 1128
rect 186497 1123 186563 1126
rect 190361 1123 190427 1126
rect 190821 1186 190887 1189
rect 191046 1186 191052 1188
rect 190821 1184 191052 1186
rect 190821 1128 190826 1184
rect 190882 1128 191052 1184
rect 190821 1126 191052 1128
rect 190821 1123 190887 1126
rect 191046 1124 191052 1126
rect 191116 1124 191122 1188
rect 191414 1186 191420 1188
rect 191238 1126 191420 1186
rect 184289 1050 184355 1053
rect 184062 1048 184355 1050
rect 184062 992 184294 1048
rect 184350 992 184355 1048
rect 184062 990 184355 992
rect 166809 987 166875 990
rect 183921 987 183987 990
rect 184289 987 184355 990
rect 184422 988 184428 1052
rect 184492 1050 184498 1052
rect 189758 1050 189764 1052
rect 184492 990 189764 1050
rect 184492 988 184498 990
rect 189758 988 189764 990
rect 189828 988 189834 1052
rect 189901 1050 189967 1053
rect 191238 1050 191298 1126
rect 191414 1124 191420 1126
rect 191484 1124 191490 1188
rect 191557 1186 191623 1189
rect 196709 1186 196775 1189
rect 191557 1184 196775 1186
rect 191557 1128 191562 1184
rect 191618 1128 196714 1184
rect 196770 1128 196775 1184
rect 191557 1126 196775 1128
rect 191557 1123 191623 1126
rect 196709 1123 196775 1126
rect 196934 1124 196940 1188
rect 197004 1186 197010 1188
rect 198089 1186 198155 1189
rect 209037 1186 209103 1189
rect 197004 1184 198155 1186
rect 197004 1128 198094 1184
rect 198150 1128 198155 1184
rect 197004 1126 198155 1128
rect 197004 1124 197010 1126
rect 198089 1123 198155 1126
rect 198230 1184 209103 1186
rect 198230 1128 209042 1184
rect 209098 1128 209103 1184
rect 198230 1126 209103 1128
rect 189901 1048 191298 1050
rect 189901 992 189906 1048
rect 189962 992 191298 1048
rect 189901 990 191298 992
rect 191373 1050 191439 1053
rect 197169 1050 197235 1053
rect 191373 1048 197235 1050
rect 191373 992 191378 1048
rect 191434 992 197174 1048
rect 197230 992 197235 1048
rect 191373 990 197235 992
rect 189901 987 189967 990
rect 191373 987 191439 990
rect 197169 987 197235 990
rect 197302 988 197308 1052
rect 197372 1050 197378 1052
rect 198230 1050 198290 1126
rect 209037 1123 209103 1126
rect 209221 1188 209287 1189
rect 209221 1184 209268 1188
rect 209332 1186 209338 1188
rect 209497 1186 209563 1189
rect 211889 1186 211955 1189
rect 209221 1128 209226 1184
rect 209221 1124 209268 1128
rect 209332 1126 209378 1186
rect 209497 1184 211955 1186
rect 209497 1128 209502 1184
rect 209558 1128 211894 1184
rect 211950 1128 211955 1184
rect 209497 1126 211955 1128
rect 209332 1124 209338 1126
rect 209221 1123 209287 1124
rect 209497 1123 209563 1126
rect 211889 1123 211955 1126
rect 212022 1124 212028 1188
rect 212092 1186 212098 1188
rect 217726 1186 217732 1188
rect 212092 1126 217732 1186
rect 212092 1124 212098 1126
rect 217726 1124 217732 1126
rect 217796 1124 217802 1188
rect 217869 1186 217935 1189
rect 224953 1186 225019 1189
rect 225137 1188 225203 1189
rect 217869 1184 225019 1186
rect 217869 1128 217874 1184
rect 217930 1128 224958 1184
rect 225014 1128 225019 1184
rect 217869 1126 225019 1128
rect 217869 1123 217935 1126
rect 224953 1123 225019 1126
rect 225086 1124 225092 1188
rect 225156 1186 225203 1188
rect 225321 1186 225387 1189
rect 226609 1186 226675 1189
rect 225156 1184 225248 1186
rect 225198 1128 225248 1184
rect 225156 1126 225248 1128
rect 225321 1184 226675 1186
rect 225321 1128 225326 1184
rect 225382 1128 226614 1184
rect 226670 1128 226675 1184
rect 225321 1126 226675 1128
rect 225156 1124 225203 1126
rect 225137 1123 225203 1124
rect 225321 1123 225387 1126
rect 226609 1123 226675 1126
rect 226742 1124 226748 1188
rect 226812 1186 226818 1188
rect 252737 1186 252803 1189
rect 226812 1184 252803 1186
rect 226812 1128 252742 1184
rect 252798 1128 252803 1184
rect 226812 1126 252803 1128
rect 226812 1124 226818 1126
rect 252737 1123 252803 1126
rect 197372 990 198290 1050
rect 198365 1050 198431 1053
rect 247401 1050 247467 1053
rect 198365 1048 247467 1050
rect 198365 992 198370 1048
rect 198426 992 247406 1048
rect 247462 992 247467 1048
rect 198365 990 247467 992
rect 197372 988 197378 990
rect 198365 987 198431 990
rect 247401 987 247467 990
rect 247534 988 247540 1052
rect 247604 1050 247610 1052
rect 247769 1050 247835 1053
rect 247604 1048 247835 1050
rect 247604 992 247774 1048
rect 247830 992 247835 1048
rect 247604 990 247835 992
rect 247604 988 247610 990
rect 247769 987 247835 990
rect 247902 988 247908 1052
rect 247972 1050 247978 1052
rect 250529 1050 250595 1053
rect 247972 1048 250595 1050
rect 247972 992 250534 1048
rect 250590 992 250595 1048
rect 247972 990 250595 992
rect 247972 988 247978 990
rect 250529 987 250595 990
rect 250713 1050 250779 1053
rect 251633 1050 251699 1053
rect 252686 1050 252692 1052
rect 250713 1048 251699 1050
rect 250713 992 250718 1048
rect 250774 992 251638 1048
rect 251694 992 251699 1048
rect 250713 990 251699 992
rect 250713 987 250779 990
rect 251633 987 251699 990
rect 251774 990 252692 1050
rect 130028 854 135730 914
rect 130028 852 130034 854
rect 135846 852 135852 916
rect 135916 914 135922 916
rect 138381 914 138447 917
rect 139393 914 139459 917
rect 135916 854 137938 914
rect 135916 852 135922 854
rect 130326 778 130332 780
rect 129782 718 130332 778
rect 129292 716 129298 718
rect 129641 715 129707 718
rect 130326 716 130332 718
rect 130396 716 130402 780
rect 130510 716 130516 780
rect 130580 778 130586 780
rect 134926 778 134932 780
rect 130580 718 134932 778
rect 130580 716 130586 718
rect 134926 716 134932 718
rect 134996 716 135002 780
rect 135294 716 135300 780
rect 135364 778 135370 780
rect 136081 778 136147 781
rect 135364 776 136147 778
rect 135364 720 136086 776
rect 136142 720 136147 776
rect 135364 718 136147 720
rect 135364 716 135370 718
rect 136081 715 136147 718
rect 136214 716 136220 780
rect 136284 778 136290 780
rect 137686 778 137692 780
rect 136284 718 137692 778
rect 136284 716 136290 718
rect 137686 716 137692 718
rect 137756 716 137762 780
rect 137878 778 137938 854
rect 138381 912 139459 914
rect 138381 856 138386 912
rect 138442 856 139398 912
rect 139454 856 139459 912
rect 138381 854 139459 856
rect 138381 851 138447 854
rect 139393 851 139459 854
rect 139577 914 139643 917
rect 150750 914 150756 916
rect 139577 912 150756 914
rect 139577 856 139582 912
rect 139638 856 150756 912
rect 139577 854 150756 856
rect 139577 851 139643 854
rect 150750 852 150756 854
rect 150820 852 150826 916
rect 150934 852 150940 916
rect 151004 914 151010 916
rect 151169 914 151235 917
rect 151004 912 151235 914
rect 151004 856 151174 912
rect 151230 856 151235 912
rect 151004 854 151235 856
rect 151004 852 151010 854
rect 151169 851 151235 854
rect 151302 852 151308 916
rect 151372 914 151378 916
rect 197721 914 197787 917
rect 151372 912 197787 914
rect 151372 856 197726 912
rect 197782 856 197787 912
rect 151372 854 197787 856
rect 151372 852 151378 854
rect 197721 851 197787 854
rect 197854 852 197860 916
rect 197924 852 197930 916
rect 198181 914 198247 917
rect 231342 914 231348 916
rect 198181 912 231348 914
rect 198181 856 198186 912
rect 198242 856 231348 912
rect 198181 854 231348 856
rect 139393 778 139459 781
rect 137878 776 139459 778
rect 137878 720 139398 776
rect 139454 720 139459 776
rect 137878 718 139459 720
rect 139393 715 139459 718
rect 139577 778 139643 781
rect 142245 778 142311 781
rect 139577 776 142311 778
rect 139577 720 139582 776
rect 139638 720 142250 776
rect 142306 720 142311 776
rect 139577 718 142311 720
rect 139577 715 139643 718
rect 142245 715 142311 718
rect 142429 778 142495 781
rect 144177 778 144243 781
rect 142429 776 144243 778
rect 142429 720 142434 776
rect 142490 720 144182 776
rect 144238 720 144243 776
rect 142429 718 144243 720
rect 142429 715 142495 718
rect 144177 715 144243 718
rect 144310 716 144316 780
rect 144380 778 144386 780
rect 145598 778 145604 780
rect 144380 718 145604 778
rect 144380 716 144386 718
rect 145598 716 145604 718
rect 145668 716 145674 780
rect 145741 778 145807 781
rect 146937 778 147003 781
rect 145741 776 147003 778
rect 145741 720 145746 776
rect 145802 720 146942 776
rect 146998 720 147003 776
rect 145741 718 147003 720
rect 145741 715 145807 718
rect 146937 715 147003 718
rect 147070 716 147076 780
rect 147140 778 147146 780
rect 161473 778 161539 781
rect 147140 718 156522 778
rect 147140 716 147146 718
rect 112345 640 114018 642
rect 112345 584 112350 640
rect 112406 584 114018 640
rect 112345 582 114018 584
rect 114093 642 114159 645
rect 115749 642 115815 645
rect 114093 640 115815 642
rect 114093 584 114098 640
rect 114154 584 115754 640
rect 115810 584 115815 640
rect 114093 582 115815 584
rect 112345 579 112411 582
rect 114093 579 114159 582
rect 115749 579 115815 582
rect 115933 642 115999 645
rect 120901 642 120967 645
rect 115933 640 120967 642
rect 115933 584 115938 640
rect 115994 584 120906 640
rect 120962 584 120967 640
rect 115933 582 120967 584
rect 115933 579 115999 582
rect 120901 579 120967 582
rect 121177 642 121243 645
rect 123753 642 123819 645
rect 121177 640 123819 642
rect 121177 584 121182 640
rect 121238 584 123758 640
rect 123814 584 123819 640
rect 121177 582 123819 584
rect 121177 579 121243 582
rect 123753 579 123819 582
rect 123937 642 124003 645
rect 124070 642 124076 644
rect 123937 640 124076 642
rect 123937 584 123942 640
rect 123998 584 124076 640
rect 123937 582 124076 584
rect 123937 579 124003 582
rect 124070 580 124076 582
rect 124140 580 124146 644
rect 124213 642 124279 645
rect 135345 642 135411 645
rect 124213 640 129520 642
rect 124213 584 124218 640
rect 124274 608 129520 640
rect 129782 640 135411 642
rect 129782 608 135350 640
rect 124274 584 135350 608
rect 135406 584 135411 640
rect 124213 582 135411 584
rect 124213 579 124279 582
rect 129460 548 129842 582
rect 135345 579 135411 582
rect 135478 580 135484 644
rect 135548 642 135554 644
rect 139894 642 139900 644
rect 135548 582 139900 642
rect 135548 580 135554 582
rect 139894 580 139900 582
rect 139964 580 139970 644
rect 140037 642 140103 645
rect 150249 642 150315 645
rect 151077 642 151143 645
rect 151302 642 151308 644
rect 140037 640 150315 642
rect 140037 584 140042 640
rect 140098 584 150254 640
rect 150310 584 150315 640
rect 140037 582 150315 584
rect 140037 579 140103 582
rect 150249 579 150315 582
rect 150574 582 151002 642
rect 102734 446 103162 506
rect 103278 444 103284 508
rect 103348 506 103354 508
rect 111742 506 111748 508
rect 103348 446 111748 506
rect 103348 444 103354 446
rect 111742 444 111748 446
rect 111812 444 111818 508
rect 111885 506 111951 509
rect 112069 506 112135 509
rect 111885 504 112135 506
rect 111885 448 111890 504
rect 111946 448 112074 504
rect 112130 448 112135 504
rect 111885 446 112135 448
rect 111885 443 111951 446
rect 112069 443 112135 446
rect 112294 444 112300 508
rect 112364 506 112370 508
rect 129273 506 129339 509
rect 112364 446 122850 506
rect 112364 444 112370 446
rect 65333 370 65399 373
rect 73337 370 73403 373
rect 65333 368 73403 370
rect 65333 312 65338 368
rect 65394 312 73342 368
rect 73398 312 73403 368
rect 65333 310 73403 312
rect 65333 307 65399 310
rect 73337 307 73403 310
rect 73797 370 73863 373
rect 92473 370 92539 373
rect 73797 368 92539 370
rect 73797 312 73802 368
rect 73858 312 92478 368
rect 92534 312 92539 368
rect 73797 310 92539 312
rect 73797 307 73863 310
rect 92473 307 92539 310
rect 92657 370 92723 373
rect 122649 370 122715 373
rect 92657 368 122715 370
rect 92657 312 92662 368
rect 92718 312 122654 368
rect 122710 312 122715 368
rect 92657 310 122715 312
rect 122790 370 122850 446
rect 123158 504 129339 506
rect 123158 448 129278 504
rect 129334 448 129339 504
rect 123158 446 129339 448
rect 123158 370 123218 446
rect 129273 443 129339 446
rect 129917 506 129983 509
rect 150574 506 150634 582
rect 150801 508 150867 509
rect 150750 506 150756 508
rect 129917 504 150634 506
rect 129917 448 129922 504
rect 129978 448 150634 504
rect 129917 446 150634 448
rect 150710 446 150756 506
rect 150820 504 150867 508
rect 150862 448 150867 504
rect 129917 443 129983 446
rect 150750 444 150756 446
rect 150820 444 150867 448
rect 150942 506 151002 582
rect 151077 640 151308 642
rect 151077 584 151082 640
rect 151138 584 151308 640
rect 151077 582 151308 584
rect 151077 579 151143 582
rect 151302 580 151308 582
rect 151372 580 151378 644
rect 151445 642 151511 645
rect 156270 642 156276 644
rect 151445 640 156276 642
rect 151445 584 151450 640
rect 151506 584 156276 640
rect 151445 582 156276 584
rect 151445 579 151511 582
rect 156270 580 156276 582
rect 156340 580 156346 644
rect 156462 642 156522 718
rect 157014 776 161539 778
rect 157014 720 161478 776
rect 161534 720 161539 776
rect 157014 718 161539 720
rect 157014 642 157074 718
rect 161473 715 161539 718
rect 161606 716 161612 780
rect 161676 716 161682 780
rect 161749 778 161815 781
rect 163129 778 163195 781
rect 161749 776 163195 778
rect 161749 720 161754 776
rect 161810 720 163134 776
rect 163190 720 163195 776
rect 161749 718 163195 720
rect 156462 582 157074 642
rect 157149 642 157215 645
rect 157609 642 157675 645
rect 157885 644 157951 645
rect 157885 642 157932 644
rect 157149 640 157675 642
rect 157149 584 157154 640
rect 157210 584 157614 640
rect 157670 584 157675 640
rect 157149 582 157675 584
rect 157840 640 157932 642
rect 157840 584 157890 640
rect 157840 582 157932 584
rect 157149 579 157215 582
rect 157609 579 157675 582
rect 157885 580 157932 582
rect 157996 580 158002 644
rect 158069 642 158135 645
rect 161614 642 161674 716
rect 161749 715 161815 718
rect 163129 715 163195 718
rect 163262 716 163268 780
rect 163332 778 163338 780
rect 163681 778 163747 781
rect 163332 776 163747 778
rect 163332 720 163686 776
rect 163742 720 163747 776
rect 163332 718 163747 720
rect 163332 716 163338 718
rect 163681 715 163747 718
rect 163865 778 163931 781
rect 176009 778 176075 781
rect 163865 776 176075 778
rect 163865 720 163870 776
rect 163926 720 176014 776
rect 176070 720 176075 776
rect 163865 718 176075 720
rect 163865 715 163931 718
rect 176009 715 176075 718
rect 176193 778 176259 781
rect 184197 778 184263 781
rect 176193 776 184263 778
rect 176193 720 176198 776
rect 176254 720 184202 776
rect 184258 720 184263 776
rect 176193 718 184263 720
rect 176193 715 176259 718
rect 184197 715 184263 718
rect 184381 778 184447 781
rect 190310 778 190316 780
rect 184381 776 190316 778
rect 184381 720 184386 776
rect 184442 720 190316 776
rect 184381 718 190316 720
rect 184381 715 184447 718
rect 190310 716 190316 718
rect 190380 716 190386 780
rect 190453 778 190519 781
rect 197537 778 197603 781
rect 190453 776 197603 778
rect 190453 720 190458 776
rect 190514 720 197542 776
rect 197598 720 197603 776
rect 190453 718 197603 720
rect 197862 778 197922 852
rect 198181 851 198247 854
rect 231342 852 231348 854
rect 231412 852 231418 916
rect 231485 914 231551 917
rect 232630 914 232636 916
rect 231485 912 232636 914
rect 231485 856 231490 912
rect 231546 856 232636 912
rect 231485 854 232636 856
rect 231485 851 231551 854
rect 232630 852 232636 854
rect 232700 852 232706 916
rect 232814 852 232820 916
rect 232884 914 232890 916
rect 233141 914 233207 917
rect 233325 916 233391 917
rect 233325 914 233372 916
rect 232884 912 233207 914
rect 232884 856 233146 912
rect 233202 856 233207 912
rect 232884 854 233207 856
rect 233280 912 233372 914
rect 233280 856 233330 912
rect 233280 854 233372 856
rect 232884 852 232890 854
rect 233141 851 233207 854
rect 233325 852 233372 854
rect 233436 852 233442 916
rect 233734 852 233740 916
rect 233804 914 233810 916
rect 246757 914 246823 917
rect 233804 912 246823 914
rect 233804 856 246762 912
rect 246818 856 246823 912
rect 233804 854 246823 856
rect 233804 852 233810 854
rect 233325 851 233391 852
rect 246757 851 246823 854
rect 246941 914 247007 917
rect 250161 914 250227 917
rect 246941 912 250227 914
rect 246941 856 246946 912
rect 247002 856 250166 912
rect 250222 856 250227 912
rect 246941 854 250227 856
rect 246941 851 247007 854
rect 250161 851 250227 854
rect 250294 852 250300 916
rect 250364 914 250370 916
rect 251774 914 251834 990
rect 252686 988 252692 990
rect 252756 988 252762 1052
rect 252878 1050 252938 1398
rect 253422 1396 253428 1398
rect 253492 1396 253498 1460
rect 253614 1458 253674 1534
rect 253790 1532 253796 1596
rect 253860 1594 253866 1596
rect 256601 1594 256667 1597
rect 258214 1594 258274 1670
rect 261702 1668 261708 1670
rect 261772 1668 261778 1732
rect 262029 1730 262095 1733
rect 268469 1730 268535 1733
rect 268694 1730 268700 1732
rect 262029 1728 268394 1730
rect 262029 1672 262034 1728
rect 262090 1672 268394 1728
rect 262029 1670 268394 1672
rect 262029 1667 262095 1670
rect 268334 1597 268394 1670
rect 268469 1728 268700 1730
rect 268469 1672 268474 1728
rect 268530 1672 268700 1728
rect 268469 1670 268700 1672
rect 268469 1667 268535 1670
rect 268694 1668 268700 1670
rect 268764 1668 268770 1732
rect 268837 1730 268903 1733
rect 268837 1728 272074 1730
rect 268837 1672 268842 1728
rect 268898 1672 272074 1728
rect 268837 1670 272074 1672
rect 268837 1667 268903 1670
rect 253860 1592 256667 1594
rect 253860 1536 256606 1592
rect 256662 1536 256667 1592
rect 253860 1534 256667 1536
rect 253860 1532 253866 1534
rect 256601 1531 256667 1534
rect 256926 1534 258274 1594
rect 254025 1458 254091 1461
rect 253614 1456 254091 1458
rect 253614 1400 254030 1456
rect 254086 1400 254091 1456
rect 253614 1398 254091 1400
rect 254025 1395 254091 1398
rect 254209 1458 254275 1461
rect 256926 1458 256986 1534
rect 258390 1532 258396 1596
rect 258460 1594 258466 1596
rect 261886 1594 261892 1596
rect 258460 1534 261892 1594
rect 258460 1532 258466 1534
rect 261886 1532 261892 1534
rect 261956 1532 261962 1596
rect 262029 1594 262095 1597
rect 262029 1592 268210 1594
rect 262029 1536 262034 1592
rect 262090 1536 268210 1592
rect 262029 1534 268210 1536
rect 268334 1592 268443 1597
rect 270953 1594 271019 1597
rect 271873 1594 271939 1597
rect 268334 1536 268382 1592
rect 268438 1536 268443 1592
rect 268334 1534 268443 1536
rect 262029 1531 262095 1534
rect 254209 1456 256986 1458
rect 254209 1400 254214 1456
rect 254270 1400 256986 1456
rect 254209 1398 256986 1400
rect 257061 1458 257127 1461
rect 258073 1458 258139 1461
rect 257061 1456 258139 1458
rect 257061 1400 257066 1456
rect 257122 1400 258078 1456
rect 258134 1400 258139 1456
rect 257061 1398 258139 1400
rect 254209 1395 254275 1398
rect 257061 1395 257127 1398
rect 258073 1395 258139 1398
rect 259085 1458 259151 1461
rect 260465 1458 260531 1461
rect 260649 1460 260715 1461
rect 259085 1456 260531 1458
rect 259085 1400 259090 1456
rect 259146 1400 260470 1456
rect 260526 1400 260531 1456
rect 259085 1398 260531 1400
rect 259085 1395 259151 1398
rect 260465 1395 260531 1398
rect 260598 1396 260604 1460
rect 260668 1458 260715 1460
rect 260668 1456 260760 1458
rect 260710 1400 260760 1456
rect 260668 1398 260760 1400
rect 260668 1396 260715 1398
rect 260966 1396 260972 1460
rect 261036 1458 261042 1460
rect 268009 1458 268075 1461
rect 261036 1456 268075 1458
rect 261036 1400 268014 1456
rect 268070 1400 268075 1456
rect 261036 1398 268075 1400
rect 268150 1458 268210 1534
rect 268377 1531 268443 1534
rect 268518 1592 271019 1594
rect 268518 1536 270958 1592
rect 271014 1536 271019 1592
rect 268518 1534 271019 1536
rect 268518 1458 268578 1534
rect 270953 1531 271019 1534
rect 271094 1592 271939 1594
rect 271094 1536 271878 1592
rect 271934 1536 271939 1592
rect 271094 1534 271939 1536
rect 272014 1594 272074 1670
rect 272190 1668 272196 1732
rect 272260 1730 272266 1732
rect 278998 1730 279004 1732
rect 272260 1670 279004 1730
rect 272260 1668 272266 1670
rect 278998 1668 279004 1670
rect 279068 1668 279074 1732
rect 279325 1730 279391 1733
rect 285622 1730 285628 1732
rect 279325 1728 285628 1730
rect 279325 1672 279330 1728
rect 279386 1672 285628 1728
rect 279325 1670 285628 1672
rect 279325 1667 279391 1670
rect 285622 1668 285628 1670
rect 285692 1668 285698 1732
rect 285765 1730 285831 1733
rect 294086 1730 294092 1766
rect 285765 1728 294092 1730
rect 285765 1672 285770 1728
rect 285826 1702 294092 1728
rect 294156 1702 294162 1766
rect 285826 1672 294154 1702
rect 285765 1670 294154 1672
rect 285765 1667 285831 1670
rect 294454 1668 294460 1732
rect 294524 1730 294530 1732
rect 294597 1730 294663 1733
rect 294524 1728 294663 1730
rect 294524 1672 294602 1728
rect 294658 1672 294663 1728
rect 294524 1670 294663 1672
rect 294524 1668 294530 1670
rect 294597 1667 294663 1670
rect 294965 1730 295031 1733
rect 309961 1730 310027 1733
rect 310462 1730 310468 1732
rect 294965 1728 309794 1730
rect 294965 1672 294970 1728
rect 295026 1672 309794 1728
rect 294965 1670 309794 1672
rect 294965 1667 295031 1670
rect 279785 1594 279851 1597
rect 272014 1592 279851 1594
rect 272014 1536 279790 1592
rect 279846 1536 279851 1592
rect 272014 1534 279851 1536
rect 268837 1460 268903 1461
rect 268837 1458 268884 1460
rect 268150 1398 268578 1458
rect 268792 1456 268884 1458
rect 268792 1400 268842 1456
rect 268792 1398 268884 1400
rect 261036 1396 261042 1398
rect 260649 1395 260715 1396
rect 268009 1395 268075 1398
rect 268837 1396 268884 1398
rect 268948 1396 268954 1460
rect 269021 1458 269087 1461
rect 271094 1458 271154 1534
rect 271873 1531 271939 1534
rect 279785 1531 279851 1534
rect 279969 1594 280035 1597
rect 280153 1594 280219 1597
rect 279969 1592 280219 1594
rect 279969 1536 279974 1592
rect 280030 1536 280158 1592
rect 280214 1536 280219 1592
rect 279969 1534 280219 1536
rect 279969 1531 280035 1534
rect 280153 1531 280219 1534
rect 280521 1594 280587 1597
rect 295609 1594 295675 1597
rect 280521 1592 285506 1594
rect 280521 1536 280526 1592
rect 280582 1536 285506 1592
rect 280521 1534 285506 1536
rect 280521 1531 280587 1534
rect 269021 1456 271154 1458
rect 269021 1400 269026 1456
rect 269082 1400 271154 1456
rect 269021 1398 271154 1400
rect 271229 1458 271295 1461
rect 273529 1460 273595 1461
rect 271229 1456 271706 1458
rect 271229 1400 271234 1456
rect 271290 1400 271706 1456
rect 271229 1398 271706 1400
rect 268837 1395 268903 1396
rect 269021 1395 269087 1398
rect 271229 1395 271295 1398
rect 253054 1260 253060 1324
rect 253124 1322 253130 1324
rect 253841 1322 253907 1325
rect 253124 1320 253907 1322
rect 253124 1264 253846 1320
rect 253902 1264 253907 1320
rect 253124 1262 253907 1264
rect 253124 1260 253130 1262
rect 253841 1259 253907 1262
rect 254025 1322 254091 1325
rect 256366 1322 256372 1324
rect 254025 1320 256372 1322
rect 254025 1264 254030 1320
rect 254086 1264 256372 1320
rect 254025 1262 256372 1264
rect 254025 1259 254091 1262
rect 256366 1260 256372 1262
rect 256436 1260 256442 1324
rect 256509 1322 256575 1325
rect 261201 1322 261267 1325
rect 256509 1320 261267 1322
rect 256509 1264 256514 1320
rect 256570 1264 261206 1320
rect 261262 1264 261267 1320
rect 256509 1262 261267 1264
rect 256509 1259 256575 1262
rect 261201 1259 261267 1262
rect 261385 1322 261451 1325
rect 262673 1322 262739 1325
rect 261385 1320 262739 1322
rect 261385 1264 261390 1320
rect 261446 1264 262678 1320
rect 262734 1264 262739 1320
rect 261385 1262 262739 1264
rect 261385 1259 261451 1262
rect 262673 1259 262739 1262
rect 262806 1260 262812 1324
rect 262876 1322 262882 1324
rect 264830 1322 264836 1324
rect 262876 1262 264836 1322
rect 262876 1260 262882 1262
rect 264830 1260 264836 1262
rect 264900 1260 264906 1324
rect 265341 1322 265407 1325
rect 271413 1322 271479 1325
rect 265341 1320 271479 1322
rect 265341 1264 265346 1320
rect 265402 1264 271418 1320
rect 271474 1264 271479 1320
rect 265341 1262 271479 1264
rect 271646 1322 271706 1398
rect 271822 1396 271828 1460
rect 271892 1458 271898 1460
rect 273294 1458 273300 1460
rect 271892 1398 273300 1458
rect 271892 1396 271898 1398
rect 273294 1396 273300 1398
rect 273364 1396 273370 1460
rect 273478 1458 273484 1460
rect 273438 1398 273484 1458
rect 273548 1456 273595 1460
rect 273590 1400 273595 1456
rect 273478 1396 273484 1398
rect 273548 1396 273595 1400
rect 273662 1396 273668 1460
rect 273732 1458 273738 1460
rect 279366 1458 279372 1460
rect 273732 1398 279372 1458
rect 273732 1396 273738 1398
rect 279366 1396 279372 1398
rect 279436 1396 279442 1460
rect 280470 1396 280476 1460
rect 280540 1458 280546 1460
rect 280540 1398 281274 1458
rect 280540 1396 280546 1398
rect 273529 1395 273595 1396
rect 280521 1322 280587 1325
rect 280981 1324 281047 1325
rect 280981 1322 281028 1324
rect 271646 1320 280587 1322
rect 271646 1264 280526 1320
rect 280582 1264 280587 1320
rect 271646 1262 280587 1264
rect 280936 1320 281028 1322
rect 280936 1264 280986 1320
rect 280936 1262 281028 1264
rect 265341 1259 265407 1262
rect 271413 1259 271479 1262
rect 280521 1259 280587 1262
rect 280981 1260 281028 1262
rect 281092 1260 281098 1324
rect 281214 1322 281274 1398
rect 281390 1396 281396 1460
rect 281460 1458 281466 1460
rect 281533 1458 281599 1461
rect 281460 1456 281599 1458
rect 281460 1400 281538 1456
rect 281594 1400 281599 1456
rect 281460 1398 281599 1400
rect 281460 1396 281466 1398
rect 281533 1395 281599 1398
rect 281717 1458 281783 1461
rect 285305 1458 285371 1461
rect 281717 1456 285371 1458
rect 281717 1400 281722 1456
rect 281778 1400 285310 1456
rect 285366 1400 285371 1456
rect 281717 1398 285371 1400
rect 285446 1458 285506 1534
rect 285814 1592 295675 1594
rect 285814 1536 295614 1592
rect 295670 1536 295675 1592
rect 285814 1534 295675 1536
rect 285814 1458 285874 1534
rect 295609 1531 295675 1534
rect 295793 1594 295859 1597
rect 296110 1594 296116 1596
rect 295793 1592 296116 1594
rect 295793 1536 295798 1592
rect 295854 1536 296116 1592
rect 295793 1534 296116 1536
rect 295793 1531 295859 1534
rect 296110 1532 296116 1534
rect 296180 1532 296186 1596
rect 296253 1594 296319 1597
rect 305637 1594 305703 1597
rect 296253 1592 305703 1594
rect 296253 1536 296258 1592
rect 296314 1536 305642 1592
rect 305698 1536 305703 1592
rect 296253 1534 305703 1536
rect 296253 1531 296319 1534
rect 305637 1531 305703 1534
rect 305821 1594 305887 1597
rect 307017 1594 307083 1597
rect 305821 1592 307083 1594
rect 305821 1536 305826 1592
rect 305882 1536 307022 1592
rect 307078 1536 307083 1592
rect 305821 1534 307083 1536
rect 305821 1531 305887 1534
rect 307017 1531 307083 1534
rect 307201 1594 307267 1597
rect 309225 1594 309291 1597
rect 307201 1592 309291 1594
rect 307201 1536 307206 1592
rect 307262 1536 309230 1592
rect 309286 1536 309291 1592
rect 307201 1534 309291 1536
rect 309734 1594 309794 1670
rect 309961 1728 310468 1730
rect 309961 1672 309966 1728
rect 310022 1672 310468 1728
rect 309961 1670 310468 1672
rect 309961 1667 310027 1670
rect 310462 1668 310468 1670
rect 310532 1668 310538 1732
rect 310646 1668 310652 1732
rect 310716 1730 310722 1732
rect 321737 1730 321803 1733
rect 310716 1728 321803 1730
rect 310716 1672 321742 1728
rect 321798 1672 321803 1728
rect 310716 1670 321803 1672
rect 310716 1668 310722 1670
rect 321737 1667 321803 1670
rect 321921 1730 321987 1733
rect 347405 1730 347471 1733
rect 321921 1728 347471 1730
rect 321921 1672 321926 1728
rect 321982 1672 347410 1728
rect 347466 1672 347471 1728
rect 321921 1670 347471 1672
rect 321921 1667 321987 1670
rect 347405 1667 347471 1670
rect 348325 1730 348391 1733
rect 373717 1730 373783 1733
rect 348325 1728 373783 1730
rect 348325 1672 348330 1728
rect 348386 1672 373722 1728
rect 373778 1672 373783 1728
rect 348325 1670 373783 1672
rect 348325 1667 348391 1670
rect 373717 1667 373783 1670
rect 373901 1730 373967 1733
rect 380157 1730 380223 1733
rect 373901 1728 380223 1730
rect 373901 1672 373906 1728
rect 373962 1672 380162 1728
rect 380218 1672 380223 1728
rect 373901 1670 380223 1672
rect 373901 1667 373967 1670
rect 380157 1667 380223 1670
rect 380341 1730 380407 1733
rect 385718 1730 385724 1732
rect 380341 1728 385724 1730
rect 380341 1672 380346 1728
rect 380402 1672 385724 1728
rect 380341 1670 385724 1672
rect 380341 1667 380407 1670
rect 385718 1668 385724 1670
rect 385788 1668 385794 1732
rect 389081 1730 389147 1733
rect 395429 1730 395495 1733
rect 389081 1728 395495 1730
rect 389081 1672 389086 1728
rect 389142 1672 395434 1728
rect 395490 1672 395495 1728
rect 389081 1670 395495 1672
rect 389081 1667 389147 1670
rect 395429 1667 395495 1670
rect 398649 1730 398715 1733
rect 399569 1730 399635 1733
rect 398649 1728 399635 1730
rect 398649 1672 398654 1728
rect 398710 1672 399574 1728
rect 399630 1672 399635 1728
rect 398649 1670 399635 1672
rect 398649 1667 398715 1670
rect 399569 1667 399635 1670
rect 403709 1730 403775 1733
rect 415669 1730 415735 1733
rect 403709 1728 415735 1730
rect 403709 1672 403714 1728
rect 403770 1672 415674 1728
rect 415730 1672 415735 1728
rect 403709 1670 415735 1672
rect 403709 1667 403775 1670
rect 415669 1667 415735 1670
rect 418797 1730 418863 1733
rect 432321 1730 432387 1733
rect 418797 1728 432387 1730
rect 418797 1672 418802 1728
rect 418858 1672 432326 1728
rect 432382 1672 432387 1728
rect 418797 1670 432387 1672
rect 418797 1667 418863 1670
rect 432321 1667 432387 1670
rect 436001 1730 436067 1733
rect 443453 1730 443519 1733
rect 436001 1728 443519 1730
rect 436001 1672 436006 1728
rect 436062 1672 443458 1728
rect 443514 1672 443519 1728
rect 436001 1670 443519 1672
rect 436001 1667 436067 1670
rect 443453 1667 443519 1670
rect 443637 1730 443703 1733
rect 453297 1730 453363 1733
rect 443637 1728 453363 1730
rect 443637 1672 443642 1728
rect 443698 1672 453302 1728
rect 453358 1672 453363 1728
rect 443637 1670 453363 1672
rect 443637 1667 443703 1670
rect 453297 1667 453363 1670
rect 462865 1730 462931 1733
rect 474917 1730 474983 1733
rect 462865 1728 474983 1730
rect 462865 1672 462870 1728
rect 462926 1672 474922 1728
rect 474978 1672 474983 1728
rect 462865 1670 474983 1672
rect 462865 1667 462931 1670
rect 474917 1667 474983 1670
rect 481265 1730 481331 1733
rect 488993 1730 489059 1733
rect 481265 1728 489059 1730
rect 481265 1672 481270 1728
rect 481326 1672 488998 1728
rect 489054 1672 489059 1728
rect 481265 1670 489059 1672
rect 481265 1667 481331 1670
rect 488993 1667 489059 1670
rect 501781 1730 501847 1733
rect 512361 1730 512427 1733
rect 501781 1728 512427 1730
rect 501781 1672 501786 1728
rect 501842 1672 512366 1728
rect 512422 1672 512427 1728
rect 501781 1670 512427 1672
rect 501781 1667 501847 1670
rect 512361 1667 512427 1670
rect 513230 1668 513236 1732
rect 513300 1730 513306 1732
rect 522573 1730 522639 1733
rect 513300 1728 522639 1730
rect 513300 1672 522578 1728
rect 522634 1672 522639 1728
rect 513300 1670 522639 1672
rect 513300 1668 513306 1670
rect 522573 1667 522639 1670
rect 529381 1730 529447 1733
rect 567142 1730 567148 1732
rect 529381 1728 567148 1730
rect 529381 1672 529386 1728
rect 529442 1672 567148 1728
rect 529381 1670 567148 1672
rect 529381 1667 529447 1670
rect 567142 1668 567148 1670
rect 567212 1668 567218 1732
rect 567285 1730 567351 1733
rect 569585 1732 569651 1733
rect 569166 1730 569172 1732
rect 567285 1728 569172 1730
rect 567285 1672 567290 1728
rect 567346 1672 569172 1728
rect 567285 1670 569172 1672
rect 567285 1667 567351 1670
rect 569166 1668 569172 1670
rect 569236 1668 569242 1732
rect 569534 1730 569540 1732
rect 569494 1670 569540 1730
rect 569604 1728 569651 1732
rect 569646 1672 569651 1728
rect 569534 1668 569540 1670
rect 569604 1668 569651 1672
rect 569585 1667 569651 1668
rect 319529 1594 319595 1597
rect 309734 1592 319595 1594
rect 309734 1536 319534 1592
rect 319590 1536 319595 1592
rect 309734 1534 319595 1536
rect 307201 1531 307267 1534
rect 309225 1531 309291 1534
rect 319529 1531 319595 1534
rect 319713 1594 319779 1597
rect 352925 1594 352991 1597
rect 319713 1592 352991 1594
rect 319713 1536 319718 1592
rect 319774 1536 352930 1592
rect 352986 1536 352991 1592
rect 319713 1534 352991 1536
rect 319713 1531 319779 1534
rect 352925 1531 352991 1534
rect 354254 1532 354260 1596
rect 354324 1594 354330 1596
rect 365989 1594 366055 1597
rect 354324 1592 366055 1594
rect 354324 1536 365994 1592
rect 366050 1536 366055 1592
rect 354324 1534 366055 1536
rect 354324 1532 354330 1534
rect 365989 1531 366055 1534
rect 366173 1594 366239 1597
rect 406837 1594 406903 1597
rect 366173 1592 406903 1594
rect 366173 1536 366178 1592
rect 366234 1536 406842 1592
rect 406898 1536 406903 1592
rect 366173 1534 406903 1536
rect 366173 1531 366239 1534
rect 406837 1531 406903 1534
rect 407021 1594 407087 1597
rect 415117 1594 415183 1597
rect 407021 1592 415183 1594
rect 407021 1536 407026 1592
rect 407082 1536 415122 1592
rect 415178 1536 415183 1592
rect 407021 1534 415183 1536
rect 407021 1531 407087 1534
rect 415117 1531 415183 1534
rect 418797 1594 418863 1597
rect 440693 1594 440759 1597
rect 418797 1592 440759 1594
rect 418797 1536 418802 1592
rect 418858 1536 440698 1592
rect 440754 1536 440759 1592
rect 418797 1534 440759 1536
rect 418797 1531 418863 1534
rect 440693 1531 440759 1534
rect 453205 1594 453271 1597
rect 462589 1594 462655 1597
rect 453205 1592 462655 1594
rect 453205 1536 453210 1592
rect 453266 1536 462594 1592
rect 462650 1536 462655 1592
rect 453205 1534 462655 1536
rect 453205 1531 453271 1534
rect 462589 1531 462655 1534
rect 471513 1594 471579 1597
rect 559097 1596 559163 1597
rect 558862 1594 558868 1596
rect 471513 1592 558868 1594
rect 471513 1536 471518 1592
rect 471574 1536 558868 1592
rect 471513 1534 558868 1536
rect 471513 1531 471579 1534
rect 558862 1532 558868 1534
rect 558932 1532 558938 1596
rect 559046 1594 559052 1596
rect 559006 1534 559052 1594
rect 559116 1592 559163 1596
rect 559158 1536 559163 1592
rect 559046 1532 559052 1534
rect 559116 1532 559163 1536
rect 559097 1531 559163 1532
rect 559373 1594 559439 1597
rect 565813 1594 565879 1597
rect 559373 1592 565879 1594
rect 559373 1536 559378 1592
rect 559434 1536 565818 1592
rect 565874 1536 565879 1592
rect 559373 1534 565879 1536
rect 559373 1531 559439 1534
rect 565813 1531 565879 1534
rect 285446 1398 285874 1458
rect 285949 1458 286015 1461
rect 556429 1458 556495 1461
rect 285949 1456 556495 1458
rect 285949 1400 285954 1456
rect 286010 1400 556434 1456
rect 556490 1400 556495 1456
rect 285949 1398 556495 1400
rect 281717 1395 281783 1398
rect 285305 1395 285371 1398
rect 285949 1395 286015 1398
rect 556429 1395 556495 1398
rect 559414 1396 559420 1460
rect 559484 1458 559490 1460
rect 560150 1458 560156 1460
rect 559484 1398 560156 1458
rect 559484 1396 559490 1398
rect 560150 1396 560156 1398
rect 560220 1396 560226 1460
rect 565813 1458 565879 1461
rect 566406 1458 566412 1460
rect 565813 1456 566412 1458
rect 565813 1400 565818 1456
rect 565874 1400 566412 1456
rect 565813 1398 566412 1400
rect 565813 1395 565879 1398
rect 566406 1396 566412 1398
rect 566476 1396 566482 1460
rect 289629 1322 289695 1325
rect 294689 1322 294755 1325
rect 281214 1262 287714 1322
rect 280981 1259 281047 1260
rect 253013 1186 253079 1189
rect 268878 1186 268884 1188
rect 253013 1184 268884 1186
rect 253013 1128 253018 1184
rect 253074 1128 268884 1184
rect 253013 1126 268884 1128
rect 253013 1123 253079 1126
rect 268878 1124 268884 1126
rect 268948 1124 268954 1188
rect 269205 1186 269271 1189
rect 273253 1186 273319 1189
rect 269205 1184 273319 1186
rect 269205 1128 269210 1184
rect 269266 1128 273258 1184
rect 273314 1128 273319 1184
rect 269205 1126 273319 1128
rect 269205 1123 269271 1126
rect 273253 1123 273319 1126
rect 273437 1186 273503 1189
rect 279417 1186 279483 1189
rect 273437 1184 279483 1186
rect 273437 1128 273442 1184
rect 273498 1128 279422 1184
rect 279478 1128 279483 1184
rect 273437 1126 279483 1128
rect 273437 1123 273503 1126
rect 279417 1123 279483 1126
rect 279550 1124 279556 1188
rect 279620 1186 279626 1188
rect 287513 1186 287579 1189
rect 279620 1184 287579 1186
rect 279620 1128 287518 1184
rect 287574 1128 287579 1184
rect 279620 1126 287579 1128
rect 279620 1124 279626 1126
rect 287513 1123 287579 1126
rect 253289 1050 253355 1053
rect 252878 1048 253355 1050
rect 252878 992 253294 1048
rect 253350 992 253355 1048
rect 252878 990 253355 992
rect 253289 987 253355 990
rect 253422 988 253428 1052
rect 253492 1050 253498 1052
rect 255865 1050 255931 1053
rect 253492 1048 255931 1050
rect 253492 992 255870 1048
rect 255926 992 255931 1048
rect 253492 990 255931 992
rect 253492 988 253498 990
rect 255865 987 255931 990
rect 255998 988 256004 1052
rect 256068 1050 256074 1052
rect 261937 1050 262003 1053
rect 262305 1052 262371 1053
rect 262254 1050 262260 1052
rect 256068 1048 262003 1050
rect 256068 992 261942 1048
rect 261998 992 262003 1048
rect 256068 990 262003 992
rect 262214 990 262260 1050
rect 262324 1048 262371 1052
rect 262366 992 262371 1048
rect 256068 988 256074 990
rect 261937 987 262003 990
rect 262254 988 262260 990
rect 262324 988 262371 992
rect 262305 987 262371 988
rect 262489 1050 262555 1053
rect 285673 1050 285739 1053
rect 262489 1048 285739 1050
rect 262489 992 262494 1048
rect 262550 992 285678 1048
rect 285734 992 285739 1048
rect 262489 990 285739 992
rect 287654 1050 287714 1262
rect 289629 1320 294755 1322
rect 289629 1264 289634 1320
rect 289690 1264 294694 1320
rect 294750 1264 294755 1320
rect 289629 1262 294755 1264
rect 289629 1259 289695 1262
rect 294689 1259 294755 1262
rect 294822 1260 294828 1324
rect 294892 1322 294898 1324
rect 294965 1322 295031 1325
rect 294892 1320 295031 1322
rect 294892 1264 294970 1320
rect 295026 1264 295031 1320
rect 294892 1262 295031 1264
rect 294892 1260 294898 1262
rect 294965 1259 295031 1262
rect 295149 1322 295215 1325
rect 317689 1322 317755 1325
rect 295149 1320 317755 1322
rect 295149 1264 295154 1320
rect 295210 1264 317694 1320
rect 317750 1264 317755 1320
rect 295149 1262 317755 1264
rect 295149 1259 295215 1262
rect 317689 1259 317755 1262
rect 317822 1260 317828 1324
rect 317892 1322 317898 1324
rect 318333 1322 318399 1325
rect 317892 1320 318399 1322
rect 317892 1264 318338 1320
rect 318394 1264 318399 1320
rect 317892 1262 318399 1264
rect 317892 1260 317898 1262
rect 318333 1259 318399 1262
rect 318609 1322 318675 1325
rect 322933 1322 322999 1325
rect 318609 1320 322999 1322
rect 318609 1264 318614 1320
rect 318670 1264 322938 1320
rect 322994 1264 322999 1320
rect 318609 1262 322999 1264
rect 318609 1259 318675 1262
rect 322933 1259 322999 1262
rect 323117 1322 323183 1325
rect 324814 1322 324820 1324
rect 323117 1320 324820 1322
rect 323117 1264 323122 1320
rect 323178 1264 324820 1320
rect 323117 1262 324820 1264
rect 323117 1259 323183 1262
rect 324814 1260 324820 1262
rect 324884 1260 324890 1324
rect 324957 1322 325023 1325
rect 327533 1322 327599 1325
rect 327717 1324 327783 1325
rect 327717 1322 327764 1324
rect 324957 1320 327599 1322
rect 324957 1264 324962 1320
rect 325018 1264 327538 1320
rect 327594 1264 327599 1320
rect 324957 1262 327599 1264
rect 327672 1320 327764 1322
rect 327672 1264 327722 1320
rect 327672 1262 327764 1264
rect 324957 1259 325023 1262
rect 327533 1259 327599 1262
rect 327717 1260 327764 1262
rect 327828 1260 327834 1324
rect 327901 1322 327967 1325
rect 364701 1322 364767 1325
rect 327901 1320 364767 1322
rect 327901 1264 327906 1320
rect 327962 1264 364706 1320
rect 364762 1264 364767 1320
rect 327901 1262 364767 1264
rect 327717 1259 327783 1260
rect 327901 1259 327967 1262
rect 364701 1259 364767 1262
rect 365989 1322 366055 1325
rect 372470 1322 372476 1324
rect 365989 1320 372476 1322
rect 365989 1264 365994 1320
rect 366050 1264 372476 1320
rect 365989 1262 372476 1264
rect 365989 1259 366055 1262
rect 372470 1260 372476 1262
rect 372540 1260 372546 1324
rect 373349 1322 373415 1325
rect 406653 1322 406719 1325
rect 373349 1320 406719 1322
rect 373349 1264 373354 1320
rect 373410 1264 406658 1320
rect 406714 1264 406719 1320
rect 373349 1262 406719 1264
rect 373349 1259 373415 1262
rect 406653 1259 406719 1262
rect 406837 1322 406903 1325
rect 418797 1322 418863 1325
rect 406837 1320 418863 1322
rect 406837 1264 406842 1320
rect 406898 1264 418802 1320
rect 418858 1264 418863 1320
rect 406837 1262 418863 1264
rect 406837 1259 406903 1262
rect 418797 1259 418863 1262
rect 419390 1260 419396 1324
rect 419460 1322 419466 1324
rect 436001 1322 436067 1325
rect 443177 1322 443243 1325
rect 419460 1320 436067 1322
rect 419460 1264 436006 1320
rect 436062 1264 436067 1320
rect 419460 1262 436067 1264
rect 419460 1260 419466 1262
rect 436001 1259 436067 1262
rect 439454 1320 443243 1322
rect 439454 1264 443182 1320
rect 443238 1264 443243 1320
rect 439454 1262 443243 1264
rect 287789 1186 287855 1189
rect 289537 1186 289603 1189
rect 290365 1188 290431 1189
rect 287789 1184 289603 1186
rect 287789 1128 287794 1184
rect 287850 1128 289542 1184
rect 289598 1128 289603 1184
rect 287789 1126 289603 1128
rect 287789 1123 287855 1126
rect 289537 1123 289603 1126
rect 289670 1124 289676 1188
rect 289740 1186 289746 1188
rect 290038 1186 290044 1188
rect 289740 1126 290044 1186
rect 289740 1124 289746 1126
rect 290038 1124 290044 1126
rect 290108 1124 290114 1188
rect 290365 1184 290412 1188
rect 290476 1186 290482 1188
rect 296713 1186 296779 1189
rect 290365 1128 290370 1184
rect 290365 1124 290412 1128
rect 290476 1126 290522 1186
rect 290598 1184 296779 1186
rect 290598 1128 296718 1184
rect 296774 1128 296779 1184
rect 290598 1126 296779 1128
rect 290476 1124 290482 1126
rect 290365 1123 290431 1124
rect 290598 1050 290658 1126
rect 296713 1123 296779 1126
rect 296846 1124 296852 1188
rect 296916 1186 296922 1188
rect 308806 1186 308812 1188
rect 296916 1126 308812 1186
rect 296916 1124 296922 1126
rect 308806 1124 308812 1126
rect 308876 1124 308882 1188
rect 308949 1186 309015 1189
rect 309961 1186 310027 1189
rect 321921 1186 321987 1189
rect 308949 1184 309794 1186
rect 308949 1128 308954 1184
rect 309010 1128 309794 1184
rect 308949 1126 309794 1128
rect 308949 1123 309015 1126
rect 287654 990 290658 1050
rect 293861 1050 293927 1053
rect 296897 1050 296963 1053
rect 293861 1048 296963 1050
rect 293861 992 293866 1048
rect 293922 992 296902 1048
rect 296958 992 296963 1048
rect 293861 990 296963 992
rect 262489 987 262555 990
rect 285673 987 285739 990
rect 293861 987 293927 990
rect 296897 987 296963 990
rect 299933 1050 299999 1053
rect 303286 1050 303292 1052
rect 299933 1048 303292 1050
rect 299933 992 299938 1048
rect 299994 992 303292 1048
rect 299933 990 303292 992
rect 299933 987 299999 990
rect 303286 988 303292 990
rect 303356 988 303362 1052
rect 303429 1050 303495 1053
rect 306925 1050 306991 1053
rect 303429 1048 306991 1050
rect 303429 992 303434 1048
rect 303490 992 306930 1048
rect 306986 992 306991 1048
rect 303429 990 306991 992
rect 303429 987 303495 990
rect 306925 987 306991 990
rect 307109 1050 307175 1053
rect 309317 1050 309383 1053
rect 307109 1048 309383 1050
rect 307109 992 307114 1048
rect 307170 992 309322 1048
rect 309378 992 309383 1048
rect 307109 990 309383 992
rect 309734 1050 309794 1126
rect 309961 1184 321987 1186
rect 309961 1128 309966 1184
rect 310022 1128 321926 1184
rect 321982 1128 321987 1184
rect 309961 1126 321987 1128
rect 309961 1123 310027 1126
rect 321921 1123 321987 1126
rect 322105 1186 322171 1189
rect 328310 1186 328316 1188
rect 322105 1184 328316 1186
rect 322105 1128 322110 1184
rect 322166 1128 328316 1184
rect 322105 1126 328316 1128
rect 322105 1123 322171 1126
rect 328310 1124 328316 1126
rect 328380 1124 328386 1188
rect 328494 1124 328500 1188
rect 328564 1186 328570 1188
rect 328821 1186 328887 1189
rect 328564 1184 328887 1186
rect 328564 1128 328826 1184
rect 328882 1128 328887 1184
rect 328564 1126 328887 1128
rect 328564 1124 328570 1126
rect 328821 1123 328887 1126
rect 329741 1186 329807 1189
rect 331765 1186 331831 1189
rect 329741 1184 331831 1186
rect 329741 1128 329746 1184
rect 329802 1128 331770 1184
rect 331826 1128 331831 1184
rect 329741 1126 331831 1128
rect 329741 1123 329807 1126
rect 331765 1123 331831 1126
rect 331949 1186 332015 1189
rect 335813 1186 335879 1189
rect 331949 1184 335879 1186
rect 331949 1128 331954 1184
rect 332010 1128 335818 1184
rect 335874 1128 335879 1184
rect 331949 1126 335879 1128
rect 331949 1123 332015 1126
rect 335813 1123 335879 1126
rect 335997 1186 336063 1189
rect 348325 1186 348391 1189
rect 335997 1184 348391 1186
rect 335997 1128 336002 1184
rect 336058 1128 348330 1184
rect 348386 1128 348391 1184
rect 335997 1126 348391 1128
rect 335997 1123 336063 1126
rect 348325 1123 348391 1126
rect 348918 1124 348924 1188
rect 348988 1186 348994 1188
rect 366173 1186 366239 1189
rect 348988 1184 366239 1186
rect 348988 1128 366178 1184
rect 366234 1128 366239 1184
rect 348988 1126 366239 1128
rect 348988 1124 348994 1126
rect 366173 1123 366239 1126
rect 370446 1124 370452 1188
rect 370516 1186 370522 1188
rect 372521 1186 372587 1189
rect 370516 1184 372587 1186
rect 370516 1128 372526 1184
rect 372582 1128 372587 1184
rect 370516 1126 372587 1128
rect 370516 1124 370522 1126
rect 372521 1123 372587 1126
rect 373717 1186 373783 1189
rect 389081 1186 389147 1189
rect 373717 1184 389147 1186
rect 373717 1128 373722 1184
rect 373778 1128 389086 1184
rect 389142 1128 389147 1184
rect 373717 1126 389147 1128
rect 373717 1123 373783 1126
rect 389081 1123 389147 1126
rect 389357 1186 389423 1189
rect 439454 1186 439514 1262
rect 443177 1259 443243 1262
rect 453297 1322 453363 1325
rect 460565 1322 460631 1325
rect 453297 1320 460631 1322
rect 453297 1264 453302 1320
rect 453358 1264 460570 1320
rect 460626 1264 460631 1320
rect 453297 1262 460631 1264
rect 453297 1259 453363 1262
rect 460565 1259 460631 1262
rect 462589 1322 462655 1325
rect 476389 1322 476455 1325
rect 462589 1320 476455 1322
rect 462589 1264 462594 1320
rect 462650 1264 476394 1320
rect 476450 1264 476455 1320
rect 462589 1262 476455 1264
rect 462589 1259 462655 1262
rect 476389 1259 476455 1262
rect 476573 1322 476639 1325
rect 482185 1322 482251 1325
rect 501321 1322 501387 1325
rect 476573 1320 482251 1322
rect 476573 1264 476578 1320
rect 476634 1264 482190 1320
rect 482246 1264 482251 1320
rect 476573 1262 482251 1264
rect 476573 1259 476639 1262
rect 482185 1259 482251 1262
rect 482326 1320 501387 1322
rect 482326 1264 501326 1320
rect 501382 1264 501387 1320
rect 482326 1262 501387 1264
rect 389357 1184 439514 1186
rect 389357 1128 389362 1184
rect 389418 1128 439514 1184
rect 389357 1126 439514 1128
rect 440693 1186 440759 1189
rect 482326 1186 482386 1262
rect 501321 1259 501387 1262
rect 504173 1322 504239 1325
rect 516685 1322 516751 1325
rect 504173 1320 516751 1322
rect 504173 1264 504178 1320
rect 504234 1264 516690 1320
rect 516746 1264 516751 1320
rect 504173 1262 516751 1264
rect 504173 1259 504239 1262
rect 516685 1259 516751 1262
rect 516869 1322 516935 1325
rect 537293 1322 537359 1325
rect 516869 1320 537359 1322
rect 516869 1264 516874 1320
rect 516930 1264 537298 1320
rect 537354 1264 537359 1320
rect 516869 1262 537359 1264
rect 516869 1259 516935 1262
rect 537293 1259 537359 1262
rect 538765 1322 538831 1325
rect 552473 1322 552539 1325
rect 559557 1322 559623 1325
rect 538765 1320 552539 1322
rect 538765 1264 538770 1320
rect 538826 1264 552478 1320
rect 552534 1264 552539 1320
rect 538765 1262 552539 1264
rect 538765 1259 538831 1262
rect 552473 1259 552539 1262
rect 552614 1320 559623 1322
rect 552614 1264 559562 1320
rect 559618 1264 559623 1320
rect 552614 1262 559623 1264
rect 440693 1184 482386 1186
rect 440693 1128 440698 1184
rect 440754 1128 482386 1184
rect 440693 1126 482386 1128
rect 389357 1123 389423 1126
rect 440693 1123 440759 1126
rect 483790 1124 483796 1188
rect 483860 1186 483866 1188
rect 514150 1186 514156 1188
rect 483860 1126 514156 1186
rect 483860 1124 483866 1126
rect 514150 1124 514156 1126
rect 514220 1124 514226 1188
rect 531773 1186 531839 1189
rect 552614 1186 552674 1262
rect 559557 1259 559623 1262
rect 564433 1322 564499 1325
rect 564934 1322 564940 1324
rect 564433 1320 564940 1322
rect 564433 1264 564438 1320
rect 564494 1264 564940 1320
rect 564433 1262 564940 1264
rect 564433 1259 564499 1262
rect 564934 1260 564940 1262
rect 565004 1260 565010 1324
rect 531773 1184 552674 1186
rect 531773 1128 531778 1184
rect 531834 1128 552674 1184
rect 531773 1126 552674 1128
rect 552749 1186 552815 1189
rect 557993 1186 558059 1189
rect 552749 1184 558059 1186
rect 552749 1128 552754 1184
rect 552810 1128 557998 1184
rect 558054 1128 558059 1184
rect 552749 1126 558059 1128
rect 531773 1123 531839 1126
rect 552749 1123 552815 1126
rect 557993 1123 558059 1126
rect 561438 1124 561444 1188
rect 561508 1186 561514 1188
rect 568389 1186 568455 1189
rect 561508 1184 568455 1186
rect 561508 1128 568394 1184
rect 568450 1128 568455 1184
rect 561508 1126 568455 1128
rect 561508 1124 561514 1126
rect 568389 1123 568455 1126
rect 326889 1050 326955 1053
rect 327073 1052 327139 1053
rect 309734 1048 326955 1050
rect 309734 992 326894 1048
rect 326950 992 326955 1048
rect 309734 990 326955 992
rect 307109 987 307175 990
rect 309317 987 309383 990
rect 326889 987 326955 990
rect 327022 988 327028 1052
rect 327092 1050 327139 1052
rect 327257 1050 327323 1053
rect 568665 1050 568731 1053
rect 327092 1048 327184 1050
rect 327134 992 327184 1048
rect 327092 990 327184 992
rect 327257 1048 568731 1050
rect 327257 992 327262 1048
rect 327318 992 568670 1048
rect 568726 992 568731 1048
rect 327257 990 568731 992
rect 327092 988 327139 990
rect 327073 987 327139 988
rect 327257 987 327323 990
rect 568665 987 568731 990
rect 250364 854 251834 914
rect 250364 852 250370 854
rect 251950 852 251956 916
rect 252020 914 252026 916
rect 252461 914 252527 917
rect 252020 912 252527 914
rect 252020 856 252466 912
rect 252522 856 252527 912
rect 252020 854 252527 856
rect 252020 852 252026 854
rect 252461 851 252527 854
rect 252921 914 252987 917
rect 253657 914 253723 917
rect 252921 912 253723 914
rect 252921 856 252926 912
rect 252982 856 253662 912
rect 253718 856 253723 912
rect 252921 854 253723 856
rect 252921 851 252987 854
rect 253657 851 253723 854
rect 253790 852 253796 916
rect 253860 914 253866 916
rect 255630 914 255636 916
rect 253860 854 255636 914
rect 253860 852 253866 854
rect 255630 852 255636 854
rect 255700 852 255706 916
rect 309777 914 309843 917
rect 255822 912 309843 914
rect 255822 856 309782 912
rect 309838 856 309843 912
rect 255822 854 309843 856
rect 198406 778 198412 780
rect 197862 718 198412 778
rect 190453 715 190519 718
rect 197537 715 197603 718
rect 198406 716 198412 718
rect 198476 716 198482 780
rect 198641 778 198707 781
rect 221089 778 221155 781
rect 224401 778 224467 781
rect 198641 776 221155 778
rect 198641 720 198646 776
rect 198702 720 221094 776
rect 221150 720 221155 776
rect 198641 718 221155 720
rect 198641 715 198707 718
rect 221089 715 221155 718
rect 221230 776 224467 778
rect 221230 720 224406 776
rect 224462 720 224467 776
rect 221230 718 224467 720
rect 158069 640 161674 642
rect 158069 584 158074 640
rect 158130 584 161674 640
rect 158069 582 161674 584
rect 161749 642 161815 645
rect 163497 642 163563 645
rect 161749 640 163563 642
rect 161749 584 161754 640
rect 161810 584 163502 640
rect 163558 584 163563 640
rect 161749 582 163563 584
rect 157885 579 157951 580
rect 158069 579 158135 582
rect 161749 579 161815 582
rect 163497 579 163563 582
rect 163630 580 163636 644
rect 163700 642 163706 644
rect 169661 642 169727 645
rect 169845 644 169911 645
rect 169845 642 169892 644
rect 163700 640 169727 642
rect 163700 584 169666 640
rect 169722 584 169727 640
rect 163700 582 169727 584
rect 169800 640 169892 642
rect 169800 584 169850 640
rect 169800 582 169892 584
rect 163700 580 163706 582
rect 169661 579 169727 582
rect 169845 580 169892 582
rect 169956 580 169962 644
rect 170029 642 170095 645
rect 175038 642 175044 644
rect 170029 640 175044 642
rect 170029 584 170034 640
rect 170090 584 175044 640
rect 170029 582 175044 584
rect 169845 579 169911 580
rect 170029 579 170095 582
rect 175038 580 175044 582
rect 175108 580 175114 644
rect 175406 580 175412 644
rect 175476 642 175482 644
rect 177246 642 177252 644
rect 175476 582 177252 642
rect 175476 580 175482 582
rect 177246 580 177252 582
rect 177316 580 177322 644
rect 177389 642 177455 645
rect 177798 642 177804 644
rect 177389 640 177804 642
rect 177389 584 177394 640
rect 177450 584 177804 640
rect 177389 582 177804 584
rect 177389 579 177455 582
rect 177798 580 177804 582
rect 177868 580 177874 644
rect 177941 642 178007 645
rect 197353 642 197419 645
rect 177941 640 197419 642
rect 177941 584 177946 640
rect 178002 584 197358 640
rect 197414 584 197419 640
rect 177941 582 197419 584
rect 177941 579 178007 582
rect 197353 579 197419 582
rect 198457 642 198523 645
rect 204110 642 204116 644
rect 198457 640 204116 642
rect 198457 584 198462 640
rect 198518 584 204116 640
rect 198457 582 204116 584
rect 198457 579 198523 582
rect 204110 580 204116 582
rect 204180 580 204186 644
rect 204253 642 204319 645
rect 204529 642 204595 645
rect 204253 640 204595 642
rect 204253 584 204258 640
rect 204314 584 204534 640
rect 204590 584 204595 640
rect 204253 582 204595 584
rect 204253 579 204319 582
rect 204529 579 204595 582
rect 204662 580 204668 644
rect 204732 642 204738 644
rect 205081 642 205147 645
rect 204732 640 205147 642
rect 204732 584 205086 640
rect 205142 584 205147 640
rect 204732 582 205147 584
rect 204732 580 204738 582
rect 205081 579 205147 582
rect 205214 580 205220 644
rect 205284 642 205290 644
rect 207841 642 207907 645
rect 205284 640 207907 642
rect 205284 584 207846 640
rect 207902 584 207907 640
rect 205284 582 207907 584
rect 205284 580 205290 582
rect 207841 579 207907 582
rect 207974 580 207980 644
rect 208044 642 208050 644
rect 210366 642 210372 644
rect 208044 582 210372 642
rect 208044 580 208050 582
rect 210366 580 210372 582
rect 210436 580 210442 644
rect 210550 580 210556 644
rect 210620 642 210626 644
rect 211286 642 211292 644
rect 210620 582 211292 642
rect 210620 580 210626 582
rect 211286 580 211292 582
rect 211356 580 211362 644
rect 211429 642 211495 645
rect 215017 642 215083 645
rect 211429 640 215083 642
rect 211429 584 211434 640
rect 211490 584 215022 640
rect 215078 584 215083 640
rect 211429 582 215083 584
rect 211429 579 211495 582
rect 215017 579 215083 582
rect 215201 642 215267 645
rect 217777 642 217843 645
rect 215201 640 217843 642
rect 215201 584 215206 640
rect 215262 584 217782 640
rect 217838 584 217843 640
rect 215201 582 217843 584
rect 215201 579 215267 582
rect 217777 579 217843 582
rect 217961 642 218027 645
rect 219198 642 219204 644
rect 217961 640 219204 642
rect 217961 584 217966 640
rect 218022 584 219204 640
rect 217961 582 219204 584
rect 217961 579 218027 582
rect 219198 580 219204 582
rect 219268 580 219274 644
rect 219341 642 219407 645
rect 221230 642 221290 718
rect 224401 715 224467 718
rect 224585 778 224651 781
rect 231158 778 231164 780
rect 224585 776 231164 778
rect 224585 720 224590 776
rect 224646 720 231164 776
rect 224585 718 231164 720
rect 224585 715 224651 718
rect 231158 716 231164 718
rect 231228 716 231234 780
rect 231301 778 231367 781
rect 238201 778 238267 781
rect 231301 776 238267 778
rect 231301 720 231306 776
rect 231362 720 238206 776
rect 238262 720 238267 776
rect 231301 718 238267 720
rect 231301 715 231367 718
rect 238201 715 238267 718
rect 238385 778 238451 781
rect 239121 778 239187 781
rect 238385 776 239187 778
rect 238385 720 238390 776
rect 238446 720 239126 776
rect 239182 720 239187 776
rect 238385 718 239187 720
rect 238385 715 238451 718
rect 239121 715 239187 718
rect 239305 778 239371 781
rect 245009 778 245075 781
rect 239305 776 245075 778
rect 239305 720 239310 776
rect 239366 720 245014 776
rect 245070 720 245075 776
rect 239305 718 245075 720
rect 239305 715 239371 718
rect 245009 715 245075 718
rect 245142 716 245148 780
rect 245212 778 245218 780
rect 246430 778 246436 780
rect 245212 718 246436 778
rect 245212 716 245218 718
rect 246430 716 246436 718
rect 246500 716 246506 780
rect 246614 716 246620 780
rect 246684 778 246690 780
rect 247861 778 247927 781
rect 252318 778 252324 780
rect 246684 718 247786 778
rect 246684 716 246690 718
rect 219341 640 221290 642
rect 219341 584 219346 640
rect 219402 584 221290 640
rect 219341 582 221290 584
rect 221365 642 221431 645
rect 232957 642 233023 645
rect 221365 640 233023 642
rect 221365 584 221370 640
rect 221426 584 232962 640
rect 233018 584 233023 640
rect 221365 582 233023 584
rect 219341 579 219407 582
rect 221365 579 221431 582
rect 232957 579 233023 582
rect 233141 642 233207 645
rect 247585 642 247651 645
rect 233141 640 247651 642
rect 233141 584 233146 640
rect 233202 584 247590 640
rect 247646 584 247651 640
rect 233141 582 247651 584
rect 247726 642 247786 718
rect 247861 776 252324 778
rect 247861 720 247866 776
rect 247922 720 252324 776
rect 247861 718 252324 720
rect 247861 715 247927 718
rect 252318 716 252324 718
rect 252388 716 252394 780
rect 252502 716 252508 780
rect 252572 778 252578 780
rect 255822 778 255882 854
rect 309777 851 309843 854
rect 309910 852 309916 916
rect 309980 914 309986 916
rect 314745 914 314811 917
rect 328545 916 328611 917
rect 309980 912 314811 914
rect 309980 856 314750 912
rect 314806 856 314811 912
rect 309980 854 314811 856
rect 309980 852 309986 854
rect 314745 851 314811 854
rect 314878 852 314884 916
rect 314948 914 314954 916
rect 328310 914 328316 916
rect 314948 854 328316 914
rect 314948 852 314954 854
rect 328310 852 328316 854
rect 328380 852 328386 916
rect 328540 852 328546 916
rect 328610 914 328616 916
rect 328610 854 328702 914
rect 328610 852 328616 854
rect 329046 852 329052 916
rect 329116 914 329122 916
rect 329649 914 329715 917
rect 329116 912 329715 914
rect 329116 856 329654 912
rect 329710 856 329715 912
rect 329116 854 329715 856
rect 329116 852 329122 854
rect 328545 851 328611 852
rect 329649 851 329715 854
rect 329833 914 329899 917
rect 335997 914 336063 917
rect 329833 912 336063 914
rect 329833 856 329838 912
rect 329894 856 336002 912
rect 336058 856 336063 912
rect 329833 854 336063 856
rect 329833 851 329899 854
rect 335997 851 336063 854
rect 336181 914 336247 917
rect 349521 914 349587 917
rect 336181 912 349587 914
rect 336181 856 336186 912
rect 336242 856 349526 912
rect 349582 856 349587 912
rect 336181 854 349587 856
rect 336181 851 336247 854
rect 349521 851 349587 854
rect 352189 914 352255 917
rect 356237 914 356303 917
rect 352189 912 356303 914
rect 352189 856 352194 912
rect 352250 856 356242 912
rect 356298 856 356303 912
rect 352189 854 356303 856
rect 352189 851 352255 854
rect 356237 851 356303 854
rect 356421 914 356487 917
rect 356421 912 357818 914
rect 356421 856 356426 912
rect 356482 856 357818 912
rect 356421 854 357818 856
rect 356421 851 356487 854
rect 252572 718 255882 778
rect 255957 778 256023 781
rect 258206 778 258212 780
rect 255957 776 258212 778
rect 255957 720 255962 776
rect 256018 720 258212 776
rect 255957 718 258212 720
rect 252572 716 252578 718
rect 255957 715 256023 718
rect 258206 716 258212 718
rect 258276 716 258282 780
rect 258349 778 258415 781
rect 260833 780 260899 781
rect 260230 778 260236 780
rect 258349 776 260236 778
rect 258349 720 258354 776
rect 258410 720 260236 776
rect 258349 718 260236 720
rect 258349 715 258415 718
rect 260230 716 260236 718
rect 260300 716 260306 780
rect 260782 778 260788 780
rect 260742 718 260788 778
rect 260852 776 260899 780
rect 260894 720 260899 776
rect 260782 716 260788 718
rect 260852 716 260899 720
rect 261150 716 261156 780
rect 261220 778 261226 780
rect 261845 778 261911 781
rect 262673 778 262739 781
rect 261220 718 261770 778
rect 261220 716 261226 718
rect 260833 715 260899 716
rect 248270 642 248276 644
rect 247726 582 248276 642
rect 233141 579 233207 582
rect 247585 579 247651 582
rect 248270 580 248276 582
rect 248340 580 248346 644
rect 248413 642 248479 645
rect 261569 642 261635 645
rect 248413 640 261635 642
rect 248413 584 248418 640
rect 248474 584 261574 640
rect 261630 584 261635 640
rect 248413 582 261635 584
rect 261710 642 261770 718
rect 261845 776 262739 778
rect 261845 720 261850 776
rect 261906 720 262678 776
rect 262734 720 262739 776
rect 261845 718 262739 720
rect 261845 715 261911 718
rect 262673 715 262739 718
rect 262857 778 262923 781
rect 265985 778 266051 781
rect 262857 776 266051 778
rect 262857 720 262862 776
rect 262918 720 265990 776
rect 266046 720 266051 776
rect 262857 718 266051 720
rect 262857 715 262923 718
rect 265985 715 266051 718
rect 266261 778 266327 781
rect 271045 778 271111 781
rect 266261 776 271111 778
rect 266261 720 266266 776
rect 266322 720 271050 776
rect 271106 720 271111 776
rect 266261 718 271111 720
rect 266261 715 266327 718
rect 271045 715 271111 718
rect 271229 778 271295 781
rect 279877 778 279943 781
rect 271229 776 279943 778
rect 271229 720 271234 776
rect 271290 720 279882 776
rect 279938 720 279943 776
rect 271229 718 279943 720
rect 271229 715 271295 718
rect 279877 715 279943 718
rect 280102 716 280108 780
rect 280172 778 280178 780
rect 280245 778 280311 781
rect 280172 776 280311 778
rect 280172 720 280250 776
rect 280306 720 280311 776
rect 280172 718 280311 720
rect 280172 716 280178 718
rect 280245 715 280311 718
rect 280654 716 280660 780
rect 280724 778 280730 780
rect 281901 778 281967 781
rect 280724 776 281967 778
rect 280724 720 281906 776
rect 281962 720 281967 776
rect 280724 718 281967 720
rect 280724 716 280730 718
rect 281901 715 281967 718
rect 282085 778 282151 781
rect 285305 778 285371 781
rect 282085 776 285371 778
rect 282085 720 282090 776
rect 282146 720 285310 776
rect 285366 720 285371 776
rect 282085 718 285371 720
rect 282085 715 282151 718
rect 285305 715 285371 718
rect 285765 778 285831 781
rect 290365 778 290431 781
rect 294781 780 294847 781
rect 294781 778 294828 780
rect 285765 776 290431 778
rect 285765 720 285770 776
rect 285826 720 290370 776
rect 290426 720 290431 776
rect 285765 718 290431 720
rect 294736 776 294828 778
rect 294736 720 294786 776
rect 294736 718 294828 720
rect 285765 715 285831 718
rect 290365 715 290431 718
rect 294781 716 294828 718
rect 294892 716 294898 780
rect 295241 778 295307 781
rect 348693 778 348759 781
rect 353886 778 353892 780
rect 295241 776 348759 778
rect 295241 720 295246 776
rect 295302 720 348698 776
rect 348754 720 348759 776
rect 295241 718 348759 720
rect 294781 715 294847 716
rect 295241 715 295307 718
rect 348693 715 348759 718
rect 349846 718 353892 778
rect 262581 642 262647 645
rect 261710 640 262647 642
rect 261710 584 262586 640
rect 262642 584 262647 640
rect 261710 582 262647 584
rect 248413 579 248479 582
rect 261569 579 261635 582
rect 262581 579 262647 582
rect 264830 580 264836 644
rect 264900 642 264906 644
rect 266813 642 266879 645
rect 264900 640 266879 642
rect 264900 584 266818 640
rect 266874 584 266879 640
rect 264900 582 266879 584
rect 264900 580 264906 582
rect 266813 579 266879 582
rect 266997 642 267063 645
rect 336181 642 336247 645
rect 266997 640 336247 642
rect 266997 584 267002 640
rect 267058 584 336186 640
rect 336242 584 336247 640
rect 266997 582 336247 584
rect 266997 579 267063 582
rect 336181 579 336247 582
rect 336365 642 336431 645
rect 338614 642 338620 644
rect 336365 640 338620 642
rect 336365 584 336370 640
rect 336426 584 338620 640
rect 336365 582 338620 584
rect 336365 579 336431 582
rect 338614 580 338620 582
rect 338684 580 338690 644
rect 338798 580 338804 644
rect 338868 642 338874 644
rect 342662 642 342668 644
rect 338868 582 342668 642
rect 338868 580 338874 582
rect 342662 580 342668 582
rect 342732 580 342738 644
rect 343081 642 343147 645
rect 349846 642 349906 718
rect 353886 716 353892 718
rect 353956 716 353962 780
rect 354029 778 354095 781
rect 357617 778 357683 781
rect 354029 776 357683 778
rect 354029 720 354034 776
rect 354090 720 357622 776
rect 357678 720 357683 776
rect 354029 718 357683 720
rect 357758 778 357818 854
rect 358118 852 358124 916
rect 358188 914 358194 916
rect 564566 914 564572 916
rect 358188 854 564572 914
rect 358188 852 358194 854
rect 564566 852 564572 854
rect 564636 852 564642 916
rect 362718 778 362724 780
rect 357758 718 362724 778
rect 354029 715 354095 718
rect 357617 715 357683 718
rect 362718 716 362724 718
rect 362788 716 362794 780
rect 364701 778 364767 781
rect 373349 778 373415 781
rect 364701 776 373415 778
rect 364701 720 364706 776
rect 364762 720 373354 776
rect 373410 720 373415 776
rect 364701 718 373415 720
rect 364701 715 364767 718
rect 373349 715 373415 718
rect 376753 778 376819 781
rect 381537 778 381603 781
rect 376753 776 381603 778
rect 376753 720 376758 776
rect 376814 720 381542 776
rect 381598 720 381603 776
rect 376753 718 381603 720
rect 376753 715 376819 718
rect 381537 715 381603 718
rect 385902 716 385908 780
rect 385972 778 385978 780
rect 406101 778 406167 781
rect 385972 776 406167 778
rect 385972 720 406106 776
rect 406162 720 406167 776
rect 385972 718 406167 720
rect 385972 716 385978 718
rect 406101 715 406167 718
rect 406377 778 406443 781
rect 434989 778 435055 781
rect 406377 776 435055 778
rect 406377 720 406382 776
rect 406438 720 434994 776
rect 435050 720 435055 776
rect 406377 718 435055 720
rect 406377 715 406443 718
rect 434989 715 435055 718
rect 440182 716 440188 780
rect 440252 778 440258 780
rect 449750 778 449756 780
rect 440252 718 449756 778
rect 440252 716 440258 718
rect 449750 716 449756 718
rect 449820 716 449826 780
rect 460565 778 460631 781
rect 476573 778 476639 781
rect 460565 776 476639 778
rect 460565 720 460570 776
rect 460626 720 476578 776
rect 476634 720 476639 776
rect 460565 718 476639 720
rect 460565 715 460631 718
rect 476573 715 476639 718
rect 482185 778 482251 781
rect 504173 778 504239 781
rect 482185 776 504239 778
rect 482185 720 482190 776
rect 482246 720 504178 776
rect 504234 720 504239 776
rect 482185 718 504239 720
rect 482185 715 482251 718
rect 504173 715 504239 718
rect 512637 778 512703 781
rect 515581 778 515647 781
rect 512637 776 515647 778
rect 512637 720 512642 776
rect 512698 720 515586 776
rect 515642 720 515647 776
rect 512637 718 515647 720
rect 512637 715 512703 718
rect 515581 715 515647 718
rect 516685 778 516751 781
rect 531773 778 531839 781
rect 516685 776 531839 778
rect 516685 720 516690 776
rect 516746 720 531778 776
rect 531834 720 531839 776
rect 516685 718 531839 720
rect 516685 715 516751 718
rect 531773 715 531839 718
rect 536925 778 536991 781
rect 539542 778 539548 780
rect 536925 776 539548 778
rect 536925 720 536930 776
rect 536986 720 539548 776
rect 536925 718 539548 720
rect 536925 715 536991 718
rect 539542 716 539548 718
rect 539612 716 539618 780
rect 559557 778 559623 781
rect 563094 778 563100 780
rect 559557 776 563100 778
rect 559557 720 559562 776
rect 559618 720 563100 776
rect 559557 718 563100 720
rect 559557 715 559623 718
rect 563094 716 563100 718
rect 563164 716 563170 780
rect 569125 778 569191 781
rect 569125 776 569234 778
rect 569125 720 569130 776
rect 569186 720 569234 776
rect 569125 715 569234 720
rect 343081 640 349906 642
rect 343081 584 343086 640
rect 343142 584 349906 640
rect 343081 582 349906 584
rect 343081 579 343147 582
rect 350022 580 350028 644
rect 350092 642 350098 644
rect 356513 642 356579 645
rect 350092 640 356579 642
rect 350092 584 356518 640
rect 356574 584 356579 640
rect 350092 582 356579 584
rect 350092 580 350098 582
rect 356513 579 356579 582
rect 356973 642 357039 645
rect 365069 642 365135 645
rect 356973 640 365135 642
rect 356973 584 356978 640
rect 357034 584 365074 640
rect 365130 584 365135 640
rect 356973 582 365135 584
rect 356973 579 357039 582
rect 365069 579 365135 582
rect 365253 642 365319 645
rect 380341 642 380407 645
rect 365253 640 380407 642
rect 365253 584 365258 640
rect 365314 584 380346 640
rect 380402 584 380407 640
rect 365253 582 380407 584
rect 365253 579 365319 582
rect 380341 579 380407 582
rect 386045 642 386111 645
rect 390502 642 390508 644
rect 386045 640 390508 642
rect 386045 584 386050 640
rect 386106 584 390508 640
rect 386045 582 390508 584
rect 386045 579 386111 582
rect 390502 580 390508 582
rect 390572 580 390578 644
rect 393405 642 393471 645
rect 411253 642 411319 645
rect 393405 640 411319 642
rect 393405 584 393410 640
rect 393466 584 411258 640
rect 411314 584 411319 640
rect 393405 582 411319 584
rect 393405 579 393471 582
rect 411253 579 411319 582
rect 415117 642 415183 645
rect 427813 642 427879 645
rect 415117 640 427879 642
rect 415117 584 415122 640
rect 415178 584 427818 640
rect 427874 584 427879 640
rect 415117 582 427879 584
rect 415117 579 415183 582
rect 427813 579 427879 582
rect 430614 580 430620 644
rect 430684 642 430690 644
rect 434478 642 434484 644
rect 430684 582 434484 642
rect 430684 580 430690 582
rect 434478 580 434484 582
rect 434548 580 434554 644
rect 442809 642 442875 645
rect 476757 642 476823 645
rect 442809 640 476823 642
rect 442809 584 442814 640
rect 442870 584 476762 640
rect 476818 584 476823 640
rect 442809 582 476823 584
rect 442809 579 442875 582
rect 476757 579 476823 582
rect 490189 642 490255 645
rect 509049 642 509115 645
rect 522573 642 522639 645
rect 536741 642 536807 645
rect 559782 642 559788 644
rect 490189 640 509115 642
rect 490189 584 490194 640
rect 490250 584 509054 640
rect 509110 584 509115 640
rect 490189 582 509115 584
rect 490189 579 490255 582
rect 509049 579 509115 582
rect 512686 582 522498 642
rect 156873 506 156939 509
rect 150942 504 156939 506
rect 150942 448 156878 504
rect 156934 448 156939 504
rect 150942 446 156939 448
rect 150801 443 150867 444
rect 156873 443 156939 446
rect 157149 506 157215 509
rect 190637 506 190703 509
rect 157149 504 190703 506
rect 157149 448 157154 504
rect 157210 448 190642 504
rect 190698 448 190703 504
rect 157149 446 190703 448
rect 157149 443 157215 446
rect 190637 443 190703 446
rect 190862 444 190868 508
rect 190932 506 190938 508
rect 191281 506 191347 509
rect 190932 504 191347 506
rect 190932 448 191286 504
rect 191342 448 191347 504
rect 190932 446 191347 448
rect 190932 444 190938 446
rect 191281 443 191347 446
rect 191414 444 191420 508
rect 191484 506 191490 508
rect 197118 506 197124 508
rect 191484 446 197124 506
rect 191484 444 191490 446
rect 197118 444 197124 446
rect 197188 444 197194 508
rect 197629 506 197695 509
rect 198181 508 198247 509
rect 197854 506 197860 508
rect 197629 504 197860 506
rect 197629 448 197634 504
rect 197690 448 197860 504
rect 197629 446 197860 448
rect 197629 443 197695 446
rect 197854 444 197860 446
rect 197924 444 197930 508
rect 198181 506 198228 508
rect 198136 504 198228 506
rect 198136 448 198186 504
rect 198136 446 198228 448
rect 198181 444 198228 446
rect 198292 444 198298 508
rect 198365 506 198431 509
rect 442717 506 442783 509
rect 198365 504 442783 506
rect 198365 448 198370 504
rect 198426 448 442722 504
rect 442778 448 442783 504
rect 198365 446 442783 448
rect 198181 443 198247 444
rect 198365 443 198431 446
rect 442717 443 442783 446
rect 462998 444 463004 508
rect 463068 506 463074 508
rect 469070 506 469076 508
rect 463068 446 469076 506
rect 463068 444 463074 446
rect 469070 444 469076 446
rect 469140 444 469146 508
rect 473486 444 473492 508
rect 473556 506 473562 508
rect 509877 506 509943 509
rect 473556 504 509943 506
rect 473556 448 509882 504
rect 509938 448 509943 504
rect 473556 446 509943 448
rect 473556 444 473562 446
rect 509877 443 509943 446
rect 122790 310 123218 370
rect 123293 370 123359 373
rect 153101 370 153167 373
rect 123293 368 153167 370
rect 123293 312 123298 368
rect 123354 312 153106 368
rect 153162 312 153167 368
rect 123293 310 153167 312
rect 92657 307 92723 310
rect 122649 307 122715 310
rect 123293 307 123359 310
rect 153101 307 153167 310
rect 153285 370 153351 373
rect 156873 370 156939 373
rect 153285 368 156939 370
rect 153285 312 153290 368
rect 153346 312 156878 368
rect 156934 312 156939 368
rect 153285 310 156939 312
rect 153285 307 153351 310
rect 156873 307 156939 310
rect 157333 370 157399 373
rect 157793 370 157859 373
rect 157333 368 157859 370
rect 157333 312 157338 368
rect 157394 312 157798 368
rect 157854 312 157859 368
rect 157333 310 157859 312
rect 157333 307 157399 310
rect 157793 307 157859 310
rect 157926 308 157932 372
rect 157996 370 158002 372
rect 161238 370 161244 372
rect 157996 310 161244 370
rect 157996 308 158002 310
rect 161238 308 161244 310
rect 161308 308 161314 372
rect 161381 370 161447 373
rect 163129 370 163195 373
rect 161381 368 163195 370
rect 161381 312 161386 368
rect 161442 312 163134 368
rect 163190 312 163195 368
rect 161381 310 163195 312
rect 161381 307 161447 310
rect 163129 307 163195 310
rect 163313 370 163379 373
rect 224309 370 224375 373
rect 163313 368 224375 370
rect 163313 312 163318 368
rect 163374 312 224314 368
rect 224370 312 224375 368
rect 163313 310 224375 312
rect 163313 307 163379 310
rect 224309 307 224375 310
rect 224677 370 224743 373
rect 248321 370 248387 373
rect 224677 368 248387 370
rect 224677 312 224682 368
rect 224738 312 248326 368
rect 248382 312 248387 368
rect 224677 310 248387 312
rect 224677 307 224743 310
rect 248321 307 248387 310
rect 248781 370 248847 373
rect 290774 370 290780 372
rect 248781 368 290780 370
rect 248781 312 248786 368
rect 248842 312 290780 368
rect 248781 310 290780 312
rect 248781 307 248847 310
rect 290774 308 290780 310
rect 290844 308 290850 372
rect 291142 308 291148 372
rect 291212 370 291218 372
rect 358169 370 358235 373
rect 291212 368 358235 370
rect 291212 312 358174 368
rect 358230 312 358235 368
rect 291212 310 358235 312
rect 291212 308 291218 310
rect 358169 307 358235 310
rect 365069 370 365135 373
rect 386045 370 386111 373
rect 365069 368 386111 370
rect 365069 312 365074 368
rect 365130 312 386050 368
rect 386106 312 386111 368
rect 365069 310 386111 312
rect 365069 307 365135 310
rect 386045 307 386111 310
rect 390502 308 390508 372
rect 390572 370 390578 372
rect 406377 370 406443 373
rect 390572 368 406443 370
rect 390572 312 406382 368
rect 406438 312 406443 368
rect 390572 310 406443 312
rect 390572 308 390578 310
rect 406377 307 406443 310
rect 406653 370 406719 373
rect 413645 370 413711 373
rect 406653 368 413711 370
rect 406653 312 406658 368
rect 406714 312 413650 368
rect 413706 312 413711 368
rect 406653 310 413711 312
rect 406653 307 406719 310
rect 413645 307 413711 310
rect 418838 308 418844 372
rect 418908 370 418914 372
rect 422150 370 422156 372
rect 418908 310 422156 370
rect 418908 308 418914 310
rect 422150 308 422156 310
rect 422220 308 422226 372
rect 425697 370 425763 373
rect 426934 370 426940 372
rect 425697 368 426940 370
rect 425697 312 425702 368
rect 425758 312 426940 368
rect 425697 310 426940 312
rect 425697 307 425763 310
rect 426934 308 426940 310
rect 427004 308 427010 372
rect 427813 370 427879 373
rect 442942 370 442948 372
rect 427813 368 442948 370
rect 427813 312 427818 368
rect 427874 312 442948 368
rect 427813 310 442948 312
rect 427813 307 427879 310
rect 442942 308 442948 310
rect 443012 308 443018 372
rect 443177 370 443243 373
rect 473118 370 473124 372
rect 443177 368 473124 370
rect 443177 312 443182 368
rect 443238 312 473124 368
rect 443177 310 473124 312
rect 443177 307 443243 310
rect 473118 308 473124 310
rect 473188 308 473194 372
rect 476798 308 476804 372
rect 476868 370 476874 372
rect 490598 370 490604 372
rect 476868 310 490604 370
rect 476868 308 476874 310
rect 490598 308 490604 310
rect 490668 308 490674 372
rect 512686 370 512746 582
rect 522246 506 522252 508
rect 504222 310 512746 370
rect 512870 446 522252 506
rect 66713 234 66779 237
rect 65198 232 66779 234
rect 65198 176 66718 232
rect 66774 176 66779 232
rect 65198 174 66779 176
rect 61377 171 61443 174
rect 64413 171 64479 174
rect 66713 171 66779 174
rect 66897 234 66963 237
rect 73521 234 73587 237
rect 73838 234 73844 236
rect 66897 232 73587 234
rect 66897 176 66902 232
rect 66958 176 73526 232
rect 73582 176 73587 232
rect 66897 174 73587 176
rect 66897 171 66963 174
rect 73521 171 73587 174
rect 73662 174 73844 234
rect 1894 36 1900 100
rect 1964 98 1970 100
rect 9857 98 9923 101
rect 1964 96 9923 98
rect 1964 40 9862 96
rect 9918 40 9923 96
rect 1964 38 9923 40
rect 1964 36 1970 38
rect 9857 35 9923 38
rect 10225 98 10291 101
rect 73662 98 73722 174
rect 73838 172 73844 174
rect 73908 172 73914 236
rect 74073 234 74139 237
rect 77661 234 77727 237
rect 74073 232 77727 234
rect 74073 176 74078 232
rect 74134 176 77666 232
rect 77722 176 77727 232
rect 74073 174 77727 176
rect 74073 171 74139 174
rect 77661 171 77727 174
rect 78213 234 78279 237
rect 82169 234 82235 237
rect 78213 232 82235 234
rect 78213 176 78218 232
rect 78274 176 82174 232
rect 82230 176 82235 232
rect 78213 174 82235 176
rect 78213 171 78279 174
rect 82169 171 82235 174
rect 82302 172 82308 236
rect 82372 234 82378 236
rect 84193 234 84259 237
rect 82372 232 84259 234
rect 82372 176 84198 232
rect 84254 176 84259 232
rect 82372 174 84259 176
rect 82372 172 82378 174
rect 84193 171 84259 174
rect 84377 234 84443 237
rect 85430 234 85436 236
rect 84377 232 85436 234
rect 84377 176 84382 232
rect 84438 176 85436 232
rect 84377 174 85436 176
rect 84377 171 84443 174
rect 85430 172 85436 174
rect 85500 172 85506 236
rect 85614 172 85620 236
rect 85684 234 85690 236
rect 87270 234 87276 236
rect 85684 174 87276 234
rect 85684 172 85690 174
rect 87270 172 87276 174
rect 87340 172 87346 236
rect 87505 234 87571 237
rect 92974 234 92980 236
rect 87505 232 92980 234
rect 87505 176 87510 232
rect 87566 176 92980 232
rect 87505 174 92980 176
rect 87505 171 87571 174
rect 92974 172 92980 174
rect 93044 172 93050 236
rect 93158 172 93164 236
rect 93228 234 93234 236
rect 93577 234 93643 237
rect 93228 232 93643 234
rect 93228 176 93582 232
rect 93638 176 93643 232
rect 93228 174 93643 176
rect 93228 172 93234 174
rect 93577 171 93643 174
rect 93761 234 93827 237
rect 93894 234 93900 236
rect 93761 232 93900 234
rect 93761 176 93766 232
rect 93822 176 93900 232
rect 93761 174 93900 176
rect 93761 171 93827 174
rect 93894 172 93900 174
rect 93964 172 93970 236
rect 94262 172 94268 236
rect 94332 234 94338 236
rect 97809 234 97875 237
rect 94332 232 97875 234
rect 94332 176 97814 232
rect 97870 176 97875 232
rect 94332 174 97875 176
rect 94332 172 94338 174
rect 97809 171 97875 174
rect 98269 234 98335 237
rect 108941 234 109007 237
rect 111701 234 111767 237
rect 116577 234 116643 237
rect 98269 232 108866 234
rect 98269 176 98274 232
rect 98330 176 108866 232
rect 98269 174 108866 176
rect 98269 171 98335 174
rect 10225 96 73722 98
rect 10225 40 10230 96
rect 10286 40 73722 96
rect 10225 38 73722 40
rect 73889 98 73955 101
rect 74206 98 74212 100
rect 73889 96 74212 98
rect 73889 40 73894 96
rect 73950 40 74212 96
rect 73889 38 74212 40
rect 10225 35 10291 38
rect 73889 35 73955 38
rect 74206 36 74212 38
rect 74276 36 74282 100
rect 74533 98 74599 101
rect 78622 98 78628 100
rect 74533 96 78628 98
rect 74533 40 74538 96
rect 74594 40 78628 96
rect 74533 38 78628 40
rect 74533 35 74599 38
rect 78622 36 78628 38
rect 78692 36 78698 100
rect 78857 98 78923 101
rect 81382 98 81388 100
rect 78857 96 81388 98
rect 78857 40 78862 96
rect 78918 40 81388 96
rect 78857 38 81388 40
rect 78857 35 78923 38
rect 81382 36 81388 38
rect 81452 36 81458 100
rect 81617 98 81683 101
rect 82905 98 82971 101
rect 81617 96 82971 98
rect 81617 40 81622 96
rect 81678 40 82910 96
rect 82966 40 82971 96
rect 81617 38 82971 40
rect 81617 35 81683 38
rect 82905 35 82971 38
rect 83038 36 83044 100
rect 83108 98 83114 100
rect 84193 98 84259 101
rect 83108 96 84259 98
rect 83108 40 84198 96
rect 84254 40 84259 96
rect 83108 38 84259 40
rect 83108 36 83114 38
rect 84193 35 84259 38
rect 84326 36 84332 100
rect 84396 98 84402 100
rect 89662 98 89668 100
rect 84396 38 89668 98
rect 84396 36 84402 38
rect 89662 36 89668 38
rect 89732 36 89738 100
rect 92606 36 92612 100
rect 92676 98 92682 100
rect 93853 98 93919 101
rect 92676 96 93919 98
rect 92676 40 93858 96
rect 93914 40 93919 96
rect 92676 38 93919 40
rect 92676 36 92682 38
rect 93853 35 93919 38
rect 94129 98 94195 101
rect 101029 98 101095 101
rect 94129 96 101095 98
rect 94129 40 94134 96
rect 94190 40 101034 96
rect 101090 40 101095 96
rect 94129 38 101095 40
rect 94129 35 94195 38
rect 101029 35 101095 38
rect 101438 36 101444 100
rect 101508 98 101514 100
rect 101765 98 101831 101
rect 101508 96 101831 98
rect 101508 40 101770 96
rect 101826 40 101831 96
rect 101508 38 101831 40
rect 101508 36 101514 38
rect 101765 35 101831 38
rect 101949 98 102015 101
rect 108573 98 108639 101
rect 101949 96 108639 98
rect 101949 40 101954 96
rect 102010 40 108578 96
rect 108634 40 108639 96
rect 101949 38 108639 40
rect 108806 98 108866 174
rect 108941 232 111767 234
rect 108941 176 108946 232
rect 109002 176 111706 232
rect 111762 176 111767 232
rect 108941 174 111767 176
rect 108941 171 109007 174
rect 111701 171 111767 174
rect 111888 232 116643 234
rect 111888 176 116582 232
rect 116638 176 116643 232
rect 111888 174 116643 176
rect 111888 98 111948 174
rect 116577 171 116643 174
rect 116710 172 116716 236
rect 116780 172 116786 236
rect 116853 234 116919 237
rect 150985 234 151051 237
rect 116853 232 151051 234
rect 116853 176 116858 232
rect 116914 176 150990 232
rect 151046 176 151051 232
rect 116853 174 151051 176
rect 108806 38 111948 98
rect 112621 98 112687 101
rect 116718 98 116778 172
rect 116853 171 116919 174
rect 150985 171 151051 174
rect 151813 234 151879 237
rect 198365 234 198431 237
rect 151813 232 198431 234
rect 151813 176 151818 232
rect 151874 176 198370 232
rect 198426 176 198431 232
rect 151813 174 198431 176
rect 151813 171 151879 174
rect 198365 171 198431 174
rect 198549 234 198615 237
rect 248413 234 248479 237
rect 198549 232 248479 234
rect 198549 176 198554 232
rect 198610 176 248418 232
rect 248474 176 248479 232
rect 198549 174 248479 176
rect 198549 171 198615 174
rect 248413 171 248479 174
rect 248689 234 248755 237
rect 265065 234 265131 237
rect 248689 232 265131 234
rect 248689 176 248694 232
rect 248750 176 265070 232
rect 265126 176 265131 232
rect 248689 174 265131 176
rect 248689 171 248755 174
rect 265065 171 265131 174
rect 265617 234 265683 237
rect 461669 234 461735 237
rect 265617 232 461735 234
rect 265617 176 265622 232
rect 265678 176 461674 232
rect 461730 176 461735 232
rect 265617 174 461735 176
rect 265617 171 265683 174
rect 461669 171 461735 174
rect 473353 234 473419 237
rect 473721 234 473787 237
rect 473353 232 473787 234
rect 473353 176 473358 232
rect 473414 176 473726 232
rect 473782 176 473787 232
rect 473353 174 473787 176
rect 473353 171 473419 174
rect 473721 171 473787 174
rect 486141 234 486207 237
rect 504222 234 504282 310
rect 486141 232 504282 234
rect 486141 176 486146 232
rect 486202 176 504282 232
rect 486141 174 504282 176
rect 486141 171 486207 174
rect 504398 172 504404 236
rect 504468 234 504474 236
rect 512870 234 512930 446
rect 522246 444 522252 446
rect 522316 444 522322 508
rect 522438 506 522498 582
rect 522573 640 536807 642
rect 522573 584 522578 640
rect 522634 584 536746 640
rect 536802 584 536807 640
rect 522573 582 536807 584
rect 522573 579 522639 582
rect 536741 579 536807 582
rect 545438 582 559788 642
rect 522438 446 528754 506
rect 504468 174 512930 234
rect 528694 234 528754 446
rect 539542 444 539548 508
rect 539612 506 539618 508
rect 545438 506 545498 582
rect 559782 580 559788 582
rect 559852 580 559858 644
rect 539612 446 545498 506
rect 545665 506 545731 509
rect 569174 506 569234 715
rect 545665 504 569234 506
rect 545665 448 545670 504
rect 545726 448 569234 504
rect 545665 446 569234 448
rect 539612 444 539618 446
rect 545665 443 545731 446
rect 528829 370 528895 373
rect 538765 370 538831 373
rect 528829 368 538831 370
rect 528829 312 528834 368
rect 528890 312 538770 368
rect 538826 312 538831 368
rect 528829 310 538831 312
rect 528829 307 528895 310
rect 538765 307 538831 310
rect 538949 370 539015 373
rect 559373 370 559439 373
rect 538949 368 559439 370
rect 538949 312 538954 368
rect 539010 312 559378 368
rect 559434 312 559439 368
rect 538949 310 559439 312
rect 538949 307 539015 310
rect 559373 307 559439 310
rect 545665 234 545731 237
rect 528694 232 545731 234
rect 528694 176 545670 232
rect 545726 176 545731 232
rect 528694 174 545731 176
rect 504468 172 504474 174
rect 545665 171 545731 174
rect 112621 96 116778 98
rect 112621 40 112626 96
rect 112682 40 116778 96
rect 112621 38 116778 40
rect 101949 35 102015 38
rect 108573 35 108639 38
rect 112621 35 112687 38
rect 116894 36 116900 100
rect 116964 98 116970 100
rect 119470 98 119476 100
rect 116964 38 119476 98
rect 116964 36 116970 38
rect 119470 36 119476 38
rect 119540 36 119546 100
rect 119613 98 119679 101
rect 569677 98 569743 101
rect 119613 96 569743 98
rect 119613 40 119618 96
rect 119674 40 569682 96
rect 569738 40 569743 96
rect 119613 38 569743 40
rect 119613 35 119679 38
rect 569677 35 569743 38
<< via3 >>
rect 550588 680988 550652 681052
rect 434668 680852 434732 680916
rect 344876 680580 344940 680644
rect 434668 680580 434732 680644
rect 550588 680580 550652 680644
rect 559788 680716 559852 680780
rect 561996 680580 562060 680644
rect 559052 680444 559116 680508
rect 561260 680444 561324 680508
rect 561628 680504 561692 680508
rect 561628 680448 561642 680504
rect 561642 680448 561692 680504
rect 561628 680444 561692 680448
rect 563100 680444 563164 680508
rect 564572 680444 564636 680508
rect 567148 680444 567212 680508
rect 559420 680308 559484 680372
rect 560708 680368 560772 680372
rect 560708 680312 560758 680368
rect 560758 680312 560772 680368
rect 560708 680308 560772 680312
rect 561076 680308 561140 680372
rect 562364 680308 562428 680372
rect 563652 680308 563716 680372
rect 566412 680368 566476 680372
rect 566412 680312 566426 680368
rect 566426 680312 566476 680368
rect 566412 680308 566476 680312
rect 3142 339688 3206 339692
rect 3142 339632 3146 339688
rect 3146 339632 3202 339688
rect 3202 339632 3206 339688
rect 3142 339628 3206 339632
rect 3142 321056 3206 321060
rect 3142 321000 3146 321056
rect 3146 321000 3202 321056
rect 3202 321000 3206 321056
rect 3142 320996 3206 321000
rect 570460 284608 570524 284612
rect 570460 284552 570510 284608
rect 570510 284552 570524 284608
rect 570460 284548 570524 284552
rect 569218 260128 569282 260132
rect 569218 260072 569222 260128
rect 569222 260072 569278 260128
rect 569278 260072 569282 260128
rect 569218 260068 569282 260072
rect 568390 248432 568454 248436
rect 568390 248376 568394 248432
rect 568394 248376 568450 248432
rect 568450 248376 568454 248432
rect 568390 248372 568454 248376
rect 568850 222320 568914 222324
rect 568850 222264 568854 222320
rect 568854 222264 568910 222320
rect 568910 222264 568914 222320
rect 568850 222260 568914 222264
rect 1348 221504 1412 221508
rect 1348 221448 1398 221504
rect 1398 221448 1412 221504
rect 1348 221444 1412 221448
rect 1348 214568 1412 214572
rect 1348 214512 1362 214568
rect 1362 214512 1412 214568
rect 1348 214508 1412 214512
rect 1532 198188 1596 198252
rect 568574 193624 568638 193628
rect 568574 193568 568578 193624
rect 568578 193568 568634 193624
rect 568634 193568 568638 193624
rect 568574 193564 568638 193568
rect 570276 193624 570340 193628
rect 570276 193568 570326 193624
rect 570326 193568 570340 193624
rect 570276 193564 570340 193568
rect 568298 193488 568362 193492
rect 568298 193432 568302 193488
rect 568302 193432 568358 193488
rect 568358 193432 568362 193488
rect 568298 193428 568362 193432
rect 570460 193428 570524 193492
rect 570644 193428 570708 193492
rect 2866 185328 2930 185332
rect 2866 185272 2870 185328
rect 2870 185272 2926 185328
rect 2926 185272 2930 185328
rect 2866 185268 2930 185272
rect 569172 178528 569236 178532
rect 569172 178472 569222 178528
rect 569222 178472 569236 178528
rect 569172 178468 569236 178472
rect 568482 174584 568546 174588
rect 568482 174528 568486 174584
rect 568486 174528 568542 174584
rect 568542 174528 568546 174584
rect 568482 174524 568546 174528
rect 1532 173088 1596 173092
rect 1532 173032 1546 173088
rect 1546 173032 1596 173088
rect 1532 173028 1596 173032
rect 1532 167588 1596 167652
rect 1532 146976 1596 146980
rect 1532 146920 1582 146976
rect 1582 146920 1596 146976
rect 1532 146916 1596 146920
rect 1532 138680 1596 138684
rect 1532 138624 1546 138680
rect 1546 138624 1596 138680
rect 1532 138620 1596 138624
rect 1348 108156 1412 108220
rect 1532 107068 1596 107132
rect 1532 99588 1596 99652
rect 570276 99376 570340 99380
rect 570276 99320 570326 99376
rect 570326 99320 570340 99376
rect 570276 99316 570340 99320
rect 3510 96112 3574 96116
rect 3510 96056 3514 96112
rect 3514 96056 3570 96112
rect 3570 96056 3574 96112
rect 3510 96052 3574 96056
rect 570460 90068 570524 90132
rect 1532 45868 1596 45932
rect 3740 40352 3804 40356
rect 3740 40296 3790 40352
rect 3790 40296 3804 40352
rect 3740 40292 3804 40296
rect 570276 34912 570340 34916
rect 570276 34856 570326 34912
rect 570326 34856 570340 34912
rect 570276 34852 570340 34856
rect 1532 33220 1596 33284
rect 612 32328 676 32332
rect 612 32272 662 32328
rect 662 32272 676 32328
rect 612 32268 676 32272
rect 1532 30288 1596 30292
rect 1532 30232 1546 30288
rect 1546 30232 1596 30288
rect 1532 30228 1596 30232
rect 1348 29744 1412 29748
rect 1348 29688 1398 29744
rect 1398 29688 1412 29744
rect 1348 29684 1412 29688
rect 1532 26964 1596 27028
rect 1348 26828 1412 26892
rect 980 25740 1044 25804
rect 1532 20028 1596 20092
rect 1348 19892 1412 19956
rect 1164 19756 1228 19820
rect 1532 17988 1596 18052
rect 20116 13288 20180 13292
rect 20116 13232 20130 13288
rect 20130 13232 20180 13288
rect 20116 13228 20180 13232
rect 980 12820 1044 12884
rect 570276 12336 570340 12340
rect 570276 12280 570326 12336
rect 570326 12280 570340 12336
rect 570276 12276 570340 12280
rect 1532 8800 1596 8804
rect 1532 8744 1582 8800
rect 1582 8744 1596 8800
rect 1532 8740 1596 8744
rect 19932 7984 19996 7988
rect 19932 7928 19982 7984
rect 19982 7928 19996 7984
rect 19932 7924 19996 7928
rect 612 7848 676 7852
rect 612 7792 626 7848
rect 626 7792 676 7848
rect 612 7788 676 7792
rect 225828 6428 225892 6492
rect 225828 5128 225892 5132
rect 225828 5072 225842 5128
rect 225842 5072 225892 5128
rect 225828 5068 225892 5072
rect 1348 4388 1412 4452
rect 570460 4388 570524 4452
rect 124306 3768 124370 3772
rect 124306 3712 124310 3768
rect 124310 3712 124366 3768
rect 124366 3712 124370 3768
rect 124306 3708 124370 3712
rect 177942 3768 178006 3772
rect 177942 3712 177946 3768
rect 177946 3712 178002 3768
rect 178002 3712 178006 3768
rect 177942 3708 178006 3712
rect 268378 3768 268442 3772
rect 268378 3712 268382 3768
rect 268382 3712 268438 3768
rect 268438 3712 268442 3768
rect 268378 3708 268442 3712
rect 91738 1804 91802 1868
rect 3004 1668 3068 1732
rect 65012 1668 65076 1732
rect 68692 1668 68756 1732
rect 72556 1668 72620 1732
rect 52316 1532 52380 1596
rect 3004 1396 3068 1460
rect 39068 1396 39132 1460
rect 56364 1396 56428 1460
rect 58572 1532 58636 1596
rect 66668 1532 66732 1596
rect 73108 1532 73172 1596
rect 73292 1532 73356 1596
rect 75316 1668 75380 1732
rect 76052 1668 76116 1732
rect 76788 1668 76852 1732
rect 75500 1532 75564 1596
rect 76420 1532 76484 1596
rect 82492 1668 82556 1732
rect 83596 1668 83660 1732
rect 85804 1668 85868 1732
rect 88012 1668 88076 1732
rect 88196 1668 88260 1732
rect 83044 1532 83108 1596
rect 92796 1668 92860 1732
rect 92980 1668 93044 1732
rect 94452 1668 94516 1732
rect 73476 1396 73540 1460
rect 83412 1456 83476 1460
rect 83412 1400 83426 1456
rect 83426 1400 83476 1456
rect 83412 1396 83476 1400
rect 95372 1668 95436 1732
rect 95556 1668 95620 1732
rect 100340 1668 100404 1732
rect 111564 1668 111628 1732
rect 120764 1668 120828 1732
rect 94820 1532 94884 1596
rect 95740 1532 95804 1596
rect 101812 1532 101876 1596
rect 103284 1532 103348 1596
rect 83044 1260 83108 1324
rect 83228 1260 83292 1324
rect 90956 1260 91020 1324
rect 101076 1456 101140 1460
rect 101076 1400 101126 1456
rect 101126 1400 101140 1456
rect 101076 1396 101140 1400
rect 102916 1396 102980 1460
rect 111196 1592 111260 1596
rect 111196 1536 111246 1592
rect 111246 1536 111260 1592
rect 111196 1532 111260 1536
rect 124444 1668 124508 1732
rect 125916 1668 125980 1732
rect 127940 1668 128004 1732
rect 128860 1668 128924 1732
rect 135300 1728 135364 1732
rect 135300 1672 135350 1728
rect 135350 1672 135364 1728
rect 135300 1668 135364 1672
rect 135668 1728 135732 1732
rect 135668 1672 135682 1728
rect 135682 1672 135732 1728
rect 135668 1668 135732 1672
rect 136082 1668 136146 1732
rect 136404 1668 136468 1732
rect 139348 1668 139412 1732
rect 141004 1668 141068 1732
rect 96476 1260 96540 1324
rect 97764 1260 97828 1324
rect 100340 1260 100404 1324
rect 101260 1260 101324 1324
rect 102180 1260 102244 1324
rect 102364 1320 102428 1324
rect 111748 1396 111812 1460
rect 128492 1532 128556 1596
rect 120764 1396 120828 1460
rect 102364 1264 102378 1320
rect 102378 1264 102428 1320
rect 102364 1260 102428 1264
rect 103284 1260 103348 1324
rect 2820 1124 2884 1188
rect 10916 1124 10980 1188
rect 39436 1124 39500 1188
rect 60596 1124 60660 1188
rect 64644 1124 64708 1188
rect 66852 1124 66916 1188
rect 82308 1124 82372 1188
rect 82676 1124 82740 1188
rect 90588 1124 90652 1188
rect 46796 1048 46860 1052
rect 46796 992 46810 1048
rect 46810 992 46860 1048
rect 46796 988 46860 992
rect 63724 988 63788 1052
rect 72924 988 72988 1052
rect 73108 988 73172 1052
rect 73476 988 73540 1052
rect 92428 1124 92492 1188
rect 101260 1124 101324 1188
rect 83228 988 83292 1052
rect 83412 988 83476 1052
rect 131436 1320 131500 1324
rect 131436 1264 131486 1320
rect 131486 1264 131500 1320
rect 131436 1260 131500 1264
rect 134380 1260 134444 1324
rect 135116 1396 135180 1460
rect 136588 1396 136652 1460
rect 141740 1668 141804 1732
rect 145788 1728 145852 1732
rect 145788 1672 145838 1728
rect 145838 1672 145852 1728
rect 145788 1668 145852 1672
rect 146156 1728 146220 1732
rect 146156 1672 146206 1728
rect 146206 1672 146220 1728
rect 146156 1668 146220 1672
rect 146340 1668 146404 1732
rect 148180 1668 148244 1732
rect 152228 1668 152292 1732
rect 138612 1396 138676 1460
rect 138796 1396 138860 1460
rect 136956 1320 137020 1324
rect 136956 1264 136970 1320
rect 136970 1264 137020 1320
rect 136956 1260 137020 1264
rect 141188 1260 141252 1324
rect 144868 1532 144932 1596
rect 145972 1532 146036 1596
rect 147260 1532 147324 1596
rect 147812 1532 147876 1596
rect 154436 1668 154500 1732
rect 156092 1668 156156 1732
rect 158484 1668 158548 1732
rect 166948 1668 167012 1732
rect 168972 1668 169036 1732
rect 157564 1396 157628 1460
rect 107148 1124 107212 1188
rect 107516 1124 107580 1188
rect 111380 1124 111444 1188
rect 111564 1184 111628 1188
rect 111564 1128 111614 1184
rect 111614 1128 111628 1184
rect 111564 1124 111628 1128
rect 111794 1124 111858 1188
rect 112484 1124 112548 1188
rect 120212 1124 120276 1188
rect 125364 1124 125428 1188
rect 126836 1124 126900 1188
rect 128308 1124 128372 1188
rect 123708 1048 123772 1052
rect 123708 992 123758 1048
rect 123758 992 123772 1048
rect 123708 988 123772 992
rect 124076 988 124140 1052
rect 128676 988 128740 1052
rect 10548 852 10612 916
rect 19196 852 19260 916
rect 28212 852 28276 916
rect 82308 852 82372 916
rect 82676 852 82740 916
rect 91324 852 91388 916
rect 91692 852 91756 916
rect 92244 852 92308 916
rect 129596 852 129660 916
rect 91876 716 91940 780
rect 102364 716 102428 780
rect 102916 716 102980 780
rect 106964 716 107028 780
rect 107700 716 107764 780
rect 111564 716 111628 780
rect 111748 716 111812 780
rect 428 308 492 372
rect 14964 308 15028 372
rect 61148 172 61212 236
rect 74212 444 74276 508
rect 76052 444 76116 508
rect 78628 444 78692 508
rect 79364 444 79428 508
rect 80284 444 80348 508
rect 102548 444 102612 508
rect 122972 716 123036 780
rect 129228 716 129292 780
rect 129964 988 130028 1052
rect 135484 988 135548 1052
rect 129964 852 130028 916
rect 139578 1124 139642 1188
rect 139900 1124 139964 1188
rect 141188 1124 141252 1188
rect 147444 1124 147508 1188
rect 147996 1260 148060 1324
rect 148180 1260 148244 1324
rect 148732 1124 148796 1188
rect 150756 1124 150820 1188
rect 151308 1124 151372 1188
rect 153884 1260 153948 1324
rect 157932 1532 157996 1596
rect 160140 1532 160204 1596
rect 161060 1532 161124 1596
rect 169340 1532 169404 1596
rect 169892 1668 169956 1732
rect 175780 1668 175844 1732
rect 175964 1668 176028 1732
rect 178172 1668 178236 1732
rect 178908 1668 178972 1732
rect 171180 1532 171244 1596
rect 171732 1532 171796 1596
rect 173020 1532 173084 1596
rect 157932 1456 157996 1460
rect 157932 1400 157982 1456
rect 157982 1400 157996 1456
rect 157932 1396 157996 1400
rect 159404 1396 159468 1460
rect 159772 1396 159836 1460
rect 161244 1396 161308 1460
rect 161612 1396 161676 1460
rect 164004 1396 164068 1460
rect 176884 1396 176948 1460
rect 177068 1396 177132 1460
rect 178172 1532 178236 1596
rect 178356 1532 178420 1596
rect 179644 1532 179708 1596
rect 181852 1532 181916 1596
rect 177988 1396 178052 1460
rect 161980 1260 162044 1324
rect 163452 1260 163516 1324
rect 169892 1260 169956 1324
rect 170076 1260 170140 1324
rect 166212 1124 166276 1188
rect 168788 1124 168852 1188
rect 173940 1260 174004 1324
rect 175964 1260 176028 1324
rect 176332 1260 176396 1324
rect 179460 1260 179524 1324
rect 180380 1260 180444 1324
rect 173388 1124 173452 1188
rect 176148 1124 176212 1188
rect 180932 1124 180996 1188
rect 183692 1260 183756 1324
rect 184060 1532 184124 1596
rect 184980 1668 185044 1732
rect 192340 1668 192404 1732
rect 194732 1668 194796 1732
rect 194916 1668 194980 1732
rect 190500 1532 190564 1596
rect 195836 1532 195900 1596
rect 197124 1532 197188 1596
rect 191052 1396 191116 1460
rect 198412 1532 198476 1596
rect 197492 1396 197556 1460
rect 198780 1396 198844 1460
rect 207980 1668 208044 1732
rect 216812 1668 216876 1732
rect 220308 1668 220372 1732
rect 200988 1532 201052 1596
rect 203196 1532 203260 1596
rect 204300 1532 204364 1596
rect 204668 1532 204732 1596
rect 204852 1592 204916 1596
rect 204852 1536 204866 1592
rect 204866 1536 204916 1592
rect 204852 1532 204916 1536
rect 200436 1396 200500 1460
rect 189764 1260 189828 1324
rect 191236 1260 191300 1324
rect 208348 1396 208412 1460
rect 209820 1396 209884 1460
rect 210188 1532 210252 1596
rect 210924 1396 210988 1460
rect 212028 1396 212092 1460
rect 210004 1260 210068 1324
rect 218284 1396 218348 1460
rect 224540 1456 224604 1460
rect 224540 1400 224554 1456
rect 224554 1400 224604 1456
rect 224540 1396 224604 1400
rect 224908 1532 224972 1596
rect 234292 1668 234356 1732
rect 237972 1668 238036 1732
rect 245332 1668 245396 1732
rect 247540 1668 247604 1732
rect 238708 1532 238772 1596
rect 239076 1532 239140 1596
rect 241836 1532 241900 1596
rect 249748 1532 249812 1596
rect 214788 1320 214852 1324
rect 214788 1264 214838 1320
rect 214838 1264 214852 1320
rect 214788 1260 214852 1264
rect 217548 1260 217612 1324
rect 243124 1396 243188 1460
rect 245148 1396 245212 1460
rect 246620 1396 246684 1460
rect 246804 1396 246868 1460
rect 248828 1396 248892 1460
rect 250116 1396 250180 1460
rect 253244 1532 253308 1596
rect 227116 1260 227180 1324
rect 227484 1320 227548 1324
rect 227484 1264 227498 1320
rect 227498 1264 227548 1320
rect 227484 1260 227548 1264
rect 227668 1260 227732 1324
rect 229140 1260 229204 1324
rect 229324 1260 229388 1324
rect 245516 1260 245580 1324
rect 245700 1260 245764 1324
rect 247908 1260 247972 1324
rect 250484 1260 250548 1324
rect 251220 1260 251284 1324
rect 163820 988 163884 1052
rect 191052 1124 191116 1188
rect 184428 988 184492 1052
rect 189764 988 189828 1052
rect 191420 1124 191484 1188
rect 196940 1124 197004 1188
rect 197308 988 197372 1052
rect 209268 1184 209332 1188
rect 209268 1128 209282 1184
rect 209282 1128 209332 1184
rect 209268 1124 209332 1128
rect 212028 1124 212092 1188
rect 217732 1124 217796 1188
rect 225092 1184 225156 1188
rect 225092 1128 225142 1184
rect 225142 1128 225156 1184
rect 225092 1124 225156 1128
rect 226748 1124 226812 1188
rect 247540 988 247604 1052
rect 247908 988 247972 1052
rect 135852 852 135916 916
rect 130332 716 130396 780
rect 130516 716 130580 780
rect 134932 716 134996 780
rect 135300 716 135364 780
rect 136220 716 136284 780
rect 137692 716 137756 780
rect 150756 852 150820 916
rect 150940 852 151004 916
rect 151308 852 151372 916
rect 197860 852 197924 916
rect 144316 716 144380 780
rect 145604 716 145668 780
rect 147076 716 147140 780
rect 124076 580 124140 644
rect 135484 580 135548 644
rect 139900 580 139964 644
rect 103284 444 103348 508
rect 111748 444 111812 508
rect 112300 444 112364 508
rect 150756 504 150820 508
rect 150756 448 150806 504
rect 150806 448 150820 504
rect 150756 444 150820 448
rect 151308 580 151372 644
rect 156276 580 156340 644
rect 161612 716 161676 780
rect 157932 640 157996 644
rect 157932 584 157946 640
rect 157946 584 157996 640
rect 157932 580 157996 584
rect 163268 716 163332 780
rect 190316 716 190380 780
rect 231348 852 231412 916
rect 232636 852 232700 916
rect 232820 852 232884 916
rect 233372 912 233436 916
rect 233372 856 233386 912
rect 233386 856 233436 912
rect 233372 852 233436 856
rect 233740 852 233804 916
rect 250300 852 250364 916
rect 252692 988 252756 1052
rect 253428 1396 253492 1460
rect 253796 1532 253860 1596
rect 261708 1668 261772 1732
rect 268700 1668 268764 1732
rect 258396 1532 258460 1596
rect 261892 1532 261956 1596
rect 260604 1456 260668 1460
rect 260604 1400 260654 1456
rect 260654 1400 260668 1456
rect 260604 1396 260668 1400
rect 260972 1396 261036 1460
rect 272196 1668 272260 1732
rect 279004 1668 279068 1732
rect 285628 1668 285692 1732
rect 294092 1702 294156 1766
rect 294460 1668 294524 1732
rect 268884 1456 268948 1460
rect 268884 1400 268898 1456
rect 268898 1400 268948 1456
rect 268884 1396 268948 1400
rect 253060 1260 253124 1324
rect 256372 1260 256436 1324
rect 262812 1260 262876 1324
rect 264836 1260 264900 1324
rect 271828 1396 271892 1460
rect 273300 1396 273364 1460
rect 273484 1456 273548 1460
rect 273484 1400 273534 1456
rect 273534 1400 273548 1456
rect 273484 1396 273548 1400
rect 273668 1396 273732 1460
rect 279372 1396 279436 1460
rect 280476 1396 280540 1460
rect 281028 1320 281092 1324
rect 281028 1264 281042 1320
rect 281042 1264 281092 1320
rect 281028 1260 281092 1264
rect 281396 1396 281460 1460
rect 296116 1532 296180 1596
rect 310468 1668 310532 1732
rect 310652 1668 310716 1732
rect 385724 1668 385788 1732
rect 513236 1668 513300 1732
rect 567148 1668 567212 1732
rect 569172 1668 569236 1732
rect 569540 1728 569604 1732
rect 569540 1672 569590 1728
rect 569590 1672 569604 1728
rect 569540 1668 569604 1672
rect 354260 1532 354324 1596
rect 558868 1532 558932 1596
rect 559052 1592 559116 1596
rect 559052 1536 559102 1592
rect 559102 1536 559116 1592
rect 559052 1532 559116 1536
rect 559420 1396 559484 1460
rect 560156 1396 560220 1460
rect 566412 1396 566476 1460
rect 268884 1124 268948 1188
rect 279556 1124 279620 1188
rect 253428 988 253492 1052
rect 256004 988 256068 1052
rect 262260 1048 262324 1052
rect 262260 992 262310 1048
rect 262310 992 262324 1048
rect 262260 988 262324 992
rect 294828 1260 294892 1324
rect 317828 1260 317892 1324
rect 324820 1260 324884 1324
rect 327764 1320 327828 1324
rect 327764 1264 327778 1320
rect 327778 1264 327828 1320
rect 327764 1260 327828 1264
rect 372476 1260 372540 1324
rect 419396 1260 419460 1324
rect 289676 1124 289740 1188
rect 290044 1124 290108 1188
rect 290412 1184 290476 1188
rect 290412 1128 290426 1184
rect 290426 1128 290476 1184
rect 290412 1124 290476 1128
rect 296852 1124 296916 1188
rect 308812 1124 308876 1188
rect 303292 988 303356 1052
rect 328316 1124 328380 1188
rect 328500 1124 328564 1188
rect 348924 1124 348988 1188
rect 370452 1124 370516 1188
rect 483796 1124 483860 1188
rect 514156 1124 514220 1188
rect 564940 1260 565004 1324
rect 561444 1124 561508 1188
rect 327028 1048 327092 1052
rect 327028 992 327078 1048
rect 327078 992 327092 1048
rect 327028 988 327092 992
rect 251956 852 252020 916
rect 253796 852 253860 916
rect 255636 852 255700 916
rect 198412 716 198476 780
rect 163636 580 163700 644
rect 169892 640 169956 644
rect 169892 584 169906 640
rect 169906 584 169956 640
rect 169892 580 169956 584
rect 175044 580 175108 644
rect 175412 580 175476 644
rect 177252 580 177316 644
rect 177804 580 177868 644
rect 204116 580 204180 644
rect 204668 580 204732 644
rect 205220 580 205284 644
rect 207980 580 208044 644
rect 210372 580 210436 644
rect 210556 580 210620 644
rect 211292 580 211356 644
rect 219204 580 219268 644
rect 231164 716 231228 780
rect 245148 716 245212 780
rect 246436 716 246500 780
rect 246620 716 246684 780
rect 252324 716 252388 780
rect 252508 716 252572 780
rect 309916 852 309980 916
rect 314884 852 314948 916
rect 328316 852 328380 916
rect 328546 912 328610 916
rect 328546 856 328550 912
rect 328550 856 328606 912
rect 328606 856 328610 912
rect 328546 852 328610 856
rect 329052 852 329116 916
rect 258212 716 258276 780
rect 260236 716 260300 780
rect 260788 776 260852 780
rect 260788 720 260838 776
rect 260838 720 260852 776
rect 260788 716 260852 720
rect 261156 716 261220 780
rect 248276 580 248340 644
rect 280108 716 280172 780
rect 280660 716 280724 780
rect 294828 776 294892 780
rect 294828 720 294842 776
rect 294842 720 294892 776
rect 294828 716 294892 720
rect 264836 580 264900 644
rect 338620 580 338684 644
rect 338804 580 338868 644
rect 342668 580 342732 644
rect 353892 716 353956 780
rect 358124 852 358188 916
rect 564572 852 564636 916
rect 362724 716 362788 780
rect 385908 716 385972 780
rect 440188 716 440252 780
rect 449756 716 449820 780
rect 539548 716 539612 780
rect 563100 716 563164 780
rect 350028 580 350092 644
rect 390508 580 390572 644
rect 430620 580 430684 644
rect 434484 580 434548 644
rect 190868 444 190932 508
rect 191420 444 191484 508
rect 197124 444 197188 508
rect 197860 444 197924 508
rect 198228 504 198292 508
rect 198228 448 198242 504
rect 198242 448 198292 504
rect 198228 444 198292 448
rect 463004 444 463068 508
rect 469076 444 469140 508
rect 473492 444 473556 508
rect 157932 308 157996 372
rect 161244 308 161308 372
rect 290780 308 290844 372
rect 291148 308 291212 372
rect 390508 308 390572 372
rect 418844 308 418908 372
rect 422156 308 422220 372
rect 426940 308 427004 372
rect 442948 308 443012 372
rect 473124 308 473188 372
rect 476804 308 476868 372
rect 490604 308 490668 372
rect 1900 36 1964 100
rect 73844 172 73908 236
rect 82308 172 82372 236
rect 85436 172 85500 236
rect 85620 172 85684 236
rect 87276 172 87340 236
rect 92980 172 93044 236
rect 93164 172 93228 236
rect 93900 172 93964 236
rect 94268 172 94332 236
rect 74212 36 74276 100
rect 78628 36 78692 100
rect 81388 36 81452 100
rect 83044 36 83108 100
rect 84332 36 84396 100
rect 89668 36 89732 100
rect 92612 36 92676 100
rect 101444 36 101508 100
rect 116716 172 116780 236
rect 504404 172 504468 236
rect 522252 444 522316 508
rect 539548 444 539612 508
rect 559788 580 559852 644
rect 116900 36 116964 100
rect 119476 36 119540 100
<< metal4 >>
rect -8436 711278 -7836 711300
rect -8436 711042 -8254 711278
rect -8018 711042 -7836 711278
rect -8436 710958 -7836 711042
rect -8436 710722 -8254 710958
rect -8018 710722 -7836 710958
rect -8436 679254 -7836 710722
rect 591760 711278 592360 711300
rect 591760 711042 591942 711278
rect 592178 711042 592360 711278
rect 591760 710958 592360 711042
rect 591760 710722 591942 710958
rect 592178 710722 592360 710958
rect -8436 679018 -8254 679254
rect -8018 679018 -7836 679254
rect -8436 678934 -7836 679018
rect -8436 678698 -8254 678934
rect -8018 678698 -7836 678934
rect -8436 643254 -7836 678698
rect -8436 643018 -8254 643254
rect -8018 643018 -7836 643254
rect -8436 642934 -7836 643018
rect -8436 642698 -8254 642934
rect -8018 642698 -7836 642934
rect -8436 607254 -7836 642698
rect -8436 607018 -8254 607254
rect -8018 607018 -7836 607254
rect -8436 606934 -7836 607018
rect -8436 606698 -8254 606934
rect -8018 606698 -7836 606934
rect -8436 571254 -7836 606698
rect -8436 571018 -8254 571254
rect -8018 571018 -7836 571254
rect -8436 570934 -7836 571018
rect -8436 570698 -8254 570934
rect -8018 570698 -7836 570934
rect -8436 535254 -7836 570698
rect -8436 535018 -8254 535254
rect -8018 535018 -7836 535254
rect -8436 534934 -7836 535018
rect -8436 534698 -8254 534934
rect -8018 534698 -7836 534934
rect -8436 499254 -7836 534698
rect -8436 499018 -8254 499254
rect -8018 499018 -7836 499254
rect -8436 498934 -7836 499018
rect -8436 498698 -8254 498934
rect -8018 498698 -7836 498934
rect -8436 463254 -7836 498698
rect -8436 463018 -8254 463254
rect -8018 463018 -7836 463254
rect -8436 462934 -7836 463018
rect -8436 462698 -8254 462934
rect -8018 462698 -7836 462934
rect -8436 427254 -7836 462698
rect -8436 427018 -8254 427254
rect -8018 427018 -7836 427254
rect -8436 426934 -7836 427018
rect -8436 426698 -8254 426934
rect -8018 426698 -7836 426934
rect -8436 391254 -7836 426698
rect -8436 391018 -8254 391254
rect -8018 391018 -7836 391254
rect -8436 390934 -7836 391018
rect -8436 390698 -8254 390934
rect -8018 390698 -7836 390934
rect -8436 355254 -7836 390698
rect -8436 355018 -8254 355254
rect -8018 355018 -7836 355254
rect -8436 354934 -7836 355018
rect -8436 354698 -8254 354934
rect -8018 354698 -7836 354934
rect -8436 319254 -7836 354698
rect -8436 319018 -8254 319254
rect -8018 319018 -7836 319254
rect -8436 318934 -7836 319018
rect -8436 318698 -8254 318934
rect -8018 318698 -7836 318934
rect -8436 283254 -7836 318698
rect -8436 283018 -8254 283254
rect -8018 283018 -7836 283254
rect -8436 282934 -7836 283018
rect -8436 282698 -8254 282934
rect -8018 282698 -7836 282934
rect -8436 247254 -7836 282698
rect -8436 247018 -8254 247254
rect -8018 247018 -7836 247254
rect -8436 246934 -7836 247018
rect -8436 246698 -8254 246934
rect -8018 246698 -7836 246934
rect -8436 211254 -7836 246698
rect -8436 211018 -8254 211254
rect -8018 211018 -7836 211254
rect -8436 210934 -7836 211018
rect -8436 210698 -8254 210934
rect -8018 210698 -7836 210934
rect -8436 175254 -7836 210698
rect -8436 175018 -8254 175254
rect -8018 175018 -7836 175254
rect -8436 174934 -7836 175018
rect -8436 174698 -8254 174934
rect -8018 174698 -7836 174934
rect -8436 139254 -7836 174698
rect -8436 139018 -8254 139254
rect -8018 139018 -7836 139254
rect -8436 138934 -7836 139018
rect -8436 138698 -8254 138934
rect -8018 138698 -7836 138934
rect -8436 103254 -7836 138698
rect -8436 103018 -8254 103254
rect -8018 103018 -7836 103254
rect -8436 102934 -7836 103018
rect -8436 102698 -8254 102934
rect -8018 102698 -7836 102934
rect -8436 67254 -7836 102698
rect -8436 67018 -8254 67254
rect -8018 67018 -7836 67254
rect -8436 66934 -7836 67018
rect -8436 66698 -8254 66934
rect -8018 66698 -7836 66934
rect -8436 31254 -7836 66698
rect -8436 31018 -8254 31254
rect -8018 31018 -7836 31254
rect -8436 30934 -7836 31018
rect -8436 30698 -8254 30934
rect -8018 30698 -7836 30934
rect -8436 -6786 -7836 30698
rect -7516 710358 -6916 710380
rect -7516 710122 -7334 710358
rect -7098 710122 -6916 710358
rect -7516 710038 -6916 710122
rect -7516 709802 -7334 710038
rect -7098 709802 -6916 710038
rect -7516 697254 -6916 709802
rect 590840 710358 591440 710380
rect 590840 710122 591022 710358
rect 591258 710122 591440 710358
rect 590840 710038 591440 710122
rect 590840 709802 591022 710038
rect 591258 709802 591440 710038
rect -7516 697018 -7334 697254
rect -7098 697018 -6916 697254
rect -7516 696934 -6916 697018
rect -7516 696698 -7334 696934
rect -7098 696698 -6916 696934
rect -7516 661254 -6916 696698
rect -7516 661018 -7334 661254
rect -7098 661018 -6916 661254
rect -7516 660934 -6916 661018
rect -7516 660698 -7334 660934
rect -7098 660698 -6916 660934
rect -7516 625254 -6916 660698
rect -7516 625018 -7334 625254
rect -7098 625018 -6916 625254
rect -7516 624934 -6916 625018
rect -7516 624698 -7334 624934
rect -7098 624698 -6916 624934
rect -7516 589254 -6916 624698
rect -7516 589018 -7334 589254
rect -7098 589018 -6916 589254
rect -7516 588934 -6916 589018
rect -7516 588698 -7334 588934
rect -7098 588698 -6916 588934
rect -7516 553254 -6916 588698
rect -7516 553018 -7334 553254
rect -7098 553018 -6916 553254
rect -7516 552934 -6916 553018
rect -7516 552698 -7334 552934
rect -7098 552698 -6916 552934
rect -7516 517254 -6916 552698
rect -7516 517018 -7334 517254
rect -7098 517018 -6916 517254
rect -7516 516934 -6916 517018
rect -7516 516698 -7334 516934
rect -7098 516698 -6916 516934
rect -7516 481254 -6916 516698
rect -7516 481018 -7334 481254
rect -7098 481018 -6916 481254
rect -7516 480934 -6916 481018
rect -7516 480698 -7334 480934
rect -7098 480698 -6916 480934
rect -7516 445254 -6916 480698
rect -7516 445018 -7334 445254
rect -7098 445018 -6916 445254
rect -7516 444934 -6916 445018
rect -7516 444698 -7334 444934
rect -7098 444698 -6916 444934
rect -7516 409254 -6916 444698
rect -7516 409018 -7334 409254
rect -7098 409018 -6916 409254
rect -7516 408934 -6916 409018
rect -7516 408698 -7334 408934
rect -7098 408698 -6916 408934
rect -7516 373254 -6916 408698
rect -7516 373018 -7334 373254
rect -7098 373018 -6916 373254
rect -7516 372934 -6916 373018
rect -7516 372698 -7334 372934
rect -7098 372698 -6916 372934
rect -7516 337254 -6916 372698
rect -7516 337018 -7334 337254
rect -7098 337018 -6916 337254
rect -7516 336934 -6916 337018
rect -7516 336698 -7334 336934
rect -7098 336698 -6916 336934
rect -7516 301254 -6916 336698
rect -7516 301018 -7334 301254
rect -7098 301018 -6916 301254
rect -7516 300934 -6916 301018
rect -7516 300698 -7334 300934
rect -7098 300698 -6916 300934
rect -7516 265254 -6916 300698
rect -7516 265018 -7334 265254
rect -7098 265018 -6916 265254
rect -7516 264934 -6916 265018
rect -7516 264698 -7334 264934
rect -7098 264698 -6916 264934
rect -7516 229254 -6916 264698
rect -7516 229018 -7334 229254
rect -7098 229018 -6916 229254
rect -7516 228934 -6916 229018
rect -7516 228698 -7334 228934
rect -7098 228698 -6916 228934
rect -7516 193254 -6916 228698
rect -7516 193018 -7334 193254
rect -7098 193018 -6916 193254
rect -7516 192934 -6916 193018
rect -7516 192698 -7334 192934
rect -7098 192698 -6916 192934
rect -7516 157254 -6916 192698
rect -7516 157018 -7334 157254
rect -7098 157018 -6916 157254
rect -7516 156934 -6916 157018
rect -7516 156698 -7334 156934
rect -7098 156698 -6916 156934
rect -7516 121254 -6916 156698
rect -7516 121018 -7334 121254
rect -7098 121018 -6916 121254
rect -7516 120934 -6916 121018
rect -7516 120698 -7334 120934
rect -7098 120698 -6916 120934
rect -7516 85254 -6916 120698
rect -7516 85018 -7334 85254
rect -7098 85018 -6916 85254
rect -7516 84934 -6916 85018
rect -7516 84698 -7334 84934
rect -7098 84698 -6916 84934
rect -7516 49254 -6916 84698
rect -7516 49018 -7334 49254
rect -7098 49018 -6916 49254
rect -7516 48934 -6916 49018
rect -7516 48698 -7334 48934
rect -7098 48698 -6916 48934
rect -7516 13254 -6916 48698
rect -7516 13018 -7334 13254
rect -7098 13018 -6916 13254
rect -7516 12934 -6916 13018
rect -7516 12698 -7334 12934
rect -7098 12698 -6916 12934
rect -7516 -5866 -6916 12698
rect -6596 709438 -5996 709460
rect -6596 709202 -6414 709438
rect -6178 709202 -5996 709438
rect -6596 709118 -5996 709202
rect -6596 708882 -6414 709118
rect -6178 708882 -5996 709118
rect -6596 675654 -5996 708882
rect 589920 709438 590520 709460
rect 589920 709202 590102 709438
rect 590338 709202 590520 709438
rect 589920 709118 590520 709202
rect 589920 708882 590102 709118
rect 590338 708882 590520 709118
rect -6596 675418 -6414 675654
rect -6178 675418 -5996 675654
rect -6596 675334 -5996 675418
rect -6596 675098 -6414 675334
rect -6178 675098 -5996 675334
rect -6596 639654 -5996 675098
rect -6596 639418 -6414 639654
rect -6178 639418 -5996 639654
rect -6596 639334 -5996 639418
rect -6596 639098 -6414 639334
rect -6178 639098 -5996 639334
rect -6596 603654 -5996 639098
rect -6596 603418 -6414 603654
rect -6178 603418 -5996 603654
rect -6596 603334 -5996 603418
rect -6596 603098 -6414 603334
rect -6178 603098 -5996 603334
rect -6596 567654 -5996 603098
rect -6596 567418 -6414 567654
rect -6178 567418 -5996 567654
rect -6596 567334 -5996 567418
rect -6596 567098 -6414 567334
rect -6178 567098 -5996 567334
rect -6596 531654 -5996 567098
rect -6596 531418 -6414 531654
rect -6178 531418 -5996 531654
rect -6596 531334 -5996 531418
rect -6596 531098 -6414 531334
rect -6178 531098 -5996 531334
rect -6596 495654 -5996 531098
rect -6596 495418 -6414 495654
rect -6178 495418 -5996 495654
rect -6596 495334 -5996 495418
rect -6596 495098 -6414 495334
rect -6178 495098 -5996 495334
rect -6596 459654 -5996 495098
rect -6596 459418 -6414 459654
rect -6178 459418 -5996 459654
rect -6596 459334 -5996 459418
rect -6596 459098 -6414 459334
rect -6178 459098 -5996 459334
rect -6596 423654 -5996 459098
rect -6596 423418 -6414 423654
rect -6178 423418 -5996 423654
rect -6596 423334 -5996 423418
rect -6596 423098 -6414 423334
rect -6178 423098 -5996 423334
rect -6596 387654 -5996 423098
rect -6596 387418 -6414 387654
rect -6178 387418 -5996 387654
rect -6596 387334 -5996 387418
rect -6596 387098 -6414 387334
rect -6178 387098 -5996 387334
rect -6596 351654 -5996 387098
rect -6596 351418 -6414 351654
rect -6178 351418 -5996 351654
rect -6596 351334 -5996 351418
rect -6596 351098 -6414 351334
rect -6178 351098 -5996 351334
rect -6596 315654 -5996 351098
rect -6596 315418 -6414 315654
rect -6178 315418 -5996 315654
rect -6596 315334 -5996 315418
rect -6596 315098 -6414 315334
rect -6178 315098 -5996 315334
rect -6596 279654 -5996 315098
rect -6596 279418 -6414 279654
rect -6178 279418 -5996 279654
rect -6596 279334 -5996 279418
rect -6596 279098 -6414 279334
rect -6178 279098 -5996 279334
rect -6596 243654 -5996 279098
rect -6596 243418 -6414 243654
rect -6178 243418 -5996 243654
rect -6596 243334 -5996 243418
rect -6596 243098 -6414 243334
rect -6178 243098 -5996 243334
rect -6596 207654 -5996 243098
rect -6596 207418 -6414 207654
rect -6178 207418 -5996 207654
rect -6596 207334 -5996 207418
rect -6596 207098 -6414 207334
rect -6178 207098 -5996 207334
rect -6596 171654 -5996 207098
rect -6596 171418 -6414 171654
rect -6178 171418 -5996 171654
rect -6596 171334 -5996 171418
rect -6596 171098 -6414 171334
rect -6178 171098 -5996 171334
rect -6596 135654 -5996 171098
rect -6596 135418 -6414 135654
rect -6178 135418 -5996 135654
rect -6596 135334 -5996 135418
rect -6596 135098 -6414 135334
rect -6178 135098 -5996 135334
rect -6596 99654 -5996 135098
rect -6596 99418 -6414 99654
rect -6178 99418 -5996 99654
rect -6596 99334 -5996 99418
rect -6596 99098 -6414 99334
rect -6178 99098 -5996 99334
rect -6596 63654 -5996 99098
rect -6596 63418 -6414 63654
rect -6178 63418 -5996 63654
rect -6596 63334 -5996 63418
rect -6596 63098 -6414 63334
rect -6178 63098 -5996 63334
rect -6596 27654 -5996 63098
rect -6596 27418 -6414 27654
rect -6178 27418 -5996 27654
rect -6596 27334 -5996 27418
rect -6596 27098 -6414 27334
rect -6178 27098 -5996 27334
rect -6596 -4946 -5996 27098
rect -5676 708518 -5076 708540
rect -5676 708282 -5494 708518
rect -5258 708282 -5076 708518
rect -5676 708198 -5076 708282
rect -5676 707962 -5494 708198
rect -5258 707962 -5076 708198
rect -5676 693654 -5076 707962
rect 589000 708518 589600 708540
rect 589000 708282 589182 708518
rect 589418 708282 589600 708518
rect 589000 708198 589600 708282
rect 589000 707962 589182 708198
rect 589418 707962 589600 708198
rect -5676 693418 -5494 693654
rect -5258 693418 -5076 693654
rect -5676 693334 -5076 693418
rect -5676 693098 -5494 693334
rect -5258 693098 -5076 693334
rect -5676 657654 -5076 693098
rect -5676 657418 -5494 657654
rect -5258 657418 -5076 657654
rect -5676 657334 -5076 657418
rect -5676 657098 -5494 657334
rect -5258 657098 -5076 657334
rect -5676 621654 -5076 657098
rect -5676 621418 -5494 621654
rect -5258 621418 -5076 621654
rect -5676 621334 -5076 621418
rect -5676 621098 -5494 621334
rect -5258 621098 -5076 621334
rect -5676 585654 -5076 621098
rect -5676 585418 -5494 585654
rect -5258 585418 -5076 585654
rect -5676 585334 -5076 585418
rect -5676 585098 -5494 585334
rect -5258 585098 -5076 585334
rect -5676 549654 -5076 585098
rect -5676 549418 -5494 549654
rect -5258 549418 -5076 549654
rect -5676 549334 -5076 549418
rect -5676 549098 -5494 549334
rect -5258 549098 -5076 549334
rect -5676 513654 -5076 549098
rect -5676 513418 -5494 513654
rect -5258 513418 -5076 513654
rect -5676 513334 -5076 513418
rect -5676 513098 -5494 513334
rect -5258 513098 -5076 513334
rect -5676 477654 -5076 513098
rect -5676 477418 -5494 477654
rect -5258 477418 -5076 477654
rect -5676 477334 -5076 477418
rect -5676 477098 -5494 477334
rect -5258 477098 -5076 477334
rect -5676 441654 -5076 477098
rect -5676 441418 -5494 441654
rect -5258 441418 -5076 441654
rect -5676 441334 -5076 441418
rect -5676 441098 -5494 441334
rect -5258 441098 -5076 441334
rect -5676 405654 -5076 441098
rect -5676 405418 -5494 405654
rect -5258 405418 -5076 405654
rect -5676 405334 -5076 405418
rect -5676 405098 -5494 405334
rect -5258 405098 -5076 405334
rect -5676 369654 -5076 405098
rect -5676 369418 -5494 369654
rect -5258 369418 -5076 369654
rect -5676 369334 -5076 369418
rect -5676 369098 -5494 369334
rect -5258 369098 -5076 369334
rect -5676 333654 -5076 369098
rect -5676 333418 -5494 333654
rect -5258 333418 -5076 333654
rect -5676 333334 -5076 333418
rect -5676 333098 -5494 333334
rect -5258 333098 -5076 333334
rect -5676 297654 -5076 333098
rect -5676 297418 -5494 297654
rect -5258 297418 -5076 297654
rect -5676 297334 -5076 297418
rect -5676 297098 -5494 297334
rect -5258 297098 -5076 297334
rect -5676 261654 -5076 297098
rect -5676 261418 -5494 261654
rect -5258 261418 -5076 261654
rect -5676 261334 -5076 261418
rect -5676 261098 -5494 261334
rect -5258 261098 -5076 261334
rect -5676 225654 -5076 261098
rect -5676 225418 -5494 225654
rect -5258 225418 -5076 225654
rect -5676 225334 -5076 225418
rect -5676 225098 -5494 225334
rect -5258 225098 -5076 225334
rect -5676 189654 -5076 225098
rect -5676 189418 -5494 189654
rect -5258 189418 -5076 189654
rect -5676 189334 -5076 189418
rect -5676 189098 -5494 189334
rect -5258 189098 -5076 189334
rect -5676 153654 -5076 189098
rect -5676 153418 -5494 153654
rect -5258 153418 -5076 153654
rect -5676 153334 -5076 153418
rect -5676 153098 -5494 153334
rect -5258 153098 -5076 153334
rect -5676 117654 -5076 153098
rect -5676 117418 -5494 117654
rect -5258 117418 -5076 117654
rect -5676 117334 -5076 117418
rect -5676 117098 -5494 117334
rect -5258 117098 -5076 117334
rect -5676 81654 -5076 117098
rect -5676 81418 -5494 81654
rect -5258 81418 -5076 81654
rect -5676 81334 -5076 81418
rect -5676 81098 -5494 81334
rect -5258 81098 -5076 81334
rect -5676 45654 -5076 81098
rect -5676 45418 -5494 45654
rect -5258 45418 -5076 45654
rect -5676 45334 -5076 45418
rect -5676 45098 -5494 45334
rect -5258 45098 -5076 45334
rect -5676 9654 -5076 45098
rect -5676 9418 -5494 9654
rect -5258 9418 -5076 9654
rect -5676 9334 -5076 9418
rect -5676 9098 -5494 9334
rect -5258 9098 -5076 9334
rect -5676 -4026 -5076 9098
rect -4756 707598 -4156 707620
rect -4756 707362 -4574 707598
rect -4338 707362 -4156 707598
rect -4756 707278 -4156 707362
rect -4756 707042 -4574 707278
rect -4338 707042 -4156 707278
rect -4756 672054 -4156 707042
rect 588080 707598 588680 707620
rect 588080 707362 588262 707598
rect 588498 707362 588680 707598
rect 588080 707278 588680 707362
rect 588080 707042 588262 707278
rect 588498 707042 588680 707278
rect -4756 671818 -4574 672054
rect -4338 671818 -4156 672054
rect -4756 671734 -4156 671818
rect -4756 671498 -4574 671734
rect -4338 671498 -4156 671734
rect -4756 636054 -4156 671498
rect -4756 635818 -4574 636054
rect -4338 635818 -4156 636054
rect -4756 635734 -4156 635818
rect -4756 635498 -4574 635734
rect -4338 635498 -4156 635734
rect -4756 600054 -4156 635498
rect -4756 599818 -4574 600054
rect -4338 599818 -4156 600054
rect -4756 599734 -4156 599818
rect -4756 599498 -4574 599734
rect -4338 599498 -4156 599734
rect -4756 564054 -4156 599498
rect -4756 563818 -4574 564054
rect -4338 563818 -4156 564054
rect -4756 563734 -4156 563818
rect -4756 563498 -4574 563734
rect -4338 563498 -4156 563734
rect -4756 528054 -4156 563498
rect -4756 527818 -4574 528054
rect -4338 527818 -4156 528054
rect -4756 527734 -4156 527818
rect -4756 527498 -4574 527734
rect -4338 527498 -4156 527734
rect -4756 492054 -4156 527498
rect -4756 491818 -4574 492054
rect -4338 491818 -4156 492054
rect -4756 491734 -4156 491818
rect -4756 491498 -4574 491734
rect -4338 491498 -4156 491734
rect -4756 456054 -4156 491498
rect -4756 455818 -4574 456054
rect -4338 455818 -4156 456054
rect -4756 455734 -4156 455818
rect -4756 455498 -4574 455734
rect -4338 455498 -4156 455734
rect -4756 420054 -4156 455498
rect -4756 419818 -4574 420054
rect -4338 419818 -4156 420054
rect -4756 419734 -4156 419818
rect -4756 419498 -4574 419734
rect -4338 419498 -4156 419734
rect -4756 384054 -4156 419498
rect -4756 383818 -4574 384054
rect -4338 383818 -4156 384054
rect -4756 383734 -4156 383818
rect -4756 383498 -4574 383734
rect -4338 383498 -4156 383734
rect -4756 348054 -4156 383498
rect -4756 347818 -4574 348054
rect -4338 347818 -4156 348054
rect -4756 347734 -4156 347818
rect -4756 347498 -4574 347734
rect -4338 347498 -4156 347734
rect -4756 312054 -4156 347498
rect -4756 311818 -4574 312054
rect -4338 311818 -4156 312054
rect -4756 311734 -4156 311818
rect -4756 311498 -4574 311734
rect -4338 311498 -4156 311734
rect -4756 276054 -4156 311498
rect -4756 275818 -4574 276054
rect -4338 275818 -4156 276054
rect -4756 275734 -4156 275818
rect -4756 275498 -4574 275734
rect -4338 275498 -4156 275734
rect -4756 240054 -4156 275498
rect -4756 239818 -4574 240054
rect -4338 239818 -4156 240054
rect -4756 239734 -4156 239818
rect -4756 239498 -4574 239734
rect -4338 239498 -4156 239734
rect -4756 204054 -4156 239498
rect -4756 203818 -4574 204054
rect -4338 203818 -4156 204054
rect -4756 203734 -4156 203818
rect -4756 203498 -4574 203734
rect -4338 203498 -4156 203734
rect -4756 168054 -4156 203498
rect -4756 167818 -4574 168054
rect -4338 167818 -4156 168054
rect -4756 167734 -4156 167818
rect -4756 167498 -4574 167734
rect -4338 167498 -4156 167734
rect -4756 132054 -4156 167498
rect -4756 131818 -4574 132054
rect -4338 131818 -4156 132054
rect -4756 131734 -4156 131818
rect -4756 131498 -4574 131734
rect -4338 131498 -4156 131734
rect -4756 96054 -4156 131498
rect -4756 95818 -4574 96054
rect -4338 95818 -4156 96054
rect -4756 95734 -4156 95818
rect -4756 95498 -4574 95734
rect -4338 95498 -4156 95734
rect -4756 60054 -4156 95498
rect -4756 59818 -4574 60054
rect -4338 59818 -4156 60054
rect -4756 59734 -4156 59818
rect -4756 59498 -4574 59734
rect -4338 59498 -4156 59734
rect -4756 24054 -4156 59498
rect -4756 23818 -4574 24054
rect -4338 23818 -4156 24054
rect -4756 23734 -4156 23818
rect -4756 23498 -4574 23734
rect -4338 23498 -4156 23734
rect -4756 -3106 -4156 23498
rect -3836 706678 -3236 706700
rect -3836 706442 -3654 706678
rect -3418 706442 -3236 706678
rect -3836 706358 -3236 706442
rect -3836 706122 -3654 706358
rect -3418 706122 -3236 706358
rect -3836 690054 -3236 706122
rect 587160 706678 587760 706700
rect 587160 706442 587342 706678
rect 587578 706442 587760 706678
rect 587160 706358 587760 706442
rect 587160 706122 587342 706358
rect 587578 706122 587760 706358
rect -3836 689818 -3654 690054
rect -3418 689818 -3236 690054
rect -3836 689734 -3236 689818
rect -3836 689498 -3654 689734
rect -3418 689498 -3236 689734
rect -3836 654054 -3236 689498
rect -3836 653818 -3654 654054
rect -3418 653818 -3236 654054
rect -3836 653734 -3236 653818
rect -3836 653498 -3654 653734
rect -3418 653498 -3236 653734
rect -3836 618054 -3236 653498
rect -3836 617818 -3654 618054
rect -3418 617818 -3236 618054
rect -3836 617734 -3236 617818
rect -3836 617498 -3654 617734
rect -3418 617498 -3236 617734
rect -3836 582054 -3236 617498
rect -3836 581818 -3654 582054
rect -3418 581818 -3236 582054
rect -3836 581734 -3236 581818
rect -3836 581498 -3654 581734
rect -3418 581498 -3236 581734
rect -3836 546054 -3236 581498
rect -3836 545818 -3654 546054
rect -3418 545818 -3236 546054
rect -3836 545734 -3236 545818
rect -3836 545498 -3654 545734
rect -3418 545498 -3236 545734
rect -3836 510054 -3236 545498
rect -3836 509818 -3654 510054
rect -3418 509818 -3236 510054
rect -3836 509734 -3236 509818
rect -3836 509498 -3654 509734
rect -3418 509498 -3236 509734
rect -3836 474054 -3236 509498
rect -3836 473818 -3654 474054
rect -3418 473818 -3236 474054
rect -3836 473734 -3236 473818
rect -3836 473498 -3654 473734
rect -3418 473498 -3236 473734
rect -3836 438054 -3236 473498
rect -3836 437818 -3654 438054
rect -3418 437818 -3236 438054
rect -3836 437734 -3236 437818
rect -3836 437498 -3654 437734
rect -3418 437498 -3236 437734
rect -3836 402054 -3236 437498
rect -3836 401818 -3654 402054
rect -3418 401818 -3236 402054
rect -3836 401734 -3236 401818
rect -3836 401498 -3654 401734
rect -3418 401498 -3236 401734
rect -3836 366054 -3236 401498
rect -3836 365818 -3654 366054
rect -3418 365818 -3236 366054
rect -3836 365734 -3236 365818
rect -3836 365498 -3654 365734
rect -3418 365498 -3236 365734
rect -3836 330054 -3236 365498
rect -3836 329818 -3654 330054
rect -3418 329818 -3236 330054
rect -3836 329734 -3236 329818
rect -3836 329498 -3654 329734
rect -3418 329498 -3236 329734
rect -3836 294054 -3236 329498
rect -3836 293818 -3654 294054
rect -3418 293818 -3236 294054
rect -3836 293734 -3236 293818
rect -3836 293498 -3654 293734
rect -3418 293498 -3236 293734
rect -3836 258054 -3236 293498
rect -3836 257818 -3654 258054
rect -3418 257818 -3236 258054
rect -3836 257734 -3236 257818
rect -3836 257498 -3654 257734
rect -3418 257498 -3236 257734
rect -3836 222054 -3236 257498
rect -3836 221818 -3654 222054
rect -3418 221818 -3236 222054
rect -3836 221734 -3236 221818
rect -3836 221498 -3654 221734
rect -3418 221498 -3236 221734
rect -3836 186054 -3236 221498
rect -3836 185818 -3654 186054
rect -3418 185818 -3236 186054
rect -3836 185734 -3236 185818
rect -3836 185498 -3654 185734
rect -3418 185498 -3236 185734
rect -3836 150054 -3236 185498
rect -3836 149818 -3654 150054
rect -3418 149818 -3236 150054
rect -3836 149734 -3236 149818
rect -3836 149498 -3654 149734
rect -3418 149498 -3236 149734
rect -3836 114054 -3236 149498
rect -3836 113818 -3654 114054
rect -3418 113818 -3236 114054
rect -3836 113734 -3236 113818
rect -3836 113498 -3654 113734
rect -3418 113498 -3236 113734
rect -3836 78054 -3236 113498
rect -3836 77818 -3654 78054
rect -3418 77818 -3236 78054
rect -3836 77734 -3236 77818
rect -3836 77498 -3654 77734
rect -3418 77498 -3236 77734
rect -3836 42054 -3236 77498
rect -3836 41818 -3654 42054
rect -3418 41818 -3236 42054
rect -3836 41734 -3236 41818
rect -3836 41498 -3654 41734
rect -3418 41498 -3236 41734
rect -3836 6054 -3236 41498
rect -3836 5818 -3654 6054
rect -3418 5818 -3236 6054
rect -3836 5734 -3236 5818
rect -3836 5498 -3654 5734
rect -3418 5498 -3236 5734
rect -3836 -2186 -3236 5498
rect -2916 705758 -2316 705780
rect -2916 705522 -2734 705758
rect -2498 705522 -2316 705758
rect -2916 705438 -2316 705522
rect -2916 705202 -2734 705438
rect -2498 705202 -2316 705438
rect -2916 668454 -2316 705202
rect 586240 705758 586840 705780
rect 586240 705522 586422 705758
rect 586658 705522 586840 705758
rect 586240 705438 586840 705522
rect 586240 705202 586422 705438
rect 586658 705202 586840 705438
rect -2916 668218 -2734 668454
rect -2498 668218 -2316 668454
rect -2916 668134 -2316 668218
rect -2916 667898 -2734 668134
rect -2498 667898 -2316 668134
rect -2916 632454 -2316 667898
rect -2916 632218 -2734 632454
rect -2498 632218 -2316 632454
rect -2916 632134 -2316 632218
rect -2916 631898 -2734 632134
rect -2498 631898 -2316 632134
rect -2916 596454 -2316 631898
rect -2916 596218 -2734 596454
rect -2498 596218 -2316 596454
rect -2916 596134 -2316 596218
rect -2916 595898 -2734 596134
rect -2498 595898 -2316 596134
rect -2916 560454 -2316 595898
rect -2916 560218 -2734 560454
rect -2498 560218 -2316 560454
rect -2916 560134 -2316 560218
rect -2916 559898 -2734 560134
rect -2498 559898 -2316 560134
rect -2916 524454 -2316 559898
rect -2916 524218 -2734 524454
rect -2498 524218 -2316 524454
rect -2916 524134 -2316 524218
rect -2916 523898 -2734 524134
rect -2498 523898 -2316 524134
rect -2916 488454 -2316 523898
rect -2916 488218 -2734 488454
rect -2498 488218 -2316 488454
rect -2916 488134 -2316 488218
rect -2916 487898 -2734 488134
rect -2498 487898 -2316 488134
rect -2916 452454 -2316 487898
rect -2916 452218 -2734 452454
rect -2498 452218 -2316 452454
rect -2916 452134 -2316 452218
rect -2916 451898 -2734 452134
rect -2498 451898 -2316 452134
rect -2916 416454 -2316 451898
rect -2916 416218 -2734 416454
rect -2498 416218 -2316 416454
rect -2916 416134 -2316 416218
rect -2916 415898 -2734 416134
rect -2498 415898 -2316 416134
rect -2916 380454 -2316 415898
rect -2916 380218 -2734 380454
rect -2498 380218 -2316 380454
rect -2916 380134 -2316 380218
rect -2916 379898 -2734 380134
rect -2498 379898 -2316 380134
rect -2916 344454 -2316 379898
rect -2916 344218 -2734 344454
rect -2498 344218 -2316 344454
rect -2916 344134 -2316 344218
rect -2916 343898 -2734 344134
rect -2498 343898 -2316 344134
rect -2916 308454 -2316 343898
rect -2916 308218 -2734 308454
rect -2498 308218 -2316 308454
rect -2916 308134 -2316 308218
rect -2916 307898 -2734 308134
rect -2498 307898 -2316 308134
rect -2916 272454 -2316 307898
rect -2916 272218 -2734 272454
rect -2498 272218 -2316 272454
rect -2916 272134 -2316 272218
rect -2916 271898 -2734 272134
rect -2498 271898 -2316 272134
rect -2916 236454 -2316 271898
rect -2916 236218 -2734 236454
rect -2498 236218 -2316 236454
rect -2916 236134 -2316 236218
rect -2916 235898 -2734 236134
rect -2498 235898 -2316 236134
rect -2916 200454 -2316 235898
rect -2916 200218 -2734 200454
rect -2498 200218 -2316 200454
rect -2916 200134 -2316 200218
rect -2916 199898 -2734 200134
rect -2498 199898 -2316 200134
rect -2916 164454 -2316 199898
rect -2916 164218 -2734 164454
rect -2498 164218 -2316 164454
rect -2916 164134 -2316 164218
rect -2916 163898 -2734 164134
rect -2498 163898 -2316 164134
rect -2916 128454 -2316 163898
rect -2916 128218 -2734 128454
rect -2498 128218 -2316 128454
rect -2916 128134 -2316 128218
rect -2916 127898 -2734 128134
rect -2498 127898 -2316 128134
rect -2916 92454 -2316 127898
rect -2916 92218 -2734 92454
rect -2498 92218 -2316 92454
rect -2916 92134 -2316 92218
rect -2916 91898 -2734 92134
rect -2498 91898 -2316 92134
rect -2916 56454 -2316 91898
rect -2916 56218 -2734 56454
rect -2498 56218 -2316 56454
rect -2916 56134 -2316 56218
rect -2916 55898 -2734 56134
rect -2498 55898 -2316 56134
rect -2916 20454 -2316 55898
rect -2916 20218 -2734 20454
rect -2498 20218 -2316 20454
rect -2916 20134 -2316 20218
rect -2916 19898 -2734 20134
rect -2498 19898 -2316 20134
rect -2916 -1266 -2316 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 550587 681052 550653 681053
rect 550587 680988 550588 681052
rect 550652 680988 550653 681052
rect 550587 680987 550653 680988
rect 434667 680916 434733 680917
rect 434667 680852 434668 680916
rect 434732 680852 434733 680916
rect 434667 680851 434733 680852
rect 434670 680645 434730 680851
rect 550590 680645 550650 680987
rect 559787 680780 559853 680781
rect 559787 680716 559788 680780
rect 559852 680716 559853 680780
rect 559787 680715 559853 680716
rect 344875 680644 344941 680645
rect 344875 680580 344876 680644
rect 344940 680580 344941 680644
rect 344875 680579 344941 680580
rect 434667 680644 434733 680645
rect 434667 680580 434668 680644
rect 434732 680580 434733 680644
rect 434667 680579 434733 680580
rect 550587 680644 550653 680645
rect 550587 680580 550588 680644
rect 550652 680580 550653 680644
rect 550587 680579 550653 680580
rect 344878 680458 344938 680579
rect 559051 680508 559117 680509
rect 559051 680444 559052 680508
rect 559116 680506 559117 680508
rect 559116 680446 559298 680506
rect 559116 680444 559117 680446
rect 559051 680443 559117 680444
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect 558870 645010 558930 676142
rect 559238 666178 559298 680446
rect 559419 680372 559485 680373
rect 559419 680308 559420 680372
rect 559484 680308 559485 680372
rect 559419 680307 559485 680308
rect 559422 674250 559482 680307
rect 559790 676378 559850 680715
rect 561995 680644 562061 680645
rect 561995 680580 561996 680644
rect 562060 680580 562061 680644
rect 561995 680579 562061 680580
rect 561259 680508 561325 680509
rect 561259 680444 561260 680508
rect 561324 680444 561325 680508
rect 561259 680443 561325 680444
rect 561627 680508 561693 680509
rect 561627 680444 561628 680508
rect 561692 680444 561693 680508
rect 561627 680443 561693 680444
rect 560707 680372 560773 680373
rect 560707 680308 560708 680372
rect 560772 680308 560773 680372
rect 560707 680307 560773 680308
rect 561075 680372 561141 680373
rect 561075 680308 561076 680372
rect 561140 680308 561141 680372
rect 561075 680307 561141 680308
rect 559422 674190 559666 674250
rect 559606 647050 559666 674190
rect 559974 666030 560254 666090
rect 559974 653170 560034 666030
rect 560710 660650 560770 680307
rect 560342 660590 560770 660650
rect 560342 653850 560402 660590
rect 560342 653790 560954 653850
rect 558686 644950 558930 645010
rect 559238 646990 559666 647050
rect 559790 653110 560034 653170
rect 558686 640250 558746 644950
rect 558686 640190 558930 640250
rect 558870 624610 558930 640190
rect 559238 638210 559298 646990
rect 559790 646370 559850 653110
rect 559790 646310 560034 646370
rect 559974 642290 560034 646310
rect 559974 642230 560402 642290
rect 560342 638210 560402 642230
rect 559238 638150 560770 638210
rect 559054 632710 560034 632770
rect 559054 627330 559114 632710
rect 559974 630730 560034 632710
rect 560342 630730 560402 638150
rect 559974 630670 560402 630730
rect 560710 629370 560770 638150
rect 559238 629310 560770 629370
rect 559238 628690 559298 629310
rect 559238 628630 559850 628690
rect 559054 627270 559298 627330
rect 558870 624550 559114 624610
rect 559054 623250 559114 624550
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect 558870 623190 559114 623250
rect 3141 339692 3207 339693
rect 3141 339628 3142 339692
rect 3206 339690 3207 339692
rect 3206 339630 3434 339690
rect 3206 339628 3207 339630
rect 3141 339627 3207 339628
rect 3374 334216 3434 339630
rect 3190 334156 3434 334216
rect 3190 326770 3250 334156
rect 3190 326710 3434 326770
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect 3374 324050 3434 326710
rect 3190 323990 3434 324050
rect 3190 323370 3250 323990
rect 3144 323310 3250 323370
rect 3144 321061 3204 323310
rect 3141 321060 3207 321061
rect 3141 320996 3142 321060
rect 3206 320996 3207 321060
rect 3141 320995 3207 320996
rect 558870 309090 558930 623190
rect 559238 540970 559298 627270
rect 559790 618490 559850 628630
rect 560894 621210 560954 653790
rect 559606 618430 559850 618490
rect 560526 621150 560954 621210
rect 559238 540910 559482 540970
rect 559422 532130 559482 540910
rect 559606 534850 559666 618430
rect 560526 615090 560586 621150
rect 560526 615030 560770 615090
rect 560710 608290 560770 615030
rect 560342 608230 560770 608290
rect 560342 604890 560402 608230
rect 560342 604830 560586 604890
rect 560526 594010 560586 604830
rect 560526 593950 560770 594010
rect 560710 579050 560770 593950
rect 560526 578990 560770 579050
rect 560526 562730 560586 578990
rect 560526 562670 560770 562730
rect 560710 553890 560770 562670
rect 560710 553830 560954 553890
rect 560894 543690 560954 553830
rect 560342 543630 560954 543690
rect 560342 534850 560402 543630
rect 559606 534790 559850 534850
rect 560342 534790 560770 534850
rect 559790 532130 559850 534790
rect 559238 532070 559482 532130
rect 559606 532070 559850 532130
rect 558870 309030 559114 309090
rect 559054 295490 559114 309030
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect 558870 295430 559114 295490
rect 1347 221508 1413 221509
rect 1347 221444 1348 221508
rect 1412 221444 1413 221508
rect 1347 221443 1413 221444
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect 1350 214573 1410 221443
rect 1347 214572 1413 214573
rect 1347 214508 1348 214572
rect 1412 214508 1413 214572
rect 1347 214507 1413 214508
rect 1531 198252 1597 198253
rect 1531 198188 1532 198252
rect 1596 198188 1597 198252
rect 1531 198187 1597 198188
rect 1534 185330 1594 198187
rect 2865 185332 2931 185333
rect 2865 185330 2866 185332
rect 1534 185270 2866 185330
rect 2865 185268 2866 185270
rect 2930 185268 2931 185332
rect 2865 185267 2931 185268
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect 1531 173092 1597 173093
rect 1531 173028 1532 173092
rect 1596 173028 1597 173092
rect 1531 173027 1597 173028
rect 1534 167653 1594 173027
rect 1531 167652 1597 167653
rect 1531 167588 1532 167652
rect 1596 167588 1597 167652
rect 1531 167587 1597 167588
rect 1531 146980 1597 146981
rect 1531 146916 1532 146980
rect 1596 146916 1597 146980
rect 1531 146915 1597 146916
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect 1534 138685 1594 146915
rect 1531 138684 1597 138685
rect 1531 138620 1532 138684
rect 1596 138620 1597 138684
rect 1531 138619 1597 138620
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect 1347 108220 1413 108221
rect 1347 108156 1348 108220
rect 1412 108156 1413 108220
rect 1347 108155 1413 108156
rect 1350 96250 1410 108155
rect 1531 107132 1597 107133
rect 1531 107068 1532 107132
rect 1596 107130 1597 107132
rect 1596 107070 3066 107130
rect 1596 107068 1597 107070
rect 1531 107067 1597 107068
rect 1531 99652 1597 99653
rect 1531 99588 1532 99652
rect 1596 99650 1597 99652
rect 3006 99650 3066 107070
rect 1596 99590 3066 99650
rect 1596 99588 1597 99590
rect 1531 99587 1597 99588
rect 1350 96190 3572 96250
rect 3512 96117 3572 96190
rect 3509 96116 3575 96117
rect 3509 96052 3510 96116
rect 3574 96052 3575 96116
rect 3509 96051 3575 96052
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect 1531 45932 1597 45933
rect 1531 45868 1532 45932
rect 1596 45868 1597 45932
rect 1531 45867 1597 45868
rect 1534 43890 1594 45867
rect 1534 43830 3802 43890
rect 3742 40357 3802 43830
rect 3739 40356 3805 40357
rect 3739 40292 3740 40356
rect 3804 40292 3805 40356
rect 3739 40291 3805 40292
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect 982 25805 1042 34222
rect 1350 29749 1410 36262
rect 1718 33690 1778 35582
rect 1534 33630 1778 33690
rect 1534 33285 1594 33630
rect 1531 33284 1597 33285
rect 1531 33220 1532 33284
rect 1596 33220 1597 33284
rect 1531 33219 1597 33220
rect 1531 30292 1597 30293
rect 1531 30228 1532 30292
rect 1596 30290 1597 30292
rect 1718 30290 1778 32862
rect 1596 30230 1778 30290
rect 1596 30228 1597 30230
rect 1531 30227 1597 30228
rect 1347 29748 1413 29749
rect 1347 29684 1348 29748
rect 1412 29684 1413 29748
rect 1347 29683 1413 29684
rect 1350 26893 1410 28782
rect 1531 27028 1597 27029
rect 1531 26964 1532 27028
rect 1596 27026 1597 27028
rect 1718 27026 1778 29462
rect 1596 26966 1778 27026
rect 1596 26964 1597 26966
rect 1531 26963 1597 26964
rect 1347 26892 1413 26893
rect 1347 26828 1348 26892
rect 1412 26828 1413 26892
rect 1347 26827 1413 26828
rect 979 25804 1045 25805
rect 979 25740 980 25804
rect 1044 25740 1045 25804
rect 979 25739 1045 25740
rect 1166 19821 1226 25382
rect 1534 20093 1594 24702
rect 1531 20092 1597 20093
rect 1531 20028 1532 20092
rect 1596 20028 1597 20092
rect 1531 20027 1597 20028
rect 1347 19956 1413 19957
rect 1347 19892 1348 19956
rect 1412 19892 1413 19956
rect 1347 19891 1413 19892
rect 1163 19820 1229 19821
rect 1163 19756 1164 19820
rect 1228 19756 1229 19820
rect 1163 19755 1229 19756
rect 1350 16010 1410 19891
rect 1531 18052 1597 18053
rect 1531 17988 1532 18052
rect 1596 18050 1597 18052
rect 1902 18050 1962 26062
rect 1596 17990 1962 18050
rect 1596 17988 1597 17990
rect 1531 17987 1597 17988
rect 558870 16098 558930 295430
rect 559238 212530 559298 532070
rect 559606 499490 559666 532070
rect 560710 530090 560770 534790
rect 560526 530030 560770 530090
rect 560526 524650 560586 530030
rect 560342 524590 560586 524650
rect 560342 519890 560402 524590
rect 560342 519830 560586 519890
rect 560526 518530 560586 519830
rect 560158 518470 560586 518530
rect 560158 509690 560218 518470
rect 560158 509630 560770 509690
rect 560710 504930 560770 509630
rect 560710 504870 560954 504930
rect 559606 499430 560034 499490
rect 559974 489970 560034 499430
rect 560894 495410 560954 504870
rect 559606 489910 560034 489970
rect 560526 495350 560954 495410
rect 559606 451210 559666 489910
rect 560526 485210 560586 495350
rect 560526 485150 560770 485210
rect 560710 480450 560770 485150
rect 560710 480390 560954 480450
rect 560894 470930 560954 480390
rect 560710 470870 560954 470930
rect 560710 451210 560770 470870
rect 559606 451150 559850 451210
rect 559790 441690 559850 451150
rect 560342 451150 560770 451210
rect 560342 445770 560402 451150
rect 560342 445710 560770 445770
rect 559606 441630 559850 441690
rect 559606 402930 559666 441630
rect 560710 436930 560770 445710
rect 560526 436870 560770 436930
rect 560526 428770 560586 436870
rect 560158 428710 560586 428770
rect 560158 418570 560218 428710
rect 560158 418510 560770 418570
rect 560710 412450 560770 418510
rect 560710 412390 560954 412450
rect 560894 407690 560954 412390
rect 560342 407630 560954 407690
rect 560342 402930 560402 407630
rect 559606 402870 560034 402930
rect 560342 402870 560586 402930
rect 559974 393410 560034 402870
rect 560526 398170 560586 402870
rect 560526 398110 560770 398170
rect 559606 393350 560034 393410
rect 559606 354650 559666 393350
rect 560710 380490 560770 398110
rect 559790 380430 560770 380490
rect 559790 379130 559850 380430
rect 559790 379070 560218 379130
rect 560158 369610 560218 379070
rect 560158 369550 560586 369610
rect 560526 360090 560586 369550
rect 560526 360030 560770 360090
rect 559606 354590 559850 354650
rect 559790 343770 559850 354590
rect 560710 345130 560770 360030
rect 560710 345070 560954 345130
rect 559606 343710 559850 343770
rect 559606 286650 559666 343710
rect 560894 334930 560954 345070
rect 560710 334870 560954 334930
rect 560710 333570 560770 334870
rect 560158 333510 560770 333570
rect 560158 325410 560218 333510
rect 560158 325350 560402 325410
rect 560342 324050 560402 325350
rect 560342 323990 560586 324050
rect 560526 323370 560586 323990
rect 560526 323310 560770 323370
rect 560710 306370 560770 323310
rect 560710 306310 560954 306370
rect 560894 290730 560954 306310
rect 559422 286590 559666 286650
rect 560526 290670 560954 290730
rect 560526 286650 560586 290670
rect 560526 286590 560770 286650
rect 559422 278490 559482 286590
rect 560710 283250 560770 286590
rect 560342 283190 560770 283250
rect 559422 278430 559666 278490
rect 559606 277130 559666 278430
rect 559606 277070 559850 277130
rect 559790 268290 559850 277070
rect 560342 272370 560402 283190
rect 560342 272310 560586 272370
rect 559606 268230 559850 268290
rect 559238 212470 559482 212530
rect 559422 207770 559482 212470
rect 559238 207710 559482 207770
rect 559238 36498 559298 207710
rect 559606 35818 559666 268230
rect 560526 264210 560586 272310
rect 560342 264150 560586 264210
rect 560342 262850 560402 264150
rect 560342 262790 560770 262850
rect 560710 254010 560770 262790
rect 560342 253950 560770 254010
rect 560342 233610 560402 253950
rect 560342 233550 560770 233610
rect 560710 228170 560770 233550
rect 560710 228110 560954 228170
rect 560894 223410 560954 228110
rect 560526 223350 560954 223410
rect 560526 215930 560586 223350
rect 560526 215870 560770 215930
rect 560710 214570 560770 215870
rect 560342 214510 560770 214570
rect 560342 207090 560402 214510
rect 560342 207030 560770 207090
rect 560710 205050 560770 207030
rect 560526 204990 560770 205050
rect 560526 196210 560586 204990
rect 561078 197570 561138 680307
rect 560342 196150 560586 196210
rect 560710 197510 561138 197570
rect 560342 190090 560402 196150
rect 560710 194170 560770 197510
rect 561262 196210 561322 680443
rect 561078 196150 561322 196210
rect 561078 194850 561138 196150
rect 561078 194790 561322 194850
rect 560710 194110 561138 194170
rect 560342 190030 560586 190090
rect 560526 187370 560586 190030
rect 560342 187310 560586 187370
rect 560342 186010 560402 187310
rect 560342 185950 560770 186010
rect 560710 176490 560770 185950
rect 560710 176430 560954 176490
rect 560894 166970 560954 176430
rect 560526 166910 560954 166970
rect 560526 156770 560586 166910
rect 560526 156710 560770 156770
rect 560710 152010 560770 156710
rect 560710 151950 560954 152010
rect 560894 142490 560954 151950
rect 560710 142430 560954 142490
rect 560710 131610 560770 142430
rect 560710 131550 560954 131610
rect 560894 128210 560954 131550
rect 560710 128150 560954 128210
rect 560710 122770 560770 128150
rect 560710 122710 560954 122770
rect 560894 113250 560954 122710
rect 560710 113190 560954 113250
rect 560710 109170 560770 113190
rect 560710 109110 560954 109170
rect 560894 104410 560954 109110
rect 560710 104350 560954 104410
rect 560710 103730 560770 104350
rect 560526 103670 560770 103730
rect 560526 99650 560586 103670
rect 560526 99590 560770 99650
rect 560710 98290 560770 99590
rect 560158 98230 560770 98290
rect 560158 90810 560218 98230
rect 560158 90750 560402 90810
rect 560342 76530 560402 90750
rect 560342 76470 560586 76530
rect 560526 69730 560586 76470
rect 560526 69670 560770 69730
rect 560710 54770 560770 69670
rect 560342 54710 560770 54770
rect 560342 50010 560402 54710
rect 560342 49950 560954 50010
rect 560894 45250 560954 49950
rect 560526 45190 560954 45250
rect 560526 40490 560586 45190
rect 560526 40430 560770 40490
rect 559790 24938 559850 34902
rect 560710 29018 560770 40430
rect 561078 33098 561138 194110
rect 561262 33690 561322 194790
rect 561262 33630 561506 33690
rect 561446 32418 561506 33630
rect 561630 33010 561690 680443
rect 561998 35138 562058 680579
rect 563099 680508 563165 680509
rect 563099 680444 563100 680508
rect 563164 680444 563165 680508
rect 563099 680443 563165 680444
rect 564571 680508 564637 680509
rect 564571 680444 564572 680508
rect 564636 680444 564637 680508
rect 567147 680508 567213 680509
rect 564571 680443 564637 680444
rect 562363 680372 562429 680373
rect 562363 680308 562364 680372
rect 562428 680308 562429 680372
rect 562363 680307 562429 680308
rect 562366 34458 562426 680307
rect 561630 32950 561874 33010
rect 561814 29698 561874 32950
rect 1350 15950 2330 16010
rect 982 12885 1042 15182
rect 979 12884 1045 12885
rect 979 12820 980 12884
rect 1044 12820 1045 12884
rect 979 12819 1045 12820
rect 1534 8805 1594 10422
rect 1531 8804 1597 8805
rect 1531 8740 1532 8804
rect 1596 8740 1597 8804
rect 1531 8739 1597 8740
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect 1902 101 1962 13822
rect 2270 9890 2330 15950
rect 4846 12018 4906 13822
rect 558686 9890 558746 11782
rect 559790 11338 559850 18582
rect 2270 9830 2882 9890
rect 558686 9830 558930 9890
rect 2822 1189 2882 9830
rect 19931 7988 19997 7989
rect 19931 7938 19932 7988
rect 19996 7938 19997 7988
rect 3003 1732 3069 1733
rect 3003 1668 3004 1732
rect 3068 1668 3069 1732
rect 3003 1667 3069 1668
rect 3006 1461 3066 1667
rect 3003 1460 3069 1461
rect 3003 1396 3004 1460
rect 3068 1396 3069 1460
rect 3003 1395 3069 1396
rect 2819 1188 2885 1189
rect 2819 1124 2820 1188
rect 2884 1124 2885 1188
rect 4846 1138 4906 7022
rect 125514 3030 125610 3090
rect 10915 1188 10981 1189
rect 2819 1123 2885 1124
rect 10915 1124 10916 1188
rect 10980 1124 10981 1188
rect 10915 1123 10981 1124
rect 10547 852 10548 902
rect 10612 852 10613 902
rect 10547 851 10613 852
rect 10918 458 10978 1123
rect 14966 373 15026 2942
rect 19195 852 19196 902
rect 19260 852 19261 902
rect 19195 851 19261 852
rect 28211 852 28212 902
rect 28276 852 28277 902
rect 28211 851 28277 852
rect 28950 458 29010 2942
rect 52318 1597 52378 2942
rect 65198 2350 67834 2410
rect 65011 1732 65077 1733
rect 65011 1730 65012 1732
rect 64646 1670 65012 1730
rect 52315 1596 52381 1597
rect 52315 1532 52316 1596
rect 52380 1532 52381 1596
rect 58571 1596 58637 1597
rect 58571 1594 58572 1596
rect 52315 1531 52381 1532
rect 56366 1534 58572 1594
rect 56366 1461 56426 1534
rect 58571 1532 58572 1534
rect 58636 1532 58637 1596
rect 58571 1531 58637 1532
rect 39067 1460 39133 1461
rect 39067 1396 39068 1460
rect 39132 1396 39133 1460
rect 39067 1395 39133 1396
rect 56363 1460 56429 1461
rect 56363 1396 56364 1460
rect 56428 1396 56429 1460
rect 56363 1395 56429 1396
rect 39070 1138 39130 1395
rect 64646 1189 64706 1670
rect 65011 1668 65012 1670
rect 65076 1668 65077 1732
rect 65011 1667 65077 1668
rect 39435 1188 39501 1189
rect 39435 1124 39436 1188
rect 39500 1124 39501 1188
rect 60595 1188 60661 1189
rect 39435 1123 39501 1124
rect 39438 458 39498 1123
rect 60595 1124 60596 1188
rect 60660 1124 60661 1188
rect 60595 1123 60661 1124
rect 64643 1188 64709 1189
rect 64643 1124 64644 1188
rect 64708 1124 64709 1188
rect 65198 1186 65258 2350
rect 67774 1866 67834 2350
rect 67774 1806 73354 1866
rect 68691 1732 68757 1733
rect 66670 1670 67282 1730
rect 66670 1597 66730 1670
rect 66667 1596 66733 1597
rect 66667 1532 66668 1596
rect 66732 1532 66733 1596
rect 66667 1531 66733 1532
rect 64643 1123 64709 1124
rect 65014 1126 65258 1186
rect 66851 1188 66917 1189
rect 66851 1138 66852 1188
rect 66916 1138 66917 1188
rect 60598 1050 60658 1123
rect 63723 1052 63789 1053
rect 63723 1050 63724 1052
rect 60598 990 63724 1050
rect 63723 988 63724 990
rect 63788 988 63789 1052
rect 63723 987 63789 988
rect 14963 372 15029 373
rect 14963 308 14964 372
rect 15028 308 15029 372
rect 14963 307 15029 308
rect 65014 370 65074 1126
rect 67222 1050 67282 1670
rect 68691 1668 68692 1732
rect 68756 1730 68757 1732
rect 72555 1732 72621 1733
rect 72555 1730 72556 1732
rect 68756 1670 72556 1730
rect 68756 1668 68757 1670
rect 68691 1667 68757 1668
rect 72555 1668 72556 1670
rect 72620 1668 72621 1732
rect 72555 1667 72621 1668
rect 73294 1597 73354 1806
rect 73107 1596 73173 1597
rect 73107 1532 73108 1596
rect 73172 1532 73173 1596
rect 73107 1531 73173 1532
rect 73291 1596 73357 1597
rect 73291 1532 73292 1596
rect 73356 1532 73357 1596
rect 74950 1594 75010 2942
rect 76422 2410 76482 2942
rect 76422 2350 76666 2410
rect 75315 1732 75381 1733
rect 75315 1668 75316 1732
rect 75380 1730 75381 1732
rect 76051 1732 76117 1733
rect 76051 1730 76052 1732
rect 75380 1670 76052 1730
rect 75380 1668 75381 1670
rect 75315 1667 75381 1668
rect 76051 1668 76052 1670
rect 76116 1668 76117 1732
rect 76051 1667 76117 1668
rect 75499 1596 75565 1597
rect 75499 1594 75500 1596
rect 74950 1534 75500 1594
rect 73291 1531 73357 1532
rect 75499 1532 75500 1534
rect 75564 1532 75565 1596
rect 76419 1596 76485 1597
rect 76419 1594 76420 1596
rect 75499 1531 75565 1532
rect 75686 1534 76420 1594
rect 67222 990 68974 1050
rect 73110 1053 73170 1531
rect 73475 1460 73541 1461
rect 73475 1396 73476 1460
rect 73540 1396 73541 1460
rect 73475 1395 73541 1396
rect 73478 1053 73538 1395
rect 72923 1052 72989 1053
rect 72923 988 72924 1052
rect 72988 988 72989 1052
rect 72923 987 72989 988
rect 73107 1052 73173 1053
rect 73107 988 73108 1052
rect 73172 988 73173 1052
rect 73107 987 73173 988
rect 73475 1052 73541 1053
rect 73475 988 73476 1052
rect 73540 988 73541 1052
rect 73475 987 73541 988
rect 72926 914 72986 987
rect 75686 914 75746 1534
rect 76419 1532 76420 1534
rect 76484 1532 76485 1596
rect 76606 1594 76666 2350
rect 76790 2350 77586 2410
rect 76790 1733 76850 2350
rect 77526 1866 77586 2350
rect 78630 1866 78690 2942
rect 82310 1866 82370 2942
rect 91510 1866 91570 2942
rect 94822 2410 94882 2942
rect 95742 2410 95802 2942
rect 92062 2350 93226 2410
rect 94822 2350 95250 2410
rect 91737 1868 91803 1869
rect 91737 1866 91738 1868
rect 77526 1806 78690 1866
rect 81758 1806 82370 1866
rect 88014 1806 88442 1866
rect 91510 1806 91738 1866
rect 76787 1732 76853 1733
rect 76787 1668 76788 1732
rect 76852 1668 76853 1732
rect 81758 1730 81818 1806
rect 88014 1733 88074 1806
rect 76787 1667 76853 1668
rect 76974 1670 81818 1730
rect 82491 1732 82557 1733
rect 76974 1594 77034 1670
rect 82491 1668 82492 1732
rect 82556 1730 82557 1732
rect 83595 1732 83661 1733
rect 82556 1670 82922 1730
rect 82556 1668 82557 1670
rect 82491 1667 82557 1668
rect 76606 1534 77034 1594
rect 82862 1594 82922 1670
rect 83595 1668 83596 1732
rect 83660 1730 83661 1732
rect 85803 1732 85869 1733
rect 85803 1730 85804 1732
rect 83660 1670 85804 1730
rect 83660 1668 83661 1670
rect 83595 1667 83661 1668
rect 85803 1668 85804 1670
rect 85868 1668 85869 1732
rect 85803 1667 85869 1668
rect 88011 1732 88077 1733
rect 88011 1668 88012 1732
rect 88076 1668 88077 1732
rect 88011 1667 88077 1668
rect 88195 1732 88261 1733
rect 88195 1668 88196 1732
rect 88260 1668 88261 1732
rect 88382 1730 88442 1806
rect 91737 1804 91738 1806
rect 91802 1804 91803 1868
rect 92062 1866 92122 2350
rect 93166 1866 93226 2350
rect 91737 1803 91803 1804
rect 91924 1806 92122 1866
rect 92614 1806 93042 1866
rect 93166 1806 95066 1866
rect 91924 1730 91984 1806
rect 88382 1670 91984 1730
rect 88195 1667 88261 1668
rect 83043 1596 83109 1597
rect 83043 1594 83044 1596
rect 82862 1534 83044 1594
rect 76419 1531 76485 1532
rect 83043 1532 83044 1534
rect 83108 1532 83109 1596
rect 83043 1531 83109 1532
rect 83414 1534 85682 1594
rect 83414 1461 83474 1534
rect 83411 1460 83477 1461
rect 72926 854 75746 914
rect 78814 1398 83290 1458
rect 73478 582 76298 642
rect 73478 458 73538 582
rect 74211 508 74277 509
rect 74211 506 74212 508
rect 63542 310 65074 370
rect 61147 236 61213 237
rect 61147 172 61148 236
rect 61212 234 61213 236
rect 63542 234 63602 310
rect 61212 174 63602 234
rect 73846 446 74212 506
rect 73846 237 73906 446
rect 74211 444 74212 446
rect 74276 444 74277 508
rect 76051 508 76117 509
rect 74211 443 74277 444
rect 73843 236 73909 237
rect 61212 172 61213 174
rect 61147 171 61213 172
rect 73843 172 73844 236
rect 73908 172 73909 236
rect 76051 444 76052 508
rect 76116 444 76117 508
rect 76238 506 76298 582
rect 78627 508 78693 509
rect 78627 506 78628 508
rect 76238 446 78628 506
rect 76051 443 76117 444
rect 78627 444 78628 446
rect 78692 444 78693 508
rect 78627 443 78693 444
rect 76054 370 76114 443
rect 78814 370 78874 1398
rect 83230 1325 83290 1398
rect 83411 1396 83412 1460
rect 83476 1396 83477 1460
rect 83411 1395 83477 1396
rect 83043 1324 83109 1325
rect 80286 1262 82922 1322
rect 80286 509 80346 1262
rect 82307 1188 82373 1189
rect 82307 1124 82308 1188
rect 82372 1186 82373 1188
rect 82675 1188 82741 1189
rect 82675 1186 82676 1188
rect 82372 1126 82676 1186
rect 82372 1124 82373 1126
rect 82307 1123 82373 1124
rect 82675 1124 82676 1126
rect 82740 1124 82741 1188
rect 82675 1123 82741 1124
rect 82310 990 82738 1050
rect 82310 917 82370 990
rect 82678 917 82738 990
rect 82307 916 82373 917
rect 82307 852 82308 916
rect 82372 852 82373 916
rect 82307 851 82373 852
rect 82675 916 82741 917
rect 82675 852 82676 916
rect 82740 852 82741 916
rect 82675 851 82741 852
rect 79363 508 79429 509
rect 79363 444 79364 508
rect 79428 444 79429 508
rect 79363 443 79429 444
rect 80283 508 80349 509
rect 80283 444 80284 508
rect 80348 444 80349 508
rect 80283 443 80349 444
rect 79366 370 79426 443
rect 76054 310 78874 370
rect 79182 310 79426 370
rect 73843 171 73909 172
rect 1899 100 1965 101
rect 1899 36 1900 100
rect 1964 36 1965 100
rect 1899 35 1965 36
rect 74211 100 74277 101
rect 74211 36 74212 100
rect 74276 98 74277 100
rect 74582 98 74642 222
rect 74276 38 74642 98
rect 78627 100 78693 101
rect 74276 36 74277 38
rect 74211 35 74277 36
rect 78627 36 78628 100
rect 78692 98 78693 100
rect 79182 98 79242 310
rect 82307 236 82373 237
rect 82307 172 82308 236
rect 82372 172 82373 236
rect 82307 171 82373 172
rect 78692 38 79242 98
rect 81387 100 81453 101
rect 78692 36 78693 38
rect 78627 35 78693 36
rect 81387 36 81388 100
rect 81452 98 81453 100
rect 82310 98 82370 171
rect 81452 38 82370 98
rect 82862 98 82922 1262
rect 83043 1260 83044 1324
rect 83108 1260 83109 1324
rect 83043 1259 83109 1260
rect 83227 1324 83293 1325
rect 83227 1260 83228 1324
rect 83292 1260 83293 1324
rect 83227 1259 83293 1260
rect 83046 1186 83106 1259
rect 83046 1126 83474 1186
rect 83414 1053 83474 1126
rect 83227 1052 83293 1053
rect 83227 988 83228 1052
rect 83292 988 83293 1052
rect 83227 987 83293 988
rect 83411 1052 83477 1053
rect 83411 988 83412 1052
rect 83476 988 83477 1052
rect 83411 987 83477 988
rect 83043 100 83109 101
rect 83043 98 83044 100
rect 82862 38 83044 98
rect 81452 36 81453 38
rect 81387 35 81453 36
rect 83043 36 83044 38
rect 83108 36 83109 100
rect 83230 98 83290 987
rect 85622 237 85682 1534
rect 88198 1138 88258 1667
rect 92614 1594 92674 1806
rect 92982 1733 93042 1806
rect 92795 1732 92861 1733
rect 92795 1668 92796 1732
rect 92860 1668 92861 1732
rect 92795 1667 92861 1668
rect 92979 1732 93045 1733
rect 92979 1668 92980 1732
rect 93044 1668 93045 1732
rect 92979 1667 93045 1668
rect 94451 1732 94517 1733
rect 94451 1668 94452 1732
rect 94516 1730 94517 1732
rect 94516 1670 94882 1730
rect 94516 1668 94517 1670
rect 94451 1667 94517 1668
rect 88750 1534 92674 1594
rect 92798 1594 92858 1667
rect 94822 1597 94882 1670
rect 94819 1596 94885 1597
rect 92798 1534 94514 1594
rect 88750 778 88810 1534
rect 90590 1398 94330 1458
rect 90590 1189 90650 1398
rect 90955 1324 91021 1325
rect 90955 1260 90956 1324
rect 91020 1260 91021 1324
rect 90955 1259 91021 1260
rect 91326 1262 92306 1322
rect 90587 1188 90653 1189
rect 90587 1124 90588 1188
rect 90652 1124 90653 1188
rect 90587 1123 90653 1124
rect 87278 718 88810 778
rect 90958 778 91018 1259
rect 91326 917 91386 1262
rect 91323 916 91389 917
rect 91323 852 91324 916
rect 91388 852 91389 916
rect 92246 917 92306 1262
rect 92427 1188 92493 1189
rect 92427 1124 92428 1188
rect 92492 1124 92493 1188
rect 92427 1123 92493 1124
rect 92243 916 92309 917
rect 91323 851 91389 852
rect 91691 852 91692 902
rect 91756 852 91757 902
rect 91691 851 91757 852
rect 92243 852 92244 916
rect 92308 852 92309 916
rect 92243 851 92309 852
rect 91875 780 91941 781
rect 91875 778 91876 780
rect 90958 718 91876 778
rect 87278 237 87338 718
rect 91875 716 91876 718
rect 91940 716 91941 780
rect 91875 715 91941 716
rect 92430 642 92490 1123
rect 87462 582 92490 642
rect 85435 236 85501 237
rect 85435 172 85436 236
rect 85500 172 85501 236
rect 85435 171 85501 172
rect 85619 236 85685 237
rect 85619 172 85620 236
rect 85684 172 85685 236
rect 85619 171 85685 172
rect 87275 236 87341 237
rect 87275 172 87276 236
rect 87340 172 87341 236
rect 87275 171 87341 172
rect 84331 100 84397 101
rect 84331 98 84332 100
rect 83230 38 84332 98
rect 83043 35 83109 36
rect 84331 36 84332 38
rect 84396 36 84397 100
rect 85438 98 85498 171
rect 87462 98 87522 582
rect 92762 310 93226 370
rect 93166 237 93226 310
rect 92979 236 93045 237
rect 92979 172 92980 236
rect 93044 172 93045 236
rect 92979 171 93045 172
rect 93163 236 93229 237
rect 93163 172 93164 236
rect 93228 172 93229 236
rect 94270 237 94330 1398
rect 94454 778 94514 1534
rect 94819 1532 94820 1596
rect 94884 1532 94885 1596
rect 94819 1531 94885 1532
rect 95006 1458 95066 1806
rect 95190 1594 95250 2350
rect 95374 2350 95802 2410
rect 95374 1733 95434 2350
rect 96846 1866 96906 2942
rect 95742 1806 96906 1866
rect 95371 1732 95437 1733
rect 95371 1668 95372 1732
rect 95436 1668 95437 1732
rect 95371 1667 95437 1668
rect 95555 1732 95621 1733
rect 95555 1668 95556 1732
rect 95620 1668 95621 1732
rect 95555 1667 95621 1668
rect 95558 1594 95618 1667
rect 95742 1597 95802 1806
rect 100339 1732 100405 1733
rect 100339 1668 100340 1732
rect 100404 1730 100405 1732
rect 100404 1670 102610 1730
rect 100404 1668 100405 1670
rect 100339 1667 100405 1668
rect 95190 1534 95618 1594
rect 95739 1596 95805 1597
rect 95739 1532 95740 1596
rect 95804 1532 95805 1596
rect 101811 1596 101877 1597
rect 101811 1594 101812 1596
rect 95739 1531 95805 1532
rect 95926 1534 101812 1594
rect 95926 1458 95986 1534
rect 101811 1532 101812 1534
rect 101876 1532 101877 1596
rect 101811 1531 101877 1532
rect 101075 1460 101141 1461
rect 101075 1458 101076 1460
rect 95006 1398 95986 1458
rect 97766 1398 101076 1458
rect 97766 1325 97826 1398
rect 101075 1396 101076 1398
rect 101140 1396 101141 1460
rect 101075 1395 101141 1396
rect 101262 1398 102426 1458
rect 101262 1325 101322 1398
rect 102366 1325 102426 1398
rect 96475 1324 96541 1325
rect 96475 1260 96476 1324
rect 96540 1260 96541 1324
rect 96475 1259 96541 1260
rect 97763 1324 97829 1325
rect 97763 1260 97764 1324
rect 97828 1260 97829 1324
rect 100339 1324 100405 1325
rect 100339 1322 100340 1324
rect 97763 1259 97829 1260
rect 97950 1262 100340 1322
rect 96478 1186 96538 1259
rect 97950 1186 98010 1262
rect 100339 1260 100340 1262
rect 100404 1260 100405 1324
rect 100339 1259 100405 1260
rect 101259 1324 101325 1325
rect 101259 1260 101260 1324
rect 101324 1260 101325 1324
rect 101259 1259 101325 1260
rect 102179 1324 102245 1325
rect 102179 1260 102180 1324
rect 102244 1260 102245 1324
rect 102179 1259 102245 1260
rect 102363 1324 102429 1325
rect 102363 1260 102364 1324
rect 102428 1260 102429 1324
rect 102550 1322 102610 1670
rect 102734 1458 102794 2942
rect 103654 2350 116042 2410
rect 103283 1596 103349 1597
rect 103283 1532 103284 1596
rect 103348 1594 103349 1596
rect 103654 1594 103714 2350
rect 115982 1866 116042 2350
rect 125550 1866 125610 3030
rect 126102 2410 126162 2942
rect 127206 2410 127266 2942
rect 126102 2350 126530 2410
rect 111198 1806 111810 1866
rect 115982 1806 124690 1866
rect 125550 1806 126162 1866
rect 126470 1818 126530 2350
rect 126700 2350 127266 2410
rect 127942 2350 134258 2410
rect 111198 1597 111258 1806
rect 111563 1732 111629 1733
rect 111563 1730 111564 1732
rect 111382 1670 111564 1730
rect 103348 1534 103714 1594
rect 111195 1596 111261 1597
rect 103348 1532 103349 1534
rect 103283 1531 103349 1532
rect 111195 1532 111196 1596
rect 111260 1532 111261 1596
rect 111195 1531 111261 1532
rect 102915 1460 102981 1461
rect 102915 1458 102916 1460
rect 102734 1398 102916 1458
rect 102915 1396 102916 1398
rect 102980 1396 102981 1460
rect 102915 1395 102981 1396
rect 103102 1398 109234 1458
rect 103102 1322 103162 1398
rect 102550 1262 103162 1322
rect 103283 1324 103349 1325
rect 102363 1259 102429 1260
rect 103283 1260 103284 1324
rect 103348 1322 103349 1324
rect 103348 1262 107762 1322
rect 103348 1260 103349 1262
rect 103283 1259 103349 1260
rect 96478 1126 98010 1186
rect 101259 1188 101325 1189
rect 101259 1124 101260 1188
rect 101324 1124 101325 1188
rect 102182 1186 102242 1259
rect 107147 1188 107213 1189
rect 107147 1186 107148 1188
rect 102182 1126 104634 1186
rect 101259 1123 101325 1124
rect 101262 1050 101322 1123
rect 101262 990 102978 1050
rect 102918 781 102978 990
rect 102363 780 102429 781
rect 102363 778 102364 780
rect 94454 718 102364 778
rect 102363 716 102364 718
rect 102428 716 102429 780
rect 102363 715 102429 716
rect 102915 780 102981 781
rect 102915 716 102916 780
rect 102980 716 102981 780
rect 102915 715 102981 716
rect 102550 582 103346 642
rect 102550 509 102610 582
rect 103286 509 103346 582
rect 102547 508 102613 509
rect 102547 444 102548 508
rect 102612 444 102613 508
rect 102547 443 102613 444
rect 103283 508 103349 509
rect 103283 444 103284 508
rect 103348 444 103349 508
rect 104574 458 104634 1126
rect 104942 1126 107148 1186
rect 104942 1050 105002 1126
rect 107147 1124 107148 1126
rect 107212 1124 107213 1188
rect 107515 1188 107581 1189
rect 107515 1186 107516 1188
rect 107147 1123 107213 1124
rect 107334 1126 107516 1186
rect 107334 1050 107394 1126
rect 107515 1124 107516 1126
rect 107580 1124 107581 1188
rect 107515 1123 107581 1124
rect 107702 1050 107762 1262
rect 104758 990 105002 1050
rect 106782 990 107394 1050
rect 107518 990 107762 1050
rect 109174 1050 109234 1398
rect 111382 1189 111442 1670
rect 111563 1668 111564 1670
rect 111628 1668 111629 1732
rect 111750 1730 111810 1806
rect 120763 1732 120829 1733
rect 120763 1730 120764 1732
rect 111750 1670 120764 1730
rect 111563 1667 111629 1668
rect 120763 1668 120764 1670
rect 120828 1668 120829 1732
rect 124443 1732 124509 1733
rect 124443 1730 124444 1732
rect 120763 1667 120829 1668
rect 122974 1670 124444 1730
rect 122974 1594 123034 1670
rect 124443 1668 124444 1670
rect 124508 1668 124509 1732
rect 124630 1730 124690 1806
rect 125915 1732 125981 1733
rect 125915 1730 125916 1732
rect 124630 1670 125916 1730
rect 124443 1667 124509 1668
rect 125915 1668 125916 1670
rect 125980 1668 125981 1732
rect 125915 1667 125981 1668
rect 111566 1534 123034 1594
rect 111566 1189 111626 1534
rect 111747 1460 111813 1461
rect 111747 1396 111748 1460
rect 111812 1458 111813 1460
rect 120763 1460 120829 1461
rect 120763 1458 120764 1460
rect 111812 1398 111994 1458
rect 111812 1396 111813 1398
rect 111747 1395 111813 1396
rect 111379 1188 111445 1189
rect 111379 1124 111380 1188
rect 111444 1124 111445 1188
rect 111379 1123 111445 1124
rect 111563 1188 111629 1189
rect 111563 1124 111564 1188
rect 111628 1124 111629 1188
rect 111793 1188 111859 1189
rect 111793 1186 111794 1188
rect 111563 1123 111629 1124
rect 111750 1124 111794 1186
rect 111858 1124 111859 1188
rect 111750 1123 111859 1124
rect 111750 1050 111810 1123
rect 109174 990 111810 1050
rect 111934 1050 111994 1398
rect 112486 1398 120764 1458
rect 112486 1189 112546 1398
rect 120763 1396 120764 1398
rect 120828 1396 120829 1460
rect 120763 1395 120829 1396
rect 124262 1262 125610 1322
rect 112483 1188 112549 1189
rect 112483 1124 112484 1188
rect 112548 1124 112549 1188
rect 112483 1123 112549 1124
rect 120211 1188 120277 1189
rect 120211 1124 120212 1188
rect 120276 1186 120277 1188
rect 120276 1126 123770 1186
rect 120276 1124 120277 1126
rect 120211 1123 120277 1124
rect 123710 1053 123770 1126
rect 123707 1052 123773 1053
rect 111934 990 112546 1050
rect 104758 642 104818 990
rect 104758 582 104864 642
rect 103283 443 103349 444
rect 94267 236 94333 237
rect 93163 171 93229 172
rect 93899 172 93900 222
rect 93964 172 93965 222
rect 93899 171 93965 172
rect 94267 172 94268 236
rect 94332 172 94333 236
rect 94267 171 94333 172
rect 85438 38 87522 98
rect 89667 100 89733 101
rect 84331 35 84397 36
rect 89667 36 89668 100
rect 89732 98 89733 100
rect 92611 100 92677 101
rect 92611 98 92612 100
rect 89732 38 92612 98
rect 89732 36 89733 38
rect 89667 35 89733 36
rect 92611 36 92612 38
rect 92676 36 92677 100
rect 92982 98 93042 171
rect 101443 100 101509 101
rect 101443 98 101444 100
rect 92982 38 101444 98
rect 92611 35 92677 36
rect 101443 36 101444 38
rect 101508 36 101509 100
rect 103838 98 103898 222
rect 104804 98 104864 582
rect 106782 458 106842 990
rect 106963 780 107029 781
rect 106963 716 106964 780
rect 107028 778 107029 780
rect 107028 718 107210 778
rect 107028 716 107029 718
rect 106963 715 107029 716
rect 107150 370 107210 718
rect 107518 642 107578 990
rect 107699 780 107765 781
rect 107699 716 107700 780
rect 107764 778 107765 780
rect 111563 780 111629 781
rect 107764 718 108130 778
rect 107764 716 107765 718
rect 107699 715 107765 716
rect 107518 582 107946 642
rect 107150 310 107430 370
rect 107886 234 107946 582
rect 108070 370 108130 718
rect 111563 716 111564 780
rect 111628 778 111629 780
rect 111747 780 111813 781
rect 111747 778 111748 780
rect 111628 718 111748 778
rect 111628 716 111629 718
rect 111563 715 111629 716
rect 111747 716 111748 718
rect 111812 716 111813 780
rect 112486 778 112546 990
rect 117454 990 123586 1050
rect 117454 778 117514 990
rect 123526 914 123586 990
rect 123707 988 123708 1052
rect 123772 988 123773 1052
rect 124075 1052 124141 1053
rect 124075 1050 124076 1052
rect 123707 987 123773 988
rect 123894 990 124076 1050
rect 123894 914 123954 990
rect 124075 988 124076 990
rect 124140 988 124141 1052
rect 124075 987 124141 988
rect 124262 914 124322 1262
rect 125363 1188 125429 1189
rect 125363 1124 125364 1188
rect 125428 1124 125429 1188
rect 125363 1123 125429 1124
rect 123526 854 123954 914
rect 124078 854 124322 914
rect 125366 914 125426 1123
rect 125550 1050 125610 1262
rect 126102 1186 126162 1806
rect 126700 1458 126760 2350
rect 127942 1733 128002 2350
rect 134198 1866 134258 2350
rect 128494 1806 134074 1866
rect 134198 1806 135546 1866
rect 127939 1732 128005 1733
rect 127939 1668 127940 1732
rect 128004 1668 128005 1732
rect 127939 1667 128005 1668
rect 128494 1597 128554 1806
rect 128859 1732 128925 1733
rect 128859 1668 128860 1732
rect 128924 1730 128925 1732
rect 134014 1730 134074 1806
rect 135299 1732 135365 1733
rect 135299 1730 135300 1732
rect 128924 1670 133890 1730
rect 134014 1670 135300 1730
rect 128924 1668 128925 1670
rect 128859 1667 128925 1668
rect 128491 1596 128557 1597
rect 127206 1458 127266 1582
rect 128491 1532 128492 1596
rect 128556 1532 128557 1596
rect 128491 1531 128557 1532
rect 126700 1398 127082 1458
rect 127206 1398 131682 1458
rect 126835 1188 126901 1189
rect 126835 1186 126836 1188
rect 126102 1126 126836 1186
rect 126835 1124 126836 1126
rect 126900 1124 126901 1188
rect 126835 1123 126901 1124
rect 127022 1050 127082 1398
rect 131435 1324 131501 1325
rect 131435 1322 131436 1324
rect 125550 990 127082 1050
rect 127206 1262 131436 1322
rect 127206 914 127266 1262
rect 131435 1260 131436 1262
rect 131500 1260 131501 1324
rect 131435 1259 131501 1260
rect 128307 1188 128373 1189
rect 128307 1124 128308 1188
rect 128372 1124 128373 1188
rect 128307 1123 128373 1124
rect 125366 854 127266 914
rect 122971 780 123037 781
rect 122971 778 122972 780
rect 112486 718 117514 778
rect 122422 718 122972 778
rect 111747 715 111813 716
rect 111747 508 111813 509
rect 111747 444 111748 508
rect 111812 506 111813 508
rect 112299 508 112365 509
rect 112299 506 112300 508
rect 111812 446 112300 506
rect 111812 444 111813 446
rect 111747 443 111813 444
rect 112299 444 112300 446
rect 112364 444 112365 508
rect 112299 443 112365 444
rect 122422 370 122482 718
rect 122971 716 122972 718
rect 123036 716 123037 780
rect 124078 778 124138 854
rect 128310 778 128370 1123
rect 128675 1052 128741 1053
rect 128675 988 128676 1052
rect 128740 1050 128741 1052
rect 129963 1052 130029 1053
rect 129963 1050 129964 1052
rect 128740 990 129964 1050
rect 128740 988 128741 990
rect 128675 987 128741 988
rect 129963 988 129964 990
rect 130028 988 130029 1052
rect 131622 1050 131682 1398
rect 133830 1186 133890 1670
rect 135299 1668 135300 1670
rect 135364 1668 135365 1732
rect 135486 1730 135546 1806
rect 135667 1732 135733 1733
rect 135667 1730 135668 1732
rect 135486 1670 135668 1730
rect 135299 1667 135365 1668
rect 135667 1668 135668 1670
rect 135732 1668 135733 1732
rect 135667 1667 135733 1668
rect 135854 1594 135914 2942
rect 136590 2410 136650 2942
rect 145974 2410 146034 2942
rect 136038 2350 136650 2410
rect 139534 2350 145482 2410
rect 145974 2350 146770 2410
rect 136038 1733 136098 2350
rect 136222 1806 136650 1866
rect 136038 1732 136147 1733
rect 136038 1670 136082 1732
rect 136081 1668 136082 1670
rect 136146 1668 136147 1732
rect 136081 1667 136147 1668
rect 135118 1534 135914 1594
rect 135118 1461 135178 1534
rect 135115 1460 135181 1461
rect 135115 1396 135116 1460
rect 135180 1396 135181 1460
rect 136222 1458 136282 1806
rect 136403 1732 136469 1733
rect 136403 1668 136404 1732
rect 136468 1668 136469 1732
rect 136590 1730 136650 1806
rect 139347 1732 139413 1733
rect 139347 1730 139348 1732
rect 136590 1670 136834 1730
rect 136403 1667 136469 1668
rect 135115 1395 135181 1396
rect 135302 1398 136282 1458
rect 134379 1324 134445 1325
rect 134379 1260 134380 1324
rect 134444 1322 134445 1324
rect 135302 1322 135362 1398
rect 134444 1262 135362 1322
rect 134444 1260 134445 1262
rect 134379 1259 134445 1260
rect 136406 1186 136466 1667
rect 136587 1460 136653 1461
rect 136587 1396 136588 1460
rect 136652 1396 136653 1460
rect 136587 1395 136653 1396
rect 133830 1126 136466 1186
rect 135483 1052 135549 1053
rect 131622 990 135362 1050
rect 129963 987 130029 988
rect 129595 916 129661 917
rect 129595 852 129596 916
rect 129660 914 129661 916
rect 129963 916 130029 917
rect 129963 914 129964 916
rect 129660 854 129964 914
rect 129660 852 129661 854
rect 129595 851 129661 852
rect 129963 852 129964 854
rect 130028 852 130029 916
rect 129963 851 130029 852
rect 130334 854 135178 914
rect 130334 781 130394 854
rect 129227 780 129293 781
rect 129227 778 129228 780
rect 122971 715 123037 716
rect 123158 718 124138 778
rect 124308 718 124506 778
rect 128310 718 129228 778
rect 108070 310 113466 370
rect 113406 234 113466 310
rect 115246 310 122482 370
rect 115246 234 115306 310
rect 107886 174 113282 234
rect 113406 174 115306 234
rect 116715 236 116781 237
rect 103838 38 104864 98
rect 113222 98 113282 174
rect 116715 172 116716 236
rect 116780 234 116781 236
rect 123158 234 123218 718
rect 124075 644 124141 645
rect 124075 580 124076 644
rect 124140 642 124141 644
rect 124308 642 124368 718
rect 124140 582 124368 642
rect 124446 642 124506 718
rect 129227 716 129228 718
rect 129292 716 129293 780
rect 129227 715 129293 716
rect 130331 780 130397 781
rect 130331 716 130332 780
rect 130396 716 130397 780
rect 130331 715 130397 716
rect 130515 780 130581 781
rect 130515 716 130516 780
rect 130580 716 130581 780
rect 130515 715 130581 716
rect 134931 780 134997 781
rect 134931 716 134932 780
rect 134996 716 134997 780
rect 134931 715 134997 716
rect 130518 642 130578 715
rect 134934 642 134994 715
rect 135118 642 135178 854
rect 135302 781 135362 990
rect 135483 988 135484 1052
rect 135548 988 135549 1052
rect 135483 987 135549 988
rect 135486 914 135546 987
rect 135851 916 135917 917
rect 135851 914 135852 916
rect 135486 854 135852 914
rect 135851 852 135852 854
rect 135916 852 135917 916
rect 135851 851 135917 852
rect 135299 780 135365 781
rect 135299 716 135300 780
rect 135364 716 135365 780
rect 136219 780 136285 781
rect 136219 778 136220 780
rect 135299 715 135365 716
rect 135670 718 136220 778
rect 135483 644 135549 645
rect 135483 642 135484 644
rect 124446 582 130578 642
rect 130702 582 134442 642
rect 134934 582 135040 642
rect 135118 582 135484 642
rect 124140 580 124141 582
rect 124075 579 124141 580
rect 116780 174 123218 234
rect 130702 370 130762 582
rect 123674 310 130762 370
rect 134382 370 134442 582
rect 134980 506 135040 582
rect 135483 580 135484 582
rect 135548 580 135549 644
rect 135483 579 135549 580
rect 135670 506 135730 718
rect 136219 716 136220 718
rect 136284 716 136285 780
rect 136219 715 136285 716
rect 136590 642 136650 1395
rect 136774 1186 136834 1670
rect 138614 1670 139348 1730
rect 138614 1461 138674 1670
rect 139347 1668 139348 1670
rect 139412 1668 139413 1732
rect 139347 1667 139413 1668
rect 138611 1460 138677 1461
rect 138611 1396 138612 1460
rect 138676 1396 138677 1460
rect 138611 1395 138677 1396
rect 138795 1460 138861 1461
rect 138795 1396 138796 1460
rect 138860 1396 138861 1460
rect 138795 1395 138861 1396
rect 136955 1324 137021 1325
rect 136955 1260 136956 1324
rect 137020 1322 137021 1324
rect 138798 1322 138858 1395
rect 139534 1322 139594 2350
rect 145422 1866 145482 2350
rect 141926 1806 145298 1866
rect 145422 1806 146034 1866
rect 141003 1732 141069 1733
rect 141003 1668 141004 1732
rect 141068 1730 141069 1732
rect 141739 1732 141805 1733
rect 141739 1730 141740 1732
rect 141068 1670 141740 1730
rect 141068 1668 141069 1670
rect 141003 1667 141069 1668
rect 141739 1668 141740 1670
rect 141804 1668 141805 1732
rect 141739 1667 141805 1668
rect 141926 1594 141986 1806
rect 145238 1730 145298 1806
rect 145787 1732 145853 1733
rect 145787 1730 145788 1732
rect 137020 1262 138858 1322
rect 139350 1262 139594 1322
rect 141006 1534 141986 1594
rect 142478 1670 145114 1730
rect 145238 1670 145788 1730
rect 137020 1260 137021 1262
rect 136955 1259 137021 1260
rect 139350 1186 139410 1262
rect 139577 1188 139643 1189
rect 139577 1186 139578 1188
rect 136774 1126 139410 1186
rect 139534 1124 139578 1186
rect 139642 1124 139643 1188
rect 139899 1188 139965 1189
rect 139899 1186 139900 1188
rect 139534 1123 139643 1124
rect 139718 1126 139900 1186
rect 139534 1050 139594 1123
rect 137878 990 139594 1050
rect 137691 780 137757 781
rect 137691 716 137692 780
rect 137756 778 137757 780
rect 137878 778 137938 990
rect 139718 914 139778 1126
rect 139899 1124 139900 1126
rect 139964 1124 139965 1188
rect 139899 1123 139965 1124
rect 137756 718 137938 778
rect 138062 854 139778 914
rect 137756 716 137757 718
rect 137691 715 137757 716
rect 138062 642 138122 854
rect 141006 778 141066 1534
rect 142478 1458 142538 1670
rect 144867 1596 144933 1597
rect 144867 1532 144868 1596
rect 144932 1532 144933 1596
rect 145054 1594 145114 1670
rect 145787 1668 145788 1670
rect 145852 1668 145853 1732
rect 145974 1730 146034 1806
rect 146155 1732 146221 1733
rect 146155 1730 146156 1732
rect 145974 1670 146156 1730
rect 145787 1667 145853 1668
rect 146155 1668 146156 1670
rect 146220 1668 146221 1732
rect 146155 1667 146221 1668
rect 146339 1732 146405 1733
rect 146339 1668 146340 1732
rect 146404 1668 146405 1732
rect 146339 1667 146405 1668
rect 145971 1596 146037 1597
rect 145971 1594 145972 1596
rect 145054 1534 145972 1594
rect 144867 1531 144933 1532
rect 145971 1532 145972 1534
rect 146036 1532 146037 1596
rect 145971 1531 146037 1532
rect 141190 1398 142538 1458
rect 144870 1458 144930 1531
rect 146342 1458 146402 1667
rect 144870 1398 146402 1458
rect 141190 1325 141250 1398
rect 141187 1324 141253 1325
rect 141187 1260 141188 1324
rect 141252 1260 141253 1324
rect 141187 1259 141253 1260
rect 141187 1188 141253 1189
rect 141187 1124 141188 1188
rect 141252 1124 141253 1188
rect 146710 1186 146770 2350
rect 153702 1866 153762 2942
rect 147078 1806 152658 1866
rect 153702 1806 154028 1866
rect 147078 1322 147138 1806
rect 148179 1732 148245 1733
rect 148179 1730 148180 1732
rect 147262 1670 148180 1730
rect 147262 1597 147322 1670
rect 148179 1668 148180 1670
rect 148244 1668 148245 1732
rect 148179 1667 148245 1668
rect 152227 1732 152293 1733
rect 152227 1668 152228 1732
rect 152292 1730 152293 1732
rect 152292 1670 152474 1730
rect 152292 1668 152293 1670
rect 152227 1667 152293 1668
rect 147259 1596 147325 1597
rect 147259 1532 147260 1596
rect 147324 1532 147325 1596
rect 147259 1531 147325 1532
rect 147811 1596 147877 1597
rect 147811 1532 147812 1596
rect 147876 1594 147877 1596
rect 147876 1534 148242 1594
rect 147876 1532 147877 1534
rect 147811 1531 147877 1532
rect 148182 1325 148242 1534
rect 148366 1534 152290 1594
rect 147995 1324 148061 1325
rect 147078 1262 147506 1322
rect 147446 1189 147506 1262
rect 147995 1260 147996 1324
rect 148060 1260 148061 1324
rect 147995 1259 148061 1260
rect 148179 1324 148245 1325
rect 148179 1260 148180 1324
rect 148244 1260 148245 1324
rect 148179 1259 148245 1260
rect 147443 1188 147509 1189
rect 141187 1123 141253 1124
rect 136590 582 138122 642
rect 139350 718 141066 778
rect 141190 778 141250 1123
rect 146710 1126 147322 1186
rect 144315 780 144381 781
rect 144315 778 144316 780
rect 141190 718 144316 778
rect 134382 310 134662 370
rect 134980 446 135730 506
rect 139350 370 139410 718
rect 144315 716 144316 718
rect 144380 716 144381 780
rect 144315 715 144381 716
rect 145603 780 145669 781
rect 145603 716 145604 780
rect 145668 716 145669 780
rect 146342 778 146402 902
rect 147075 780 147141 781
rect 147075 778 147076 780
rect 146342 718 147076 778
rect 145603 715 145669 716
rect 147075 716 147076 718
rect 147140 716 147141 780
rect 147262 778 147322 1126
rect 147443 1124 147444 1188
rect 147508 1124 147509 1188
rect 147998 1138 148058 1259
rect 147443 1123 147509 1124
rect 148366 778 148426 1534
rect 149102 1398 152106 1458
rect 147262 718 148426 778
rect 148550 1262 148978 1322
rect 147075 715 147141 716
rect 139899 644 139965 645
rect 139899 580 139900 644
rect 139964 580 139965 644
rect 145606 642 145666 715
rect 148550 642 148610 1262
rect 148731 1188 148797 1189
rect 148731 1124 148732 1188
rect 148796 1124 148797 1188
rect 148731 1123 148797 1124
rect 145606 582 148610 642
rect 139899 579 139965 580
rect 139902 506 139962 579
rect 148734 506 148794 1123
rect 148918 642 148978 1262
rect 149102 642 149162 1398
rect 150758 1262 151922 1322
rect 150758 1189 150818 1262
rect 150755 1188 150821 1189
rect 150755 1124 150756 1188
rect 150820 1124 150821 1188
rect 150755 1123 150821 1124
rect 151307 1188 151373 1189
rect 151307 1124 151308 1188
rect 151372 1124 151373 1188
rect 151307 1123 151373 1124
rect 151310 1050 151370 1123
rect 150758 990 151186 1050
rect 151310 990 151452 1050
rect 150758 917 150818 990
rect 150755 916 150821 917
rect 150390 778 150450 902
rect 150755 852 150756 916
rect 150820 852 150821 916
rect 150755 851 150821 852
rect 150939 916 151005 917
rect 150939 852 150940 916
rect 151004 852 151005 916
rect 151126 914 151186 990
rect 151307 916 151373 917
rect 151307 914 151308 916
rect 151126 854 151308 914
rect 150939 851 151005 852
rect 151307 852 151308 854
rect 151372 852 151373 916
rect 151307 851 151373 852
rect 150942 778 151002 851
rect 150390 718 151002 778
rect 148918 582 149162 642
rect 151307 644 151373 645
rect 151307 580 151308 644
rect 151372 642 151373 644
rect 151372 582 151554 642
rect 151372 580 151373 582
rect 151307 579 151373 580
rect 139902 446 148794 506
rect 150755 508 150821 509
rect 150755 458 150756 508
rect 150820 458 150821 508
rect 151494 458 151554 582
rect 135118 310 139410 370
rect 116780 172 116781 174
rect 116715 171 116781 172
rect 116899 100 116965 101
rect 116899 98 116900 100
rect 113222 38 116900 98
rect 101443 35 101509 36
rect 116899 36 116900 38
rect 116964 36 116965 100
rect 116899 35 116965 36
rect 119475 100 119541 101
rect 119475 36 119476 100
rect 119540 98 119541 100
rect 135118 98 135178 310
rect 151862 370 151922 1262
rect 152046 914 152106 1398
rect 152230 1186 152290 1534
rect 152414 1458 152474 1670
rect 152598 1594 152658 1806
rect 154438 1733 154498 2942
rect 154435 1732 154501 1733
rect 154435 1668 154436 1732
rect 154500 1668 154501 1732
rect 155358 1730 155418 2942
rect 156094 1733 156154 2942
rect 154435 1667 154501 1668
rect 154806 1670 155418 1730
rect 156091 1732 156157 1733
rect 154806 1594 154866 1670
rect 156091 1668 156092 1732
rect 156156 1668 156157 1732
rect 156091 1667 156157 1668
rect 157931 1596 157997 1597
rect 157931 1594 157932 1596
rect 152598 1534 154866 1594
rect 155174 1534 157932 1594
rect 155174 1458 155234 1534
rect 157931 1532 157932 1534
rect 157996 1532 157997 1596
rect 157931 1531 157997 1532
rect 152414 1398 155234 1458
rect 157563 1460 157629 1461
rect 157563 1396 157564 1460
rect 157628 1458 157629 1460
rect 157931 1460 157997 1461
rect 157931 1458 157932 1460
rect 157628 1398 157932 1458
rect 157628 1396 157629 1398
rect 157563 1395 157629 1396
rect 157931 1396 157932 1398
rect 157996 1396 157997 1460
rect 157931 1395 157997 1396
rect 153883 1324 153949 1325
rect 153883 1260 153884 1324
rect 153948 1322 153949 1324
rect 158118 1322 158178 2942
rect 158670 2350 170322 2410
rect 158483 1732 158549 1733
rect 158483 1668 158484 1732
rect 158548 1668 158549 1732
rect 158483 1667 158549 1668
rect 153948 1262 158178 1322
rect 153948 1260 153949 1262
rect 153883 1259 153949 1260
rect 158486 1186 158546 1667
rect 152230 1126 158546 1186
rect 158670 1050 158730 2350
rect 170262 1866 170322 2350
rect 169342 1806 170138 1866
rect 170262 1806 171426 1866
rect 166947 1732 167013 1733
rect 166947 1730 166948 1732
rect 159186 1718 160018 1730
rect 159038 1670 160018 1718
rect 159403 1460 159469 1461
rect 159403 1396 159404 1460
rect 159468 1396 159469 1460
rect 159403 1395 159469 1396
rect 159771 1460 159837 1461
rect 159771 1396 159772 1460
rect 159836 1396 159837 1460
rect 159958 1458 160018 1670
rect 160142 1670 166948 1730
rect 160142 1597 160202 1670
rect 166947 1668 166948 1670
rect 167012 1668 167013 1732
rect 166947 1667 167013 1668
rect 168971 1732 169037 1733
rect 168971 1668 168972 1732
rect 169036 1668 169037 1732
rect 168971 1667 169037 1668
rect 160139 1596 160205 1597
rect 160139 1532 160140 1596
rect 160204 1532 160205 1596
rect 160139 1531 160205 1532
rect 161059 1596 161125 1597
rect 161059 1532 161060 1596
rect 161124 1594 161125 1596
rect 161124 1534 166642 1594
rect 161124 1532 161125 1534
rect 161059 1531 161125 1532
rect 161243 1460 161309 1461
rect 159958 1398 160202 1458
rect 159771 1395 159837 1396
rect 159406 1138 159466 1395
rect 152598 990 158730 1050
rect 152598 914 152658 990
rect 152046 854 152658 914
rect 159774 778 159834 1395
rect 160142 1138 160202 1398
rect 161243 1396 161244 1460
rect 161308 1396 161309 1460
rect 161611 1460 161677 1461
rect 161611 1410 161612 1460
rect 161676 1410 161677 1460
rect 164003 1460 164069 1461
rect 161243 1395 161309 1396
rect 161246 1050 161306 1395
rect 164003 1396 164004 1460
rect 164068 1458 164069 1460
rect 164068 1398 166458 1458
rect 164068 1396 164069 1398
rect 164003 1395 164069 1396
rect 161979 1324 162045 1325
rect 161979 1260 161980 1324
rect 162044 1260 162045 1324
rect 161979 1259 162045 1260
rect 163451 1324 163517 1325
rect 163451 1260 163452 1324
rect 163516 1260 163517 1324
rect 163451 1259 163517 1260
rect 161982 1050 162042 1259
rect 163454 1186 163514 1259
rect 166211 1188 166277 1189
rect 161246 990 162042 1050
rect 161614 902 162262 914
rect 163454 1126 164618 1186
rect 163819 1052 163885 1053
rect 163819 988 163820 1052
rect 163884 988 163885 1052
rect 163819 987 163885 988
rect 161614 854 162410 902
rect 161614 781 161674 854
rect 156278 718 159834 778
rect 161611 780 161677 781
rect 156278 645 156338 718
rect 161611 716 161612 780
rect 161676 716 161677 780
rect 163267 780 163333 781
rect 163267 778 163268 780
rect 161611 715 161677 716
rect 161798 718 163268 778
rect 156275 644 156341 645
rect 156275 580 156276 644
rect 156340 580 156341 644
rect 156275 579 156341 580
rect 157931 644 157997 645
rect 157931 580 157932 644
rect 157996 642 157997 644
rect 161798 642 161858 718
rect 163267 716 163268 718
rect 163332 716 163333 780
rect 163267 715 163333 716
rect 163635 644 163701 645
rect 163635 642 163636 644
rect 157996 582 161858 642
rect 161982 582 163636 642
rect 157996 580 157997 582
rect 157931 579 157997 580
rect 157931 372 157997 373
rect 157931 370 157932 372
rect 151862 310 157932 370
rect 157931 308 157932 310
rect 157996 308 157997 372
rect 157931 307 157997 308
rect 161243 372 161309 373
rect 161243 308 161244 372
rect 161308 370 161309 372
rect 161982 370 162042 582
rect 163635 580 163636 582
rect 163700 580 163701 644
rect 163635 579 163701 580
rect 163822 458 163882 987
rect 164558 458 164618 1126
rect 166211 1124 166212 1188
rect 166276 1124 166277 1188
rect 166211 1123 166277 1124
rect 166214 914 166274 1123
rect 166398 1050 166458 1398
rect 166582 1186 166642 1534
rect 168787 1188 168853 1189
rect 168787 1186 168788 1188
rect 166582 1126 168788 1186
rect 168787 1124 168788 1126
rect 168852 1124 168853 1188
rect 168974 1186 169034 1667
rect 169342 1597 169402 1806
rect 169891 1732 169957 1733
rect 169891 1668 169892 1732
rect 169956 1668 169957 1732
rect 169891 1667 169957 1668
rect 169339 1596 169405 1597
rect 169339 1532 169340 1596
rect 169404 1532 169405 1596
rect 169339 1531 169405 1532
rect 169894 1325 169954 1667
rect 170078 1594 170138 1806
rect 171179 1596 171245 1597
rect 171179 1594 171180 1596
rect 170078 1534 171180 1594
rect 171179 1532 171180 1534
rect 171244 1532 171245 1596
rect 171366 1594 171426 1806
rect 175782 1806 176210 1866
rect 175782 1733 175842 1806
rect 175779 1732 175845 1733
rect 171918 1670 173266 1730
rect 171731 1596 171797 1597
rect 171731 1594 171732 1596
rect 171366 1534 171732 1594
rect 171179 1531 171245 1532
rect 171731 1532 171732 1534
rect 171796 1532 171797 1596
rect 171731 1531 171797 1532
rect 169891 1324 169957 1325
rect 169891 1260 169892 1324
rect 169956 1260 169957 1324
rect 169891 1259 169957 1260
rect 170075 1324 170141 1325
rect 170075 1260 170076 1324
rect 170140 1260 170141 1324
rect 171918 1322 171978 1670
rect 173019 1596 173085 1597
rect 173019 1532 173020 1596
rect 173084 1532 173085 1596
rect 173206 1594 173266 1670
rect 175779 1668 175780 1732
rect 175844 1668 175845 1732
rect 175779 1667 175845 1668
rect 175963 1732 176029 1733
rect 175963 1668 175964 1732
rect 176028 1668 176029 1732
rect 176150 1730 176210 1806
rect 185166 1806 187802 1866
rect 178171 1732 178237 1733
rect 176150 1670 177314 1730
rect 175963 1667 176029 1668
rect 173206 1534 175658 1594
rect 173019 1531 173085 1532
rect 170075 1259 170141 1260
rect 170262 1262 171978 1322
rect 173022 1322 173082 1531
rect 173939 1324 174005 1325
rect 173939 1322 173940 1324
rect 173022 1262 173940 1322
rect 170078 1186 170138 1259
rect 168974 1126 170138 1186
rect 168787 1123 168853 1124
rect 170262 1050 170322 1262
rect 173939 1260 173940 1262
rect 174004 1260 174005 1324
rect 173939 1259 174005 1260
rect 173387 1188 173453 1189
rect 173387 1186 173388 1188
rect 171182 1126 173388 1186
rect 171182 1050 171242 1126
rect 173387 1124 173388 1126
rect 173452 1124 173453 1188
rect 173387 1123 173453 1124
rect 175598 1050 175658 1534
rect 175966 1325 176026 1667
rect 176518 1534 177130 1594
rect 176518 1458 176578 1534
rect 177070 1461 177130 1534
rect 176150 1398 176578 1458
rect 176883 1460 176949 1461
rect 175963 1324 176029 1325
rect 175963 1260 175964 1324
rect 176028 1260 176029 1324
rect 175963 1259 176029 1260
rect 176150 1189 176210 1398
rect 176883 1396 176884 1460
rect 176948 1396 176949 1460
rect 176883 1395 176949 1396
rect 177067 1460 177133 1461
rect 177067 1396 177068 1460
rect 177132 1396 177133 1460
rect 177254 1458 177314 1670
rect 178171 1668 178172 1732
rect 178236 1730 178237 1732
rect 178907 1732 178973 1733
rect 178236 1670 178418 1730
rect 178236 1668 178237 1670
rect 178171 1667 178237 1668
rect 178358 1597 178418 1670
rect 178907 1668 178908 1732
rect 178972 1730 178973 1732
rect 184979 1732 185045 1733
rect 184979 1730 184980 1732
rect 178972 1670 184980 1730
rect 178972 1668 178973 1670
rect 178907 1667 178973 1668
rect 184979 1668 184980 1670
rect 185044 1668 185045 1732
rect 184979 1667 185045 1668
rect 178171 1596 178237 1597
rect 178171 1532 178172 1596
rect 178236 1532 178237 1596
rect 178171 1531 178237 1532
rect 178355 1596 178421 1597
rect 178355 1532 178356 1596
rect 178420 1532 178421 1596
rect 178355 1531 178421 1532
rect 179643 1596 179709 1597
rect 179643 1532 179644 1596
rect 179708 1594 179709 1596
rect 181851 1596 181917 1597
rect 181851 1594 181852 1596
rect 179708 1534 181852 1594
rect 179708 1532 179709 1534
rect 179643 1531 179709 1532
rect 181851 1532 181852 1534
rect 181916 1532 181917 1596
rect 184059 1596 184125 1597
rect 184059 1594 184060 1596
rect 181851 1531 181917 1532
rect 182038 1534 184060 1594
rect 177987 1460 178053 1461
rect 177987 1458 177988 1460
rect 177254 1398 177988 1458
rect 177067 1395 177133 1396
rect 177987 1396 177988 1398
rect 178052 1396 178053 1460
rect 178174 1458 178234 1531
rect 182038 1458 182098 1534
rect 184059 1532 184060 1534
rect 184124 1532 184125 1596
rect 184059 1531 184125 1532
rect 185166 1458 185226 1806
rect 187742 1730 187802 1806
rect 192339 1732 192405 1733
rect 192339 1730 192340 1732
rect 187742 1670 192340 1730
rect 192339 1668 192340 1670
rect 192404 1668 192405 1732
rect 192339 1667 192405 1668
rect 190499 1596 190565 1597
rect 190499 1532 190500 1596
rect 190564 1532 190565 1596
rect 190499 1531 190565 1532
rect 178174 1398 182098 1458
rect 183694 1398 185226 1458
rect 190502 1458 190562 1531
rect 191051 1460 191117 1461
rect 191051 1458 191052 1460
rect 190502 1398 191052 1458
rect 177987 1395 178053 1396
rect 176331 1324 176397 1325
rect 176331 1260 176332 1324
rect 176396 1260 176397 1324
rect 176331 1259 176397 1260
rect 176147 1188 176213 1189
rect 176147 1124 176148 1188
rect 176212 1124 176213 1188
rect 176147 1123 176213 1124
rect 176334 1050 176394 1259
rect 176886 1186 176946 1395
rect 183694 1325 183754 1398
rect 191051 1396 191052 1398
rect 191116 1396 191117 1460
rect 191051 1395 191117 1396
rect 179459 1324 179525 1325
rect 179459 1260 179460 1324
rect 179524 1322 179525 1324
rect 180379 1324 180445 1325
rect 180379 1322 180380 1324
rect 179524 1262 180380 1322
rect 179524 1260 179525 1262
rect 179459 1259 179525 1260
rect 180379 1260 180380 1262
rect 180444 1260 180445 1324
rect 180379 1259 180445 1260
rect 183691 1324 183757 1325
rect 183691 1260 183692 1324
rect 183756 1260 183757 1324
rect 189763 1324 189829 1325
rect 189763 1322 189764 1324
rect 183691 1259 183757 1260
rect 183878 1262 189764 1322
rect 180931 1188 180997 1189
rect 180931 1186 180932 1188
rect 176886 1126 180932 1186
rect 180931 1124 180932 1126
rect 180996 1124 180997 1188
rect 183878 1186 183938 1262
rect 189763 1260 189764 1262
rect 189828 1260 189829 1324
rect 191235 1324 191301 1325
rect 191235 1322 191236 1324
rect 189763 1259 189829 1260
rect 189950 1262 191236 1322
rect 189950 1186 190010 1262
rect 191235 1260 191236 1262
rect 191300 1260 191301 1324
rect 194182 1322 194242 2942
rect 194918 1733 194978 2262
rect 194731 1732 194797 1733
rect 194731 1668 194732 1732
rect 194796 1668 194797 1732
rect 194731 1667 194797 1668
rect 194915 1732 194981 1733
rect 194915 1668 194916 1732
rect 194980 1668 194981 1732
rect 195654 1730 195714 2942
rect 194915 1667 194981 1668
rect 195102 1670 195714 1730
rect 197126 1670 200682 1730
rect 194734 1594 194794 1667
rect 195102 1594 195162 1670
rect 197126 1597 197186 1670
rect 194734 1534 195162 1594
rect 195835 1596 195901 1597
rect 195835 1532 195836 1596
rect 195900 1532 195901 1596
rect 195835 1531 195901 1532
rect 197123 1596 197189 1597
rect 197123 1532 197124 1596
rect 197188 1532 197189 1596
rect 197123 1531 197189 1532
rect 198411 1596 198477 1597
rect 198411 1532 198412 1596
rect 198476 1594 198477 1596
rect 198476 1534 200498 1594
rect 198476 1532 198477 1534
rect 198411 1531 198477 1532
rect 195838 1458 195898 1531
rect 200438 1461 200498 1534
rect 197491 1460 197557 1461
rect 197491 1458 197492 1460
rect 195838 1398 197492 1458
rect 197491 1396 197492 1398
rect 197556 1396 197557 1460
rect 197491 1395 197557 1396
rect 198779 1460 198845 1461
rect 198779 1396 198780 1460
rect 198844 1396 198845 1460
rect 198779 1395 198845 1396
rect 200435 1460 200501 1461
rect 200435 1396 200436 1460
rect 200500 1396 200501 1460
rect 200622 1458 200682 1670
rect 200990 1597 201050 2942
rect 224174 2410 224234 2942
rect 225094 2410 225154 2942
rect 211294 2350 215402 2410
rect 224174 2350 224602 2410
rect 225094 2350 225706 2410
rect 207979 1732 208045 1733
rect 204670 1670 205098 1730
rect 204670 1597 204730 1670
rect 200987 1596 201053 1597
rect 200987 1532 200988 1596
rect 201052 1532 201053 1596
rect 200987 1531 201053 1532
rect 203195 1596 203261 1597
rect 203195 1532 203196 1596
rect 203260 1532 203261 1596
rect 203195 1531 203261 1532
rect 204299 1596 204365 1597
rect 204299 1532 204300 1596
rect 204364 1532 204365 1596
rect 204299 1531 204365 1532
rect 204667 1596 204733 1597
rect 204667 1532 204668 1596
rect 204732 1532 204733 1596
rect 204667 1531 204733 1532
rect 204851 1596 204917 1597
rect 204851 1532 204852 1596
rect 204916 1532 204917 1596
rect 204851 1531 204917 1532
rect 203198 1458 203258 1531
rect 200622 1398 203258 1458
rect 204302 1458 204362 1531
rect 204854 1458 204914 1531
rect 204302 1398 204914 1458
rect 205038 1458 205098 1670
rect 207979 1668 207980 1732
rect 208044 1668 208045 1732
rect 211294 1730 211354 2350
rect 215342 1866 215402 2350
rect 215342 1806 216138 1866
rect 216078 1730 216138 1806
rect 220310 1806 223902 1866
rect 220310 1733 220370 1806
rect 216811 1732 216877 1733
rect 216811 1730 216812 1732
rect 207979 1667 208045 1668
rect 210926 1670 211354 1730
rect 211478 1670 215954 1730
rect 216078 1670 216812 1730
rect 207982 1594 208042 1667
rect 210187 1596 210253 1597
rect 210187 1594 210188 1596
rect 207982 1534 210188 1594
rect 210187 1532 210188 1534
rect 210252 1532 210253 1596
rect 210187 1531 210253 1532
rect 210926 1461 210986 1670
rect 208347 1460 208413 1461
rect 208347 1458 208348 1460
rect 205038 1398 208348 1458
rect 200435 1395 200501 1396
rect 208347 1396 208348 1398
rect 208412 1396 208413 1460
rect 208347 1395 208413 1396
rect 209819 1460 209885 1461
rect 209819 1396 209820 1460
rect 209884 1458 209885 1460
rect 210923 1460 210989 1461
rect 209884 1398 210066 1458
rect 209884 1396 209885 1398
rect 209819 1395 209885 1396
rect 198782 1322 198842 1395
rect 210006 1325 210066 1398
rect 210923 1396 210924 1460
rect 210988 1396 210989 1460
rect 210923 1395 210989 1396
rect 210003 1324 210069 1325
rect 194182 1262 197738 1322
rect 198782 1262 209514 1322
rect 191235 1259 191301 1260
rect 180931 1123 180997 1124
rect 181118 1126 183938 1186
rect 184614 1126 190010 1186
rect 191051 1188 191117 1189
rect 181118 1050 181178 1126
rect 166398 990 170322 1050
rect 170446 990 171242 1050
rect 175046 990 175474 1050
rect 175598 990 176394 1050
rect 176518 990 181178 1050
rect 184427 1052 184493 1053
rect 170446 914 170506 990
rect 166214 854 170506 914
rect 169158 718 170322 778
rect 169158 458 169218 718
rect 169891 644 169957 645
rect 169891 580 169892 644
rect 169956 580 169957 644
rect 169891 579 169957 580
rect 169894 458 169954 579
rect 161308 310 162042 370
rect 161308 308 161309 310
rect 161243 307 161309 308
rect 170262 370 170322 718
rect 175046 645 175106 990
rect 175414 914 175474 990
rect 176518 914 176578 990
rect 184427 988 184428 1052
rect 184492 988 184493 1052
rect 184427 987 184493 988
rect 184430 914 184490 987
rect 175414 854 176578 914
rect 177806 854 184490 914
rect 175043 644 175109 645
rect 175043 580 175044 644
rect 175108 580 175109 644
rect 175043 579 175109 580
rect 177806 645 177866 854
rect 184614 778 184674 1126
rect 191051 1124 191052 1188
rect 191116 1124 191117 1188
rect 191051 1123 191117 1124
rect 191419 1188 191485 1189
rect 191419 1124 191420 1188
rect 191484 1186 191485 1188
rect 196939 1188 197005 1189
rect 196939 1186 196940 1188
rect 191484 1126 196940 1186
rect 191484 1124 191485 1126
rect 191419 1123 191485 1124
rect 196939 1124 196940 1126
rect 197004 1124 197005 1188
rect 196939 1123 197005 1124
rect 189763 1052 189829 1053
rect 189763 988 189764 1052
rect 189828 1050 189829 1052
rect 191054 1050 191114 1123
rect 197307 1052 197373 1053
rect 197307 1050 197308 1052
rect 189828 990 190562 1050
rect 191054 990 197308 1050
rect 189828 988 189829 990
rect 189763 987 189829 988
rect 177990 718 184674 778
rect 190315 780 190381 781
rect 177251 644 177317 645
rect 177251 580 177252 644
rect 177316 580 177317 644
rect 177251 579 177317 580
rect 177803 644 177869 645
rect 177803 580 177804 644
rect 177868 580 177869 644
rect 177803 579 177869 580
rect 170262 310 176246 370
rect 177254 370 177314 579
rect 177990 370 178050 718
rect 190315 716 190316 780
rect 190380 716 190381 780
rect 190315 715 190381 716
rect 190318 506 190378 715
rect 190502 642 190562 990
rect 197307 988 197308 990
rect 197372 988 197373 1052
rect 197307 987 197373 988
rect 197678 914 197738 1262
rect 209267 1188 209333 1189
rect 209267 1186 209268 1188
rect 198552 1126 206018 1186
rect 198552 1050 198612 1126
rect 198230 990 198612 1050
rect 197859 916 197925 917
rect 197859 914 197860 916
rect 197678 854 197860 914
rect 197859 852 197860 854
rect 197924 852 197925 916
rect 198230 914 198290 990
rect 197859 851 197925 852
rect 198092 854 198290 914
rect 198414 854 204868 914
rect 198092 778 198152 854
rect 198414 781 198474 854
rect 196758 718 198152 778
rect 198411 780 198477 781
rect 190502 582 191482 642
rect 191422 509 191482 582
rect 190867 508 190933 509
rect 190867 506 190868 508
rect 190318 446 190868 506
rect 190867 444 190868 446
rect 190932 444 190933 508
rect 190867 443 190933 444
rect 191419 508 191485 509
rect 191419 444 191420 508
rect 191484 444 191485 508
rect 196758 458 196818 718
rect 198411 716 198412 780
rect 198476 716 198477 780
rect 198411 715 198477 716
rect 204115 644 204181 645
rect 197126 582 198428 642
rect 197126 509 197186 582
rect 197123 508 197189 509
rect 191419 443 191485 444
rect 177254 310 178050 370
rect 197123 444 197124 508
rect 197188 444 197189 508
rect 197859 508 197925 509
rect 197859 458 197860 508
rect 197924 458 197925 508
rect 198227 508 198293 509
rect 197123 443 197189 444
rect 198227 444 198228 508
rect 198292 444 198293 508
rect 198368 506 198428 582
rect 204115 580 204116 644
rect 204180 642 204181 644
rect 204667 644 204733 645
rect 204667 642 204668 644
rect 204180 582 204668 642
rect 204180 580 204181 582
rect 204115 579 204181 580
rect 204667 580 204668 582
rect 204732 580 204733 644
rect 204808 642 204868 854
rect 205958 778 206018 1126
rect 208718 1126 209268 1186
rect 208718 778 208778 1126
rect 209267 1124 209268 1126
rect 209332 1124 209333 1188
rect 209267 1123 209333 1124
rect 205958 718 208778 778
rect 205219 644 205285 645
rect 205219 642 205220 644
rect 204808 582 205220 642
rect 204667 579 204733 580
rect 205219 580 205220 582
rect 205284 580 205285 644
rect 205219 579 205285 580
rect 207979 644 208045 645
rect 207979 580 207980 644
rect 208044 580 208045 644
rect 207979 579 208045 580
rect 207982 506 208042 579
rect 198368 446 208042 506
rect 209454 506 209514 1262
rect 210003 1260 210004 1324
rect 210068 1260 210069 1324
rect 211478 1322 211538 1670
rect 215894 1594 215954 1670
rect 216811 1668 216812 1670
rect 216876 1668 216877 1732
rect 220307 1732 220373 1733
rect 216811 1667 216877 1668
rect 216998 1670 218714 1730
rect 216998 1594 217058 1670
rect 215894 1534 217058 1594
rect 218102 1534 218530 1594
rect 212027 1460 212093 1461
rect 212027 1396 212028 1460
rect 212092 1396 212093 1460
rect 218102 1458 218162 1534
rect 212027 1395 212093 1396
rect 217366 1398 218162 1458
rect 218283 1460 218349 1461
rect 210003 1259 210069 1260
rect 210374 1262 211538 1322
rect 210374 645 210434 1262
rect 212030 1189 212090 1395
rect 214787 1324 214853 1325
rect 214787 1322 214788 1324
rect 213870 1262 214788 1322
rect 212027 1188 212093 1189
rect 210742 1126 211722 1186
rect 210371 644 210437 645
rect 210371 580 210372 644
rect 210436 580 210437 644
rect 210371 579 210437 580
rect 210555 644 210621 645
rect 210555 580 210556 644
rect 210620 580 210621 644
rect 210555 579 210621 580
rect 210558 506 210618 579
rect 209454 446 210618 506
rect 198227 443 198293 444
rect 198230 370 198290 443
rect 210742 370 210802 1126
rect 211291 644 211357 645
rect 211291 580 211292 644
rect 211356 580 211357 644
rect 211291 579 211357 580
rect 211294 506 211354 579
rect 211662 506 211722 1126
rect 212027 1124 212028 1188
rect 212092 1124 212093 1188
rect 212027 1123 212093 1124
rect 213870 506 213930 1262
rect 214787 1260 214788 1262
rect 214852 1260 214853 1324
rect 214787 1259 214853 1260
rect 217366 506 217426 1398
rect 218283 1396 218284 1460
rect 218348 1396 218349 1460
rect 218283 1395 218349 1396
rect 217547 1324 217613 1325
rect 217547 1260 217548 1324
rect 217612 1260 217613 1324
rect 218286 1322 218346 1395
rect 217547 1259 217613 1260
rect 217734 1262 218346 1322
rect 217550 1050 217610 1259
rect 217734 1189 217794 1262
rect 217731 1188 217797 1189
rect 217731 1124 217732 1188
rect 217796 1124 217797 1188
rect 217731 1123 217797 1124
rect 217550 990 217794 1050
rect 217734 642 217794 990
rect 218470 778 218530 1534
rect 218654 1050 218714 1670
rect 220307 1668 220308 1732
rect 220372 1668 220373 1732
rect 224542 1866 224602 2350
rect 224542 1806 225154 1866
rect 220307 1667 220373 1668
rect 224907 1596 224973 1597
rect 224907 1594 224908 1596
rect 220862 1534 224908 1594
rect 220862 1050 220922 1534
rect 224907 1532 224908 1534
rect 224972 1532 224973 1596
rect 224907 1531 224973 1532
rect 224539 1460 224605 1461
rect 224539 1396 224540 1460
rect 224604 1458 224605 1460
rect 225094 1458 225154 1806
rect 224604 1398 225154 1458
rect 224604 1396 224605 1398
rect 224539 1395 224605 1396
rect 218654 990 220922 1050
rect 221046 1262 225338 1322
rect 221046 778 221106 1262
rect 225091 1188 225157 1189
rect 225091 1124 225092 1188
rect 225156 1124 225157 1188
rect 225091 1123 225157 1124
rect 218470 718 221106 778
rect 219203 644 219269 645
rect 217734 582 217840 642
rect 211294 446 211492 506
rect 211662 446 213930 506
rect 214054 446 217426 506
rect 217780 458 217840 582
rect 219203 580 219204 644
rect 219268 642 219269 644
rect 225094 642 225154 1123
rect 225278 1050 225338 1262
rect 225646 1050 225706 2350
rect 225830 1186 225890 2642
rect 226934 2410 226994 2942
rect 226198 2350 226994 2410
rect 226198 1322 226258 2350
rect 227854 1866 227914 2942
rect 226566 1818 227914 1866
rect 226714 1806 227914 1818
rect 228774 1730 228834 2942
rect 253430 2410 253490 2942
rect 227118 1670 228834 1730
rect 229510 2350 234170 2410
rect 227118 1325 227178 1670
rect 227486 1534 227730 1594
rect 227486 1325 227546 1534
rect 227670 1325 227730 1534
rect 229510 1458 229570 2350
rect 234110 1730 234170 2350
rect 245150 2350 245762 2410
rect 234291 1732 234357 1733
rect 234291 1730 234292 1732
rect 229142 1398 229570 1458
rect 231166 1670 233986 1730
rect 234110 1670 234292 1730
rect 229142 1325 229202 1398
rect 227115 1324 227181 1325
rect 226198 1262 226994 1322
rect 226747 1188 226813 1189
rect 226747 1186 226748 1188
rect 225830 1126 226748 1186
rect 226747 1124 226748 1126
rect 226812 1124 226813 1188
rect 226747 1123 226813 1124
rect 226934 1050 226994 1262
rect 227115 1260 227116 1324
rect 227180 1260 227181 1324
rect 227115 1259 227181 1260
rect 227483 1324 227549 1325
rect 227483 1260 227484 1324
rect 227548 1260 227549 1324
rect 227483 1259 227549 1260
rect 227667 1324 227733 1325
rect 227667 1260 227668 1324
rect 227732 1260 227733 1324
rect 227667 1259 227733 1260
rect 229139 1324 229205 1325
rect 229139 1260 229140 1324
rect 229204 1260 229205 1324
rect 229139 1259 229205 1260
rect 229323 1324 229389 1325
rect 229323 1260 229324 1324
rect 229388 1260 229389 1324
rect 229323 1259 229389 1260
rect 225278 990 226994 1050
rect 225646 778 225706 990
rect 229326 778 229386 1259
rect 231166 781 231226 1670
rect 233926 1594 233986 1670
rect 234291 1668 234292 1670
rect 234356 1668 234357 1732
rect 234291 1667 234357 1668
rect 237971 1732 238037 1733
rect 237971 1668 237972 1732
rect 238036 1668 238037 1732
rect 237971 1667 238037 1668
rect 237974 1594 238034 1667
rect 238707 1596 238773 1597
rect 238707 1594 238708 1596
rect 231350 1534 233802 1594
rect 233926 1534 234170 1594
rect 237974 1534 238708 1594
rect 231350 917 231410 1534
rect 231534 1262 233618 1322
rect 231347 916 231413 917
rect 231347 852 231348 916
rect 231412 852 231413 916
rect 231347 851 231413 852
rect 225646 718 229386 778
rect 231163 780 231229 781
rect 231163 716 231164 780
rect 231228 716 231229 780
rect 231163 715 231229 716
rect 231534 642 231594 1262
rect 219268 582 221290 642
rect 225094 582 231594 642
rect 232454 990 232882 1050
rect 219268 580 219269 582
rect 219203 579 219269 580
rect 198230 310 210802 370
rect 211432 370 211492 446
rect 214054 370 214114 446
rect 211432 310 214114 370
rect 221230 370 221290 582
rect 232454 458 232514 990
rect 232822 917 232882 990
rect 232635 916 232701 917
rect 232635 852 232636 916
rect 232700 852 232701 916
rect 232635 851 232701 852
rect 232819 916 232885 917
rect 232819 852 232820 916
rect 232884 852 232885 916
rect 232819 851 232885 852
rect 233371 916 233437 917
rect 233371 852 233372 916
rect 233436 852 233437 916
rect 233371 851 233437 852
rect 232638 778 232698 851
rect 232638 718 233250 778
rect 233190 458 233250 718
rect 233374 642 233434 851
rect 233558 778 233618 1262
rect 233742 917 233802 1534
rect 234110 1458 234170 1534
rect 238707 1532 238708 1534
rect 238772 1532 238773 1596
rect 238707 1531 238773 1532
rect 239075 1596 239141 1597
rect 239075 1532 239076 1596
rect 239140 1532 239141 1596
rect 239075 1531 239141 1532
rect 241835 1596 241901 1597
rect 241835 1532 241836 1596
rect 241900 1532 241901 1596
rect 241835 1531 241901 1532
rect 239078 1458 239138 1531
rect 234110 1398 239138 1458
rect 241838 1458 241898 1531
rect 245150 1461 245210 2350
rect 245702 1866 245762 2350
rect 253246 2350 253490 2410
rect 260238 2410 260298 2942
rect 260238 2350 261402 2410
rect 245702 1806 249258 1866
rect 245331 1732 245397 1733
rect 245331 1668 245332 1732
rect 245396 1730 245397 1732
rect 247539 1732 247605 1733
rect 245396 1670 247418 1730
rect 245396 1668 245397 1670
rect 245331 1667 245397 1668
rect 247358 1594 247418 1670
rect 247539 1668 247540 1732
rect 247604 1730 247605 1732
rect 247604 1670 248154 1730
rect 247604 1668 247605 1670
rect 247539 1667 247605 1668
rect 245334 1534 246866 1594
rect 247358 1534 247970 1594
rect 243123 1460 243189 1461
rect 243123 1458 243124 1460
rect 241838 1398 243124 1458
rect 243123 1396 243124 1398
rect 243188 1396 243189 1460
rect 243123 1395 243189 1396
rect 245147 1460 245213 1461
rect 245147 1396 245148 1460
rect 245212 1396 245213 1460
rect 245147 1395 245213 1396
rect 245334 1322 245394 1534
rect 246806 1461 246866 1534
rect 246619 1460 246685 1461
rect 245518 1398 246314 1458
rect 245518 1325 245578 1398
rect 234110 1262 245394 1322
rect 245515 1324 245581 1325
rect 233739 916 233805 917
rect 233739 852 233740 916
rect 233804 852 233805 916
rect 233739 851 233805 852
rect 234110 778 234170 1262
rect 245515 1260 245516 1324
rect 245580 1260 245581 1324
rect 245515 1259 245581 1260
rect 245699 1324 245765 1325
rect 245699 1260 245700 1324
rect 245764 1260 245765 1324
rect 245699 1259 245765 1260
rect 241250 990 242118 1050
rect 233558 718 234170 778
rect 245147 780 245213 781
rect 245147 716 245148 780
rect 245212 716 245213 780
rect 245147 715 245213 716
rect 233374 582 233618 642
rect 221230 310 224638 370
rect 233558 370 233618 582
rect 245150 370 245210 715
rect 245702 458 245762 1259
rect 233558 310 245210 370
rect 246254 370 246314 1398
rect 246619 1396 246620 1460
rect 246684 1396 246685 1460
rect 246619 1395 246685 1396
rect 246803 1460 246869 1461
rect 246803 1396 246804 1460
rect 246868 1396 246869 1460
rect 246803 1395 246869 1396
rect 246622 781 246682 1395
rect 247910 1325 247970 1534
rect 247907 1324 247973 1325
rect 247907 1260 247908 1324
rect 247972 1260 247973 1324
rect 247907 1259 247973 1260
rect 246806 1126 247786 1186
rect 246435 780 246501 781
rect 246435 716 246436 780
rect 246500 716 246501 780
rect 246435 715 246501 716
rect 246619 780 246685 781
rect 246619 716 246620 780
rect 246684 716 246685 780
rect 246619 715 246685 716
rect 246438 642 246498 715
rect 246806 642 246866 1126
rect 247539 1052 247605 1053
rect 247539 1050 247540 1052
rect 246438 582 246866 642
rect 246990 990 247540 1050
rect 246990 370 247050 990
rect 247539 988 247540 990
rect 247604 988 247605 1052
rect 247726 1050 247786 1126
rect 247907 1052 247973 1053
rect 247907 1050 247908 1052
rect 247726 990 247908 1050
rect 247539 987 247605 988
rect 247907 988 247908 990
rect 247972 988 247973 1052
rect 247907 987 247973 988
rect 248094 458 248154 1670
rect 248278 1534 249074 1594
rect 248278 645 248338 1534
rect 248827 1460 248893 1461
rect 248827 1396 248828 1460
rect 248892 1396 248893 1460
rect 248827 1395 248893 1396
rect 248275 644 248341 645
rect 248275 580 248276 644
rect 248340 580 248341 644
rect 248830 642 248890 1395
rect 249014 778 249074 1534
rect 249198 914 249258 1806
rect 253246 1597 253306 2350
rect 249747 1596 249813 1597
rect 249747 1532 249748 1596
rect 249812 1594 249813 1596
rect 253243 1596 253309 1597
rect 249812 1534 250178 1594
rect 249812 1532 249813 1534
rect 249747 1531 249813 1532
rect 250118 1461 250178 1534
rect 253243 1532 253244 1596
rect 253308 1532 253309 1596
rect 253795 1596 253861 1597
rect 253795 1594 253796 1596
rect 253243 1531 253309 1532
rect 253430 1534 253796 1594
rect 253430 1461 253490 1534
rect 253795 1532 253796 1534
rect 253860 1532 253861 1596
rect 258395 1596 258461 1597
rect 258395 1594 258396 1596
rect 253795 1531 253861 1532
rect 253982 1534 258396 1594
rect 250115 1460 250181 1461
rect 250115 1396 250116 1460
rect 250180 1396 250181 1460
rect 250115 1395 250181 1396
rect 253427 1460 253493 1461
rect 253427 1396 253428 1460
rect 253492 1396 253493 1460
rect 253427 1395 253493 1396
rect 250483 1324 250549 1325
rect 250483 1260 250484 1324
rect 250548 1260 250549 1324
rect 250483 1259 250549 1260
rect 251219 1324 251285 1325
rect 251219 1260 251220 1324
rect 251284 1322 251285 1324
rect 253059 1324 253125 1325
rect 253059 1322 253060 1324
rect 251284 1262 253060 1322
rect 251284 1260 251285 1262
rect 251219 1259 251285 1260
rect 253059 1260 253060 1262
rect 253124 1260 253125 1324
rect 253059 1259 253125 1260
rect 250486 1186 250546 1259
rect 250486 1126 252938 1186
rect 252691 1052 252757 1053
rect 252691 988 252692 1052
rect 252756 988 252757 1052
rect 252878 1050 252938 1126
rect 253427 1052 253493 1053
rect 253427 1050 253428 1052
rect 252878 990 253428 1050
rect 252691 987 252757 988
rect 253427 988 253428 990
rect 253492 988 253493 1052
rect 253427 987 253493 988
rect 250299 916 250365 917
rect 250299 914 250300 916
rect 249198 854 250300 914
rect 250299 852 250300 854
rect 250364 852 250365 916
rect 250299 851 250365 852
rect 251955 916 252021 917
rect 251955 852 251956 916
rect 252020 852 252021 916
rect 252694 914 252754 987
rect 253795 916 253861 917
rect 253795 914 253796 916
rect 252694 854 253796 914
rect 251955 851 252021 852
rect 253795 852 253796 854
rect 253860 852 253861 916
rect 253795 851 253861 852
rect 251958 778 252018 851
rect 249014 718 252018 778
rect 252323 780 252389 781
rect 252323 716 252324 780
rect 252388 778 252389 780
rect 252507 780 252573 781
rect 252507 778 252508 780
rect 252388 718 252508 778
rect 252388 716 252389 718
rect 252323 715 252389 716
rect 252507 716 252508 718
rect 252572 716 252573 780
rect 253982 778 254042 1534
rect 258395 1532 258396 1534
rect 258460 1532 258461 1596
rect 258395 1531 258461 1532
rect 260606 1534 261034 1594
rect 260606 1461 260666 1534
rect 260974 1461 261034 1534
rect 260603 1460 260669 1461
rect 260603 1396 260604 1460
rect 260668 1396 260669 1460
rect 260603 1395 260669 1396
rect 260971 1460 261037 1461
rect 260971 1396 260972 1460
rect 261036 1396 261037 1460
rect 260971 1395 261037 1396
rect 256371 1324 256437 1325
rect 256371 1260 256372 1324
rect 256436 1260 256437 1324
rect 261342 1322 261402 2350
rect 279006 2350 280538 2410
rect 262262 1806 266554 1866
rect 261707 1732 261773 1733
rect 261707 1668 261708 1732
rect 261772 1668 261773 1732
rect 261707 1667 261773 1668
rect 261710 1458 261770 1667
rect 261891 1596 261957 1597
rect 261891 1532 261892 1596
rect 261956 1594 261957 1596
rect 262262 1594 262322 1806
rect 266494 1730 266554 1806
rect 267782 1806 272258 1866
rect 267782 1730 267842 1806
rect 272198 1733 272258 1806
rect 279006 1733 279066 2350
rect 280478 1866 280538 2350
rect 279742 1806 280354 1866
rect 280478 1806 281274 1866
rect 266494 1670 267842 1730
rect 268699 1732 268765 1733
rect 268699 1668 268700 1732
rect 268764 1730 268765 1732
rect 272195 1732 272261 1733
rect 268764 1670 272074 1730
rect 268764 1668 268765 1670
rect 268699 1667 268765 1668
rect 261956 1534 262322 1594
rect 268886 1534 271890 1594
rect 261956 1532 261957 1534
rect 261891 1531 261957 1532
rect 268886 1461 268946 1534
rect 271830 1461 271890 1534
rect 268883 1460 268949 1461
rect 261710 1398 263058 1458
rect 262811 1324 262877 1325
rect 262811 1322 262812 1324
rect 256371 1259 256437 1260
rect 258214 1262 261218 1322
rect 261342 1262 262812 1322
rect 256374 1138 256434 1259
rect 256003 1052 256069 1053
rect 256003 1050 256004 1052
rect 255050 990 256004 1050
rect 256003 988 256004 990
rect 256068 988 256069 1052
rect 256003 987 256069 988
rect 255635 916 255701 917
rect 255635 852 255636 916
rect 255700 852 255701 916
rect 258214 1050 258274 1262
rect 258030 990 258274 1050
rect 260238 990 261034 1050
rect 255635 851 255701 852
rect 252507 715 252573 716
rect 252694 718 254042 778
rect 252694 642 252754 718
rect 248830 582 252754 642
rect 255638 642 255698 851
rect 258030 642 258090 990
rect 260238 781 260298 990
rect 260422 854 260850 914
rect 258211 780 258277 781
rect 258211 716 258212 780
rect 258276 778 258277 780
rect 260235 780 260301 781
rect 258276 718 259378 778
rect 258276 716 258277 718
rect 258211 715 258277 716
rect 255638 582 258090 642
rect 259318 642 259378 718
rect 260235 716 260236 780
rect 260300 716 260301 780
rect 260235 715 260301 716
rect 260422 642 260482 854
rect 260790 781 260850 854
rect 260787 780 260853 781
rect 260787 716 260788 780
rect 260852 716 260853 780
rect 260787 715 260853 716
rect 259318 582 260482 642
rect 248275 579 248341 580
rect 246254 310 247050 370
rect 260974 370 261034 990
rect 261158 781 261218 1262
rect 262811 1260 262812 1262
rect 262876 1260 262877 1324
rect 262811 1259 262877 1260
rect 262259 1052 262325 1053
rect 262259 988 262260 1052
rect 262324 1050 262325 1052
rect 262998 1050 263058 1398
rect 262324 990 263058 1050
rect 263182 1398 267474 1458
rect 262324 988 262325 990
rect 262259 987 262325 988
rect 261155 780 261221 781
rect 261155 716 261156 780
rect 261220 716 261221 780
rect 261155 715 261221 716
rect 263182 370 263242 1398
rect 264835 1324 264901 1325
rect 264835 1260 264836 1324
rect 264900 1260 264901 1324
rect 264835 1259 264901 1260
rect 264838 778 264898 1259
rect 265354 990 266958 1050
rect 264838 718 265266 778
rect 264835 644 264901 645
rect 264835 580 264836 644
rect 264900 580 264901 644
rect 264835 579 264901 580
rect 264838 458 264898 579
rect 260974 310 263242 370
rect 265206 370 265266 718
rect 267414 642 267474 1398
rect 268883 1396 268884 1460
rect 268948 1396 268949 1460
rect 268883 1395 268949 1396
rect 271827 1460 271893 1461
rect 271827 1396 271828 1460
rect 271892 1396 271893 1460
rect 272014 1458 272074 1670
rect 272195 1668 272196 1732
rect 272260 1668 272261 1732
rect 272195 1667 272261 1668
rect 279003 1732 279069 1733
rect 279003 1668 279004 1732
rect 279068 1668 279069 1732
rect 279003 1667 279069 1668
rect 272566 1534 273546 1594
rect 272566 1458 272626 1534
rect 273486 1461 273546 1534
rect 272014 1398 272626 1458
rect 273299 1460 273365 1461
rect 271827 1395 271893 1396
rect 273299 1396 273300 1460
rect 273364 1396 273365 1460
rect 273299 1395 273365 1396
rect 273483 1460 273549 1461
rect 273483 1396 273484 1460
rect 273548 1396 273549 1460
rect 273483 1395 273549 1396
rect 273667 1460 273733 1461
rect 273667 1396 273668 1460
rect 273732 1396 273733 1460
rect 273667 1395 273733 1396
rect 279371 1460 279437 1461
rect 279371 1396 279372 1460
rect 279436 1458 279437 1460
rect 279742 1458 279802 1806
rect 280294 1730 280354 1806
rect 280294 1670 280722 1730
rect 280475 1460 280541 1461
rect 279436 1398 279802 1458
rect 279926 1398 280170 1458
rect 279436 1396 279437 1398
rect 279371 1395 279437 1396
rect 268883 1188 268949 1189
rect 268883 1124 268884 1188
rect 268948 1124 268949 1188
rect 268883 1123 268949 1124
rect 266458 582 267474 642
rect 268886 642 268946 1123
rect 273302 1050 273362 1395
rect 273670 1050 273730 1395
rect 279555 1188 279621 1189
rect 279555 1124 279556 1188
rect 279620 1124 279621 1188
rect 279555 1123 279621 1124
rect 279558 1050 279618 1123
rect 273302 990 273730 1050
rect 273854 990 279618 1050
rect 273854 642 273914 990
rect 279926 642 279986 1398
rect 280110 1322 280170 1398
rect 280475 1396 280476 1460
rect 280540 1396 280541 1460
rect 280475 1395 280541 1396
rect 280478 1322 280538 1395
rect 280110 1262 280538 1322
rect 280662 781 280722 1670
rect 281214 1458 281274 1806
rect 294091 1766 294157 1767
rect 285627 1732 285693 1733
rect 285627 1668 285628 1732
rect 285692 1668 285693 1732
rect 294091 1702 294092 1766
rect 294156 1702 294157 1766
rect 294462 1733 294522 2942
rect 296118 2350 297282 2410
rect 294091 1701 294157 1702
rect 294459 1732 294525 1733
rect 285627 1667 285693 1668
rect 281395 1460 281461 1461
rect 281395 1458 281396 1460
rect 281214 1398 281396 1458
rect 281395 1396 281396 1398
rect 281460 1396 281461 1460
rect 285630 1458 285690 1667
rect 294094 1594 294154 1701
rect 294459 1668 294460 1732
rect 294524 1668 294525 1732
rect 294459 1667 294525 1668
rect 296118 1597 296178 2350
rect 296115 1596 296181 1597
rect 294094 1534 295810 1594
rect 285630 1398 289738 1458
rect 281395 1395 281461 1396
rect 281027 1324 281093 1325
rect 281027 1260 281028 1324
rect 281092 1322 281093 1324
rect 281092 1262 281642 1322
rect 281092 1260 281093 1262
rect 281027 1259 281093 1260
rect 280107 780 280173 781
rect 280107 716 280108 780
rect 280172 716 280173 780
rect 280107 715 280173 716
rect 280659 780 280725 781
rect 280659 716 280660 780
rect 280724 716 280725 780
rect 280659 715 280725 716
rect 268886 582 273914 642
rect 274038 582 279986 642
rect 274038 370 274098 582
rect 280110 458 280170 715
rect 281582 458 281642 1262
rect 289678 1189 289738 1398
rect 290046 1398 290842 1458
rect 290046 1189 290106 1398
rect 290782 1322 290842 1398
rect 294827 1324 294893 1325
rect 294827 1322 294828 1324
rect 290782 1262 291026 1322
rect 289675 1188 289741 1189
rect 289675 1124 289676 1188
rect 289740 1124 289741 1188
rect 289675 1123 289741 1124
rect 290043 1188 290109 1189
rect 290043 1124 290044 1188
rect 290108 1124 290109 1188
rect 290043 1123 290109 1124
rect 290411 1188 290477 1189
rect 290411 1124 290412 1188
rect 290476 1124 290477 1188
rect 290411 1123 290477 1124
rect 290414 458 290474 1123
rect 290966 778 291026 1262
rect 293910 1262 294828 1322
rect 293910 778 293970 1262
rect 294827 1260 294828 1262
rect 294892 1260 294893 1324
rect 294827 1259 294893 1260
rect 295750 1186 295810 1534
rect 296115 1532 296116 1596
rect 296180 1532 296181 1596
rect 296115 1531 296181 1532
rect 296851 1188 296917 1189
rect 296851 1186 296852 1188
rect 295750 1126 296852 1186
rect 296851 1124 296852 1126
rect 296916 1124 296917 1188
rect 296851 1123 296917 1124
rect 290966 718 293970 778
rect 294827 780 294893 781
rect 294827 716 294828 780
rect 294892 716 294893 780
rect 294827 715 294893 716
rect 294830 458 294890 715
rect 265206 310 274098 370
rect 290779 372 290845 373
rect 290779 308 290780 372
rect 290844 370 290845 372
rect 291147 372 291213 373
rect 291147 370 291148 372
rect 290844 310 291148 370
rect 290844 308 290845 310
rect 290779 307 290845 308
rect 291147 308 291148 310
rect 291212 308 291213 372
rect 291147 307 291213 308
rect 297222 370 297282 2350
rect 310102 1594 310162 2942
rect 311206 2410 311266 2942
rect 310470 2350 311266 2410
rect 325006 2350 328378 2410
rect 310470 1733 310530 2350
rect 310467 1732 310533 1733
rect 310467 1668 310468 1732
rect 310532 1668 310533 1732
rect 310467 1667 310533 1668
rect 310651 1732 310717 1733
rect 310651 1668 310652 1732
rect 310716 1668 310717 1732
rect 325006 1730 325066 2350
rect 310651 1667 310717 1668
rect 324822 1670 325066 1730
rect 328318 1730 328378 2350
rect 328318 1670 328746 1730
rect 310654 1594 310714 1667
rect 310102 1534 310714 1594
rect 324822 1325 324882 1670
rect 317827 1324 317893 1325
rect 317827 1322 317828 1324
rect 299982 1262 303906 1322
rect 299982 370 300042 1262
rect 303294 1126 303722 1186
rect 303294 1053 303354 1126
rect 303291 1052 303357 1053
rect 303291 988 303292 1052
rect 303356 988 303357 1052
rect 303291 987 303357 988
rect 297222 310 300042 370
rect 303662 370 303722 1126
rect 303846 1050 303906 1262
rect 317462 1262 317828 1322
rect 308811 1188 308877 1189
rect 308811 1124 308812 1188
rect 308876 1186 308877 1188
rect 308876 1126 310162 1186
rect 308876 1124 308877 1126
rect 308811 1123 308877 1124
rect 303846 990 309978 1050
rect 309918 917 309978 990
rect 309915 916 309981 917
rect 309915 852 309916 916
rect 309980 852 309981 916
rect 310102 914 310162 1126
rect 314883 916 314949 917
rect 314883 914 314884 916
rect 310102 854 314884 914
rect 309915 851 309981 852
rect 314883 852 314884 854
rect 314948 852 314949 916
rect 317462 914 317522 1262
rect 317827 1260 317828 1262
rect 317892 1260 317893 1324
rect 317827 1259 317893 1260
rect 324819 1324 324885 1325
rect 324819 1260 324820 1324
rect 324884 1260 324885 1324
rect 324819 1259 324885 1260
rect 327763 1324 327829 1325
rect 327763 1260 327764 1324
rect 327828 1260 327829 1324
rect 327763 1259 327829 1260
rect 327766 1138 327826 1259
rect 328315 1188 328381 1189
rect 314883 851 314949 852
rect 315070 854 317522 914
rect 328315 1124 328316 1188
rect 328380 1186 328381 1188
rect 328499 1188 328565 1189
rect 328499 1186 328500 1188
rect 328380 1126 328500 1186
rect 328380 1124 328381 1126
rect 328315 1123 328381 1124
rect 328499 1124 328500 1126
rect 328564 1124 328565 1188
rect 328686 1186 328746 1670
rect 328686 1126 329114 1186
rect 328499 1123 328565 1124
rect 329054 917 329114 1126
rect 328315 916 328381 917
rect 315070 370 315130 854
rect 328315 852 328316 916
rect 328380 852 328381 916
rect 328315 851 328381 852
rect 328545 916 328611 917
rect 328545 852 328546 916
rect 328610 852 328611 916
rect 328545 851 328611 852
rect 329051 916 329117 917
rect 329051 852 329052 916
rect 329116 852 329117 916
rect 329051 851 329117 852
rect 328318 642 328378 851
rect 328548 642 328608 851
rect 328318 582 328608 642
rect 336782 458 336842 2942
rect 348926 1189 348986 2942
rect 354262 1597 354322 2942
rect 354259 1596 354325 1597
rect 354259 1532 354260 1596
rect 354324 1532 354325 1596
rect 354259 1531 354325 1532
rect 372478 1325 372538 2942
rect 385723 1732 385789 1733
rect 385723 1668 385724 1732
rect 385788 1730 385789 1732
rect 385788 1670 385970 1730
rect 385788 1668 385789 1670
rect 385723 1667 385789 1668
rect 372475 1324 372541 1325
rect 372475 1260 372476 1324
rect 372540 1260 372541 1324
rect 372475 1259 372541 1260
rect 348923 1188 348989 1189
rect 348923 1124 348924 1188
rect 348988 1124 348989 1188
rect 370451 1188 370517 1189
rect 370451 1138 370452 1188
rect 370516 1138 370517 1188
rect 348923 1123 348989 1124
rect 362726 990 363154 1050
rect 358123 916 358189 917
rect 338806 645 338866 902
rect 338619 644 338685 645
rect 338619 580 338620 644
rect 338684 580 338685 644
rect 338619 579 338685 580
rect 338803 644 338869 645
rect 338803 580 338804 644
rect 338868 580 338869 644
rect 338803 579 338869 580
rect 303662 310 315130 370
rect 338622 370 338682 579
rect 339542 370 339602 902
rect 350030 645 350090 902
rect 353894 781 353954 902
rect 358123 852 358124 916
rect 358188 852 358189 916
rect 358123 851 358189 852
rect 353891 780 353957 781
rect 353891 716 353892 780
rect 353956 716 353957 780
rect 353891 715 353957 716
rect 342667 644 342733 645
rect 342667 580 342668 644
rect 342732 580 342733 644
rect 342667 579 342733 580
rect 350027 644 350093 645
rect 350027 580 350028 644
rect 350092 580 350093 644
rect 350027 579 350093 580
rect 338622 310 339602 370
rect 342670 370 342730 579
rect 358126 458 358186 851
rect 362726 781 362786 990
rect 362723 780 362789 781
rect 362723 716 362724 780
rect 362788 716 362789 780
rect 362723 715 362789 716
rect 363094 458 363154 990
rect 385910 781 385970 1670
rect 419398 1325 419458 2942
rect 419395 1324 419461 1325
rect 419395 1260 419396 1324
rect 419460 1260 419461 1324
rect 419395 1259 419461 1260
rect 385907 780 385973 781
rect 385907 716 385908 780
rect 385972 716 385973 780
rect 385907 715 385973 716
rect 390507 644 390573 645
rect 390507 580 390508 644
rect 390572 580 390573 644
rect 390507 579 390573 580
rect 342670 310 343502 370
rect 390510 373 390570 579
rect 390507 372 390573 373
rect 390507 308 390508 372
rect 390572 308 390573 372
rect 390507 307 390573 308
rect 414614 370 414674 902
rect 418846 373 418906 902
rect 414210 310 414674 370
rect 418843 372 418909 373
rect 418843 308 418844 372
rect 418908 308 418909 372
rect 418843 307 418909 308
rect 426942 373 427002 2942
rect 440190 781 440250 902
rect 440187 780 440253 781
rect 440187 716 440188 780
rect 440252 716 440253 780
rect 440187 715 440253 716
rect 430619 644 430685 645
rect 430619 580 430620 644
rect 430684 580 430685 644
rect 430619 579 430685 580
rect 434483 644 434549 645
rect 434483 580 434484 644
rect 434548 580 434549 644
rect 434483 579 434549 580
rect 430622 458 430682 579
rect 434486 458 434546 579
rect 426939 372 427005 373
rect 426939 308 426940 372
rect 427004 308 427005 372
rect 426939 307 427005 308
rect 442950 373 443010 2942
rect 473126 2350 473416 2410
rect 449755 780 449821 781
rect 449755 716 449756 780
rect 449820 716 449821 780
rect 449755 715 449821 716
rect 449758 458 449818 715
rect 463006 509 463066 902
rect 463003 508 463069 509
rect 442947 372 443013 373
rect 442947 308 442948 372
rect 443012 308 443013 372
rect 442947 307 443013 308
rect 463003 444 463004 508
rect 463068 444 463069 508
rect 469075 508 469141 509
rect 469075 458 469076 508
rect 469140 458 469141 508
rect 463003 443 463069 444
rect 473126 373 473186 2350
rect 473356 1730 473416 2350
rect 473356 1670 473554 1730
rect 473494 509 473554 1670
rect 483798 1189 483858 2942
rect 513238 1733 513298 2942
rect 514526 2410 514586 2942
rect 514158 2350 514586 2410
rect 513235 1732 513301 1733
rect 513235 1668 513236 1732
rect 513300 1668 513301 1732
rect 513235 1667 513301 1668
rect 514158 1189 514218 2350
rect 558870 1597 558930 9830
rect 559054 1597 559114 11102
rect 559790 4390 560070 4450
rect 558867 1596 558933 1597
rect 558867 1532 558868 1596
rect 558932 1532 558933 1596
rect 558867 1531 558933 1532
rect 559051 1596 559117 1597
rect 559051 1532 559052 1596
rect 559116 1532 559117 1596
rect 559051 1531 559117 1532
rect 559422 1461 559482 3622
rect 559419 1460 559485 1461
rect 559419 1396 559420 1460
rect 559484 1396 559485 1460
rect 559419 1395 559485 1396
rect 483795 1188 483861 1189
rect 483795 1124 483796 1188
rect 483860 1124 483861 1188
rect 483795 1123 483861 1124
rect 514155 1188 514221 1189
rect 514155 1124 514156 1188
rect 514220 1124 514221 1188
rect 514155 1123 514221 1124
rect 522254 509 522314 902
rect 539547 780 539613 781
rect 539547 716 539548 780
rect 539612 716 539613 780
rect 539547 715 539613 716
rect 539550 509 539610 715
rect 559790 645 559850 4390
rect 560158 1461 560218 3622
rect 560155 1460 560221 1461
rect 560155 1396 560156 1460
rect 560220 1396 560221 1460
rect 560155 1395 560221 1396
rect 561446 1189 561506 26062
rect 562182 25618 562242 32182
rect 561443 1188 561509 1189
rect 561443 1124 561444 1188
rect 561508 1124 561509 1188
rect 561443 1123 561509 1124
rect 563102 781 563162 680443
rect 563651 680372 563717 680373
rect 563651 680308 563652 680372
rect 563716 680308 563717 680372
rect 563651 680307 563717 680308
rect 563654 1138 563714 680307
rect 564574 917 564634 680443
rect 567147 680444 567148 680508
rect 567212 680444 567213 680508
rect 567147 680443 567213 680444
rect 566411 680372 566477 680373
rect 566411 680308 566412 680372
rect 566476 680308 566477 680372
rect 566411 680307 566477 680308
rect 564942 1325 565002 680222
rect 566414 1461 566474 680307
rect 567150 1733 567210 680443
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 570459 284612 570525 284613
rect 570459 284610 570460 284612
rect 569910 284550 570460 284610
rect 569910 283930 569970 284550
rect 570459 284548 570460 284550
rect 570524 284548 570525 284612
rect 570459 284547 570525 284548
rect 569358 283870 569970 283930
rect 569358 273730 569418 283870
rect 569358 273670 569786 273730
rect 569726 267610 569786 273670
rect 569726 267550 570338 267610
rect 569217 260132 569283 260133
rect 569217 260130 569218 260132
rect 568806 260070 569218 260130
rect 568806 252650 568866 260070
rect 569217 260068 569218 260070
rect 569282 260068 569283 260132
rect 569217 260067 569283 260068
rect 570278 258090 570338 267550
rect 569910 258030 570338 258090
rect 569910 256730 569970 258030
rect 568622 252590 568866 252650
rect 569358 256670 569970 256730
rect 568622 248570 568682 252590
rect 568392 248510 568682 248570
rect 568392 248437 568452 248510
rect 568389 248436 568455 248437
rect 568389 248372 568390 248436
rect 568454 248372 568455 248436
rect 568389 248371 568455 248372
rect 568849 222324 568915 222325
rect 568849 222260 568850 222324
rect 568914 222260 568915 222324
rect 568849 222259 568915 222260
rect 568852 222050 568912 222259
rect 568254 221990 568912 222050
rect 568254 209810 568314 221990
rect 568254 209750 568498 209810
rect 568438 194850 568498 209750
rect 569358 194850 569418 256670
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 568438 194790 568866 194850
rect 569358 194790 570706 194850
rect 568573 193628 568639 193629
rect 568573 193564 568574 193628
rect 568638 193626 568639 193628
rect 568638 193564 568682 193626
rect 568573 193563 568682 193564
rect 568297 193492 568363 193493
rect 568297 193490 568298 193492
rect 568254 193428 568298 193490
rect 568362 193428 568363 193492
rect 568254 193427 568363 193428
rect 568254 174450 568314 193427
rect 568622 192810 568682 193563
rect 568806 193490 568866 194790
rect 570275 193628 570341 193629
rect 570275 193626 570276 193628
rect 569174 193566 570276 193626
rect 569174 193490 569234 193566
rect 570275 193564 570276 193566
rect 570340 193564 570341 193628
rect 570275 193563 570341 193564
rect 570646 193493 570706 194790
rect 570459 193492 570525 193493
rect 570459 193490 570460 193492
rect 568806 193430 569234 193490
rect 569358 193430 570460 193490
rect 568622 192750 568866 192810
rect 568806 178530 568866 192750
rect 569171 178532 569237 178533
rect 569171 178530 569172 178532
rect 568806 178470 569172 178530
rect 569171 178468 569172 178470
rect 569236 178468 569237 178532
rect 569171 178467 569237 178468
rect 568481 174588 568547 174589
rect 568481 174524 568482 174588
rect 568546 174524 568547 174588
rect 568481 174523 568547 174524
rect 568484 174450 568544 174523
rect 568254 174390 568544 174450
rect 569358 166290 569418 193430
rect 570459 193428 570460 193430
rect 570524 193428 570525 193492
rect 570459 193427 570525 193428
rect 570643 193492 570709 193493
rect 570643 193428 570644 193492
rect 570708 193428 570709 193492
rect 570643 193427 570709 193428
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 569358 166230 569786 166290
rect 569726 124810 569786 166230
rect 569358 124750 569786 124810
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 569358 100330 569418 124750
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 569358 100270 570338 100330
rect 570278 99381 570338 100270
rect 570275 99380 570341 99381
rect 570275 99316 570276 99380
rect 570340 99316 570341 99380
rect 570275 99315 570341 99316
rect 570459 90132 570525 90133
rect 570459 90130 570460 90132
rect 569542 90070 570460 90130
rect 569542 50690 569602 90070
rect 570459 90068 570460 90070
rect 570524 90068 570525 90132
rect 570459 90067 570525 90068
rect 569358 50630 569602 50690
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 569358 43210 569418 50630
rect 569358 43150 570522 43210
rect 570462 36410 570522 43150
rect 569174 36350 570522 36410
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 569174 1733 569234 36350
rect 570275 34916 570341 34917
rect 570275 34852 570276 34916
rect 570340 34852 570341 34916
rect 570275 34851 570341 34852
rect 570278 32418 570338 34851
rect 570275 12340 570341 12341
rect 570275 12276 570276 12340
rect 570340 12276 570341 12340
rect 570275 12275 570341 12276
rect 570278 11338 570338 12275
rect 569542 1733 569602 3622
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 567147 1732 567213 1733
rect 567147 1668 567148 1732
rect 567212 1668 567213 1732
rect 567147 1667 567213 1668
rect 569171 1732 569237 1733
rect 569171 1668 569172 1732
rect 569236 1668 569237 1732
rect 569171 1667 569237 1668
rect 569539 1732 569605 1733
rect 569539 1668 569540 1732
rect 569604 1668 569605 1732
rect 569539 1667 569605 1668
rect 566411 1460 566477 1461
rect 566411 1396 566412 1460
rect 566476 1396 566477 1460
rect 566411 1395 566477 1396
rect 564939 1324 565005 1325
rect 564939 1260 564940 1324
rect 565004 1260 565005 1324
rect 564939 1259 565005 1260
rect 564571 916 564637 917
rect 564571 852 564572 916
rect 564636 852 564637 916
rect 564571 851 564637 852
rect 563099 780 563165 781
rect 563099 716 563100 780
rect 563164 716 563165 780
rect 563099 715 563165 716
rect 559787 644 559853 645
rect 559787 580 559788 644
rect 559852 580 559853 644
rect 559787 579 559853 580
rect 473491 508 473557 509
rect 473491 444 473492 508
rect 473556 444 473557 508
rect 522251 508 522317 509
rect 473491 443 473557 444
rect 473123 372 473189 373
rect 473123 308 473124 372
rect 473188 308 473189 372
rect 473123 307 473189 308
rect 522251 444 522252 508
rect 522316 444 522317 508
rect 522251 443 522317 444
rect 539547 508 539613 509
rect 539547 444 539548 508
rect 539612 444 539613 508
rect 539547 443 539613 444
rect 504403 172 504404 222
rect 504468 172 504469 222
rect 504403 171 504469 172
rect 119540 38 135178 98
rect 119540 36 119541 38
rect 119475 35 119541 36
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586240 668454 586840 705202
rect 586240 668218 586422 668454
rect 586658 668218 586840 668454
rect 586240 668134 586840 668218
rect 586240 667898 586422 668134
rect 586658 667898 586840 668134
rect 586240 632454 586840 667898
rect 586240 632218 586422 632454
rect 586658 632218 586840 632454
rect 586240 632134 586840 632218
rect 586240 631898 586422 632134
rect 586658 631898 586840 632134
rect 586240 596454 586840 631898
rect 586240 596218 586422 596454
rect 586658 596218 586840 596454
rect 586240 596134 586840 596218
rect 586240 595898 586422 596134
rect 586658 595898 586840 596134
rect 586240 560454 586840 595898
rect 586240 560218 586422 560454
rect 586658 560218 586840 560454
rect 586240 560134 586840 560218
rect 586240 559898 586422 560134
rect 586658 559898 586840 560134
rect 586240 524454 586840 559898
rect 586240 524218 586422 524454
rect 586658 524218 586840 524454
rect 586240 524134 586840 524218
rect 586240 523898 586422 524134
rect 586658 523898 586840 524134
rect 586240 488454 586840 523898
rect 586240 488218 586422 488454
rect 586658 488218 586840 488454
rect 586240 488134 586840 488218
rect 586240 487898 586422 488134
rect 586658 487898 586840 488134
rect 586240 452454 586840 487898
rect 586240 452218 586422 452454
rect 586658 452218 586840 452454
rect 586240 452134 586840 452218
rect 586240 451898 586422 452134
rect 586658 451898 586840 452134
rect 586240 416454 586840 451898
rect 586240 416218 586422 416454
rect 586658 416218 586840 416454
rect 586240 416134 586840 416218
rect 586240 415898 586422 416134
rect 586658 415898 586840 416134
rect 586240 380454 586840 415898
rect 586240 380218 586422 380454
rect 586658 380218 586840 380454
rect 586240 380134 586840 380218
rect 586240 379898 586422 380134
rect 586658 379898 586840 380134
rect 586240 344454 586840 379898
rect 586240 344218 586422 344454
rect 586658 344218 586840 344454
rect 586240 344134 586840 344218
rect 586240 343898 586422 344134
rect 586658 343898 586840 344134
rect 586240 308454 586840 343898
rect 586240 308218 586422 308454
rect 586658 308218 586840 308454
rect 586240 308134 586840 308218
rect 586240 307898 586422 308134
rect 586658 307898 586840 308134
rect 586240 272454 586840 307898
rect 586240 272218 586422 272454
rect 586658 272218 586840 272454
rect 586240 272134 586840 272218
rect 586240 271898 586422 272134
rect 586658 271898 586840 272134
rect 586240 236454 586840 271898
rect 586240 236218 586422 236454
rect 586658 236218 586840 236454
rect 586240 236134 586840 236218
rect 586240 235898 586422 236134
rect 586658 235898 586840 236134
rect 586240 200454 586840 235898
rect 586240 200218 586422 200454
rect 586658 200218 586840 200454
rect 586240 200134 586840 200218
rect 586240 199898 586422 200134
rect 586658 199898 586840 200134
rect 586240 164454 586840 199898
rect 586240 164218 586422 164454
rect 586658 164218 586840 164454
rect 586240 164134 586840 164218
rect 586240 163898 586422 164134
rect 586658 163898 586840 164134
rect 586240 128454 586840 163898
rect 586240 128218 586422 128454
rect 586658 128218 586840 128454
rect 586240 128134 586840 128218
rect 586240 127898 586422 128134
rect 586658 127898 586840 128134
rect 586240 92454 586840 127898
rect 586240 92218 586422 92454
rect 586658 92218 586840 92454
rect 586240 92134 586840 92218
rect 586240 91898 586422 92134
rect 586658 91898 586840 92134
rect 586240 56454 586840 91898
rect 586240 56218 586422 56454
rect 586658 56218 586840 56454
rect 586240 56134 586840 56218
rect 586240 55898 586422 56134
rect 586658 55898 586840 56134
rect 586240 20454 586840 55898
rect 586240 20218 586422 20454
rect 586658 20218 586840 20454
rect 586240 20134 586840 20218
rect 586240 19898 586422 20134
rect 586658 19898 586840 20134
rect -2916 -1502 -2734 -1266
rect -2498 -1502 -2316 -1266
rect -2916 -1586 -2316 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 -2316 -1586
rect -2916 -1844 -2316 -1822
rect 586240 -1266 586840 19898
rect 586240 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect 586240 -1586 586840 -1502
rect 586240 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect 586240 -1844 586840 -1822
rect 587160 690054 587760 706122
rect 587160 689818 587342 690054
rect 587578 689818 587760 690054
rect 587160 689734 587760 689818
rect 587160 689498 587342 689734
rect 587578 689498 587760 689734
rect 587160 654054 587760 689498
rect 587160 653818 587342 654054
rect 587578 653818 587760 654054
rect 587160 653734 587760 653818
rect 587160 653498 587342 653734
rect 587578 653498 587760 653734
rect 587160 618054 587760 653498
rect 587160 617818 587342 618054
rect 587578 617818 587760 618054
rect 587160 617734 587760 617818
rect 587160 617498 587342 617734
rect 587578 617498 587760 617734
rect 587160 582054 587760 617498
rect 587160 581818 587342 582054
rect 587578 581818 587760 582054
rect 587160 581734 587760 581818
rect 587160 581498 587342 581734
rect 587578 581498 587760 581734
rect 587160 546054 587760 581498
rect 587160 545818 587342 546054
rect 587578 545818 587760 546054
rect 587160 545734 587760 545818
rect 587160 545498 587342 545734
rect 587578 545498 587760 545734
rect 587160 510054 587760 545498
rect 587160 509818 587342 510054
rect 587578 509818 587760 510054
rect 587160 509734 587760 509818
rect 587160 509498 587342 509734
rect 587578 509498 587760 509734
rect 587160 474054 587760 509498
rect 587160 473818 587342 474054
rect 587578 473818 587760 474054
rect 587160 473734 587760 473818
rect 587160 473498 587342 473734
rect 587578 473498 587760 473734
rect 587160 438054 587760 473498
rect 587160 437818 587342 438054
rect 587578 437818 587760 438054
rect 587160 437734 587760 437818
rect 587160 437498 587342 437734
rect 587578 437498 587760 437734
rect 587160 402054 587760 437498
rect 587160 401818 587342 402054
rect 587578 401818 587760 402054
rect 587160 401734 587760 401818
rect 587160 401498 587342 401734
rect 587578 401498 587760 401734
rect 587160 366054 587760 401498
rect 587160 365818 587342 366054
rect 587578 365818 587760 366054
rect 587160 365734 587760 365818
rect 587160 365498 587342 365734
rect 587578 365498 587760 365734
rect 587160 330054 587760 365498
rect 587160 329818 587342 330054
rect 587578 329818 587760 330054
rect 587160 329734 587760 329818
rect 587160 329498 587342 329734
rect 587578 329498 587760 329734
rect 587160 294054 587760 329498
rect 587160 293818 587342 294054
rect 587578 293818 587760 294054
rect 587160 293734 587760 293818
rect 587160 293498 587342 293734
rect 587578 293498 587760 293734
rect 587160 258054 587760 293498
rect 587160 257818 587342 258054
rect 587578 257818 587760 258054
rect 587160 257734 587760 257818
rect 587160 257498 587342 257734
rect 587578 257498 587760 257734
rect 587160 222054 587760 257498
rect 587160 221818 587342 222054
rect 587578 221818 587760 222054
rect 587160 221734 587760 221818
rect 587160 221498 587342 221734
rect 587578 221498 587760 221734
rect 587160 186054 587760 221498
rect 587160 185818 587342 186054
rect 587578 185818 587760 186054
rect 587160 185734 587760 185818
rect 587160 185498 587342 185734
rect 587578 185498 587760 185734
rect 587160 150054 587760 185498
rect 587160 149818 587342 150054
rect 587578 149818 587760 150054
rect 587160 149734 587760 149818
rect 587160 149498 587342 149734
rect 587578 149498 587760 149734
rect 587160 114054 587760 149498
rect 587160 113818 587342 114054
rect 587578 113818 587760 114054
rect 587160 113734 587760 113818
rect 587160 113498 587342 113734
rect 587578 113498 587760 113734
rect 587160 78054 587760 113498
rect 587160 77818 587342 78054
rect 587578 77818 587760 78054
rect 587160 77734 587760 77818
rect 587160 77498 587342 77734
rect 587578 77498 587760 77734
rect 587160 42054 587760 77498
rect 587160 41818 587342 42054
rect 587578 41818 587760 42054
rect 587160 41734 587760 41818
rect 587160 41498 587342 41734
rect 587578 41498 587760 41734
rect 587160 6054 587760 41498
rect 587160 5818 587342 6054
rect 587578 5818 587760 6054
rect 587160 5734 587760 5818
rect 587160 5498 587342 5734
rect 587578 5498 587760 5734
rect -3836 -2422 -3654 -2186
rect -3418 -2422 -3236 -2186
rect -3836 -2506 -3236 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 -3236 -2506
rect -3836 -2764 -3236 -2742
rect 587160 -2186 587760 5498
rect 587160 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect 587160 -2506 587760 -2422
rect 587160 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect 587160 -2764 587760 -2742
rect 588080 672054 588680 707042
rect 588080 671818 588262 672054
rect 588498 671818 588680 672054
rect 588080 671734 588680 671818
rect 588080 671498 588262 671734
rect 588498 671498 588680 671734
rect 588080 636054 588680 671498
rect 588080 635818 588262 636054
rect 588498 635818 588680 636054
rect 588080 635734 588680 635818
rect 588080 635498 588262 635734
rect 588498 635498 588680 635734
rect 588080 600054 588680 635498
rect 588080 599818 588262 600054
rect 588498 599818 588680 600054
rect 588080 599734 588680 599818
rect 588080 599498 588262 599734
rect 588498 599498 588680 599734
rect 588080 564054 588680 599498
rect 588080 563818 588262 564054
rect 588498 563818 588680 564054
rect 588080 563734 588680 563818
rect 588080 563498 588262 563734
rect 588498 563498 588680 563734
rect 588080 528054 588680 563498
rect 588080 527818 588262 528054
rect 588498 527818 588680 528054
rect 588080 527734 588680 527818
rect 588080 527498 588262 527734
rect 588498 527498 588680 527734
rect 588080 492054 588680 527498
rect 588080 491818 588262 492054
rect 588498 491818 588680 492054
rect 588080 491734 588680 491818
rect 588080 491498 588262 491734
rect 588498 491498 588680 491734
rect 588080 456054 588680 491498
rect 588080 455818 588262 456054
rect 588498 455818 588680 456054
rect 588080 455734 588680 455818
rect 588080 455498 588262 455734
rect 588498 455498 588680 455734
rect 588080 420054 588680 455498
rect 588080 419818 588262 420054
rect 588498 419818 588680 420054
rect 588080 419734 588680 419818
rect 588080 419498 588262 419734
rect 588498 419498 588680 419734
rect 588080 384054 588680 419498
rect 588080 383818 588262 384054
rect 588498 383818 588680 384054
rect 588080 383734 588680 383818
rect 588080 383498 588262 383734
rect 588498 383498 588680 383734
rect 588080 348054 588680 383498
rect 588080 347818 588262 348054
rect 588498 347818 588680 348054
rect 588080 347734 588680 347818
rect 588080 347498 588262 347734
rect 588498 347498 588680 347734
rect 588080 312054 588680 347498
rect 588080 311818 588262 312054
rect 588498 311818 588680 312054
rect 588080 311734 588680 311818
rect 588080 311498 588262 311734
rect 588498 311498 588680 311734
rect 588080 276054 588680 311498
rect 588080 275818 588262 276054
rect 588498 275818 588680 276054
rect 588080 275734 588680 275818
rect 588080 275498 588262 275734
rect 588498 275498 588680 275734
rect 588080 240054 588680 275498
rect 588080 239818 588262 240054
rect 588498 239818 588680 240054
rect 588080 239734 588680 239818
rect 588080 239498 588262 239734
rect 588498 239498 588680 239734
rect 588080 204054 588680 239498
rect 588080 203818 588262 204054
rect 588498 203818 588680 204054
rect 588080 203734 588680 203818
rect 588080 203498 588262 203734
rect 588498 203498 588680 203734
rect 588080 168054 588680 203498
rect 588080 167818 588262 168054
rect 588498 167818 588680 168054
rect 588080 167734 588680 167818
rect 588080 167498 588262 167734
rect 588498 167498 588680 167734
rect 588080 132054 588680 167498
rect 588080 131818 588262 132054
rect 588498 131818 588680 132054
rect 588080 131734 588680 131818
rect 588080 131498 588262 131734
rect 588498 131498 588680 131734
rect 588080 96054 588680 131498
rect 588080 95818 588262 96054
rect 588498 95818 588680 96054
rect 588080 95734 588680 95818
rect 588080 95498 588262 95734
rect 588498 95498 588680 95734
rect 588080 60054 588680 95498
rect 588080 59818 588262 60054
rect 588498 59818 588680 60054
rect 588080 59734 588680 59818
rect 588080 59498 588262 59734
rect 588498 59498 588680 59734
rect 588080 24054 588680 59498
rect 588080 23818 588262 24054
rect 588498 23818 588680 24054
rect 588080 23734 588680 23818
rect 588080 23498 588262 23734
rect 588498 23498 588680 23734
rect -4756 -3342 -4574 -3106
rect -4338 -3342 -4156 -3106
rect -4756 -3426 -4156 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 -4156 -3426
rect -4756 -3684 -4156 -3662
rect 588080 -3106 588680 23498
rect 588080 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect 588080 -3426 588680 -3342
rect 588080 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect 588080 -3684 588680 -3662
rect 589000 693654 589600 707962
rect 589000 693418 589182 693654
rect 589418 693418 589600 693654
rect 589000 693334 589600 693418
rect 589000 693098 589182 693334
rect 589418 693098 589600 693334
rect 589000 657654 589600 693098
rect 589000 657418 589182 657654
rect 589418 657418 589600 657654
rect 589000 657334 589600 657418
rect 589000 657098 589182 657334
rect 589418 657098 589600 657334
rect 589000 621654 589600 657098
rect 589000 621418 589182 621654
rect 589418 621418 589600 621654
rect 589000 621334 589600 621418
rect 589000 621098 589182 621334
rect 589418 621098 589600 621334
rect 589000 585654 589600 621098
rect 589000 585418 589182 585654
rect 589418 585418 589600 585654
rect 589000 585334 589600 585418
rect 589000 585098 589182 585334
rect 589418 585098 589600 585334
rect 589000 549654 589600 585098
rect 589000 549418 589182 549654
rect 589418 549418 589600 549654
rect 589000 549334 589600 549418
rect 589000 549098 589182 549334
rect 589418 549098 589600 549334
rect 589000 513654 589600 549098
rect 589000 513418 589182 513654
rect 589418 513418 589600 513654
rect 589000 513334 589600 513418
rect 589000 513098 589182 513334
rect 589418 513098 589600 513334
rect 589000 477654 589600 513098
rect 589000 477418 589182 477654
rect 589418 477418 589600 477654
rect 589000 477334 589600 477418
rect 589000 477098 589182 477334
rect 589418 477098 589600 477334
rect 589000 441654 589600 477098
rect 589000 441418 589182 441654
rect 589418 441418 589600 441654
rect 589000 441334 589600 441418
rect 589000 441098 589182 441334
rect 589418 441098 589600 441334
rect 589000 405654 589600 441098
rect 589000 405418 589182 405654
rect 589418 405418 589600 405654
rect 589000 405334 589600 405418
rect 589000 405098 589182 405334
rect 589418 405098 589600 405334
rect 589000 369654 589600 405098
rect 589000 369418 589182 369654
rect 589418 369418 589600 369654
rect 589000 369334 589600 369418
rect 589000 369098 589182 369334
rect 589418 369098 589600 369334
rect 589000 333654 589600 369098
rect 589000 333418 589182 333654
rect 589418 333418 589600 333654
rect 589000 333334 589600 333418
rect 589000 333098 589182 333334
rect 589418 333098 589600 333334
rect 589000 297654 589600 333098
rect 589000 297418 589182 297654
rect 589418 297418 589600 297654
rect 589000 297334 589600 297418
rect 589000 297098 589182 297334
rect 589418 297098 589600 297334
rect 589000 261654 589600 297098
rect 589000 261418 589182 261654
rect 589418 261418 589600 261654
rect 589000 261334 589600 261418
rect 589000 261098 589182 261334
rect 589418 261098 589600 261334
rect 589000 225654 589600 261098
rect 589000 225418 589182 225654
rect 589418 225418 589600 225654
rect 589000 225334 589600 225418
rect 589000 225098 589182 225334
rect 589418 225098 589600 225334
rect 589000 189654 589600 225098
rect 589000 189418 589182 189654
rect 589418 189418 589600 189654
rect 589000 189334 589600 189418
rect 589000 189098 589182 189334
rect 589418 189098 589600 189334
rect 589000 153654 589600 189098
rect 589000 153418 589182 153654
rect 589418 153418 589600 153654
rect 589000 153334 589600 153418
rect 589000 153098 589182 153334
rect 589418 153098 589600 153334
rect 589000 117654 589600 153098
rect 589000 117418 589182 117654
rect 589418 117418 589600 117654
rect 589000 117334 589600 117418
rect 589000 117098 589182 117334
rect 589418 117098 589600 117334
rect 589000 81654 589600 117098
rect 589000 81418 589182 81654
rect 589418 81418 589600 81654
rect 589000 81334 589600 81418
rect 589000 81098 589182 81334
rect 589418 81098 589600 81334
rect 589000 45654 589600 81098
rect 589000 45418 589182 45654
rect 589418 45418 589600 45654
rect 589000 45334 589600 45418
rect 589000 45098 589182 45334
rect 589418 45098 589600 45334
rect 589000 9654 589600 45098
rect 589000 9418 589182 9654
rect 589418 9418 589600 9654
rect 589000 9334 589600 9418
rect 589000 9098 589182 9334
rect 589418 9098 589600 9334
rect -5676 -4262 -5494 -4026
rect -5258 -4262 -5076 -4026
rect -5676 -4346 -5076 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 -5076 -4346
rect -5676 -4604 -5076 -4582
rect 589000 -4026 589600 9098
rect 589000 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect 589000 -4346 589600 -4262
rect 589000 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect 589000 -4604 589600 -4582
rect 589920 675654 590520 708882
rect 589920 675418 590102 675654
rect 590338 675418 590520 675654
rect 589920 675334 590520 675418
rect 589920 675098 590102 675334
rect 590338 675098 590520 675334
rect 589920 639654 590520 675098
rect 589920 639418 590102 639654
rect 590338 639418 590520 639654
rect 589920 639334 590520 639418
rect 589920 639098 590102 639334
rect 590338 639098 590520 639334
rect 589920 603654 590520 639098
rect 589920 603418 590102 603654
rect 590338 603418 590520 603654
rect 589920 603334 590520 603418
rect 589920 603098 590102 603334
rect 590338 603098 590520 603334
rect 589920 567654 590520 603098
rect 589920 567418 590102 567654
rect 590338 567418 590520 567654
rect 589920 567334 590520 567418
rect 589920 567098 590102 567334
rect 590338 567098 590520 567334
rect 589920 531654 590520 567098
rect 589920 531418 590102 531654
rect 590338 531418 590520 531654
rect 589920 531334 590520 531418
rect 589920 531098 590102 531334
rect 590338 531098 590520 531334
rect 589920 495654 590520 531098
rect 589920 495418 590102 495654
rect 590338 495418 590520 495654
rect 589920 495334 590520 495418
rect 589920 495098 590102 495334
rect 590338 495098 590520 495334
rect 589920 459654 590520 495098
rect 589920 459418 590102 459654
rect 590338 459418 590520 459654
rect 589920 459334 590520 459418
rect 589920 459098 590102 459334
rect 590338 459098 590520 459334
rect 589920 423654 590520 459098
rect 589920 423418 590102 423654
rect 590338 423418 590520 423654
rect 589920 423334 590520 423418
rect 589920 423098 590102 423334
rect 590338 423098 590520 423334
rect 589920 387654 590520 423098
rect 589920 387418 590102 387654
rect 590338 387418 590520 387654
rect 589920 387334 590520 387418
rect 589920 387098 590102 387334
rect 590338 387098 590520 387334
rect 589920 351654 590520 387098
rect 589920 351418 590102 351654
rect 590338 351418 590520 351654
rect 589920 351334 590520 351418
rect 589920 351098 590102 351334
rect 590338 351098 590520 351334
rect 589920 315654 590520 351098
rect 589920 315418 590102 315654
rect 590338 315418 590520 315654
rect 589920 315334 590520 315418
rect 589920 315098 590102 315334
rect 590338 315098 590520 315334
rect 589920 279654 590520 315098
rect 589920 279418 590102 279654
rect 590338 279418 590520 279654
rect 589920 279334 590520 279418
rect 589920 279098 590102 279334
rect 590338 279098 590520 279334
rect 589920 243654 590520 279098
rect 589920 243418 590102 243654
rect 590338 243418 590520 243654
rect 589920 243334 590520 243418
rect 589920 243098 590102 243334
rect 590338 243098 590520 243334
rect 589920 207654 590520 243098
rect 589920 207418 590102 207654
rect 590338 207418 590520 207654
rect 589920 207334 590520 207418
rect 589920 207098 590102 207334
rect 590338 207098 590520 207334
rect 589920 171654 590520 207098
rect 589920 171418 590102 171654
rect 590338 171418 590520 171654
rect 589920 171334 590520 171418
rect 589920 171098 590102 171334
rect 590338 171098 590520 171334
rect 589920 135654 590520 171098
rect 589920 135418 590102 135654
rect 590338 135418 590520 135654
rect 589920 135334 590520 135418
rect 589920 135098 590102 135334
rect 590338 135098 590520 135334
rect 589920 99654 590520 135098
rect 589920 99418 590102 99654
rect 590338 99418 590520 99654
rect 589920 99334 590520 99418
rect 589920 99098 590102 99334
rect 590338 99098 590520 99334
rect 589920 63654 590520 99098
rect 589920 63418 590102 63654
rect 590338 63418 590520 63654
rect 589920 63334 590520 63418
rect 589920 63098 590102 63334
rect 590338 63098 590520 63334
rect 589920 27654 590520 63098
rect 589920 27418 590102 27654
rect 590338 27418 590520 27654
rect 589920 27334 590520 27418
rect 589920 27098 590102 27334
rect 590338 27098 590520 27334
rect -6596 -5182 -6414 -4946
rect -6178 -5182 -5996 -4946
rect -6596 -5266 -5996 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 -5996 -5266
rect -6596 -5524 -5996 -5502
rect 589920 -4946 590520 27098
rect 589920 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect 589920 -5266 590520 -5182
rect 589920 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect 589920 -5524 590520 -5502
rect 590840 697254 591440 709802
rect 590840 697018 591022 697254
rect 591258 697018 591440 697254
rect 590840 696934 591440 697018
rect 590840 696698 591022 696934
rect 591258 696698 591440 696934
rect 590840 661254 591440 696698
rect 590840 661018 591022 661254
rect 591258 661018 591440 661254
rect 590840 660934 591440 661018
rect 590840 660698 591022 660934
rect 591258 660698 591440 660934
rect 590840 625254 591440 660698
rect 590840 625018 591022 625254
rect 591258 625018 591440 625254
rect 590840 624934 591440 625018
rect 590840 624698 591022 624934
rect 591258 624698 591440 624934
rect 590840 589254 591440 624698
rect 590840 589018 591022 589254
rect 591258 589018 591440 589254
rect 590840 588934 591440 589018
rect 590840 588698 591022 588934
rect 591258 588698 591440 588934
rect 590840 553254 591440 588698
rect 590840 553018 591022 553254
rect 591258 553018 591440 553254
rect 590840 552934 591440 553018
rect 590840 552698 591022 552934
rect 591258 552698 591440 552934
rect 590840 517254 591440 552698
rect 590840 517018 591022 517254
rect 591258 517018 591440 517254
rect 590840 516934 591440 517018
rect 590840 516698 591022 516934
rect 591258 516698 591440 516934
rect 590840 481254 591440 516698
rect 590840 481018 591022 481254
rect 591258 481018 591440 481254
rect 590840 480934 591440 481018
rect 590840 480698 591022 480934
rect 591258 480698 591440 480934
rect 590840 445254 591440 480698
rect 590840 445018 591022 445254
rect 591258 445018 591440 445254
rect 590840 444934 591440 445018
rect 590840 444698 591022 444934
rect 591258 444698 591440 444934
rect 590840 409254 591440 444698
rect 590840 409018 591022 409254
rect 591258 409018 591440 409254
rect 590840 408934 591440 409018
rect 590840 408698 591022 408934
rect 591258 408698 591440 408934
rect 590840 373254 591440 408698
rect 590840 373018 591022 373254
rect 591258 373018 591440 373254
rect 590840 372934 591440 373018
rect 590840 372698 591022 372934
rect 591258 372698 591440 372934
rect 590840 337254 591440 372698
rect 590840 337018 591022 337254
rect 591258 337018 591440 337254
rect 590840 336934 591440 337018
rect 590840 336698 591022 336934
rect 591258 336698 591440 336934
rect 590840 301254 591440 336698
rect 590840 301018 591022 301254
rect 591258 301018 591440 301254
rect 590840 300934 591440 301018
rect 590840 300698 591022 300934
rect 591258 300698 591440 300934
rect 590840 265254 591440 300698
rect 590840 265018 591022 265254
rect 591258 265018 591440 265254
rect 590840 264934 591440 265018
rect 590840 264698 591022 264934
rect 591258 264698 591440 264934
rect 590840 229254 591440 264698
rect 590840 229018 591022 229254
rect 591258 229018 591440 229254
rect 590840 228934 591440 229018
rect 590840 228698 591022 228934
rect 591258 228698 591440 228934
rect 590840 193254 591440 228698
rect 590840 193018 591022 193254
rect 591258 193018 591440 193254
rect 590840 192934 591440 193018
rect 590840 192698 591022 192934
rect 591258 192698 591440 192934
rect 590840 157254 591440 192698
rect 590840 157018 591022 157254
rect 591258 157018 591440 157254
rect 590840 156934 591440 157018
rect 590840 156698 591022 156934
rect 591258 156698 591440 156934
rect 590840 121254 591440 156698
rect 590840 121018 591022 121254
rect 591258 121018 591440 121254
rect 590840 120934 591440 121018
rect 590840 120698 591022 120934
rect 591258 120698 591440 120934
rect 590840 85254 591440 120698
rect 590840 85018 591022 85254
rect 591258 85018 591440 85254
rect 590840 84934 591440 85018
rect 590840 84698 591022 84934
rect 591258 84698 591440 84934
rect 590840 49254 591440 84698
rect 590840 49018 591022 49254
rect 591258 49018 591440 49254
rect 590840 48934 591440 49018
rect 590840 48698 591022 48934
rect 591258 48698 591440 48934
rect 590840 13254 591440 48698
rect 590840 13018 591022 13254
rect 591258 13018 591440 13254
rect 590840 12934 591440 13018
rect 590840 12698 591022 12934
rect 591258 12698 591440 12934
rect -7516 -6102 -7334 -5866
rect -7098 -6102 -6916 -5866
rect -7516 -6186 -6916 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 -6916 -6186
rect -7516 -6444 -6916 -6422
rect 590840 -5866 591440 12698
rect 590840 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect 590840 -6186 591440 -6102
rect 590840 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect 590840 -6444 591440 -6422
rect 591760 679254 592360 710722
rect 591760 679018 591942 679254
rect 592178 679018 592360 679254
rect 591760 678934 592360 679018
rect 591760 678698 591942 678934
rect 592178 678698 592360 678934
rect 591760 643254 592360 678698
rect 591760 643018 591942 643254
rect 592178 643018 592360 643254
rect 591760 642934 592360 643018
rect 591760 642698 591942 642934
rect 592178 642698 592360 642934
rect 591760 607254 592360 642698
rect 591760 607018 591942 607254
rect 592178 607018 592360 607254
rect 591760 606934 592360 607018
rect 591760 606698 591942 606934
rect 592178 606698 592360 606934
rect 591760 571254 592360 606698
rect 591760 571018 591942 571254
rect 592178 571018 592360 571254
rect 591760 570934 592360 571018
rect 591760 570698 591942 570934
rect 592178 570698 592360 570934
rect 591760 535254 592360 570698
rect 591760 535018 591942 535254
rect 592178 535018 592360 535254
rect 591760 534934 592360 535018
rect 591760 534698 591942 534934
rect 592178 534698 592360 534934
rect 591760 499254 592360 534698
rect 591760 499018 591942 499254
rect 592178 499018 592360 499254
rect 591760 498934 592360 499018
rect 591760 498698 591942 498934
rect 592178 498698 592360 498934
rect 591760 463254 592360 498698
rect 591760 463018 591942 463254
rect 592178 463018 592360 463254
rect 591760 462934 592360 463018
rect 591760 462698 591942 462934
rect 592178 462698 592360 462934
rect 591760 427254 592360 462698
rect 591760 427018 591942 427254
rect 592178 427018 592360 427254
rect 591760 426934 592360 427018
rect 591760 426698 591942 426934
rect 592178 426698 592360 426934
rect 591760 391254 592360 426698
rect 591760 391018 591942 391254
rect 592178 391018 592360 391254
rect 591760 390934 592360 391018
rect 591760 390698 591942 390934
rect 592178 390698 592360 390934
rect 591760 355254 592360 390698
rect 591760 355018 591942 355254
rect 592178 355018 592360 355254
rect 591760 354934 592360 355018
rect 591760 354698 591942 354934
rect 592178 354698 592360 354934
rect 591760 319254 592360 354698
rect 591760 319018 591942 319254
rect 592178 319018 592360 319254
rect 591760 318934 592360 319018
rect 591760 318698 591942 318934
rect 592178 318698 592360 318934
rect 591760 283254 592360 318698
rect 591760 283018 591942 283254
rect 592178 283018 592360 283254
rect 591760 282934 592360 283018
rect 591760 282698 591942 282934
rect 592178 282698 592360 282934
rect 591760 247254 592360 282698
rect 591760 247018 591942 247254
rect 592178 247018 592360 247254
rect 591760 246934 592360 247018
rect 591760 246698 591942 246934
rect 592178 246698 592360 246934
rect 591760 211254 592360 246698
rect 591760 211018 591942 211254
rect 592178 211018 592360 211254
rect 591760 210934 592360 211018
rect 591760 210698 591942 210934
rect 592178 210698 592360 210934
rect 591760 175254 592360 210698
rect 591760 175018 591942 175254
rect 592178 175018 592360 175254
rect 591760 174934 592360 175018
rect 591760 174698 591942 174934
rect 592178 174698 592360 174934
rect 591760 139254 592360 174698
rect 591760 139018 591942 139254
rect 592178 139018 592360 139254
rect 591760 138934 592360 139018
rect 591760 138698 591942 138934
rect 592178 138698 592360 138934
rect 591760 103254 592360 138698
rect 591760 103018 591942 103254
rect 592178 103018 592360 103254
rect 591760 102934 592360 103018
rect 591760 102698 591942 102934
rect 592178 102698 592360 102934
rect 591760 67254 592360 102698
rect 591760 67018 591942 67254
rect 592178 67018 592360 67254
rect 591760 66934 592360 67018
rect 591760 66698 591942 66934
rect 592178 66698 592360 66934
rect 591760 31254 592360 66698
rect 591760 31018 591942 31254
rect 592178 31018 592360 31254
rect 591760 30934 592360 31018
rect 591760 30698 591942 30934
rect 592178 30698 592360 30934
rect -8436 -7022 -8254 -6786
rect -8018 -7022 -7836 -6786
rect -8436 -7106 -7836 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 -7836 -7106
rect -8436 -7364 -7836 -7342
rect 591760 -6786 592360 30698
rect 591760 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect 591760 -7106 592360 -7022
rect 591760 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect 591760 -7364 592360 -7342
<< via4 >>
rect -8254 711042 -8018 711278
rect -8254 710722 -8018 710958
rect 591942 711042 592178 711278
rect 591942 710722 592178 710958
rect -8254 679018 -8018 679254
rect -8254 678698 -8018 678934
rect -8254 643018 -8018 643254
rect -8254 642698 -8018 642934
rect -8254 607018 -8018 607254
rect -8254 606698 -8018 606934
rect -8254 571018 -8018 571254
rect -8254 570698 -8018 570934
rect -8254 535018 -8018 535254
rect -8254 534698 -8018 534934
rect -8254 499018 -8018 499254
rect -8254 498698 -8018 498934
rect -8254 463018 -8018 463254
rect -8254 462698 -8018 462934
rect -8254 427018 -8018 427254
rect -8254 426698 -8018 426934
rect -8254 391018 -8018 391254
rect -8254 390698 -8018 390934
rect -8254 355018 -8018 355254
rect -8254 354698 -8018 354934
rect -8254 319018 -8018 319254
rect -8254 318698 -8018 318934
rect -8254 283018 -8018 283254
rect -8254 282698 -8018 282934
rect -8254 247018 -8018 247254
rect -8254 246698 -8018 246934
rect -8254 211018 -8018 211254
rect -8254 210698 -8018 210934
rect -8254 175018 -8018 175254
rect -8254 174698 -8018 174934
rect -8254 139018 -8018 139254
rect -8254 138698 -8018 138934
rect -8254 103018 -8018 103254
rect -8254 102698 -8018 102934
rect -8254 67018 -8018 67254
rect -8254 66698 -8018 66934
rect -8254 31018 -8018 31254
rect -8254 30698 -8018 30934
rect -7334 710122 -7098 710358
rect -7334 709802 -7098 710038
rect 591022 710122 591258 710358
rect 591022 709802 591258 710038
rect -7334 697018 -7098 697254
rect -7334 696698 -7098 696934
rect -7334 661018 -7098 661254
rect -7334 660698 -7098 660934
rect -7334 625018 -7098 625254
rect -7334 624698 -7098 624934
rect -7334 589018 -7098 589254
rect -7334 588698 -7098 588934
rect -7334 553018 -7098 553254
rect -7334 552698 -7098 552934
rect -7334 517018 -7098 517254
rect -7334 516698 -7098 516934
rect -7334 481018 -7098 481254
rect -7334 480698 -7098 480934
rect -7334 445018 -7098 445254
rect -7334 444698 -7098 444934
rect -7334 409018 -7098 409254
rect -7334 408698 -7098 408934
rect -7334 373018 -7098 373254
rect -7334 372698 -7098 372934
rect -7334 337018 -7098 337254
rect -7334 336698 -7098 336934
rect -7334 301018 -7098 301254
rect -7334 300698 -7098 300934
rect -7334 265018 -7098 265254
rect -7334 264698 -7098 264934
rect -7334 229018 -7098 229254
rect -7334 228698 -7098 228934
rect -7334 193018 -7098 193254
rect -7334 192698 -7098 192934
rect -7334 157018 -7098 157254
rect -7334 156698 -7098 156934
rect -7334 121018 -7098 121254
rect -7334 120698 -7098 120934
rect -7334 85018 -7098 85254
rect -7334 84698 -7098 84934
rect -7334 49018 -7098 49254
rect -7334 48698 -7098 48934
rect -7334 13018 -7098 13254
rect -7334 12698 -7098 12934
rect -6414 709202 -6178 709438
rect -6414 708882 -6178 709118
rect 590102 709202 590338 709438
rect 590102 708882 590338 709118
rect -6414 675418 -6178 675654
rect -6414 675098 -6178 675334
rect -6414 639418 -6178 639654
rect -6414 639098 -6178 639334
rect -6414 603418 -6178 603654
rect -6414 603098 -6178 603334
rect -6414 567418 -6178 567654
rect -6414 567098 -6178 567334
rect -6414 531418 -6178 531654
rect -6414 531098 -6178 531334
rect -6414 495418 -6178 495654
rect -6414 495098 -6178 495334
rect -6414 459418 -6178 459654
rect -6414 459098 -6178 459334
rect -6414 423418 -6178 423654
rect -6414 423098 -6178 423334
rect -6414 387418 -6178 387654
rect -6414 387098 -6178 387334
rect -6414 351418 -6178 351654
rect -6414 351098 -6178 351334
rect -6414 315418 -6178 315654
rect -6414 315098 -6178 315334
rect -6414 279418 -6178 279654
rect -6414 279098 -6178 279334
rect -6414 243418 -6178 243654
rect -6414 243098 -6178 243334
rect -6414 207418 -6178 207654
rect -6414 207098 -6178 207334
rect -6414 171418 -6178 171654
rect -6414 171098 -6178 171334
rect -6414 135418 -6178 135654
rect -6414 135098 -6178 135334
rect -6414 99418 -6178 99654
rect -6414 99098 -6178 99334
rect -6414 63418 -6178 63654
rect -6414 63098 -6178 63334
rect -6414 27418 -6178 27654
rect -6414 27098 -6178 27334
rect -5494 708282 -5258 708518
rect -5494 707962 -5258 708198
rect 589182 708282 589418 708518
rect 589182 707962 589418 708198
rect -5494 693418 -5258 693654
rect -5494 693098 -5258 693334
rect -5494 657418 -5258 657654
rect -5494 657098 -5258 657334
rect -5494 621418 -5258 621654
rect -5494 621098 -5258 621334
rect -5494 585418 -5258 585654
rect -5494 585098 -5258 585334
rect -5494 549418 -5258 549654
rect -5494 549098 -5258 549334
rect -5494 513418 -5258 513654
rect -5494 513098 -5258 513334
rect -5494 477418 -5258 477654
rect -5494 477098 -5258 477334
rect -5494 441418 -5258 441654
rect -5494 441098 -5258 441334
rect -5494 405418 -5258 405654
rect -5494 405098 -5258 405334
rect -5494 369418 -5258 369654
rect -5494 369098 -5258 369334
rect -5494 333418 -5258 333654
rect -5494 333098 -5258 333334
rect -5494 297418 -5258 297654
rect -5494 297098 -5258 297334
rect -5494 261418 -5258 261654
rect -5494 261098 -5258 261334
rect -5494 225418 -5258 225654
rect -5494 225098 -5258 225334
rect -5494 189418 -5258 189654
rect -5494 189098 -5258 189334
rect -5494 153418 -5258 153654
rect -5494 153098 -5258 153334
rect -5494 117418 -5258 117654
rect -5494 117098 -5258 117334
rect -5494 81418 -5258 81654
rect -5494 81098 -5258 81334
rect -5494 45418 -5258 45654
rect -5494 45098 -5258 45334
rect -5494 9418 -5258 9654
rect -5494 9098 -5258 9334
rect -4574 707362 -4338 707598
rect -4574 707042 -4338 707278
rect 588262 707362 588498 707598
rect 588262 707042 588498 707278
rect -4574 671818 -4338 672054
rect -4574 671498 -4338 671734
rect -4574 635818 -4338 636054
rect -4574 635498 -4338 635734
rect -4574 599818 -4338 600054
rect -4574 599498 -4338 599734
rect -4574 563818 -4338 564054
rect -4574 563498 -4338 563734
rect -4574 527818 -4338 528054
rect -4574 527498 -4338 527734
rect -4574 491818 -4338 492054
rect -4574 491498 -4338 491734
rect -4574 455818 -4338 456054
rect -4574 455498 -4338 455734
rect -4574 419818 -4338 420054
rect -4574 419498 -4338 419734
rect -4574 383818 -4338 384054
rect -4574 383498 -4338 383734
rect -4574 347818 -4338 348054
rect -4574 347498 -4338 347734
rect -4574 311818 -4338 312054
rect -4574 311498 -4338 311734
rect -4574 275818 -4338 276054
rect -4574 275498 -4338 275734
rect -4574 239818 -4338 240054
rect -4574 239498 -4338 239734
rect -4574 203818 -4338 204054
rect -4574 203498 -4338 203734
rect -4574 167818 -4338 168054
rect -4574 167498 -4338 167734
rect -4574 131818 -4338 132054
rect -4574 131498 -4338 131734
rect -4574 95818 -4338 96054
rect -4574 95498 -4338 95734
rect -4574 59818 -4338 60054
rect -4574 59498 -4338 59734
rect -4574 23818 -4338 24054
rect -4574 23498 -4338 23734
rect -3654 706442 -3418 706678
rect -3654 706122 -3418 706358
rect 587342 706442 587578 706678
rect 587342 706122 587578 706358
rect -3654 689818 -3418 690054
rect -3654 689498 -3418 689734
rect -3654 653818 -3418 654054
rect -3654 653498 -3418 653734
rect -3654 617818 -3418 618054
rect -3654 617498 -3418 617734
rect -3654 581818 -3418 582054
rect -3654 581498 -3418 581734
rect -3654 545818 -3418 546054
rect -3654 545498 -3418 545734
rect -3654 509818 -3418 510054
rect -3654 509498 -3418 509734
rect -3654 473818 -3418 474054
rect -3654 473498 -3418 473734
rect -3654 437818 -3418 438054
rect -3654 437498 -3418 437734
rect -3654 401818 -3418 402054
rect -3654 401498 -3418 401734
rect -3654 365818 -3418 366054
rect -3654 365498 -3418 365734
rect -3654 329818 -3418 330054
rect -3654 329498 -3418 329734
rect -3654 293818 -3418 294054
rect -3654 293498 -3418 293734
rect -3654 257818 -3418 258054
rect -3654 257498 -3418 257734
rect -3654 221818 -3418 222054
rect -3654 221498 -3418 221734
rect -3654 185818 -3418 186054
rect -3654 185498 -3418 185734
rect -3654 149818 -3418 150054
rect -3654 149498 -3418 149734
rect -3654 113818 -3418 114054
rect -3654 113498 -3418 113734
rect -3654 77818 -3418 78054
rect -3654 77498 -3418 77734
rect -3654 41818 -3418 42054
rect -3654 41498 -3418 41734
rect -3654 5818 -3418 6054
rect -3654 5498 -3418 5734
rect -2734 705522 -2498 705758
rect -2734 705202 -2498 705438
rect 586422 705522 586658 705758
rect 586422 705202 586658 705438
rect -2734 668218 -2498 668454
rect -2734 667898 -2498 668134
rect -2734 632218 -2498 632454
rect -2734 631898 -2498 632134
rect -2734 596218 -2498 596454
rect -2734 595898 -2498 596134
rect -2734 560218 -2498 560454
rect -2734 559898 -2498 560134
rect -2734 524218 -2498 524454
rect -2734 523898 -2498 524134
rect -2734 488218 -2498 488454
rect -2734 487898 -2498 488134
rect -2734 452218 -2498 452454
rect -2734 451898 -2498 452134
rect -2734 416218 -2498 416454
rect -2734 415898 -2498 416134
rect -2734 380218 -2498 380454
rect -2734 379898 -2498 380134
rect -2734 344218 -2498 344454
rect -2734 343898 -2498 344134
rect -2734 308218 -2498 308454
rect -2734 307898 -2498 308134
rect -2734 272218 -2498 272454
rect -2734 271898 -2498 272134
rect -2734 236218 -2498 236454
rect -2734 235898 -2498 236134
rect -2734 200218 -2498 200454
rect -2734 199898 -2498 200134
rect -2734 164218 -2498 164454
rect -2734 163898 -2498 164134
rect -2734 128218 -2498 128454
rect -2734 127898 -2498 128134
rect -2734 92218 -2498 92454
rect -2734 91898 -2498 92134
rect -2734 56218 -2498 56454
rect -2734 55898 -2498 56134
rect -2734 20218 -2498 20454
rect -2734 19898 -2498 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 344790 680222 345026 680458
rect 558782 676142 559018 676378
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect 559702 676142 559938 676378
rect 559150 665942 559386 666178
rect 560254 665942 560490 666178
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect 1262 36262 1498 36498
rect 894 34222 1130 34458
rect 526 32332 762 32418
rect 526 32268 612 32332
rect 612 32268 676 32332
rect 676 32268 762 32332
rect 526 32182 762 32268
rect 1630 35582 1866 35818
rect 1630 32862 1866 33098
rect 1630 29462 1866 29698
rect 1262 28782 1498 29018
rect 1814 26062 2050 26298
rect 1078 25382 1314 25618
rect 1446 24702 1682 24938
rect 559150 36262 559386 36498
rect 559518 35582 559754 35818
rect 559702 34902 559938 35138
rect 560990 32862 561226 33098
rect 561910 34902 562146 35138
rect 562278 34222 562514 34458
rect 561358 32182 561594 32418
rect 562094 32182 562330 32418
rect 561726 29462 561962 29698
rect 560622 28782 560858 29018
rect 561358 26062 561594 26298
rect 559702 24702 559938 24938
rect 559702 18582 559938 18818
rect 894 15182 1130 15418
rect 1814 13822 2050 14058
rect 1446 10422 1682 10658
rect 526 7852 762 7938
rect 526 7788 612 7852
rect 612 7788 676 7852
rect 676 7788 762 7852
rect 526 7702 762 7788
rect 1262 4452 1498 4538
rect 1262 4388 1348 4452
rect 1348 4388 1412 4452
rect 1412 4388 1498 4452
rect 1262 4302 1498 4388
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect 342 372 578 458
rect 342 308 428 372
rect 428 308 492 372
rect 492 308 578 372
rect 342 222 578 308
rect 558782 15862 559018 16098
rect 4758 13822 4994 14058
rect 20030 13292 20266 13378
rect 20030 13228 20116 13292
rect 20116 13228 20180 13292
rect 20180 13228 20266 13292
rect 20030 13142 20266 13228
rect 4758 11782 4994 12018
rect 558598 11782 558834 12018
rect 558966 11102 559202 11338
rect 559702 11102 559938 11338
rect 19846 7924 19932 7938
rect 19932 7924 19996 7938
rect 19996 7924 20082 7938
rect 19846 7702 20082 7924
rect 4758 7022 4994 7258
rect 225742 6492 225978 6578
rect 225742 6428 225828 6492
rect 225828 6428 225892 6492
rect 225892 6428 225978 6492
rect 225742 6342 225978 6428
rect 225742 5132 225978 5218
rect 225742 5068 225828 5132
rect 225828 5068 225892 5132
rect 225892 5068 225978 5132
rect 225742 4982 225978 5068
rect 124220 3772 124456 3858
rect 124220 3708 124306 3772
rect 124306 3708 124370 3772
rect 124370 3708 124456 3772
rect 124220 3622 124456 3708
rect 177856 3772 178092 3858
rect 177856 3708 177942 3772
rect 177942 3708 178006 3772
rect 178006 3708 178092 3772
rect 177856 3622 178092 3708
rect 268292 3772 268528 3858
rect 268292 3708 268378 3772
rect 268378 3708 268442 3772
rect 268442 3708 268528 3772
rect 268292 3622 268528 3708
rect 14878 2942 15114 3178
rect 28862 2942 29098 3178
rect 52230 2942 52466 3178
rect 74862 2942 75098 3178
rect 76334 2942 76570 3178
rect 78542 2942 78778 3178
rect 82222 2942 82458 3178
rect 91422 2942 91658 3178
rect 94734 2942 94970 3178
rect 95654 2942 95890 3178
rect 96758 2942 96994 3178
rect 102646 2942 102882 3178
rect 125278 2942 125514 3178
rect 4758 902 4994 1138
rect 10462 916 10698 1138
rect 10462 902 10548 916
rect 10548 902 10612 916
rect 10612 902 10698 916
rect 10830 222 11066 458
rect 19110 916 19346 1138
rect 19110 902 19196 916
rect 19196 902 19260 916
rect 19260 902 19346 916
rect 28126 916 28362 1138
rect 28126 902 28212 916
rect 28212 902 28276 916
rect 28276 902 28362 916
rect 38982 902 39218 1138
rect 46710 1052 46946 1138
rect 46710 988 46796 1052
rect 46796 988 46860 1052
rect 46860 988 46946 1052
rect 46710 902 46946 988
rect 28862 222 29098 458
rect 39350 222 39586 458
rect 66766 1124 66852 1138
rect 66852 1124 66916 1138
rect 66916 1124 67002 1138
rect 66766 902 67002 1124
rect 68974 902 69210 1138
rect 73390 222 73626 458
rect 74494 222 74730 458
rect 88110 902 88346 1138
rect 91606 916 91842 1138
rect 91606 902 91692 916
rect 91692 902 91756 916
rect 91756 902 91842 916
rect 92526 222 92762 458
rect 93814 236 94050 458
rect 126014 2942 126250 3178
rect 127118 2942 127354 3178
rect 135766 2942 136002 3178
rect 136502 2942 136738 3178
rect 145886 2942 146122 3178
rect 153614 2942 153850 3178
rect 154350 2942 154586 3178
rect 155270 2942 155506 3178
rect 156006 2942 156242 3178
rect 158030 2942 158266 3178
rect 194094 2942 194330 3178
rect 195566 2942 195802 3178
rect 200902 2942 201138 3178
rect 224086 2942 224322 3178
rect 225006 2942 225242 3178
rect 226846 2942 227082 3178
rect 227766 2942 228002 3178
rect 228686 2942 228922 3178
rect 253342 2942 253578 3178
rect 260150 2942 260386 3178
rect 294374 2942 294610 3178
rect 310014 2942 310250 3178
rect 311118 2942 311354 3178
rect 336694 2942 336930 3178
rect 348838 2942 349074 3178
rect 354174 2942 354410 3178
rect 372436 2942 372672 3178
rect 419310 2942 419546 3178
rect 426854 2942 427090 3178
rect 442862 2942 443098 3178
rect 483710 2942 483946 3178
rect 513150 2942 513386 3178
rect 514438 2942 514674 3178
rect 93814 222 93900 236
rect 93900 222 93964 236
rect 93964 222 94050 236
rect 103750 222 103986 458
rect 104486 222 104722 458
rect 106694 222 106930 458
rect 107430 222 107666 458
rect 126382 1582 126618 1818
rect 127118 1582 127354 1818
rect 123438 222 123674 458
rect 146254 902 146490 1138
rect 134662 222 134898 458
rect 147910 902 148146 1138
rect 150302 902 150538 1138
rect 151452 902 151688 1138
rect 150670 444 150756 458
rect 150756 444 150820 458
rect 150820 444 150906 458
rect 150670 222 150906 444
rect 151406 222 151642 458
rect 154028 1718 154264 1954
rect 158950 1718 159186 1954
rect 159318 902 159554 1138
rect 161526 1396 161612 1410
rect 161612 1396 161676 1410
rect 161676 1396 161762 1410
rect 160054 902 160290 1138
rect 161526 1174 161762 1396
rect 162262 902 162498 1138
rect 194830 2262 195066 2498
rect 225742 2642 225978 2878
rect 163734 222 163970 458
rect 164470 222 164706 458
rect 169070 222 169306 458
rect 169806 222 170042 458
rect 175326 644 175562 730
rect 175326 580 175412 644
rect 175412 580 175476 644
rect 175476 580 175562 644
rect 175326 494 175562 580
rect 176246 222 176482 458
rect 196670 222 196906 458
rect 197774 444 197860 458
rect 197860 444 197924 458
rect 197924 444 198010 458
rect 197774 222 198010 444
rect 223902 1718 224138 1954
rect 226478 1582 226714 1818
rect 217646 222 217882 458
rect 241014 902 241250 1138
rect 242118 902 242354 1138
rect 224638 222 224874 458
rect 232366 222 232602 458
rect 233102 222 233338 458
rect 245614 222 245850 458
rect 254814 902 255050 1138
rect 256286 902 256522 1138
rect 248006 222 248242 458
rect 265118 902 265354 1138
rect 266958 902 267194 1138
rect 264750 222 264986 458
rect 266222 494 266458 730
rect 280022 222 280258 458
rect 281494 222 281730 458
rect 290326 222 290562 458
rect 294742 222 294978 458
rect 326942 1052 327178 1138
rect 326942 988 327028 1052
rect 327028 988 327092 1052
rect 327092 988 327178 1052
rect 326942 902 327178 988
rect 327678 902 327914 1138
rect 338718 902 338954 1138
rect 339454 902 339690 1138
rect 349942 902 350178 1138
rect 353806 902 354042 1138
rect 370366 1124 370452 1138
rect 370452 1124 370516 1138
rect 370516 1124 370602 1138
rect 336694 222 336930 458
rect 370366 902 370602 1124
rect 414526 902 414762 1138
rect 418758 902 418994 1138
rect 343502 222 343738 458
rect 358038 222 358274 458
rect 363006 222 363242 458
rect 413974 222 414210 458
rect 422070 372 422306 458
rect 440102 902 440338 1138
rect 422070 308 422156 372
rect 422156 308 422220 372
rect 422220 308 422306 372
rect 422070 222 422306 308
rect 430534 222 430770 458
rect 434398 222 434634 458
rect 462918 902 463154 1138
rect 449670 222 449906 458
rect 468990 444 469076 458
rect 469076 444 469140 458
rect 469140 444 469226 458
rect 468990 222 469226 444
rect 559334 3622 559570 3858
rect 522166 902 522402 1138
rect 560070 4302 560306 4538
rect 560070 3622 560306 3858
rect 562094 25382 562330 25618
rect 563566 902 563802 1138
rect 564854 680222 565090 680458
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 570190 32182 570426 32418
rect 570190 11102 570426 11338
rect 570374 4452 570610 4538
rect 570374 4388 570460 4452
rect 570460 4388 570524 4452
rect 570524 4388 570610 4452
rect 570374 4302 570610 4388
rect 569454 3622 569690 3858
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 476718 372 476954 458
rect 476718 308 476804 372
rect 476804 308 476868 372
rect 476868 308 476954 372
rect 476718 222 476954 308
rect 490518 372 490754 458
rect 490518 308 490604 372
rect 490604 308 490668 372
rect 490668 308 490754 372
rect 490518 222 490754 308
rect 504318 236 504554 458
rect 504318 222 504404 236
rect 504404 222 504468 236
rect 504468 222 504554 236
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586422 668218 586658 668454
rect 586422 667898 586658 668134
rect 586422 632218 586658 632454
rect 586422 631898 586658 632134
rect 586422 596218 586658 596454
rect 586422 595898 586658 596134
rect 586422 560218 586658 560454
rect 586422 559898 586658 560134
rect 586422 524218 586658 524454
rect 586422 523898 586658 524134
rect 586422 488218 586658 488454
rect 586422 487898 586658 488134
rect 586422 452218 586658 452454
rect 586422 451898 586658 452134
rect 586422 416218 586658 416454
rect 586422 415898 586658 416134
rect 586422 380218 586658 380454
rect 586422 379898 586658 380134
rect 586422 344218 586658 344454
rect 586422 343898 586658 344134
rect 586422 308218 586658 308454
rect 586422 307898 586658 308134
rect 586422 272218 586658 272454
rect 586422 271898 586658 272134
rect 586422 236218 586658 236454
rect 586422 235898 586658 236134
rect 586422 200218 586658 200454
rect 586422 199898 586658 200134
rect 586422 164218 586658 164454
rect 586422 163898 586658 164134
rect 586422 128218 586658 128454
rect 586422 127898 586658 128134
rect 586422 92218 586658 92454
rect 586422 91898 586658 92134
rect 586422 56218 586658 56454
rect 586422 55898 586658 56134
rect 586422 20218 586658 20454
rect 586422 19898 586658 20134
rect -2734 -1502 -2498 -1266
rect -2734 -1822 -2498 -1586
rect 586422 -1502 586658 -1266
rect 586422 -1822 586658 -1586
rect 587342 689818 587578 690054
rect 587342 689498 587578 689734
rect 587342 653818 587578 654054
rect 587342 653498 587578 653734
rect 587342 617818 587578 618054
rect 587342 617498 587578 617734
rect 587342 581818 587578 582054
rect 587342 581498 587578 581734
rect 587342 545818 587578 546054
rect 587342 545498 587578 545734
rect 587342 509818 587578 510054
rect 587342 509498 587578 509734
rect 587342 473818 587578 474054
rect 587342 473498 587578 473734
rect 587342 437818 587578 438054
rect 587342 437498 587578 437734
rect 587342 401818 587578 402054
rect 587342 401498 587578 401734
rect 587342 365818 587578 366054
rect 587342 365498 587578 365734
rect 587342 329818 587578 330054
rect 587342 329498 587578 329734
rect 587342 293818 587578 294054
rect 587342 293498 587578 293734
rect 587342 257818 587578 258054
rect 587342 257498 587578 257734
rect 587342 221818 587578 222054
rect 587342 221498 587578 221734
rect 587342 185818 587578 186054
rect 587342 185498 587578 185734
rect 587342 149818 587578 150054
rect 587342 149498 587578 149734
rect 587342 113818 587578 114054
rect 587342 113498 587578 113734
rect 587342 77818 587578 78054
rect 587342 77498 587578 77734
rect 587342 41818 587578 42054
rect 587342 41498 587578 41734
rect 587342 5818 587578 6054
rect 587342 5498 587578 5734
rect -3654 -2422 -3418 -2186
rect -3654 -2742 -3418 -2506
rect 587342 -2422 587578 -2186
rect 587342 -2742 587578 -2506
rect 588262 671818 588498 672054
rect 588262 671498 588498 671734
rect 588262 635818 588498 636054
rect 588262 635498 588498 635734
rect 588262 599818 588498 600054
rect 588262 599498 588498 599734
rect 588262 563818 588498 564054
rect 588262 563498 588498 563734
rect 588262 527818 588498 528054
rect 588262 527498 588498 527734
rect 588262 491818 588498 492054
rect 588262 491498 588498 491734
rect 588262 455818 588498 456054
rect 588262 455498 588498 455734
rect 588262 419818 588498 420054
rect 588262 419498 588498 419734
rect 588262 383818 588498 384054
rect 588262 383498 588498 383734
rect 588262 347818 588498 348054
rect 588262 347498 588498 347734
rect 588262 311818 588498 312054
rect 588262 311498 588498 311734
rect 588262 275818 588498 276054
rect 588262 275498 588498 275734
rect 588262 239818 588498 240054
rect 588262 239498 588498 239734
rect 588262 203818 588498 204054
rect 588262 203498 588498 203734
rect 588262 167818 588498 168054
rect 588262 167498 588498 167734
rect 588262 131818 588498 132054
rect 588262 131498 588498 131734
rect 588262 95818 588498 96054
rect 588262 95498 588498 95734
rect 588262 59818 588498 60054
rect 588262 59498 588498 59734
rect 588262 23818 588498 24054
rect 588262 23498 588498 23734
rect -4574 -3342 -4338 -3106
rect -4574 -3662 -4338 -3426
rect 588262 -3342 588498 -3106
rect 588262 -3662 588498 -3426
rect 589182 693418 589418 693654
rect 589182 693098 589418 693334
rect 589182 657418 589418 657654
rect 589182 657098 589418 657334
rect 589182 621418 589418 621654
rect 589182 621098 589418 621334
rect 589182 585418 589418 585654
rect 589182 585098 589418 585334
rect 589182 549418 589418 549654
rect 589182 549098 589418 549334
rect 589182 513418 589418 513654
rect 589182 513098 589418 513334
rect 589182 477418 589418 477654
rect 589182 477098 589418 477334
rect 589182 441418 589418 441654
rect 589182 441098 589418 441334
rect 589182 405418 589418 405654
rect 589182 405098 589418 405334
rect 589182 369418 589418 369654
rect 589182 369098 589418 369334
rect 589182 333418 589418 333654
rect 589182 333098 589418 333334
rect 589182 297418 589418 297654
rect 589182 297098 589418 297334
rect 589182 261418 589418 261654
rect 589182 261098 589418 261334
rect 589182 225418 589418 225654
rect 589182 225098 589418 225334
rect 589182 189418 589418 189654
rect 589182 189098 589418 189334
rect 589182 153418 589418 153654
rect 589182 153098 589418 153334
rect 589182 117418 589418 117654
rect 589182 117098 589418 117334
rect 589182 81418 589418 81654
rect 589182 81098 589418 81334
rect 589182 45418 589418 45654
rect 589182 45098 589418 45334
rect 589182 9418 589418 9654
rect 589182 9098 589418 9334
rect -5494 -4262 -5258 -4026
rect -5494 -4582 -5258 -4346
rect 589182 -4262 589418 -4026
rect 589182 -4582 589418 -4346
rect 590102 675418 590338 675654
rect 590102 675098 590338 675334
rect 590102 639418 590338 639654
rect 590102 639098 590338 639334
rect 590102 603418 590338 603654
rect 590102 603098 590338 603334
rect 590102 567418 590338 567654
rect 590102 567098 590338 567334
rect 590102 531418 590338 531654
rect 590102 531098 590338 531334
rect 590102 495418 590338 495654
rect 590102 495098 590338 495334
rect 590102 459418 590338 459654
rect 590102 459098 590338 459334
rect 590102 423418 590338 423654
rect 590102 423098 590338 423334
rect 590102 387418 590338 387654
rect 590102 387098 590338 387334
rect 590102 351418 590338 351654
rect 590102 351098 590338 351334
rect 590102 315418 590338 315654
rect 590102 315098 590338 315334
rect 590102 279418 590338 279654
rect 590102 279098 590338 279334
rect 590102 243418 590338 243654
rect 590102 243098 590338 243334
rect 590102 207418 590338 207654
rect 590102 207098 590338 207334
rect 590102 171418 590338 171654
rect 590102 171098 590338 171334
rect 590102 135418 590338 135654
rect 590102 135098 590338 135334
rect 590102 99418 590338 99654
rect 590102 99098 590338 99334
rect 590102 63418 590338 63654
rect 590102 63098 590338 63334
rect 590102 27418 590338 27654
rect 590102 27098 590338 27334
rect -6414 -5182 -6178 -4946
rect -6414 -5502 -6178 -5266
rect 590102 -5182 590338 -4946
rect 590102 -5502 590338 -5266
rect 591022 697018 591258 697254
rect 591022 696698 591258 696934
rect 591022 661018 591258 661254
rect 591022 660698 591258 660934
rect 591022 625018 591258 625254
rect 591022 624698 591258 624934
rect 591022 589018 591258 589254
rect 591022 588698 591258 588934
rect 591022 553018 591258 553254
rect 591022 552698 591258 552934
rect 591022 517018 591258 517254
rect 591022 516698 591258 516934
rect 591022 481018 591258 481254
rect 591022 480698 591258 480934
rect 591022 445018 591258 445254
rect 591022 444698 591258 444934
rect 591022 409018 591258 409254
rect 591022 408698 591258 408934
rect 591022 373018 591258 373254
rect 591022 372698 591258 372934
rect 591022 337018 591258 337254
rect 591022 336698 591258 336934
rect 591022 301018 591258 301254
rect 591022 300698 591258 300934
rect 591022 265018 591258 265254
rect 591022 264698 591258 264934
rect 591022 229018 591258 229254
rect 591022 228698 591258 228934
rect 591022 193018 591258 193254
rect 591022 192698 591258 192934
rect 591022 157018 591258 157254
rect 591022 156698 591258 156934
rect 591022 121018 591258 121254
rect 591022 120698 591258 120934
rect 591022 85018 591258 85254
rect 591022 84698 591258 84934
rect 591022 49018 591258 49254
rect 591022 48698 591258 48934
rect 591022 13018 591258 13254
rect 591022 12698 591258 12934
rect -7334 -6102 -7098 -5866
rect -7334 -6422 -7098 -6186
rect 591022 -6102 591258 -5866
rect 591022 -6422 591258 -6186
rect 591942 679018 592178 679254
rect 591942 678698 592178 678934
rect 591942 643018 592178 643254
rect 591942 642698 592178 642934
rect 591942 607018 592178 607254
rect 591942 606698 592178 606934
rect 591942 571018 592178 571254
rect 591942 570698 592178 570934
rect 591942 535018 592178 535254
rect 591942 534698 592178 534934
rect 591942 499018 592178 499254
rect 591942 498698 592178 498934
rect 591942 463018 592178 463254
rect 591942 462698 592178 462934
rect 591942 427018 592178 427254
rect 591942 426698 592178 426934
rect 591942 391018 592178 391254
rect 591942 390698 592178 390934
rect 591942 355018 592178 355254
rect 591942 354698 592178 354934
rect 591942 319018 592178 319254
rect 591942 318698 592178 318934
rect 591942 283018 592178 283254
rect 591942 282698 592178 282934
rect 591942 247018 592178 247254
rect 591942 246698 592178 246934
rect 591942 211018 592178 211254
rect 591942 210698 592178 210934
rect 591942 175018 592178 175254
rect 591942 174698 592178 174934
rect 591942 139018 592178 139254
rect 591942 138698 592178 138934
rect 591942 103018 592178 103254
rect 591942 102698 592178 102934
rect 591942 67018 592178 67254
rect 591942 66698 592178 66934
rect 591942 31018 592178 31254
rect 591942 30698 592178 30934
rect -8254 -7022 -8018 -6786
rect -8254 -7342 -8018 -7106
rect 591942 -7022 592178 -6786
rect 591942 -7342 592178 -7106
<< metal5 >>
rect -8436 711300 -7836 711302
rect 591760 711300 592360 711302
rect -8436 711278 592360 711300
rect -8436 711042 -8254 711278
rect -8018 711042 591942 711278
rect 592178 711042 592360 711278
rect -8436 710958 592360 711042
rect -8436 710722 -8254 710958
rect -8018 710722 591942 710958
rect 592178 710722 592360 710958
rect -8436 710700 592360 710722
rect -8436 710698 -7836 710700
rect 591760 710698 592360 710700
rect -7516 710380 -6916 710382
rect 590840 710380 591440 710382
rect -7516 710358 591440 710380
rect -7516 710122 -7334 710358
rect -7098 710122 591022 710358
rect 591258 710122 591440 710358
rect -7516 710038 591440 710122
rect -7516 709802 -7334 710038
rect -7098 709802 591022 710038
rect 591258 709802 591440 710038
rect -7516 709780 591440 709802
rect -7516 709778 -6916 709780
rect 590840 709778 591440 709780
rect -6596 709460 -5996 709462
rect 589920 709460 590520 709462
rect -6596 709438 590520 709460
rect -6596 709202 -6414 709438
rect -6178 709202 590102 709438
rect 590338 709202 590520 709438
rect -6596 709118 590520 709202
rect -6596 708882 -6414 709118
rect -6178 708882 590102 709118
rect 590338 708882 590520 709118
rect -6596 708860 590520 708882
rect -6596 708858 -5996 708860
rect 589920 708858 590520 708860
rect -5676 708540 -5076 708542
rect 589000 708540 589600 708542
rect -5676 708518 589600 708540
rect -5676 708282 -5494 708518
rect -5258 708282 589182 708518
rect 589418 708282 589600 708518
rect -5676 708198 589600 708282
rect -5676 707962 -5494 708198
rect -5258 707962 589182 708198
rect 589418 707962 589600 708198
rect -5676 707940 589600 707962
rect -5676 707938 -5076 707940
rect 589000 707938 589600 707940
rect -4756 707620 -4156 707622
rect 588080 707620 588680 707622
rect -4756 707598 588680 707620
rect -4756 707362 -4574 707598
rect -4338 707362 588262 707598
rect 588498 707362 588680 707598
rect -4756 707278 588680 707362
rect -4756 707042 -4574 707278
rect -4338 707042 588262 707278
rect 588498 707042 588680 707278
rect -4756 707020 588680 707042
rect -4756 707018 -4156 707020
rect 588080 707018 588680 707020
rect -3836 706700 -3236 706702
rect 587160 706700 587760 706702
rect -3836 706678 587760 706700
rect -3836 706442 -3654 706678
rect -3418 706442 587342 706678
rect 587578 706442 587760 706678
rect -3836 706358 587760 706442
rect -3836 706122 -3654 706358
rect -3418 706122 587342 706358
rect 587578 706122 587760 706358
rect -3836 706100 587760 706122
rect -3836 706098 -3236 706100
rect 587160 706098 587760 706100
rect -2916 705780 -2316 705782
rect 586240 705780 586840 705782
rect -2916 705758 586840 705780
rect -2916 705522 -2734 705758
rect -2498 705522 586422 705758
rect 586658 705522 586840 705758
rect -2916 705438 586840 705522
rect -2916 705202 -2734 705438
rect -2498 705202 586422 705438
rect 586658 705202 586840 705438
rect -2916 705180 586840 705202
rect -2916 705178 -2316 705180
rect 586240 705178 586840 705180
rect -1996 704860 -1396 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 585320 704258 585920 704260
rect -7516 697276 -6916 697278
rect 590840 697276 591440 697278
rect -8436 697254 592360 697276
rect -8436 697018 -7334 697254
rect -7098 697018 591022 697254
rect 591258 697018 592360 697254
rect -8436 696934 592360 697018
rect -8436 696698 -7334 696934
rect -7098 696698 591022 696934
rect 591258 696698 592360 696934
rect -8436 696676 592360 696698
rect -7516 696674 -6916 696676
rect 590840 696674 591440 696676
rect -5676 693676 -5076 693678
rect 589000 693676 589600 693678
rect -6596 693654 590520 693676
rect -6596 693418 -5494 693654
rect -5258 693418 589182 693654
rect 589418 693418 590520 693654
rect -6596 693334 590520 693418
rect -6596 693098 -5494 693334
rect -5258 693098 589182 693334
rect 589418 693098 590520 693334
rect -6596 693076 590520 693098
rect -5676 693074 -5076 693076
rect 589000 693074 589600 693076
rect -3836 690076 -3236 690078
rect 587160 690076 587760 690078
rect -4756 690054 588680 690076
rect -4756 689818 -3654 690054
rect -3418 689818 587342 690054
rect 587578 689818 588680 690054
rect -4756 689734 588680 689818
rect -4756 689498 -3654 689734
rect -3418 689498 587342 689734
rect 587578 689498 588680 689734
rect -4756 689476 588680 689498
rect -3836 689474 -3236 689476
rect 587160 689474 587760 689476
rect -1996 686476 -1396 686478
rect 585320 686476 585920 686478
rect -2916 686454 586840 686476
rect -2916 686218 -1814 686454
rect -1578 686218 585502 686454
rect 585738 686218 586840 686454
rect -2916 686134 586840 686218
rect -2916 685898 -1814 686134
rect -1578 685898 585502 686134
rect 585738 685898 586840 686134
rect -2916 685876 586840 685898
rect -1996 685874 -1396 685876
rect 585320 685874 585920 685876
rect 364252 681540 370092 681860
rect 364252 680500 364572 681540
rect 369772 681180 370092 681540
rect 466188 681540 467244 681860
rect 466188 681180 466508 681540
rect 369772 680860 379476 681180
rect 344748 680458 364572 680500
rect 344748 680222 344790 680458
rect 345026 680222 364572 680458
rect 344748 680180 364572 680222
rect 379156 680500 379476 680860
rect 456620 680860 466508 681180
rect 466924 681180 467244 681540
rect 475940 681540 486564 681860
rect 475940 681180 476260 681540
rect 466924 680860 476260 681180
rect 486244 681180 486564 681540
rect 495260 681540 505700 681860
rect 495260 681180 495580 681540
rect 486244 680860 495580 681180
rect 505380 681180 505700 681540
rect 505380 680860 514716 681180
rect 456620 680500 456940 680860
rect 379156 680180 456940 680500
rect 514396 680500 514716 680860
rect 514396 680458 565132 680500
rect 514396 680222 564854 680458
rect 565090 680222 565132 680458
rect 514396 680180 565132 680222
rect -8436 679276 -7836 679278
rect 591760 679276 592360 679278
rect -8436 679254 592360 679276
rect -8436 679018 -8254 679254
rect -8018 679018 591942 679254
rect 592178 679018 592360 679254
rect -8436 678934 592360 679018
rect -8436 678698 -8254 678934
rect -8018 678698 591942 678934
rect 592178 678698 592360 678934
rect -8436 678676 592360 678698
rect -8436 678674 -7836 678676
rect 591760 678674 592360 678676
rect 558740 676378 559980 676420
rect 558740 676142 558782 676378
rect 559018 676142 559702 676378
rect 559938 676142 559980 676378
rect 558740 676100 559980 676142
rect -6596 675676 -5996 675678
rect 589920 675676 590520 675678
rect -6596 675654 590520 675676
rect -6596 675418 -6414 675654
rect -6178 675418 590102 675654
rect 590338 675418 590520 675654
rect -6596 675334 590520 675418
rect -6596 675098 -6414 675334
rect -6178 675098 590102 675334
rect 590338 675098 590520 675334
rect -6596 675076 590520 675098
rect -6596 675074 -5996 675076
rect 589920 675074 590520 675076
rect -4756 672076 -4156 672078
rect 588080 672076 588680 672078
rect -4756 672054 588680 672076
rect -4756 671818 -4574 672054
rect -4338 671818 588262 672054
rect 588498 671818 588680 672054
rect -4756 671734 588680 671818
rect -4756 671498 -4574 671734
rect -4338 671498 588262 671734
rect 588498 671498 588680 671734
rect -4756 671476 588680 671498
rect -4756 671474 -4156 671476
rect 588080 671474 588680 671476
rect -2916 668476 -2316 668478
rect 586240 668476 586840 668478
rect -2916 668454 586840 668476
rect -2916 668218 -2734 668454
rect -2498 668218 586422 668454
rect 586658 668218 586840 668454
rect -2916 668134 586840 668218
rect -2916 667898 -2734 668134
rect -2498 667898 586422 668134
rect 586658 667898 586840 668134
rect -2916 667876 586840 667898
rect -2916 667874 -2316 667876
rect 586240 667874 586840 667876
rect 559108 666178 560532 666220
rect 559108 665942 559150 666178
rect 559386 665942 560254 666178
rect 560490 665942 560532 666178
rect 559108 665900 560532 665942
rect -7516 661276 -6916 661278
rect 590840 661276 591440 661278
rect -8436 661254 592360 661276
rect -8436 661018 -7334 661254
rect -7098 661018 591022 661254
rect 591258 661018 592360 661254
rect -8436 660934 592360 661018
rect -8436 660698 -7334 660934
rect -7098 660698 591022 660934
rect 591258 660698 592360 660934
rect -8436 660676 592360 660698
rect -7516 660674 -6916 660676
rect 590840 660674 591440 660676
rect -5676 657676 -5076 657678
rect 589000 657676 589600 657678
rect -6596 657654 590520 657676
rect -6596 657418 -5494 657654
rect -5258 657418 589182 657654
rect 589418 657418 590520 657654
rect -6596 657334 590520 657418
rect -6596 657098 -5494 657334
rect -5258 657098 589182 657334
rect 589418 657098 590520 657334
rect -6596 657076 590520 657098
rect -5676 657074 -5076 657076
rect 589000 657074 589600 657076
rect -3836 654076 -3236 654078
rect 587160 654076 587760 654078
rect -4756 654054 588680 654076
rect -4756 653818 -3654 654054
rect -3418 653818 587342 654054
rect 587578 653818 588680 654054
rect -4756 653734 588680 653818
rect -4756 653498 -3654 653734
rect -3418 653498 587342 653734
rect 587578 653498 588680 653734
rect -4756 653476 588680 653498
rect -3836 653474 -3236 653476
rect 587160 653474 587760 653476
rect -1996 650476 -1396 650478
rect 585320 650476 585920 650478
rect -2916 650454 586840 650476
rect -2916 650218 -1814 650454
rect -1578 650218 585502 650454
rect 585738 650218 586840 650454
rect -2916 650134 586840 650218
rect -2916 649898 -1814 650134
rect -1578 649898 585502 650134
rect 585738 649898 586840 650134
rect -2916 649876 586840 649898
rect -1996 649874 -1396 649876
rect 585320 649874 585920 649876
rect -8436 643276 -7836 643278
rect 591760 643276 592360 643278
rect -8436 643254 592360 643276
rect -8436 643018 -8254 643254
rect -8018 643018 591942 643254
rect 592178 643018 592360 643254
rect -8436 642934 592360 643018
rect -8436 642698 -8254 642934
rect -8018 642698 591942 642934
rect 592178 642698 592360 642934
rect -8436 642676 592360 642698
rect -8436 642674 -7836 642676
rect 591760 642674 592360 642676
rect -6596 639676 -5996 639678
rect 589920 639676 590520 639678
rect -6596 639654 590520 639676
rect -6596 639418 -6414 639654
rect -6178 639418 590102 639654
rect 590338 639418 590520 639654
rect -6596 639334 590520 639418
rect -6596 639098 -6414 639334
rect -6178 639098 590102 639334
rect 590338 639098 590520 639334
rect -6596 639076 590520 639098
rect -6596 639074 -5996 639076
rect 589920 639074 590520 639076
rect -4756 636076 -4156 636078
rect 588080 636076 588680 636078
rect -4756 636054 588680 636076
rect -4756 635818 -4574 636054
rect -4338 635818 588262 636054
rect 588498 635818 588680 636054
rect -4756 635734 588680 635818
rect -4756 635498 -4574 635734
rect -4338 635498 588262 635734
rect 588498 635498 588680 635734
rect -4756 635476 588680 635498
rect -4756 635474 -4156 635476
rect 588080 635474 588680 635476
rect -2916 632476 -2316 632478
rect 586240 632476 586840 632478
rect -2916 632454 586840 632476
rect -2916 632218 -2734 632454
rect -2498 632218 586422 632454
rect 586658 632218 586840 632454
rect -2916 632134 586840 632218
rect -2916 631898 -2734 632134
rect -2498 631898 586422 632134
rect 586658 631898 586840 632134
rect -2916 631876 586840 631898
rect -2916 631874 -2316 631876
rect 586240 631874 586840 631876
rect -7516 625276 -6916 625278
rect 590840 625276 591440 625278
rect -8436 625254 592360 625276
rect -8436 625018 -7334 625254
rect -7098 625018 591022 625254
rect 591258 625018 592360 625254
rect -8436 624934 592360 625018
rect -8436 624698 -7334 624934
rect -7098 624698 591022 624934
rect 591258 624698 592360 624934
rect -8436 624676 592360 624698
rect -7516 624674 -6916 624676
rect 590840 624674 591440 624676
rect -5676 621676 -5076 621678
rect 589000 621676 589600 621678
rect -6596 621654 590520 621676
rect -6596 621418 -5494 621654
rect -5258 621418 589182 621654
rect 589418 621418 590520 621654
rect -6596 621334 590520 621418
rect -6596 621098 -5494 621334
rect -5258 621098 589182 621334
rect 589418 621098 590520 621334
rect -6596 621076 590520 621098
rect -5676 621074 -5076 621076
rect 589000 621074 589600 621076
rect -3836 618076 -3236 618078
rect 587160 618076 587760 618078
rect -4756 618054 588680 618076
rect -4756 617818 -3654 618054
rect -3418 617818 587342 618054
rect 587578 617818 588680 618054
rect -4756 617734 588680 617818
rect -4756 617498 -3654 617734
rect -3418 617498 587342 617734
rect 587578 617498 588680 617734
rect -4756 617476 588680 617498
rect -3836 617474 -3236 617476
rect 587160 617474 587760 617476
rect -1996 614476 -1396 614478
rect 585320 614476 585920 614478
rect -2916 614454 586840 614476
rect -2916 614218 -1814 614454
rect -1578 614218 585502 614454
rect 585738 614218 586840 614454
rect -2916 614134 586840 614218
rect -2916 613898 -1814 614134
rect -1578 613898 585502 614134
rect 585738 613898 586840 614134
rect -2916 613876 586840 613898
rect -1996 613874 -1396 613876
rect 585320 613874 585920 613876
rect -8436 607276 -7836 607278
rect 591760 607276 592360 607278
rect -8436 607254 592360 607276
rect -8436 607018 -8254 607254
rect -8018 607018 591942 607254
rect 592178 607018 592360 607254
rect -8436 606934 592360 607018
rect -8436 606698 -8254 606934
rect -8018 606698 591942 606934
rect 592178 606698 592360 606934
rect -8436 606676 592360 606698
rect -8436 606674 -7836 606676
rect 591760 606674 592360 606676
rect -6596 603676 -5996 603678
rect 589920 603676 590520 603678
rect -6596 603654 590520 603676
rect -6596 603418 -6414 603654
rect -6178 603418 590102 603654
rect 590338 603418 590520 603654
rect -6596 603334 590520 603418
rect -6596 603098 -6414 603334
rect -6178 603098 590102 603334
rect 590338 603098 590520 603334
rect -6596 603076 590520 603098
rect -6596 603074 -5996 603076
rect 589920 603074 590520 603076
rect -4756 600076 -4156 600078
rect 588080 600076 588680 600078
rect -4756 600054 588680 600076
rect -4756 599818 -4574 600054
rect -4338 599818 588262 600054
rect 588498 599818 588680 600054
rect -4756 599734 588680 599818
rect -4756 599498 -4574 599734
rect -4338 599498 588262 599734
rect 588498 599498 588680 599734
rect -4756 599476 588680 599498
rect -4756 599474 -4156 599476
rect 588080 599474 588680 599476
rect -2916 596476 -2316 596478
rect 586240 596476 586840 596478
rect -2916 596454 586840 596476
rect -2916 596218 -2734 596454
rect -2498 596218 586422 596454
rect 586658 596218 586840 596454
rect -2916 596134 586840 596218
rect -2916 595898 -2734 596134
rect -2498 595898 586422 596134
rect 586658 595898 586840 596134
rect -2916 595876 586840 595898
rect -2916 595874 -2316 595876
rect 586240 595874 586840 595876
rect -7516 589276 -6916 589278
rect 590840 589276 591440 589278
rect -8436 589254 592360 589276
rect -8436 589018 -7334 589254
rect -7098 589018 591022 589254
rect 591258 589018 592360 589254
rect -8436 588934 592360 589018
rect -8436 588698 -7334 588934
rect -7098 588698 591022 588934
rect 591258 588698 592360 588934
rect -8436 588676 592360 588698
rect -7516 588674 -6916 588676
rect 590840 588674 591440 588676
rect -5676 585676 -5076 585678
rect 589000 585676 589600 585678
rect -6596 585654 590520 585676
rect -6596 585418 -5494 585654
rect -5258 585418 589182 585654
rect 589418 585418 590520 585654
rect -6596 585334 590520 585418
rect -6596 585098 -5494 585334
rect -5258 585098 589182 585334
rect 589418 585098 590520 585334
rect -6596 585076 590520 585098
rect -5676 585074 -5076 585076
rect 589000 585074 589600 585076
rect -3836 582076 -3236 582078
rect 587160 582076 587760 582078
rect -4756 582054 588680 582076
rect -4756 581818 -3654 582054
rect -3418 581818 587342 582054
rect 587578 581818 588680 582054
rect -4756 581734 588680 581818
rect -4756 581498 -3654 581734
rect -3418 581498 587342 581734
rect 587578 581498 588680 581734
rect -4756 581476 588680 581498
rect -3836 581474 -3236 581476
rect 587160 581474 587760 581476
rect -1996 578476 -1396 578478
rect 585320 578476 585920 578478
rect -2916 578454 586840 578476
rect -2916 578218 -1814 578454
rect -1578 578218 585502 578454
rect 585738 578218 586840 578454
rect -2916 578134 586840 578218
rect -2916 577898 -1814 578134
rect -1578 577898 585502 578134
rect 585738 577898 586840 578134
rect -2916 577876 586840 577898
rect -1996 577874 -1396 577876
rect 585320 577874 585920 577876
rect -8436 571276 -7836 571278
rect 591760 571276 592360 571278
rect -8436 571254 592360 571276
rect -8436 571018 -8254 571254
rect -8018 571018 591942 571254
rect 592178 571018 592360 571254
rect -8436 570934 592360 571018
rect -8436 570698 -8254 570934
rect -8018 570698 591942 570934
rect 592178 570698 592360 570934
rect -8436 570676 592360 570698
rect -8436 570674 -7836 570676
rect 591760 570674 592360 570676
rect -6596 567676 -5996 567678
rect 589920 567676 590520 567678
rect -6596 567654 590520 567676
rect -6596 567418 -6414 567654
rect -6178 567418 590102 567654
rect 590338 567418 590520 567654
rect -6596 567334 590520 567418
rect -6596 567098 -6414 567334
rect -6178 567098 590102 567334
rect 590338 567098 590520 567334
rect -6596 567076 590520 567098
rect -6596 567074 -5996 567076
rect 589920 567074 590520 567076
rect -4756 564076 -4156 564078
rect 588080 564076 588680 564078
rect -4756 564054 588680 564076
rect -4756 563818 -4574 564054
rect -4338 563818 588262 564054
rect 588498 563818 588680 564054
rect -4756 563734 588680 563818
rect -4756 563498 -4574 563734
rect -4338 563498 588262 563734
rect 588498 563498 588680 563734
rect -4756 563476 588680 563498
rect -4756 563474 -4156 563476
rect 588080 563474 588680 563476
rect -2916 560476 -2316 560478
rect 586240 560476 586840 560478
rect -2916 560454 586840 560476
rect -2916 560218 -2734 560454
rect -2498 560218 586422 560454
rect 586658 560218 586840 560454
rect -2916 560134 586840 560218
rect -2916 559898 -2734 560134
rect -2498 559898 586422 560134
rect 586658 559898 586840 560134
rect -2916 559876 586840 559898
rect -2916 559874 -2316 559876
rect 586240 559874 586840 559876
rect -7516 553276 -6916 553278
rect 590840 553276 591440 553278
rect -8436 553254 592360 553276
rect -8436 553018 -7334 553254
rect -7098 553018 591022 553254
rect 591258 553018 592360 553254
rect -8436 552934 592360 553018
rect -8436 552698 -7334 552934
rect -7098 552698 591022 552934
rect 591258 552698 592360 552934
rect -8436 552676 592360 552698
rect -7516 552674 -6916 552676
rect 590840 552674 591440 552676
rect -5676 549676 -5076 549678
rect 589000 549676 589600 549678
rect -6596 549654 590520 549676
rect -6596 549418 -5494 549654
rect -5258 549418 589182 549654
rect 589418 549418 590520 549654
rect -6596 549334 590520 549418
rect -6596 549098 -5494 549334
rect -5258 549098 589182 549334
rect 589418 549098 590520 549334
rect -6596 549076 590520 549098
rect -5676 549074 -5076 549076
rect 589000 549074 589600 549076
rect -3836 546076 -3236 546078
rect 587160 546076 587760 546078
rect -4756 546054 588680 546076
rect -4756 545818 -3654 546054
rect -3418 545818 587342 546054
rect 587578 545818 588680 546054
rect -4756 545734 588680 545818
rect -4756 545498 -3654 545734
rect -3418 545498 587342 545734
rect 587578 545498 588680 545734
rect -4756 545476 588680 545498
rect -3836 545474 -3236 545476
rect 587160 545474 587760 545476
rect -1996 542476 -1396 542478
rect 585320 542476 585920 542478
rect -2916 542454 586840 542476
rect -2916 542218 -1814 542454
rect -1578 542218 585502 542454
rect 585738 542218 586840 542454
rect -2916 542134 586840 542218
rect -2916 541898 -1814 542134
rect -1578 541898 585502 542134
rect 585738 541898 586840 542134
rect -2916 541876 586840 541898
rect -1996 541874 -1396 541876
rect 585320 541874 585920 541876
rect -8436 535276 -7836 535278
rect 591760 535276 592360 535278
rect -8436 535254 592360 535276
rect -8436 535018 -8254 535254
rect -8018 535018 591942 535254
rect 592178 535018 592360 535254
rect -8436 534934 592360 535018
rect -8436 534698 -8254 534934
rect -8018 534698 591942 534934
rect 592178 534698 592360 534934
rect -8436 534676 592360 534698
rect -8436 534674 -7836 534676
rect 591760 534674 592360 534676
rect -6596 531676 -5996 531678
rect 589920 531676 590520 531678
rect -6596 531654 590520 531676
rect -6596 531418 -6414 531654
rect -6178 531418 590102 531654
rect 590338 531418 590520 531654
rect -6596 531334 590520 531418
rect -6596 531098 -6414 531334
rect -6178 531098 590102 531334
rect 590338 531098 590520 531334
rect -6596 531076 590520 531098
rect -6596 531074 -5996 531076
rect 589920 531074 590520 531076
rect -4756 528076 -4156 528078
rect 588080 528076 588680 528078
rect -4756 528054 588680 528076
rect -4756 527818 -4574 528054
rect -4338 527818 588262 528054
rect 588498 527818 588680 528054
rect -4756 527734 588680 527818
rect -4756 527498 -4574 527734
rect -4338 527498 588262 527734
rect 588498 527498 588680 527734
rect -4756 527476 588680 527498
rect -4756 527474 -4156 527476
rect 588080 527474 588680 527476
rect -2916 524476 -2316 524478
rect 586240 524476 586840 524478
rect -2916 524454 586840 524476
rect -2916 524218 -2734 524454
rect -2498 524218 586422 524454
rect 586658 524218 586840 524454
rect -2916 524134 586840 524218
rect -2916 523898 -2734 524134
rect -2498 523898 586422 524134
rect 586658 523898 586840 524134
rect -2916 523876 586840 523898
rect -2916 523874 -2316 523876
rect 586240 523874 586840 523876
rect -7516 517276 -6916 517278
rect 590840 517276 591440 517278
rect -8436 517254 592360 517276
rect -8436 517018 -7334 517254
rect -7098 517018 591022 517254
rect 591258 517018 592360 517254
rect -8436 516934 592360 517018
rect -8436 516698 -7334 516934
rect -7098 516698 591022 516934
rect 591258 516698 592360 516934
rect -8436 516676 592360 516698
rect -7516 516674 -6916 516676
rect 590840 516674 591440 516676
rect -5676 513676 -5076 513678
rect 589000 513676 589600 513678
rect -6596 513654 590520 513676
rect -6596 513418 -5494 513654
rect -5258 513418 589182 513654
rect 589418 513418 590520 513654
rect -6596 513334 590520 513418
rect -6596 513098 -5494 513334
rect -5258 513098 589182 513334
rect 589418 513098 590520 513334
rect -6596 513076 590520 513098
rect -5676 513074 -5076 513076
rect 589000 513074 589600 513076
rect -3836 510076 -3236 510078
rect 587160 510076 587760 510078
rect -4756 510054 588680 510076
rect -4756 509818 -3654 510054
rect -3418 509818 587342 510054
rect 587578 509818 588680 510054
rect -4756 509734 588680 509818
rect -4756 509498 -3654 509734
rect -3418 509498 587342 509734
rect 587578 509498 588680 509734
rect -4756 509476 588680 509498
rect -3836 509474 -3236 509476
rect 587160 509474 587760 509476
rect -1996 506476 -1396 506478
rect 585320 506476 585920 506478
rect -2916 506454 586840 506476
rect -2916 506218 -1814 506454
rect -1578 506218 585502 506454
rect 585738 506218 586840 506454
rect -2916 506134 586840 506218
rect -2916 505898 -1814 506134
rect -1578 505898 585502 506134
rect 585738 505898 586840 506134
rect -2916 505876 586840 505898
rect -1996 505874 -1396 505876
rect 585320 505874 585920 505876
rect -8436 499276 -7836 499278
rect 591760 499276 592360 499278
rect -8436 499254 592360 499276
rect -8436 499018 -8254 499254
rect -8018 499018 591942 499254
rect 592178 499018 592360 499254
rect -8436 498934 592360 499018
rect -8436 498698 -8254 498934
rect -8018 498698 591942 498934
rect 592178 498698 592360 498934
rect -8436 498676 592360 498698
rect -8436 498674 -7836 498676
rect 591760 498674 592360 498676
rect -6596 495676 -5996 495678
rect 589920 495676 590520 495678
rect -6596 495654 590520 495676
rect -6596 495418 -6414 495654
rect -6178 495418 590102 495654
rect 590338 495418 590520 495654
rect -6596 495334 590520 495418
rect -6596 495098 -6414 495334
rect -6178 495098 590102 495334
rect 590338 495098 590520 495334
rect -6596 495076 590520 495098
rect -6596 495074 -5996 495076
rect 589920 495074 590520 495076
rect -4756 492076 -4156 492078
rect 588080 492076 588680 492078
rect -4756 492054 588680 492076
rect -4756 491818 -4574 492054
rect -4338 491818 588262 492054
rect 588498 491818 588680 492054
rect -4756 491734 588680 491818
rect -4756 491498 -4574 491734
rect -4338 491498 588262 491734
rect 588498 491498 588680 491734
rect -4756 491476 588680 491498
rect -4756 491474 -4156 491476
rect 588080 491474 588680 491476
rect -2916 488476 -2316 488478
rect 586240 488476 586840 488478
rect -2916 488454 586840 488476
rect -2916 488218 -2734 488454
rect -2498 488218 586422 488454
rect 586658 488218 586840 488454
rect -2916 488134 586840 488218
rect -2916 487898 -2734 488134
rect -2498 487898 586422 488134
rect 586658 487898 586840 488134
rect -2916 487876 586840 487898
rect -2916 487874 -2316 487876
rect 586240 487874 586840 487876
rect -7516 481276 -6916 481278
rect 590840 481276 591440 481278
rect -8436 481254 592360 481276
rect -8436 481018 -7334 481254
rect -7098 481018 591022 481254
rect 591258 481018 592360 481254
rect -8436 480934 592360 481018
rect -8436 480698 -7334 480934
rect -7098 480698 591022 480934
rect 591258 480698 592360 480934
rect -8436 480676 592360 480698
rect -7516 480674 -6916 480676
rect 590840 480674 591440 480676
rect -5676 477676 -5076 477678
rect 589000 477676 589600 477678
rect -6596 477654 590520 477676
rect -6596 477418 -5494 477654
rect -5258 477418 589182 477654
rect 589418 477418 590520 477654
rect -6596 477334 590520 477418
rect -6596 477098 -5494 477334
rect -5258 477098 589182 477334
rect 589418 477098 590520 477334
rect -6596 477076 590520 477098
rect -5676 477074 -5076 477076
rect 589000 477074 589600 477076
rect -3836 474076 -3236 474078
rect 587160 474076 587760 474078
rect -4756 474054 588680 474076
rect -4756 473818 -3654 474054
rect -3418 473818 587342 474054
rect 587578 473818 588680 474054
rect -4756 473734 588680 473818
rect -4756 473498 -3654 473734
rect -3418 473498 587342 473734
rect 587578 473498 588680 473734
rect -4756 473476 588680 473498
rect -3836 473474 -3236 473476
rect 587160 473474 587760 473476
rect -1996 470476 -1396 470478
rect 585320 470476 585920 470478
rect -2916 470454 586840 470476
rect -2916 470218 -1814 470454
rect -1578 470218 585502 470454
rect 585738 470218 586840 470454
rect -2916 470134 586840 470218
rect -2916 469898 -1814 470134
rect -1578 469898 585502 470134
rect 585738 469898 586840 470134
rect -2916 469876 586840 469898
rect -1996 469874 -1396 469876
rect 585320 469874 585920 469876
rect -8436 463276 -7836 463278
rect 591760 463276 592360 463278
rect -8436 463254 592360 463276
rect -8436 463018 -8254 463254
rect -8018 463018 591942 463254
rect 592178 463018 592360 463254
rect -8436 462934 592360 463018
rect -8436 462698 -8254 462934
rect -8018 462698 591942 462934
rect 592178 462698 592360 462934
rect -8436 462676 592360 462698
rect -8436 462674 -7836 462676
rect 591760 462674 592360 462676
rect -6596 459676 -5996 459678
rect 589920 459676 590520 459678
rect -6596 459654 590520 459676
rect -6596 459418 -6414 459654
rect -6178 459418 590102 459654
rect 590338 459418 590520 459654
rect -6596 459334 590520 459418
rect -6596 459098 -6414 459334
rect -6178 459098 590102 459334
rect 590338 459098 590520 459334
rect -6596 459076 590520 459098
rect -6596 459074 -5996 459076
rect 589920 459074 590520 459076
rect -4756 456076 -4156 456078
rect 588080 456076 588680 456078
rect -4756 456054 588680 456076
rect -4756 455818 -4574 456054
rect -4338 455818 588262 456054
rect 588498 455818 588680 456054
rect -4756 455734 588680 455818
rect -4756 455498 -4574 455734
rect -4338 455498 588262 455734
rect 588498 455498 588680 455734
rect -4756 455476 588680 455498
rect -4756 455474 -4156 455476
rect 588080 455474 588680 455476
rect -2916 452476 -2316 452478
rect 586240 452476 586840 452478
rect -2916 452454 586840 452476
rect -2916 452218 -2734 452454
rect -2498 452218 586422 452454
rect 586658 452218 586840 452454
rect -2916 452134 586840 452218
rect -2916 451898 -2734 452134
rect -2498 451898 586422 452134
rect 586658 451898 586840 452134
rect -2916 451876 586840 451898
rect -2916 451874 -2316 451876
rect 586240 451874 586840 451876
rect -7516 445276 -6916 445278
rect 590840 445276 591440 445278
rect -8436 445254 592360 445276
rect -8436 445018 -7334 445254
rect -7098 445018 591022 445254
rect 591258 445018 592360 445254
rect -8436 444934 592360 445018
rect -8436 444698 -7334 444934
rect -7098 444698 591022 444934
rect 591258 444698 592360 444934
rect -8436 444676 592360 444698
rect -7516 444674 -6916 444676
rect 590840 444674 591440 444676
rect -5676 441676 -5076 441678
rect 589000 441676 589600 441678
rect -6596 441654 590520 441676
rect -6596 441418 -5494 441654
rect -5258 441418 589182 441654
rect 589418 441418 590520 441654
rect -6596 441334 590520 441418
rect -6596 441098 -5494 441334
rect -5258 441098 589182 441334
rect 589418 441098 590520 441334
rect -6596 441076 590520 441098
rect -5676 441074 -5076 441076
rect 589000 441074 589600 441076
rect -3836 438076 -3236 438078
rect 587160 438076 587760 438078
rect -4756 438054 588680 438076
rect -4756 437818 -3654 438054
rect -3418 437818 587342 438054
rect 587578 437818 588680 438054
rect -4756 437734 588680 437818
rect -4756 437498 -3654 437734
rect -3418 437498 587342 437734
rect 587578 437498 588680 437734
rect -4756 437476 588680 437498
rect -3836 437474 -3236 437476
rect 587160 437474 587760 437476
rect -1996 434476 -1396 434478
rect 585320 434476 585920 434478
rect -2916 434454 586840 434476
rect -2916 434218 -1814 434454
rect -1578 434218 585502 434454
rect 585738 434218 586840 434454
rect -2916 434134 586840 434218
rect -2916 433898 -1814 434134
rect -1578 433898 585502 434134
rect 585738 433898 586840 434134
rect -2916 433876 586840 433898
rect -1996 433874 -1396 433876
rect 585320 433874 585920 433876
rect -8436 427276 -7836 427278
rect 591760 427276 592360 427278
rect -8436 427254 592360 427276
rect -8436 427018 -8254 427254
rect -8018 427018 591942 427254
rect 592178 427018 592360 427254
rect -8436 426934 592360 427018
rect -8436 426698 -8254 426934
rect -8018 426698 591942 426934
rect 592178 426698 592360 426934
rect -8436 426676 592360 426698
rect -8436 426674 -7836 426676
rect 591760 426674 592360 426676
rect -6596 423676 -5996 423678
rect 589920 423676 590520 423678
rect -6596 423654 590520 423676
rect -6596 423418 -6414 423654
rect -6178 423418 590102 423654
rect 590338 423418 590520 423654
rect -6596 423334 590520 423418
rect -6596 423098 -6414 423334
rect -6178 423098 590102 423334
rect 590338 423098 590520 423334
rect -6596 423076 590520 423098
rect -6596 423074 -5996 423076
rect 589920 423074 590520 423076
rect -4756 420076 -4156 420078
rect 588080 420076 588680 420078
rect -4756 420054 588680 420076
rect -4756 419818 -4574 420054
rect -4338 419818 588262 420054
rect 588498 419818 588680 420054
rect -4756 419734 588680 419818
rect -4756 419498 -4574 419734
rect -4338 419498 588262 419734
rect 588498 419498 588680 419734
rect -4756 419476 588680 419498
rect -4756 419474 -4156 419476
rect 588080 419474 588680 419476
rect -2916 416476 -2316 416478
rect 586240 416476 586840 416478
rect -2916 416454 586840 416476
rect -2916 416218 -2734 416454
rect -2498 416218 586422 416454
rect 586658 416218 586840 416454
rect -2916 416134 586840 416218
rect -2916 415898 -2734 416134
rect -2498 415898 586422 416134
rect 586658 415898 586840 416134
rect -2916 415876 586840 415898
rect -2916 415874 -2316 415876
rect 586240 415874 586840 415876
rect -7516 409276 -6916 409278
rect 590840 409276 591440 409278
rect -8436 409254 592360 409276
rect -8436 409018 -7334 409254
rect -7098 409018 591022 409254
rect 591258 409018 592360 409254
rect -8436 408934 592360 409018
rect -8436 408698 -7334 408934
rect -7098 408698 591022 408934
rect 591258 408698 592360 408934
rect -8436 408676 592360 408698
rect -7516 408674 -6916 408676
rect 590840 408674 591440 408676
rect -5676 405676 -5076 405678
rect 589000 405676 589600 405678
rect -6596 405654 590520 405676
rect -6596 405418 -5494 405654
rect -5258 405418 589182 405654
rect 589418 405418 590520 405654
rect -6596 405334 590520 405418
rect -6596 405098 -5494 405334
rect -5258 405098 589182 405334
rect 589418 405098 590520 405334
rect -6596 405076 590520 405098
rect -5676 405074 -5076 405076
rect 589000 405074 589600 405076
rect -3836 402076 -3236 402078
rect 587160 402076 587760 402078
rect -4756 402054 588680 402076
rect -4756 401818 -3654 402054
rect -3418 401818 587342 402054
rect 587578 401818 588680 402054
rect -4756 401734 588680 401818
rect -4756 401498 -3654 401734
rect -3418 401498 587342 401734
rect 587578 401498 588680 401734
rect -4756 401476 588680 401498
rect -3836 401474 -3236 401476
rect 587160 401474 587760 401476
rect -1996 398476 -1396 398478
rect 585320 398476 585920 398478
rect -2916 398454 586840 398476
rect -2916 398218 -1814 398454
rect -1578 398218 585502 398454
rect 585738 398218 586840 398454
rect -2916 398134 586840 398218
rect -2916 397898 -1814 398134
rect -1578 397898 585502 398134
rect 585738 397898 586840 398134
rect -2916 397876 586840 397898
rect -1996 397874 -1396 397876
rect 585320 397874 585920 397876
rect -8436 391276 -7836 391278
rect 591760 391276 592360 391278
rect -8436 391254 592360 391276
rect -8436 391018 -8254 391254
rect -8018 391018 591942 391254
rect 592178 391018 592360 391254
rect -8436 390934 592360 391018
rect -8436 390698 -8254 390934
rect -8018 390698 591942 390934
rect 592178 390698 592360 390934
rect -8436 390676 592360 390698
rect -8436 390674 -7836 390676
rect 591760 390674 592360 390676
rect -6596 387676 -5996 387678
rect 589920 387676 590520 387678
rect -6596 387654 590520 387676
rect -6596 387418 -6414 387654
rect -6178 387418 590102 387654
rect 590338 387418 590520 387654
rect -6596 387334 590520 387418
rect -6596 387098 -6414 387334
rect -6178 387098 590102 387334
rect 590338 387098 590520 387334
rect -6596 387076 590520 387098
rect -6596 387074 -5996 387076
rect 589920 387074 590520 387076
rect -4756 384076 -4156 384078
rect 588080 384076 588680 384078
rect -4756 384054 588680 384076
rect -4756 383818 -4574 384054
rect -4338 383818 588262 384054
rect 588498 383818 588680 384054
rect -4756 383734 588680 383818
rect -4756 383498 -4574 383734
rect -4338 383498 588262 383734
rect 588498 383498 588680 383734
rect -4756 383476 588680 383498
rect -4756 383474 -4156 383476
rect 588080 383474 588680 383476
rect -2916 380476 -2316 380478
rect 586240 380476 586840 380478
rect -2916 380454 586840 380476
rect -2916 380218 -2734 380454
rect -2498 380218 586422 380454
rect 586658 380218 586840 380454
rect -2916 380134 586840 380218
rect -2916 379898 -2734 380134
rect -2498 379898 586422 380134
rect 586658 379898 586840 380134
rect -2916 379876 586840 379898
rect -2916 379874 -2316 379876
rect 586240 379874 586840 379876
rect -7516 373276 -6916 373278
rect 590840 373276 591440 373278
rect -8436 373254 592360 373276
rect -8436 373018 -7334 373254
rect -7098 373018 591022 373254
rect 591258 373018 592360 373254
rect -8436 372934 592360 373018
rect -8436 372698 -7334 372934
rect -7098 372698 591022 372934
rect 591258 372698 592360 372934
rect -8436 372676 592360 372698
rect -7516 372674 -6916 372676
rect 590840 372674 591440 372676
rect -5676 369676 -5076 369678
rect 589000 369676 589600 369678
rect -6596 369654 590520 369676
rect -6596 369418 -5494 369654
rect -5258 369418 589182 369654
rect 589418 369418 590520 369654
rect -6596 369334 590520 369418
rect -6596 369098 -5494 369334
rect -5258 369098 589182 369334
rect 589418 369098 590520 369334
rect -6596 369076 590520 369098
rect -5676 369074 -5076 369076
rect 589000 369074 589600 369076
rect -3836 366076 -3236 366078
rect 587160 366076 587760 366078
rect -4756 366054 588680 366076
rect -4756 365818 -3654 366054
rect -3418 365818 587342 366054
rect 587578 365818 588680 366054
rect -4756 365734 588680 365818
rect -4756 365498 -3654 365734
rect -3418 365498 587342 365734
rect 587578 365498 588680 365734
rect -4756 365476 588680 365498
rect -3836 365474 -3236 365476
rect 587160 365474 587760 365476
rect -1996 362476 -1396 362478
rect 585320 362476 585920 362478
rect -2916 362454 586840 362476
rect -2916 362218 -1814 362454
rect -1578 362218 585502 362454
rect 585738 362218 586840 362454
rect -2916 362134 586840 362218
rect -2916 361898 -1814 362134
rect -1578 361898 585502 362134
rect 585738 361898 586840 362134
rect -2916 361876 586840 361898
rect -1996 361874 -1396 361876
rect 585320 361874 585920 361876
rect -8436 355276 -7836 355278
rect 591760 355276 592360 355278
rect -8436 355254 592360 355276
rect -8436 355018 -8254 355254
rect -8018 355018 591942 355254
rect 592178 355018 592360 355254
rect -8436 354934 592360 355018
rect -8436 354698 -8254 354934
rect -8018 354698 591942 354934
rect 592178 354698 592360 354934
rect -8436 354676 592360 354698
rect -8436 354674 -7836 354676
rect 591760 354674 592360 354676
rect -6596 351676 -5996 351678
rect 589920 351676 590520 351678
rect -6596 351654 590520 351676
rect -6596 351418 -6414 351654
rect -6178 351418 590102 351654
rect 590338 351418 590520 351654
rect -6596 351334 590520 351418
rect -6596 351098 -6414 351334
rect -6178 351098 590102 351334
rect 590338 351098 590520 351334
rect -6596 351076 590520 351098
rect -6596 351074 -5996 351076
rect 589920 351074 590520 351076
rect -4756 348076 -4156 348078
rect 588080 348076 588680 348078
rect -4756 348054 588680 348076
rect -4756 347818 -4574 348054
rect -4338 347818 588262 348054
rect 588498 347818 588680 348054
rect -4756 347734 588680 347818
rect -4756 347498 -4574 347734
rect -4338 347498 588262 347734
rect 588498 347498 588680 347734
rect -4756 347476 588680 347498
rect -4756 347474 -4156 347476
rect 588080 347474 588680 347476
rect -2916 344476 -2316 344478
rect 586240 344476 586840 344478
rect -2916 344454 586840 344476
rect -2916 344218 -2734 344454
rect -2498 344218 586422 344454
rect 586658 344218 586840 344454
rect -2916 344134 586840 344218
rect -2916 343898 -2734 344134
rect -2498 343898 586422 344134
rect 586658 343898 586840 344134
rect -2916 343876 586840 343898
rect -2916 343874 -2316 343876
rect 586240 343874 586840 343876
rect -7516 337276 -6916 337278
rect 590840 337276 591440 337278
rect -8436 337254 592360 337276
rect -8436 337018 -7334 337254
rect -7098 337018 591022 337254
rect 591258 337018 592360 337254
rect -8436 336934 592360 337018
rect -8436 336698 -7334 336934
rect -7098 336698 591022 336934
rect 591258 336698 592360 336934
rect -8436 336676 592360 336698
rect -7516 336674 -6916 336676
rect 590840 336674 591440 336676
rect -5676 333676 -5076 333678
rect 589000 333676 589600 333678
rect -6596 333654 590520 333676
rect -6596 333418 -5494 333654
rect -5258 333418 589182 333654
rect 589418 333418 590520 333654
rect -6596 333334 590520 333418
rect -6596 333098 -5494 333334
rect -5258 333098 589182 333334
rect 589418 333098 590520 333334
rect -6596 333076 590520 333098
rect -5676 333074 -5076 333076
rect 589000 333074 589600 333076
rect -3836 330076 -3236 330078
rect 587160 330076 587760 330078
rect -4756 330054 588680 330076
rect -4756 329818 -3654 330054
rect -3418 329818 587342 330054
rect 587578 329818 588680 330054
rect -4756 329734 588680 329818
rect -4756 329498 -3654 329734
rect -3418 329498 587342 329734
rect 587578 329498 588680 329734
rect -4756 329476 588680 329498
rect -3836 329474 -3236 329476
rect 587160 329474 587760 329476
rect -1996 326476 -1396 326478
rect 585320 326476 585920 326478
rect -2916 326454 586840 326476
rect -2916 326218 -1814 326454
rect -1578 326218 585502 326454
rect 585738 326218 586840 326454
rect -2916 326134 586840 326218
rect -2916 325898 -1814 326134
rect -1578 325898 585502 326134
rect 585738 325898 586840 326134
rect -2916 325876 586840 325898
rect -1996 325874 -1396 325876
rect 585320 325874 585920 325876
rect -8436 319276 -7836 319278
rect 591760 319276 592360 319278
rect -8436 319254 592360 319276
rect -8436 319018 -8254 319254
rect -8018 319018 591942 319254
rect 592178 319018 592360 319254
rect -8436 318934 592360 319018
rect -8436 318698 -8254 318934
rect -8018 318698 591942 318934
rect 592178 318698 592360 318934
rect -8436 318676 592360 318698
rect -8436 318674 -7836 318676
rect 591760 318674 592360 318676
rect -6596 315676 -5996 315678
rect 589920 315676 590520 315678
rect -6596 315654 590520 315676
rect -6596 315418 -6414 315654
rect -6178 315418 590102 315654
rect 590338 315418 590520 315654
rect -6596 315334 590520 315418
rect -6596 315098 -6414 315334
rect -6178 315098 590102 315334
rect 590338 315098 590520 315334
rect -6596 315076 590520 315098
rect -6596 315074 -5996 315076
rect 589920 315074 590520 315076
rect -4756 312076 -4156 312078
rect 588080 312076 588680 312078
rect -4756 312054 588680 312076
rect -4756 311818 -4574 312054
rect -4338 311818 588262 312054
rect 588498 311818 588680 312054
rect -4756 311734 588680 311818
rect -4756 311498 -4574 311734
rect -4338 311498 588262 311734
rect 588498 311498 588680 311734
rect -4756 311476 588680 311498
rect -4756 311474 -4156 311476
rect 588080 311474 588680 311476
rect -2916 308476 -2316 308478
rect 586240 308476 586840 308478
rect -2916 308454 586840 308476
rect -2916 308218 -2734 308454
rect -2498 308218 586422 308454
rect 586658 308218 586840 308454
rect -2916 308134 586840 308218
rect -2916 307898 -2734 308134
rect -2498 307898 586422 308134
rect 586658 307898 586840 308134
rect -2916 307876 586840 307898
rect -2916 307874 -2316 307876
rect 586240 307874 586840 307876
rect -7516 301276 -6916 301278
rect 590840 301276 591440 301278
rect -8436 301254 592360 301276
rect -8436 301018 -7334 301254
rect -7098 301018 591022 301254
rect 591258 301018 592360 301254
rect -8436 300934 592360 301018
rect -8436 300698 -7334 300934
rect -7098 300698 591022 300934
rect 591258 300698 592360 300934
rect -8436 300676 592360 300698
rect -7516 300674 -6916 300676
rect 590840 300674 591440 300676
rect -5676 297676 -5076 297678
rect 589000 297676 589600 297678
rect -6596 297654 590520 297676
rect -6596 297418 -5494 297654
rect -5258 297418 589182 297654
rect 589418 297418 590520 297654
rect -6596 297334 590520 297418
rect -6596 297098 -5494 297334
rect -5258 297098 589182 297334
rect 589418 297098 590520 297334
rect -6596 297076 590520 297098
rect -5676 297074 -5076 297076
rect 589000 297074 589600 297076
rect -3836 294076 -3236 294078
rect 587160 294076 587760 294078
rect -4756 294054 588680 294076
rect -4756 293818 -3654 294054
rect -3418 293818 587342 294054
rect 587578 293818 588680 294054
rect -4756 293734 588680 293818
rect -4756 293498 -3654 293734
rect -3418 293498 587342 293734
rect 587578 293498 588680 293734
rect -4756 293476 588680 293498
rect -3836 293474 -3236 293476
rect 587160 293474 587760 293476
rect -1996 290476 -1396 290478
rect 585320 290476 585920 290478
rect -2916 290454 586840 290476
rect -2916 290218 -1814 290454
rect -1578 290218 585502 290454
rect 585738 290218 586840 290454
rect -2916 290134 586840 290218
rect -2916 289898 -1814 290134
rect -1578 289898 585502 290134
rect 585738 289898 586840 290134
rect -2916 289876 586840 289898
rect -1996 289874 -1396 289876
rect 585320 289874 585920 289876
rect -8436 283276 -7836 283278
rect 591760 283276 592360 283278
rect -8436 283254 592360 283276
rect -8436 283018 -8254 283254
rect -8018 283018 591942 283254
rect 592178 283018 592360 283254
rect -8436 282934 592360 283018
rect -8436 282698 -8254 282934
rect -8018 282698 591942 282934
rect 592178 282698 592360 282934
rect -8436 282676 592360 282698
rect -8436 282674 -7836 282676
rect 591760 282674 592360 282676
rect -6596 279676 -5996 279678
rect 589920 279676 590520 279678
rect -6596 279654 590520 279676
rect -6596 279418 -6414 279654
rect -6178 279418 590102 279654
rect 590338 279418 590520 279654
rect -6596 279334 590520 279418
rect -6596 279098 -6414 279334
rect -6178 279098 590102 279334
rect 590338 279098 590520 279334
rect -6596 279076 590520 279098
rect -6596 279074 -5996 279076
rect 589920 279074 590520 279076
rect -4756 276076 -4156 276078
rect 588080 276076 588680 276078
rect -4756 276054 588680 276076
rect -4756 275818 -4574 276054
rect -4338 275818 588262 276054
rect 588498 275818 588680 276054
rect -4756 275734 588680 275818
rect -4756 275498 -4574 275734
rect -4338 275498 588262 275734
rect 588498 275498 588680 275734
rect -4756 275476 588680 275498
rect -4756 275474 -4156 275476
rect 588080 275474 588680 275476
rect -2916 272476 -2316 272478
rect 586240 272476 586840 272478
rect -2916 272454 586840 272476
rect -2916 272218 -2734 272454
rect -2498 272218 586422 272454
rect 586658 272218 586840 272454
rect -2916 272134 586840 272218
rect -2916 271898 -2734 272134
rect -2498 271898 586422 272134
rect 586658 271898 586840 272134
rect -2916 271876 586840 271898
rect -2916 271874 -2316 271876
rect 586240 271874 586840 271876
rect -7516 265276 -6916 265278
rect 590840 265276 591440 265278
rect -8436 265254 592360 265276
rect -8436 265018 -7334 265254
rect -7098 265018 591022 265254
rect 591258 265018 592360 265254
rect -8436 264934 592360 265018
rect -8436 264698 -7334 264934
rect -7098 264698 591022 264934
rect 591258 264698 592360 264934
rect -8436 264676 592360 264698
rect -7516 264674 -6916 264676
rect 590840 264674 591440 264676
rect -5676 261676 -5076 261678
rect 589000 261676 589600 261678
rect -6596 261654 590520 261676
rect -6596 261418 -5494 261654
rect -5258 261418 589182 261654
rect 589418 261418 590520 261654
rect -6596 261334 590520 261418
rect -6596 261098 -5494 261334
rect -5258 261098 589182 261334
rect 589418 261098 590520 261334
rect -6596 261076 590520 261098
rect -5676 261074 -5076 261076
rect 589000 261074 589600 261076
rect -3836 258076 -3236 258078
rect 587160 258076 587760 258078
rect -4756 258054 588680 258076
rect -4756 257818 -3654 258054
rect -3418 257818 587342 258054
rect 587578 257818 588680 258054
rect -4756 257734 588680 257818
rect -4756 257498 -3654 257734
rect -3418 257498 587342 257734
rect 587578 257498 588680 257734
rect -4756 257476 588680 257498
rect -3836 257474 -3236 257476
rect 587160 257474 587760 257476
rect -1996 254476 -1396 254478
rect 585320 254476 585920 254478
rect -2916 254454 586840 254476
rect -2916 254218 -1814 254454
rect -1578 254218 585502 254454
rect 585738 254218 586840 254454
rect -2916 254134 586840 254218
rect -2916 253898 -1814 254134
rect -1578 253898 585502 254134
rect 585738 253898 586840 254134
rect -2916 253876 586840 253898
rect -1996 253874 -1396 253876
rect 585320 253874 585920 253876
rect -8436 247276 -7836 247278
rect 591760 247276 592360 247278
rect -8436 247254 592360 247276
rect -8436 247018 -8254 247254
rect -8018 247018 591942 247254
rect 592178 247018 592360 247254
rect -8436 246934 592360 247018
rect -8436 246698 -8254 246934
rect -8018 246698 591942 246934
rect 592178 246698 592360 246934
rect -8436 246676 592360 246698
rect -8436 246674 -7836 246676
rect 591760 246674 592360 246676
rect -6596 243676 -5996 243678
rect 589920 243676 590520 243678
rect -6596 243654 590520 243676
rect -6596 243418 -6414 243654
rect -6178 243418 590102 243654
rect 590338 243418 590520 243654
rect -6596 243334 590520 243418
rect -6596 243098 -6414 243334
rect -6178 243098 590102 243334
rect 590338 243098 590520 243334
rect -6596 243076 590520 243098
rect -6596 243074 -5996 243076
rect 589920 243074 590520 243076
rect -4756 240076 -4156 240078
rect 588080 240076 588680 240078
rect -4756 240054 588680 240076
rect -4756 239818 -4574 240054
rect -4338 239818 588262 240054
rect 588498 239818 588680 240054
rect -4756 239734 588680 239818
rect -4756 239498 -4574 239734
rect -4338 239498 588262 239734
rect 588498 239498 588680 239734
rect -4756 239476 588680 239498
rect -4756 239474 -4156 239476
rect 588080 239474 588680 239476
rect -2916 236476 -2316 236478
rect 586240 236476 586840 236478
rect -2916 236454 586840 236476
rect -2916 236218 -2734 236454
rect -2498 236218 586422 236454
rect 586658 236218 586840 236454
rect -2916 236134 586840 236218
rect -2916 235898 -2734 236134
rect -2498 235898 586422 236134
rect 586658 235898 586840 236134
rect -2916 235876 586840 235898
rect -2916 235874 -2316 235876
rect 586240 235874 586840 235876
rect -7516 229276 -6916 229278
rect 590840 229276 591440 229278
rect -8436 229254 592360 229276
rect -8436 229018 -7334 229254
rect -7098 229018 591022 229254
rect 591258 229018 592360 229254
rect -8436 228934 592360 229018
rect -8436 228698 -7334 228934
rect -7098 228698 591022 228934
rect 591258 228698 592360 228934
rect -8436 228676 592360 228698
rect -7516 228674 -6916 228676
rect 590840 228674 591440 228676
rect -5676 225676 -5076 225678
rect 589000 225676 589600 225678
rect -6596 225654 590520 225676
rect -6596 225418 -5494 225654
rect -5258 225418 589182 225654
rect 589418 225418 590520 225654
rect -6596 225334 590520 225418
rect -6596 225098 -5494 225334
rect -5258 225098 589182 225334
rect 589418 225098 590520 225334
rect -6596 225076 590520 225098
rect -5676 225074 -5076 225076
rect 589000 225074 589600 225076
rect -3836 222076 -3236 222078
rect 587160 222076 587760 222078
rect -4756 222054 588680 222076
rect -4756 221818 -3654 222054
rect -3418 221818 587342 222054
rect 587578 221818 588680 222054
rect -4756 221734 588680 221818
rect -4756 221498 -3654 221734
rect -3418 221498 587342 221734
rect 587578 221498 588680 221734
rect -4756 221476 588680 221498
rect -3836 221474 -3236 221476
rect 587160 221474 587760 221476
rect -1996 218476 -1396 218478
rect 585320 218476 585920 218478
rect -2916 218454 586840 218476
rect -2916 218218 -1814 218454
rect -1578 218218 585502 218454
rect 585738 218218 586840 218454
rect -2916 218134 586840 218218
rect -2916 217898 -1814 218134
rect -1578 217898 585502 218134
rect 585738 217898 586840 218134
rect -2916 217876 586840 217898
rect -1996 217874 -1396 217876
rect 585320 217874 585920 217876
rect -8436 211276 -7836 211278
rect 591760 211276 592360 211278
rect -8436 211254 592360 211276
rect -8436 211018 -8254 211254
rect -8018 211018 591942 211254
rect 592178 211018 592360 211254
rect -8436 210934 592360 211018
rect -8436 210698 -8254 210934
rect -8018 210698 591942 210934
rect 592178 210698 592360 210934
rect -8436 210676 592360 210698
rect -8436 210674 -7836 210676
rect 591760 210674 592360 210676
rect -6596 207676 -5996 207678
rect 589920 207676 590520 207678
rect -6596 207654 590520 207676
rect -6596 207418 -6414 207654
rect -6178 207418 590102 207654
rect 590338 207418 590520 207654
rect -6596 207334 590520 207418
rect -6596 207098 -6414 207334
rect -6178 207098 590102 207334
rect 590338 207098 590520 207334
rect -6596 207076 590520 207098
rect -6596 207074 -5996 207076
rect 589920 207074 590520 207076
rect -4756 204076 -4156 204078
rect 588080 204076 588680 204078
rect -4756 204054 588680 204076
rect -4756 203818 -4574 204054
rect -4338 203818 588262 204054
rect 588498 203818 588680 204054
rect -4756 203734 588680 203818
rect -4756 203498 -4574 203734
rect -4338 203498 588262 203734
rect 588498 203498 588680 203734
rect -4756 203476 588680 203498
rect -4756 203474 -4156 203476
rect 588080 203474 588680 203476
rect -2916 200476 -2316 200478
rect 586240 200476 586840 200478
rect -2916 200454 586840 200476
rect -2916 200218 -2734 200454
rect -2498 200218 586422 200454
rect 586658 200218 586840 200454
rect -2916 200134 586840 200218
rect -2916 199898 -2734 200134
rect -2498 199898 586422 200134
rect 586658 199898 586840 200134
rect -2916 199876 586840 199898
rect -2916 199874 -2316 199876
rect 586240 199874 586840 199876
rect -7516 193276 -6916 193278
rect 590840 193276 591440 193278
rect -8436 193254 592360 193276
rect -8436 193018 -7334 193254
rect -7098 193018 591022 193254
rect 591258 193018 592360 193254
rect -8436 192934 592360 193018
rect -8436 192698 -7334 192934
rect -7098 192698 591022 192934
rect 591258 192698 592360 192934
rect -8436 192676 592360 192698
rect -7516 192674 -6916 192676
rect 590840 192674 591440 192676
rect -5676 189676 -5076 189678
rect 589000 189676 589600 189678
rect -6596 189654 590520 189676
rect -6596 189418 -5494 189654
rect -5258 189418 589182 189654
rect 589418 189418 590520 189654
rect -6596 189334 590520 189418
rect -6596 189098 -5494 189334
rect -5258 189098 589182 189334
rect 589418 189098 590520 189334
rect -6596 189076 590520 189098
rect -5676 189074 -5076 189076
rect 589000 189074 589600 189076
rect -3836 186076 -3236 186078
rect 587160 186076 587760 186078
rect -4756 186054 588680 186076
rect -4756 185818 -3654 186054
rect -3418 185818 587342 186054
rect 587578 185818 588680 186054
rect -4756 185734 588680 185818
rect -4756 185498 -3654 185734
rect -3418 185498 587342 185734
rect 587578 185498 588680 185734
rect -4756 185476 588680 185498
rect -3836 185474 -3236 185476
rect 587160 185474 587760 185476
rect -1996 182476 -1396 182478
rect 585320 182476 585920 182478
rect -2916 182454 586840 182476
rect -2916 182218 -1814 182454
rect -1578 182218 585502 182454
rect 585738 182218 586840 182454
rect -2916 182134 586840 182218
rect -2916 181898 -1814 182134
rect -1578 181898 585502 182134
rect 585738 181898 586840 182134
rect -2916 181876 586840 181898
rect -1996 181874 -1396 181876
rect 585320 181874 585920 181876
rect -8436 175276 -7836 175278
rect 591760 175276 592360 175278
rect -8436 175254 592360 175276
rect -8436 175018 -8254 175254
rect -8018 175018 591942 175254
rect 592178 175018 592360 175254
rect -8436 174934 592360 175018
rect -8436 174698 -8254 174934
rect -8018 174698 591942 174934
rect 592178 174698 592360 174934
rect -8436 174676 592360 174698
rect -8436 174674 -7836 174676
rect 591760 174674 592360 174676
rect -6596 171676 -5996 171678
rect 589920 171676 590520 171678
rect -6596 171654 590520 171676
rect -6596 171418 -6414 171654
rect -6178 171418 590102 171654
rect 590338 171418 590520 171654
rect -6596 171334 590520 171418
rect -6596 171098 -6414 171334
rect -6178 171098 590102 171334
rect 590338 171098 590520 171334
rect -6596 171076 590520 171098
rect -6596 171074 -5996 171076
rect 589920 171074 590520 171076
rect -4756 168076 -4156 168078
rect 588080 168076 588680 168078
rect -4756 168054 588680 168076
rect -4756 167818 -4574 168054
rect -4338 167818 588262 168054
rect 588498 167818 588680 168054
rect -4756 167734 588680 167818
rect -4756 167498 -4574 167734
rect -4338 167498 588262 167734
rect 588498 167498 588680 167734
rect -4756 167476 588680 167498
rect -4756 167474 -4156 167476
rect 588080 167474 588680 167476
rect -2916 164476 -2316 164478
rect 586240 164476 586840 164478
rect -2916 164454 586840 164476
rect -2916 164218 -2734 164454
rect -2498 164218 586422 164454
rect 586658 164218 586840 164454
rect -2916 164134 586840 164218
rect -2916 163898 -2734 164134
rect -2498 163898 586422 164134
rect 586658 163898 586840 164134
rect -2916 163876 586840 163898
rect -2916 163874 -2316 163876
rect 586240 163874 586840 163876
rect -7516 157276 -6916 157278
rect 590840 157276 591440 157278
rect -8436 157254 592360 157276
rect -8436 157018 -7334 157254
rect -7098 157018 591022 157254
rect 591258 157018 592360 157254
rect -8436 156934 592360 157018
rect -8436 156698 -7334 156934
rect -7098 156698 591022 156934
rect 591258 156698 592360 156934
rect -8436 156676 592360 156698
rect -7516 156674 -6916 156676
rect 590840 156674 591440 156676
rect -5676 153676 -5076 153678
rect 589000 153676 589600 153678
rect -6596 153654 590520 153676
rect -6596 153418 -5494 153654
rect -5258 153418 589182 153654
rect 589418 153418 590520 153654
rect -6596 153334 590520 153418
rect -6596 153098 -5494 153334
rect -5258 153098 589182 153334
rect 589418 153098 590520 153334
rect -6596 153076 590520 153098
rect -5676 153074 -5076 153076
rect 589000 153074 589600 153076
rect -3836 150076 -3236 150078
rect 587160 150076 587760 150078
rect -4756 150054 588680 150076
rect -4756 149818 -3654 150054
rect -3418 149818 587342 150054
rect 587578 149818 588680 150054
rect -4756 149734 588680 149818
rect -4756 149498 -3654 149734
rect -3418 149498 587342 149734
rect 587578 149498 588680 149734
rect -4756 149476 588680 149498
rect -3836 149474 -3236 149476
rect 587160 149474 587760 149476
rect -1996 146476 -1396 146478
rect 585320 146476 585920 146478
rect -2916 146454 586840 146476
rect -2916 146218 -1814 146454
rect -1578 146218 585502 146454
rect 585738 146218 586840 146454
rect -2916 146134 586840 146218
rect -2916 145898 -1814 146134
rect -1578 145898 585502 146134
rect 585738 145898 586840 146134
rect -2916 145876 586840 145898
rect -1996 145874 -1396 145876
rect 585320 145874 585920 145876
rect -8436 139276 -7836 139278
rect 591760 139276 592360 139278
rect -8436 139254 592360 139276
rect -8436 139018 -8254 139254
rect -8018 139018 591942 139254
rect 592178 139018 592360 139254
rect -8436 138934 592360 139018
rect -8436 138698 -8254 138934
rect -8018 138698 591942 138934
rect 592178 138698 592360 138934
rect -8436 138676 592360 138698
rect -8436 138674 -7836 138676
rect 591760 138674 592360 138676
rect -6596 135676 -5996 135678
rect 589920 135676 590520 135678
rect -6596 135654 590520 135676
rect -6596 135418 -6414 135654
rect -6178 135418 590102 135654
rect 590338 135418 590520 135654
rect -6596 135334 590520 135418
rect -6596 135098 -6414 135334
rect -6178 135098 590102 135334
rect 590338 135098 590520 135334
rect -6596 135076 590520 135098
rect -6596 135074 -5996 135076
rect 589920 135074 590520 135076
rect -4756 132076 -4156 132078
rect 588080 132076 588680 132078
rect -4756 132054 588680 132076
rect -4756 131818 -4574 132054
rect -4338 131818 588262 132054
rect 588498 131818 588680 132054
rect -4756 131734 588680 131818
rect -4756 131498 -4574 131734
rect -4338 131498 588262 131734
rect 588498 131498 588680 131734
rect -4756 131476 588680 131498
rect -4756 131474 -4156 131476
rect 588080 131474 588680 131476
rect -2916 128476 -2316 128478
rect 586240 128476 586840 128478
rect -2916 128454 586840 128476
rect -2916 128218 -2734 128454
rect -2498 128218 586422 128454
rect 586658 128218 586840 128454
rect -2916 128134 586840 128218
rect -2916 127898 -2734 128134
rect -2498 127898 586422 128134
rect 586658 127898 586840 128134
rect -2916 127876 586840 127898
rect -2916 127874 -2316 127876
rect 586240 127874 586840 127876
rect -7516 121276 -6916 121278
rect 590840 121276 591440 121278
rect -8436 121254 592360 121276
rect -8436 121018 -7334 121254
rect -7098 121018 591022 121254
rect 591258 121018 592360 121254
rect -8436 120934 592360 121018
rect -8436 120698 -7334 120934
rect -7098 120698 591022 120934
rect 591258 120698 592360 120934
rect -8436 120676 592360 120698
rect -7516 120674 -6916 120676
rect 590840 120674 591440 120676
rect -5676 117676 -5076 117678
rect 589000 117676 589600 117678
rect -6596 117654 590520 117676
rect -6596 117418 -5494 117654
rect -5258 117418 589182 117654
rect 589418 117418 590520 117654
rect -6596 117334 590520 117418
rect -6596 117098 -5494 117334
rect -5258 117098 589182 117334
rect 589418 117098 590520 117334
rect -6596 117076 590520 117098
rect -5676 117074 -5076 117076
rect 589000 117074 589600 117076
rect -3836 114076 -3236 114078
rect 587160 114076 587760 114078
rect -4756 114054 588680 114076
rect -4756 113818 -3654 114054
rect -3418 113818 587342 114054
rect 587578 113818 588680 114054
rect -4756 113734 588680 113818
rect -4756 113498 -3654 113734
rect -3418 113498 587342 113734
rect 587578 113498 588680 113734
rect -4756 113476 588680 113498
rect -3836 113474 -3236 113476
rect 587160 113474 587760 113476
rect -1996 110476 -1396 110478
rect 585320 110476 585920 110478
rect -2916 110454 586840 110476
rect -2916 110218 -1814 110454
rect -1578 110218 585502 110454
rect 585738 110218 586840 110454
rect -2916 110134 586840 110218
rect -2916 109898 -1814 110134
rect -1578 109898 585502 110134
rect 585738 109898 586840 110134
rect -2916 109876 586840 109898
rect -1996 109874 -1396 109876
rect 585320 109874 585920 109876
rect -8436 103276 -7836 103278
rect 591760 103276 592360 103278
rect -8436 103254 592360 103276
rect -8436 103018 -8254 103254
rect -8018 103018 591942 103254
rect 592178 103018 592360 103254
rect -8436 102934 592360 103018
rect -8436 102698 -8254 102934
rect -8018 102698 591942 102934
rect 592178 102698 592360 102934
rect -8436 102676 592360 102698
rect -8436 102674 -7836 102676
rect 591760 102674 592360 102676
rect -6596 99676 -5996 99678
rect 589920 99676 590520 99678
rect -6596 99654 590520 99676
rect -6596 99418 -6414 99654
rect -6178 99418 590102 99654
rect 590338 99418 590520 99654
rect -6596 99334 590520 99418
rect -6596 99098 -6414 99334
rect -6178 99098 590102 99334
rect 590338 99098 590520 99334
rect -6596 99076 590520 99098
rect -6596 99074 -5996 99076
rect 589920 99074 590520 99076
rect -4756 96076 -4156 96078
rect 588080 96076 588680 96078
rect -4756 96054 588680 96076
rect -4756 95818 -4574 96054
rect -4338 95818 588262 96054
rect 588498 95818 588680 96054
rect -4756 95734 588680 95818
rect -4756 95498 -4574 95734
rect -4338 95498 588262 95734
rect 588498 95498 588680 95734
rect -4756 95476 588680 95498
rect -4756 95474 -4156 95476
rect 588080 95474 588680 95476
rect -2916 92476 -2316 92478
rect 586240 92476 586840 92478
rect -2916 92454 586840 92476
rect -2916 92218 -2734 92454
rect -2498 92218 586422 92454
rect 586658 92218 586840 92454
rect -2916 92134 586840 92218
rect -2916 91898 -2734 92134
rect -2498 91898 586422 92134
rect 586658 91898 586840 92134
rect -2916 91876 586840 91898
rect -2916 91874 -2316 91876
rect 586240 91874 586840 91876
rect -7516 85276 -6916 85278
rect 590840 85276 591440 85278
rect -8436 85254 592360 85276
rect -8436 85018 -7334 85254
rect -7098 85018 591022 85254
rect 591258 85018 592360 85254
rect -8436 84934 592360 85018
rect -8436 84698 -7334 84934
rect -7098 84698 591022 84934
rect 591258 84698 592360 84934
rect -8436 84676 592360 84698
rect -7516 84674 -6916 84676
rect 590840 84674 591440 84676
rect -5676 81676 -5076 81678
rect 589000 81676 589600 81678
rect -6596 81654 590520 81676
rect -6596 81418 -5494 81654
rect -5258 81418 589182 81654
rect 589418 81418 590520 81654
rect -6596 81334 590520 81418
rect -6596 81098 -5494 81334
rect -5258 81098 589182 81334
rect 589418 81098 590520 81334
rect -6596 81076 590520 81098
rect -5676 81074 -5076 81076
rect 589000 81074 589600 81076
rect -3836 78076 -3236 78078
rect 587160 78076 587760 78078
rect -4756 78054 588680 78076
rect -4756 77818 -3654 78054
rect -3418 77818 587342 78054
rect 587578 77818 588680 78054
rect -4756 77734 588680 77818
rect -4756 77498 -3654 77734
rect -3418 77498 587342 77734
rect 587578 77498 588680 77734
rect -4756 77476 588680 77498
rect -3836 77474 -3236 77476
rect 587160 77474 587760 77476
rect -1996 74476 -1396 74478
rect 585320 74476 585920 74478
rect -2916 74454 586840 74476
rect -2916 74218 -1814 74454
rect -1578 74218 585502 74454
rect 585738 74218 586840 74454
rect -2916 74134 586840 74218
rect -2916 73898 -1814 74134
rect -1578 73898 585502 74134
rect 585738 73898 586840 74134
rect -2916 73876 586840 73898
rect -1996 73874 -1396 73876
rect 585320 73874 585920 73876
rect -8436 67276 -7836 67278
rect 591760 67276 592360 67278
rect -8436 67254 592360 67276
rect -8436 67018 -8254 67254
rect -8018 67018 591942 67254
rect 592178 67018 592360 67254
rect -8436 66934 592360 67018
rect -8436 66698 -8254 66934
rect -8018 66698 591942 66934
rect 592178 66698 592360 66934
rect -8436 66676 592360 66698
rect -8436 66674 -7836 66676
rect 591760 66674 592360 66676
rect -6596 63676 -5996 63678
rect 589920 63676 590520 63678
rect -6596 63654 590520 63676
rect -6596 63418 -6414 63654
rect -6178 63418 590102 63654
rect 590338 63418 590520 63654
rect -6596 63334 590520 63418
rect -6596 63098 -6414 63334
rect -6178 63098 590102 63334
rect 590338 63098 590520 63334
rect -6596 63076 590520 63098
rect -6596 63074 -5996 63076
rect 589920 63074 590520 63076
rect -4756 60076 -4156 60078
rect 588080 60076 588680 60078
rect -4756 60054 588680 60076
rect -4756 59818 -4574 60054
rect -4338 59818 588262 60054
rect 588498 59818 588680 60054
rect -4756 59734 588680 59818
rect -4756 59498 -4574 59734
rect -4338 59498 588262 59734
rect 588498 59498 588680 59734
rect -4756 59476 588680 59498
rect -4756 59474 -4156 59476
rect 588080 59474 588680 59476
rect -2916 56476 -2316 56478
rect 586240 56476 586840 56478
rect -2916 56454 586840 56476
rect -2916 56218 -2734 56454
rect -2498 56218 586422 56454
rect 586658 56218 586840 56454
rect -2916 56134 586840 56218
rect -2916 55898 -2734 56134
rect -2498 55898 586422 56134
rect 586658 55898 586840 56134
rect -2916 55876 586840 55898
rect -2916 55874 -2316 55876
rect 586240 55874 586840 55876
rect -7516 49276 -6916 49278
rect 590840 49276 591440 49278
rect -8436 49254 592360 49276
rect -8436 49018 -7334 49254
rect -7098 49018 591022 49254
rect 591258 49018 592360 49254
rect -8436 48934 592360 49018
rect -8436 48698 -7334 48934
rect -7098 48698 591022 48934
rect 591258 48698 592360 48934
rect -8436 48676 592360 48698
rect -7516 48674 -6916 48676
rect 590840 48674 591440 48676
rect -5676 45676 -5076 45678
rect 589000 45676 589600 45678
rect -6596 45654 590520 45676
rect -6596 45418 -5494 45654
rect -5258 45418 589182 45654
rect 589418 45418 590520 45654
rect -6596 45334 590520 45418
rect -6596 45098 -5494 45334
rect -5258 45098 589182 45334
rect 589418 45098 590520 45334
rect -6596 45076 590520 45098
rect -5676 45074 -5076 45076
rect 589000 45074 589600 45076
rect -3836 42076 -3236 42078
rect 587160 42076 587760 42078
rect -4756 42054 588680 42076
rect -4756 41818 -3654 42054
rect -3418 41818 587342 42054
rect 587578 41818 588680 42054
rect -4756 41734 588680 41818
rect -4756 41498 -3654 41734
rect -3418 41498 587342 41734
rect 587578 41498 588680 41734
rect -4756 41476 588680 41498
rect -3836 41474 -3236 41476
rect 587160 41474 587760 41476
rect -1996 38476 -1396 38478
rect 585320 38476 585920 38478
rect -2916 38454 586840 38476
rect -2916 38218 -1814 38454
rect -1578 38218 585502 38454
rect 585738 38218 586840 38454
rect -2916 38134 586840 38218
rect -2916 37898 -1814 38134
rect -1578 37898 585502 38134
rect 585738 37898 586840 38134
rect -2916 37876 586840 37898
rect -1996 37874 -1396 37876
rect 585320 37874 585920 37876
rect 1220 36498 559428 36540
rect 1220 36262 1262 36498
rect 1498 36262 559150 36498
rect 559386 36262 559428 36498
rect 1220 36220 559428 36262
rect 1588 35818 559796 35860
rect 1588 35582 1630 35818
rect 1866 35582 559518 35818
rect 559754 35582 559796 35818
rect 1588 35540 559796 35582
rect 559660 35138 562188 35180
rect 559660 34902 559702 35138
rect 559938 34902 561910 35138
rect 562146 34902 562188 35138
rect 559660 34860 562188 34902
rect 852 34458 562556 34500
rect 852 34222 894 34458
rect 1130 34222 562278 34458
rect 562514 34222 562556 34458
rect 852 34180 562556 34222
rect 1588 33098 561268 33140
rect 1588 32862 1630 33098
rect 1866 32862 560990 33098
rect 561226 32862 561268 33098
rect 1588 32820 561268 32862
rect 484 32418 561636 32460
rect 484 32182 526 32418
rect 762 32182 561358 32418
rect 561594 32182 561636 32418
rect 484 32140 561636 32182
rect 562052 32418 570468 32460
rect 562052 32182 562094 32418
rect 562330 32182 570190 32418
rect 570426 32182 570468 32418
rect 562052 32140 570468 32182
rect -8436 31276 -7836 31278
rect 591760 31276 592360 31278
rect -8436 31254 592360 31276
rect -8436 31018 -8254 31254
rect -8018 31018 591942 31254
rect 592178 31018 592360 31254
rect -8436 30934 592360 31018
rect -8436 30698 -8254 30934
rect -8018 30698 591942 30934
rect 592178 30698 592360 30934
rect -8436 30676 592360 30698
rect -8436 30674 -7836 30676
rect 591760 30674 592360 30676
rect 1588 29698 562004 29740
rect 1588 29462 1630 29698
rect 1866 29462 561726 29698
rect 561962 29462 562004 29698
rect 1588 29420 562004 29462
rect 1220 29018 560900 29060
rect 1220 28782 1262 29018
rect 1498 28782 560622 29018
rect 560858 28782 560900 29018
rect 1220 28740 560900 28782
rect -6596 27676 -5996 27678
rect 589920 27676 590520 27678
rect -6596 27654 590520 27676
rect -6596 27418 -6414 27654
rect -6178 27418 590102 27654
rect 590338 27418 590520 27654
rect -6596 27334 590520 27418
rect -6596 27098 -6414 27334
rect -6178 27098 590102 27334
rect 590338 27098 590520 27334
rect -6596 27076 590520 27098
rect -6596 27074 -5996 27076
rect 589920 27074 590520 27076
rect 1772 26298 561636 26340
rect 1772 26062 1814 26298
rect 2050 26062 561358 26298
rect 561594 26062 561636 26298
rect 1772 26020 561636 26062
rect 1036 25618 562372 25660
rect 1036 25382 1078 25618
rect 1314 25382 562094 25618
rect 562330 25382 562372 25618
rect 1036 25340 562372 25382
rect 1404 24938 559980 24980
rect 1404 24702 1446 24938
rect 1682 24702 559702 24938
rect 559938 24702 559980 24938
rect 1404 24660 559980 24702
rect -4756 24076 -4156 24078
rect 588080 24076 588680 24078
rect -4756 24054 588680 24076
rect -4756 23818 -4574 24054
rect -4338 23818 588262 24054
rect 588498 23818 588680 24054
rect -4756 23734 588680 23818
rect -4756 23498 -4574 23734
rect -4338 23498 588262 23734
rect 588498 23498 588680 23734
rect -4756 23476 588680 23498
rect -4756 23474 -4156 23476
rect 588080 23474 588680 23476
rect -2916 20476 -2316 20478
rect 586240 20476 586840 20478
rect -2916 20454 586840 20476
rect -2916 20218 -2734 20454
rect -2498 20218 586422 20454
rect 586658 20218 586840 20454
rect -2916 20134 586840 20218
rect -2916 19898 -2734 20134
rect -2498 19898 586422 20134
rect 586658 19898 586840 20134
rect -2916 19876 586840 19898
rect -2916 19874 -2316 19876
rect 586240 19874 586840 19876
rect 199388 19220 206148 19540
rect 199388 18860 199708 19220
rect 56236 18540 63364 18860
rect 26060 17180 42388 17500
rect 26060 16140 26380 17180
rect 20908 15820 26380 16140
rect 26796 15820 37236 16140
rect 20908 15460 21228 15820
rect 852 15418 21228 15460
rect 852 15182 894 15418
rect 1130 15182 21228 15418
rect 852 15140 21228 15182
rect 26796 14780 27116 15820
rect 23300 14460 27116 14780
rect 36916 14780 37236 15820
rect 42068 15460 42388 17180
rect 56236 16820 56556 18540
rect 52372 16500 56556 16820
rect 52372 15460 52692 16500
rect 63044 16140 63364 18540
rect 199020 18540 199708 18860
rect 200308 18540 204676 18860
rect 121188 16820 121692 17500
rect 140508 16820 141012 17500
rect 159828 16820 160332 17500
rect 199020 16820 199340 18540
rect 98004 16500 107524 16820
rect 63044 15820 93908 16140
rect 42068 15140 52692 15460
rect 93588 15460 93908 15820
rect 98004 15460 98324 16500
rect 93588 15140 98324 15460
rect 107204 15460 107524 16500
rect 114196 16500 121692 16820
rect 114196 15460 114516 16500
rect 121372 16140 121692 16500
rect 133516 16500 141012 16820
rect 121372 15820 124452 16140
rect 107204 15140 114516 15460
rect 124132 15460 124452 15820
rect 133516 15460 133836 16500
rect 140692 16140 141012 16500
rect 145476 16500 149108 16820
rect 145476 16140 145796 16500
rect 140692 15820 145796 16140
rect 148788 16140 149108 16500
rect 149524 16500 173396 16820
rect 149524 16140 149844 16500
rect 148788 15820 149844 16140
rect 173076 16140 173396 16500
rect 194420 16500 199340 16820
rect 173076 15820 186092 16140
rect 124132 15140 133836 15460
rect 148788 15140 149292 15820
rect 185772 15460 186092 15820
rect 194420 15460 194740 16500
rect 200308 16140 200628 18540
rect 185772 15140 194740 15460
rect 199020 15820 200628 16140
rect 199020 14780 199340 15820
rect 36916 14460 38156 14780
rect 23300 14100 23620 14460
rect 1772 14058 5036 14100
rect 1772 13822 1814 14058
rect 2050 13822 4758 14058
rect 4994 13822 5036 14058
rect 20724 13960 23620 14100
rect 1772 13780 5036 13822
rect 19988 13780 23620 13960
rect 37836 14100 38156 14460
rect 48876 14460 52692 14780
rect 48876 14100 49196 14460
rect 37836 13780 49196 14100
rect 52372 14100 52692 14460
rect 64884 14460 73484 14780
rect 64884 14100 65204 14460
rect 52372 13780 65204 14100
rect 73164 14100 73484 14460
rect 91932 14460 199340 14780
rect 204356 14780 204676 18540
rect 205828 17500 206148 19220
rect 547516 19220 551332 19540
rect 266364 17860 276068 18180
rect 205828 17180 206700 17500
rect 206380 16140 206700 17180
rect 212452 16500 226388 16820
rect 212452 16140 212772 16500
rect 206380 15820 212772 16140
rect 226068 15460 226388 16500
rect 226804 16500 236140 16820
rect 226804 15460 227124 16500
rect 235820 16140 236140 16500
rect 246124 16500 254908 16820
rect 226068 15140 227124 15460
rect 227540 15820 234852 16140
rect 235820 15820 245708 16140
rect 227540 14780 227860 15820
rect 234532 15460 234852 15820
rect 245388 15460 245708 15820
rect 246124 15460 246444 16500
rect 254588 16140 254908 16500
rect 256980 16500 263004 16820
rect 254588 15820 255092 16140
rect 234532 15140 235404 15460
rect 245388 15140 246444 15460
rect 254772 15460 255092 15820
rect 256980 15460 257300 16500
rect 254772 15140 257300 15460
rect 262684 15460 263004 16500
rect 266364 15460 266684 17860
rect 262684 15140 266684 15460
rect 275748 15460 276068 17860
rect 547516 17500 547836 19220
rect 551012 18860 551332 19220
rect 551012 18818 559980 18860
rect 551012 18582 559702 18818
rect 559938 18582 559980 18818
rect 551012 18540 559980 18582
rect 545676 17180 547836 17500
rect 288996 15820 293364 16140
rect 288996 15460 289316 15820
rect 275748 15140 289316 15460
rect 293044 15460 293364 15820
rect 308316 15820 312684 16140
rect 308316 15460 308636 15820
rect 293044 15140 308636 15460
rect 312364 15460 312684 15820
rect 327636 15820 332004 16140
rect 327636 15460 327956 15820
rect 312364 15140 327956 15460
rect 331684 15460 332004 15820
rect 346956 15820 351324 16140
rect 346956 15460 347276 15820
rect 331684 15140 347276 15460
rect 351004 15460 351324 15820
rect 366276 15820 370644 16140
rect 366276 15460 366596 15820
rect 351004 15140 366596 15460
rect 370324 15460 370644 15820
rect 385596 15820 389964 16140
rect 385596 15460 385916 15820
rect 370324 15140 385916 15460
rect 389644 15460 389964 15820
rect 404916 15820 409284 16140
rect 404916 15460 405236 15820
rect 389644 15140 405236 15460
rect 408964 15460 409284 15820
rect 424236 15820 428604 16140
rect 424236 15460 424556 15820
rect 408964 15140 424556 15460
rect 428284 15460 428604 15820
rect 443556 15820 447924 16140
rect 443556 15460 443876 15820
rect 428284 15140 443876 15460
rect 447604 15460 447924 15820
rect 462876 15820 467244 16140
rect 462876 15460 463196 15820
rect 447604 15140 463196 15460
rect 466924 15460 467244 15820
rect 482196 15820 486564 16140
rect 482196 15460 482516 15820
rect 466924 15140 482516 15460
rect 486244 15460 486564 15820
rect 501516 15820 505884 16140
rect 501516 15460 501836 15820
rect 486244 15140 501836 15460
rect 505564 15460 505884 15820
rect 520836 15820 525204 16140
rect 520836 15460 521156 15820
rect 505564 15140 521156 15460
rect 524884 15460 525204 15820
rect 545676 15460 545996 17180
rect 548988 16098 559060 16140
rect 548988 15862 558782 16098
rect 559018 15862 559060 16098
rect 548988 15820 559060 15862
rect 548988 15460 549308 15820
rect 524884 15140 545996 15460
rect 548620 15140 549308 15460
rect 204356 14460 227860 14780
rect 91932 14100 92252 14460
rect 73164 13780 92252 14100
rect 235084 14100 235404 15140
rect 237292 14460 538268 14780
rect 237292 14100 237612 14460
rect 235084 13780 237612 14100
rect 456436 13780 456940 14460
rect 475756 13780 476260 14460
rect 495076 13780 495580 14460
rect 514396 13780 514900 14460
rect 537948 14100 538268 14460
rect 548620 14100 548940 15140
rect 537948 13780 548940 14100
rect 19988 13640 21044 13780
rect 19988 13378 20308 13640
rect -7516 13276 -6916 13278
rect 19988 13276 20030 13378
rect -8436 13254 20030 13276
rect -8436 13018 -7334 13254
rect -7098 13142 20030 13254
rect 20266 13276 20308 13378
rect 590840 13276 591440 13278
rect 20266 13254 592360 13276
rect 20266 13142 591022 13254
rect -7098 13018 591022 13142
rect 591258 13018 592360 13254
rect -8436 12934 592360 13018
rect -8436 12698 -7334 12934
rect -7098 12698 591022 12934
rect 591258 12698 592360 12934
rect -8436 12676 592360 12698
rect -7516 12674 -6916 12676
rect 78316 12420 81212 12676
rect 590840 12674 591440 12676
rect 78316 12060 78636 12420
rect 4716 12018 10556 12060
rect 4716 11782 4758 12018
rect 4994 11782 10556 12018
rect 4716 11740 10556 11782
rect 10236 11380 10556 11740
rect 11340 11740 30428 12060
rect 11340 11380 11660 11740
rect 30108 11380 30428 11740
rect 33972 11740 46988 12060
rect 10236 11060 11660 11380
rect 12628 11060 28588 11380
rect 12628 10700 12948 11060
rect 1404 10658 12948 10700
rect 1404 10422 1446 10658
rect 1682 10422 12948 10658
rect 1404 10380 12948 10422
rect 28268 10700 28588 11060
rect 29004 11060 31164 11380
rect 29004 10700 29324 11060
rect 28268 10380 29324 10700
rect 30108 10020 30428 11060
rect 30844 10700 31164 11060
rect 33972 10700 34292 11740
rect 46668 11380 46988 11740
rect 62124 11740 64836 12060
rect 62124 11380 62444 11740
rect 64516 11380 64836 11740
rect 65804 11740 78636 12060
rect 80892 12060 81212 12420
rect 80892 11740 83236 12060
rect 65804 11380 66124 11740
rect 82916 11380 83236 11740
rect 91932 11740 105684 12060
rect 91932 11380 92252 11740
rect 105364 11380 105684 11740
rect 111988 11740 117828 12060
rect 111988 11380 112308 11740
rect 30844 10380 34292 10700
rect 34892 11060 62444 11380
rect 63044 11060 66124 11380
rect 67276 11060 72564 11380
rect 82916 11060 92252 11380
rect 92668 11060 104028 11380
rect 105364 11060 112308 11380
rect 117508 11380 117828 11740
rect 118428 11740 150396 12060
rect 118428 11380 118748 11740
rect 150076 11380 150396 11740
rect 150996 11740 152972 12060
rect 150996 11380 151316 11740
rect 152652 11380 152972 11740
rect 153388 11740 154628 12060
rect 153388 11380 153708 11740
rect 117508 11060 118748 11380
rect 119716 11060 128868 11380
rect 34892 10020 35212 11060
rect 46668 10700 46988 11060
rect 63044 10700 63364 11060
rect 46668 10380 63364 10700
rect 64516 10700 64836 11060
rect 67276 10700 67596 11060
rect 64516 10380 67596 10700
rect 72244 10700 72564 11060
rect 92668 10700 92988 11060
rect 72244 10380 92988 10700
rect 103708 10700 104028 11060
rect 119716 10700 120036 11060
rect 103708 10380 120036 10700
rect 128548 10700 128868 11060
rect 130940 11060 132732 11380
rect 150076 11060 151684 11380
rect 152652 11060 153708 11380
rect 154308 11380 154628 11740
rect 178780 11740 182228 12060
rect 178780 11380 179100 11740
rect 181908 11380 182228 11740
rect 184852 11740 187012 12060
rect 184852 11380 185172 11740
rect 154308 11060 179836 11380
rect 181908 11060 185172 11380
rect 186692 11380 187012 11740
rect 187428 11380 187932 12060
rect 201964 11740 218292 12060
rect 201964 11380 202284 11740
rect 217972 11380 218292 11740
rect 225516 11740 229332 12060
rect 225516 11380 225836 11740
rect 186692 11060 202284 11380
rect 207484 11060 216820 11380
rect 217972 11060 225836 11380
rect 229012 11380 229332 11740
rect 247044 11740 249756 12060
rect 247044 11380 247364 11740
rect 249436 11380 249756 11740
rect 250356 11740 262084 12060
rect 250356 11380 250676 11740
rect 229012 11060 247364 11380
rect 247780 11060 249020 11380
rect 249436 11060 250676 11380
rect 261764 11380 262084 11740
rect 265996 11740 315260 12060
rect 265996 11380 266316 11740
rect 314940 11380 315260 11740
rect 323956 11740 334212 12060
rect 323956 11380 324276 11740
rect 333892 11380 334212 11740
rect 339964 11740 344884 12060
rect 339964 11380 340284 11740
rect 344564 11380 344884 11740
rect 345668 11740 373956 12060
rect 345668 11380 345988 11740
rect 373636 11380 373956 11740
rect 380812 12018 558876 12060
rect 380812 11782 558598 12018
rect 558834 11782 558876 12018
rect 380812 11740 558876 11782
rect 380812 11380 381132 11740
rect 261764 11060 266316 11380
rect 269676 11060 288764 11380
rect 314940 11060 324276 11380
rect 328924 11060 331636 11380
rect 333892 11060 340284 11380
rect 342724 11060 343964 11380
rect 344564 11060 345988 11380
rect 347324 11060 373220 11380
rect 373636 11060 381132 11380
rect 381548 11060 432284 11380
rect 130940 10700 131260 11060
rect 128548 10380 131260 10700
rect 132412 10700 132732 11060
rect 150444 10700 150764 11060
rect 132412 10380 150764 10700
rect 151364 10700 151684 11060
rect 178780 10700 179100 11060
rect 151364 10380 179100 10700
rect 179516 10700 179836 11060
rect 207484 10700 207804 11060
rect 179516 10380 207804 10700
rect 216500 10700 216820 11060
rect 247780 10700 248100 11060
rect 216500 10380 248100 10700
rect 248700 10700 249020 11060
rect 269676 10700 269996 11060
rect 248700 10380 269996 10700
rect 288444 10700 288764 11060
rect 328924 10700 329244 11060
rect 288444 10380 329244 10700
rect 331316 10700 331636 11060
rect 342724 10700 343044 11060
rect 331316 10380 343044 10700
rect 343644 10700 343964 11060
rect 347324 10700 347644 11060
rect 343644 10380 347644 10700
rect 372900 10700 373220 11060
rect 381548 10700 381868 11060
rect 372900 10380 381868 10700
rect 431964 10700 432284 11060
rect 443556 11060 444612 11380
rect 443556 10700 443876 11060
rect 431964 10380 443876 10700
rect 444292 10700 444612 11060
rect 453676 11060 454732 11380
rect 453676 10700 453996 11060
rect 444292 10380 453996 10700
rect 454412 10700 454732 11060
rect 462876 11060 463932 11380
rect 462876 10700 463196 11060
rect 454412 10380 463196 10700
rect 463612 10700 463932 11060
rect 472996 11060 474052 11380
rect 472996 10700 473316 11060
rect 463612 10380 473316 10700
rect 473732 10700 474052 11060
rect 482196 11060 483252 11380
rect 482196 10700 482516 11060
rect 473732 10380 482516 10700
rect 482932 10700 483252 11060
rect 492316 11060 493372 11380
rect 492316 10700 492636 11060
rect 482932 10380 492636 10700
rect 493052 10700 493372 11060
rect 501516 11060 502572 11380
rect 501516 10700 501836 11060
rect 493052 10380 501836 10700
rect 502252 10700 502572 11060
rect 511636 11060 530908 11380
rect 511636 10700 511956 11060
rect 502252 10380 511956 10700
rect 530588 10700 530908 11060
rect 540340 11338 559244 11380
rect 540340 11102 558966 11338
rect 559202 11102 559244 11338
rect 540340 11060 559244 11102
rect 559660 11338 570468 11380
rect 559660 11102 559702 11338
rect 559938 11102 570190 11338
rect 570426 11102 570468 11338
rect 559660 11060 570468 11102
rect 540340 10700 540660 11060
rect 530588 10380 540660 10700
rect 30108 9700 35212 10020
rect -5676 9676 -5076 9678
rect 589000 9676 589600 9678
rect -6596 9654 590520 9676
rect -6596 9418 -5494 9654
rect -5258 9418 589182 9654
rect 589418 9418 590520 9654
rect -6596 9334 590520 9418
rect -6596 9098 -5494 9334
rect -5258 9098 589182 9334
rect 589418 9098 590520 9334
rect -6596 9076 590520 9098
rect -5676 9074 -5076 9076
rect 589000 9074 589600 9076
rect 13916 8340 21780 8660
rect 13916 7980 14236 8340
rect 21460 7980 21780 8340
rect 38434 8340 60972 8660
rect 38434 7980 38754 8340
rect 484 7938 14236 7980
rect 484 7702 526 7938
rect 762 7702 14236 7938
rect 484 7660 14236 7702
rect 19804 7938 20124 7980
rect 19804 7702 19846 7938
rect 20082 7702 20124 7938
rect 19804 7300 20124 7702
rect 21460 7660 38754 7980
rect 60652 7980 60972 8340
rect 79788 8340 84340 8660
rect 79788 7980 80108 8340
rect 60652 7660 64836 7980
rect 4716 7258 20124 7300
rect 4716 7022 4758 7258
rect 4994 7022 20124 7258
rect 4716 6980 20124 7022
rect 64516 7300 64836 7660
rect 72980 7660 80108 7980
rect 72980 7300 73300 7660
rect 64516 6980 73300 7300
rect 84020 7300 84340 8340
rect 97084 8340 111940 8660
rect 97084 7300 97404 8340
rect 84020 6980 97404 7300
rect 111620 7300 111940 8340
rect 121188 8340 127212 8660
rect 121188 7980 121508 8340
rect 114380 7660 121508 7980
rect 126892 7980 127212 8340
rect 135724 8340 167140 8660
rect 135724 7980 136044 8340
rect 126892 7660 128638 7980
rect 114380 7300 114700 7660
rect 111620 6980 114700 7300
rect 128318 7300 128638 7660
rect 135172 7660 136044 7980
rect 166820 7980 167140 8340
rect 179332 8340 189220 8660
rect 179332 7980 179652 8340
rect 166820 7660 170084 7980
rect 135172 7300 135492 7660
rect 128318 6980 135492 7300
rect 169764 7300 170084 7660
rect 176572 7660 179652 7980
rect 176572 7300 176892 7660
rect 169764 6980 176892 7300
rect 188900 7300 189220 8340
rect 212636 8340 221420 8660
rect 212636 7300 212956 8340
rect 221100 7980 221420 8340
rect 221100 7660 226020 7980
rect 188900 6980 212956 7300
rect 225700 6578 226020 7660
rect 225700 6342 225742 6578
rect 225978 6342 226020 6578
rect 225700 6300 226020 6342
rect -3836 6076 -3236 6078
rect 587160 6076 587760 6078
rect -4756 6054 588680 6076
rect -4756 5818 -3654 6054
rect -3418 5818 587342 6054
rect 587578 5818 588680 6054
rect -4756 5734 588680 5818
rect -4756 5498 -3654 5734
rect -3418 5498 587342 5734
rect 587578 5498 588680 5734
rect -4756 5476 588680 5498
rect -3836 5474 -3236 5476
rect 587160 5474 587760 5476
rect 225700 5218 226020 5260
rect 225700 4982 225742 5218
rect 225978 4982 226020 5218
rect 1220 4538 33878 4580
rect 1220 4302 1262 4538
rect 1498 4302 33878 4538
rect 1220 4260 33878 4302
rect 33558 3900 33878 4260
rect 35444 4260 76612 4580
rect 35444 3900 35764 4260
rect 14836 3580 29140 3900
rect 33558 3580 35764 3900
rect 14836 3178 15156 3580
rect 14836 2942 14878 3178
rect 15114 2942 15156 3178
rect 14836 2900 15156 2942
rect 28820 3178 29140 3580
rect 28820 2942 28862 3178
rect 29098 2942 29140 3178
rect 28820 2900 29140 2942
rect 52188 3178 75140 3220
rect 52188 2942 52230 3178
rect 52466 2942 74862 3178
rect 75098 2942 75140 3178
rect 52188 2900 75140 2942
rect 76292 3178 76612 4260
rect 76292 2942 76334 3178
rect 76570 2942 76612 3178
rect 76292 2900 76612 2942
rect 78500 4260 80108 4580
rect 78500 3178 78820 4260
rect 79788 3900 80108 4260
rect 95980 4260 126292 4580
rect 95980 3900 96300 4260
rect 79788 3580 95012 3900
rect 78500 2942 78542 3178
rect 78778 2942 78820 3178
rect 78500 2900 78820 2942
rect 82180 3178 91700 3220
rect 82180 2942 82222 3178
rect 82458 2942 91422 3178
rect 91658 2942 91700 3178
rect 82180 2900 91700 2942
rect 94692 3178 95012 3580
rect 95796 3580 96300 3900
rect 96716 3858 124498 3900
rect 96716 3622 124220 3858
rect 124456 3622 124498 3858
rect 96716 3580 124498 3622
rect 95796 3220 96116 3580
rect 94692 2942 94734 3178
rect 94970 2942 95012 3178
rect 94692 2900 95012 2942
rect 95612 3178 96116 3220
rect 95612 2942 95654 3178
rect 95890 2942 96116 3178
rect 95612 2900 96116 2942
rect 96716 3178 97036 3580
rect 96716 2942 96758 3178
rect 96994 2942 97036 3178
rect 96716 2900 97036 2942
rect 102604 3178 125556 3220
rect 102604 2942 102646 3178
rect 102882 2942 125278 3178
rect 125514 2942 125556 3178
rect 102604 2900 125556 2942
rect 125972 3178 126292 4260
rect 134988 4260 152742 4580
rect 134988 3220 135308 4260
rect 152422 3900 152742 4260
rect 155228 4260 195108 4580
rect 125972 2942 126014 3178
rect 126250 2942 126292 3178
rect 125972 2900 126292 2942
rect 127076 3178 135308 3220
rect 127076 2942 127118 3178
rect 127354 2942 135308 3178
rect 127076 2900 135308 2942
rect 135724 3580 147130 3900
rect 152422 3580 154628 3900
rect 135724 3178 136044 3580
rect 146810 3220 147130 3580
rect 135724 2942 135766 3178
rect 136002 2942 136044 3178
rect 135724 2900 136044 2942
rect 136460 3178 146164 3220
rect 136460 2942 136502 3178
rect 136738 2942 145886 3178
rect 146122 2942 146164 3178
rect 136460 2900 146164 2942
rect 146810 3178 153892 3220
rect 146810 2942 153614 3178
rect 153850 2942 153892 3178
rect 146810 2900 153892 2942
rect 154308 3178 154628 3580
rect 154308 2942 154350 3178
rect 154586 2942 154628 3178
rect 154308 2900 154628 2942
rect 155228 3178 155548 4260
rect 155228 2942 155270 3178
rect 155506 2942 155548 3178
rect 155228 2900 155548 2942
rect 155964 3858 178134 3900
rect 155964 3622 177856 3858
rect 178092 3622 178134 3858
rect 155964 3580 178134 3622
rect 178550 3580 194372 3900
rect 155964 3178 156284 3580
rect 178550 3220 178870 3580
rect 155964 2942 156006 3178
rect 156242 2942 156284 3178
rect 155964 2900 156284 2942
rect 157988 3178 178870 3220
rect 157988 2942 158030 3178
rect 158266 2942 178870 3178
rect 157988 2900 178870 2942
rect 194052 3178 194372 3580
rect 194052 2942 194094 3178
rect 194330 2942 194372 3178
rect 194052 2900 194372 2942
rect 194788 2498 195108 4260
rect 202884 4260 221236 4580
rect 202884 3900 203204 4260
rect 195708 3580 203204 3900
rect 220916 3900 221236 4260
rect 220916 3580 225284 3900
rect 195708 3220 196028 3580
rect 195524 3178 196028 3220
rect 195524 2942 195566 3178
rect 195802 2942 196028 3178
rect 195524 2900 196028 2942
rect 200860 3178 224364 3220
rect 200860 2942 200902 3178
rect 201138 2942 224086 3178
rect 224322 2942 224364 3178
rect 200860 2900 224364 2942
rect 224964 3178 225284 3580
rect 224964 2942 225006 3178
rect 225242 2942 225284 3178
rect 224964 2900 225284 2942
rect 225700 2878 226020 4982
rect 226988 4260 259508 4580
rect 226988 3900 227308 4260
rect 259188 3900 259508 4260
rect 276116 4260 279748 4580
rect 276116 3900 276436 4260
rect 226804 3580 227308 3900
rect 227724 3580 257116 3900
rect 259188 3580 261762 3900
rect 268250 3858 276436 3900
rect 268250 3622 268292 3858
rect 268528 3622 276436 3858
rect 268250 3580 276436 3622
rect 279428 3900 279748 4260
rect 333156 4260 354452 4580
rect 279428 3580 310292 3900
rect 226804 3178 227124 3580
rect 226804 2942 226846 3178
rect 227082 2942 227124 3178
rect 226804 2900 227124 2942
rect 227724 3178 228044 3580
rect 256796 3220 257116 3580
rect 261442 3220 261762 3580
rect 227724 2942 227766 3178
rect 228002 2942 228044 3178
rect 227724 2900 228044 2942
rect 228644 3178 253620 3220
rect 228644 2942 228686 3178
rect 228922 2942 253342 3178
rect 253578 2942 253620 3178
rect 228644 2900 253620 2942
rect 256796 3178 260428 3220
rect 256796 2942 260150 3178
rect 260386 2942 260428 3178
rect 256796 2900 260428 2942
rect 261442 3178 294652 3220
rect 261442 2942 294374 3178
rect 294610 2942 294652 3178
rect 261442 2900 294652 2942
rect 309972 3178 310292 3580
rect 309972 2942 310014 3178
rect 310250 2942 310292 3178
rect 309972 2900 310292 2942
rect 311076 3580 328692 3900
rect 311076 3178 311396 3580
rect 311076 2942 311118 3178
rect 311354 2942 311396 3178
rect 311076 2900 311396 2942
rect 328372 3220 328692 3580
rect 333156 3220 333476 4260
rect 328372 2900 333476 3220
rect 336652 3580 349116 3900
rect 336652 3178 336972 3580
rect 336652 2942 336694 3178
rect 336930 2942 336972 3178
rect 336652 2900 336972 2942
rect 348796 3178 349116 3580
rect 348796 2942 348838 3178
rect 349074 2942 349116 3178
rect 348796 2900 349116 2942
rect 354132 3178 354452 4260
rect 389644 4260 403212 4580
rect 389644 3900 389964 4260
rect 354132 2942 354174 3178
rect 354410 2942 354452 3178
rect 354132 2900 354452 2942
rect 372394 3580 388676 3900
rect 372394 3178 372714 3580
rect 372394 2942 372436 3178
rect 372672 2942 372714 3178
rect 372394 2900 372714 2942
rect 388356 3220 388676 3580
rect 389460 3580 389964 3900
rect 402892 3900 403212 4260
rect 457724 4260 488726 4580
rect 457724 3900 458044 4260
rect 488406 3900 488726 4260
rect 489188 4260 490382 4580
rect 489188 3900 489508 4260
rect 402892 3580 419588 3900
rect 389460 3220 389780 3580
rect 388356 2900 389780 3220
rect 419268 3178 419588 3580
rect 419268 2942 419310 3178
rect 419546 2942 419588 3178
rect 419268 2900 419588 2942
rect 426812 3580 458044 3900
rect 472812 3580 483988 3900
rect 488406 3580 489508 3900
rect 490062 3900 490382 4260
rect 490844 4260 499444 4580
rect 490062 3580 490428 3900
rect 426812 3178 427132 3580
rect 472812 3220 473132 3580
rect 426812 2942 426854 3178
rect 427090 2942 427132 3178
rect 426812 2900 427132 2942
rect 442820 3178 473132 3220
rect 442820 2942 442862 3178
rect 443098 2942 473132 3178
rect 442820 2900 473132 2942
rect 483668 3178 483988 3580
rect 483668 2942 483710 3178
rect 483946 2942 483988 3178
rect 483668 2900 483988 2942
rect 490108 3220 490428 3580
rect 490844 3220 491164 4260
rect 499124 3900 499444 4260
rect 530956 4260 532932 4580
rect 499124 3580 513428 3900
rect 490108 2900 491164 3220
rect 513108 3178 513428 3580
rect 530956 3220 531276 4260
rect 513108 2942 513150 3178
rect 513386 2942 513428 3178
rect 513108 2900 513428 2942
rect 514396 3178 531276 3220
rect 514396 2942 514438 3178
rect 514674 2942 531276 3178
rect 514396 2900 531276 2942
rect 532612 3220 532932 4260
rect 536476 4260 541212 4580
rect 536476 3220 536796 4260
rect 532612 2900 536796 3220
rect 540892 3220 541212 4260
rect 544756 4260 549492 4580
rect 544756 3220 545076 4260
rect 540892 2900 545076 3220
rect 549172 3220 549492 4260
rect 553036 4260 558324 4580
rect 560028 4538 570652 4580
rect 560028 4302 560070 4538
rect 560306 4302 570374 4538
rect 570610 4302 570652 4538
rect 560028 4260 570652 4302
rect 553036 3220 553356 4260
rect 558004 3900 558324 4260
rect 558004 3858 559612 3900
rect 558004 3622 559334 3858
rect 559570 3622 559612 3858
rect 558004 3580 559612 3622
rect 560028 3858 569732 3900
rect 560028 3622 560070 3858
rect 560306 3622 569454 3858
rect 569690 3622 569732 3858
rect 560028 3580 569732 3622
rect 549172 2900 553356 3220
rect 225700 2642 225742 2878
rect 225978 2642 226020 2878
rect 225700 2600 226020 2642
rect -1996 2476 -1396 2478
rect 194788 2476 194830 2498
rect -2916 2454 194830 2476
rect -2916 2218 -1814 2454
rect -1578 2262 194830 2454
rect 195066 2476 195108 2498
rect 585320 2476 585920 2478
rect 195066 2454 586840 2476
rect 195066 2262 585502 2454
rect -1578 2218 585502 2262
rect 585738 2218 586840 2454
rect -2916 2134 586840 2218
rect -2916 1898 -1814 2134
rect -1578 1954 585502 2134
rect -1578 1898 154028 1954
rect -2916 1876 154028 1898
rect -1996 1874 -1396 1876
rect 126340 1818 127396 1860
rect 126340 1582 126382 1818
rect 126618 1582 127118 1818
rect 127354 1582 127396 1818
rect 153986 1718 154028 1876
rect 154264 1718 158950 1954
rect 159186 1876 223902 1954
rect 159186 1718 159228 1876
rect 153986 1676 159228 1718
rect 223860 1718 223902 1876
rect 224138 1898 585502 1954
rect 585738 1898 586840 2134
rect 224138 1876 586840 1898
rect 224138 1860 224180 1876
rect 585320 1874 585920 1876
rect 224138 1818 226756 1860
rect 224138 1718 226478 1818
rect 126340 1540 127396 1582
rect 223860 1582 226478 1718
rect 226714 1582 226756 1818
rect 223860 1540 226756 1582
rect 161484 1410 161804 1452
rect 161484 1180 161526 1410
rect 4716 1138 10740 1180
rect 4716 902 4758 1138
rect 4994 902 10462 1138
rect 10698 902 10740 1138
rect 4716 860 10740 902
rect 19068 1138 28404 1180
rect 19068 902 19110 1138
rect 19346 902 28126 1138
rect 28362 902 28404 1138
rect 19068 860 28404 902
rect 38940 1138 46252 1180
rect 38940 902 38982 1138
rect 39218 902 46252 1138
rect 38940 860 46252 902
rect 46668 1138 67044 1180
rect 46668 902 46710 1138
rect 46946 902 66766 1138
rect 67002 902 67044 1138
rect 46668 860 67044 902
rect 68932 1138 88388 1180
rect 68932 902 68974 1138
rect 69210 902 88110 1138
rect 88346 902 88388 1138
rect 68932 860 88388 902
rect 91564 1138 146532 1180
rect 91564 902 91606 1138
rect 91842 902 146254 1138
rect 146490 902 146532 1138
rect 91564 860 146532 902
rect 147868 1138 150580 1180
rect 147868 902 147910 1138
rect 148146 902 150302 1138
rect 150538 902 150580 1138
rect 147868 860 150580 902
rect 151410 1138 159596 1180
rect 151410 902 151452 1138
rect 151688 902 159318 1138
rect 159554 902 159596 1138
rect 151410 860 159596 902
rect 160012 1174 161526 1180
rect 161762 1174 161804 1410
rect 174180 1180 176294 1452
rect 201044 1180 203020 1316
rect 160012 1138 161804 1174
rect 160012 902 160054 1138
rect 160290 902 161804 1138
rect 160012 860 161804 902
rect 162220 1138 241292 1180
rect 162220 902 162262 1138
rect 162498 1132 241014 1138
rect 162498 902 174500 1132
rect 162220 860 174500 902
rect 175974 996 241014 1132
rect 175974 860 201364 996
rect 202700 902 241014 996
rect 241250 902 241292 1138
rect 202700 860 241292 902
rect 242076 1138 255092 1316
rect 242076 902 242118 1138
rect 242354 996 254814 1138
rect 242354 902 242396 996
rect 242076 860 242396 902
rect 254772 902 254814 996
rect 255050 902 255092 1138
rect 254772 860 255092 902
rect 256244 1138 265396 1180
rect 256244 902 256286 1138
rect 256522 902 265118 1138
rect 265354 902 265396 1138
rect 256244 860 265396 902
rect 266916 1138 327220 1180
rect 266916 902 266958 1138
rect 267194 902 326942 1138
rect 327178 902 327220 1138
rect 266916 860 327220 902
rect 327636 1138 338996 1180
rect 327636 902 327678 1138
rect 327914 902 338718 1138
rect 338954 902 338996 1138
rect 327636 860 338996 902
rect 339412 1138 350220 1180
rect 339412 902 339454 1138
rect 339690 902 349942 1138
rect 350178 902 350220 1138
rect 339412 860 350220 902
rect 353764 1138 370644 1180
rect 353764 902 353806 1138
rect 354042 902 370366 1138
rect 370602 902 370644 1138
rect 353764 860 370644 902
rect 384124 860 389412 1180
rect 45932 500 46252 860
rect 174916 730 175604 772
rect 174916 500 175326 730
rect 300 458 11108 500
rect 300 222 342 458
rect 578 222 10830 458
rect 11066 222 11108 458
rect 300 180 11108 222
rect 28820 458 39628 500
rect 28820 222 28862 458
rect 29098 222 39350 458
rect 39586 222 39628 458
rect 28820 180 39628 222
rect 45932 458 73668 500
rect 45932 222 73390 458
rect 73626 222 73668 458
rect 45932 180 73668 222
rect 74452 458 92804 500
rect 74452 222 74494 458
rect 74730 222 92526 458
rect 92762 222 92804 458
rect 74452 180 92804 222
rect 93772 458 104028 500
rect 93772 222 93814 458
rect 94050 222 103750 458
rect 103986 222 104028 458
rect 93772 180 104028 222
rect 104444 458 106972 500
rect 104444 222 104486 458
rect 104722 222 106694 458
rect 106930 222 106972 458
rect 104444 180 106972 222
rect 107388 458 123716 500
rect 107388 222 107430 458
rect 107666 222 123438 458
rect 123674 222 123716 458
rect 107388 180 123716 222
rect 134620 458 150948 500
rect 134620 222 134662 458
rect 134898 222 150670 458
rect 150906 222 150948 458
rect 134620 180 150948 222
rect 151364 458 164012 500
rect 151364 222 151406 458
rect 151642 222 163734 458
rect 163970 222 164012 458
rect 151364 180 164012 222
rect 164428 458 169348 500
rect 164428 222 164470 458
rect 164706 222 169070 458
rect 169306 222 169348 458
rect 164428 180 169348 222
rect 169764 494 175326 500
rect 175562 494 175604 730
rect 266180 730 266500 772
rect 169764 458 175604 494
rect 169764 222 169806 458
rect 170042 452 175604 458
rect 176204 458 196948 500
rect 170042 222 175236 452
rect 169764 180 175236 222
rect 176204 222 176246 458
rect 176482 222 196670 458
rect 196906 222 196948 458
rect 176204 180 196948 222
rect 197732 458 217924 500
rect 197732 222 197774 458
rect 198010 222 217646 458
rect 217882 222 217924 458
rect 197732 180 217924 222
rect 224596 458 232644 500
rect 224596 222 224638 458
rect 224874 222 232366 458
rect 232602 222 232644 458
rect 224596 180 232644 222
rect 233060 458 245892 500
rect 233060 222 233102 458
rect 233338 222 245614 458
rect 245850 222 245892 458
rect 233060 180 245892 222
rect 247964 458 265028 500
rect 247964 222 248006 458
rect 248242 222 264750 458
rect 264986 222 265028 458
rect 247964 180 265028 222
rect 266180 494 266222 730
rect 266458 500 266500 730
rect 384124 500 384444 860
rect 266458 494 280300 500
rect 266180 458 280300 494
rect 266180 222 280022 458
rect 280258 222 280300 458
rect 266180 180 280300 222
rect 281452 458 290604 500
rect 281452 222 281494 458
rect 281730 222 290326 458
rect 290562 222 290604 458
rect 281452 180 290604 222
rect 294700 458 336972 500
rect 294700 222 294742 458
rect 294978 222 336694 458
rect 336930 222 336972 458
rect 294700 180 336972 222
rect 343460 458 358316 500
rect 343460 222 343502 458
rect 343738 222 358038 458
rect 358274 222 358316 458
rect 343460 180 358316 222
rect 362964 458 384444 500
rect 362964 222 363006 458
rect 363242 222 384444 458
rect 362964 180 384444 222
rect 389092 500 389412 860
rect 398844 860 411308 1180
rect 414484 1138 419036 1180
rect 414484 902 414526 1138
rect 414762 902 418758 1138
rect 418994 902 419036 1138
rect 414484 860 419036 902
rect 434356 1138 440380 1180
rect 434356 902 440102 1138
rect 440338 902 440380 1138
rect 434356 860 440380 902
rect 450364 1138 463196 1180
rect 450364 902 462918 1138
rect 463154 902 463196 1138
rect 450364 860 463196 902
rect 522124 1138 563844 1180
rect 522124 902 522166 1138
rect 522402 902 563566 1138
rect 563802 902 563844 1138
rect 522124 860 563844 902
rect 398844 500 399164 860
rect 389092 180 399164 500
rect 410988 500 411308 860
rect 410988 458 414252 500
rect 410988 222 413974 458
rect 414210 222 414252 458
rect 410988 180 414252 222
rect 422028 458 430812 500
rect 422028 222 422070 458
rect 422306 222 430534 458
rect 430770 222 430812 458
rect 422028 180 430812 222
rect 434356 458 434676 860
rect 450364 636 450684 860
rect 449812 500 450684 636
rect 434356 222 434398 458
rect 434634 222 434676 458
rect 434356 180 434676 222
rect 449628 458 450684 500
rect 449628 222 449670 458
rect 449906 316 450684 458
rect 468948 458 476996 500
rect 449906 222 450132 316
rect 449628 180 450132 222
rect 468948 222 468990 458
rect 469226 222 476718 458
rect 476954 222 476996 458
rect 468948 180 476996 222
rect 490476 458 504596 500
rect 490476 222 490518 458
rect 490754 222 504318 458
rect 504554 222 504596 458
rect 490476 180 504596 222
rect -1996 -324 -1396 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 585320 -926 585920 -924
rect -2916 -1244 -2316 -1242
rect 586240 -1244 586840 -1242
rect -2916 -1266 586840 -1244
rect -2916 -1502 -2734 -1266
rect -2498 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect -2916 -1586 586840 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect -2916 -1844 586840 -1822
rect -2916 -1846 -2316 -1844
rect 586240 -1846 586840 -1844
rect -3836 -2164 -3236 -2162
rect 587160 -2164 587760 -2162
rect -3836 -2186 587760 -2164
rect -3836 -2422 -3654 -2186
rect -3418 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect -3836 -2506 587760 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect -3836 -2764 587760 -2742
rect -3836 -2766 -3236 -2764
rect 587160 -2766 587760 -2764
rect -4756 -3084 -4156 -3082
rect 588080 -3084 588680 -3082
rect -4756 -3106 588680 -3084
rect -4756 -3342 -4574 -3106
rect -4338 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect -4756 -3426 588680 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect -4756 -3684 588680 -3662
rect -4756 -3686 -4156 -3684
rect 588080 -3686 588680 -3684
rect -5676 -4004 -5076 -4002
rect 589000 -4004 589600 -4002
rect -5676 -4026 589600 -4004
rect -5676 -4262 -5494 -4026
rect -5258 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect -5676 -4346 589600 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect -5676 -4604 589600 -4582
rect -5676 -4606 -5076 -4604
rect 589000 -4606 589600 -4604
rect -6596 -4924 -5996 -4922
rect 589920 -4924 590520 -4922
rect -6596 -4946 590520 -4924
rect -6596 -5182 -6414 -4946
rect -6178 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect -6596 -5266 590520 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect -6596 -5524 590520 -5502
rect -6596 -5526 -5996 -5524
rect 589920 -5526 590520 -5524
rect -7516 -5844 -6916 -5842
rect 590840 -5844 591440 -5842
rect -7516 -5866 591440 -5844
rect -7516 -6102 -7334 -5866
rect -7098 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect -7516 -6186 591440 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect -7516 -6444 591440 -6422
rect -7516 -6446 -6916 -6444
rect 590840 -6446 591440 -6444
rect -8436 -6764 -7836 -6762
rect 591760 -6764 592360 -6762
rect -8436 -6786 592360 -6764
rect -8436 -7022 -8254 -6786
rect -8018 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect -8436 -7106 592360 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect -8436 -7364 592360 -7342
rect -8436 -7366 -7836 -7364
rect 591760 -7366 592360 -7364
use fpga  fpga250
timestamp 1607933928
transform 1 0 1000 0 1 1000
box 0 0 570000 680000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2916 -1844 586840 -1244 8 vssd1
port 637 nsew default input
rlabel metal5 s -3836 -2764 587760 -2164 8 vccd2
port 638 nsew default input
rlabel metal5 s -4756 -3684 588680 -3084 8 vssd2
port 639 nsew default input
rlabel metal5 s -5676 -4604 589600 -4004 8 vdda1
port 640 nsew default input
rlabel metal5 s -6596 -5524 590520 -4924 8 vssa1
port 641 nsew default input
rlabel metal5 s -7516 -6444 591440 -5844 8 vdda2
port 642 nsew default input
rlabel metal5 s -8436 -7364 592360 -6764 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga
  CLASS BLOCK ;
  FOREIGN fpga ;
  ORIGIN 0.000 0.000 ;
  SIZE 2850.000 BY 3400.000 ;
  PIN gpio_east[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 54.440 2850.000 55.040 ;
    END
  END gpio_east[0]
  PIN gpio_east[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 163.920 2850.000 164.520 ;
    END
  END gpio_east[1]
  PIN gpio_east[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 273.400 2850.000 274.000 ;
    END
  END gpio_east[2]
  PIN gpio_east[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 382.880 2850.000 383.480 ;
    END
  END gpio_east[3]
  PIN gpio_east[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 493.040 2850.000 493.640 ;
    END
  END gpio_east[4]
  PIN gpio_east[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 602.520 2850.000 603.120 ;
    END
  END gpio_east[5]
  PIN gpio_east[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 712.000 2850.000 712.600 ;
    END
  END gpio_east[6]
  PIN gpio_east[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 822.160 2850.000 822.760 ;
    END
  END gpio_east[7]
  PIN gpio_east[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 931.640 2850.000 932.240 ;
    END
  END gpio_east[8]
  PIN gpio_east[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1041.120 2850.000 1041.720 ;
    END
  END gpio_east[9]
  PIN gpio_north[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 54.830 3396.000 55.110 3400.000 ;
    END
  END gpio_north[0]
  PIN gpio_north[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 164.310 3396.000 164.590 3400.000 ;
    END
  END gpio_north[1]
  PIN gpio_north[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 273.790 3396.000 274.070 3400.000 ;
    END
  END gpio_north[2]
  PIN gpio_north[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 383.270 3396.000 383.550 3400.000 ;
    END
  END gpio_north[3]
  PIN gpio_north[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 493.210 3396.000 493.490 3400.000 ;
    END
  END gpio_north[4]
  PIN gpio_north[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 602.690 3396.000 602.970 3400.000 ;
    END
  END gpio_north[5]
  PIN gpio_north[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 712.170 3396.000 712.450 3400.000 ;
    END
  END gpio_north[6]
  PIN gpio_north[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 822.110 3396.000 822.390 3400.000 ;
    END
  END gpio_north[7]
  PIN gpio_north[8]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 931.590 3396.000 931.870 3400.000 ;
    END
  END gpio_north[8]
  PIN gpio_north[9]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1041.070 3396.000 1041.350 3400.000 ;
    END
  END gpio_north[9]
  PIN gpio_south[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END gpio_south[0]
  PIN gpio_south[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END gpio_south[1]
  PIN gpio_south[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END gpio_south[2]
  PIN gpio_south[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 177.650 0.000 177.930 4.000 ;
    END
  END gpio_south[3]
  PIN gpio_south[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END gpio_south[4]
  PIN gpio_south[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END gpio_south[5]
  PIN gpio_south[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 330.370 0.000 330.650 4.000 ;
    END
  END gpio_south[6]
  PIN gpio_south[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 381.430 0.000 381.710 4.000 ;
    END
  END gpio_south[7]
  PIN gpio_west[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END gpio_west[0]
  PIN gpio_west[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.920 4.000 164.520 ;
    END
  END gpio_west[1]
  PIN gpio_west[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END gpio_west[2]
  PIN gpio_west[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.880 4.000 383.480 ;
    END
  END gpio_west[3]
  PIN gpio_west[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END gpio_west[4]
  PIN gpio_west[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 602.520 4.000 603.120 ;
    END
  END gpio_west[5]
  PIN gpio_west[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 712.000 4.000 712.600 ;
    END
  END gpio_west[6]
  PIN gpio_west[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 822.160 4.000 822.760 ;
    END
  END gpio_west[7]
  PIN gpio_west[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 931.640 4.000 932.240 ;
    END
  END gpio_west[8]
  PIN gpio_west[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1041.120 4.000 1041.720 ;
    END
  END gpio_west[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1150.600 2850.000 1151.200 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1260.760 2850.000 1261.360 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1151.010 3396.000 1151.290 3400.000 ;
    END
  END wbs_ack_o
  PIN wbs_addr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1260.490 3396.000 1260.770 3400.000 ;
    END
  END wbs_addr_i[0]
  PIN wbs_addr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1479.910 3396.000 1480.190 3400.000 ;
    END
  END wbs_addr_i[10]
  PIN wbs_addr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2163.010 0.000 2163.290 4.000 ;
    END
  END wbs_addr_i[11]
  PIN wbs_addr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2213.610 0.000 2213.890 4.000 ;
    END
  END wbs_addr_i[12]
  PIN wbs_addr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1589.880 2850.000 1590.480 ;
    END
  END wbs_addr_i[13]
  PIN wbs_addr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2264.670 0.000 2264.950 4.000 ;
    END
  END wbs_addr_i[14]
  PIN wbs_addr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1589.880 4.000 1590.480 ;
    END
  END wbs_addr_i[15]
  PIN wbs_addr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1699.360 2850.000 1699.960 ;
    END
  END wbs_addr_i[16]
  PIN wbs_addr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1808.840 2850.000 1809.440 ;
    END
  END wbs_addr_i[17]
  PIN wbs_addr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2315.270 0.000 2315.550 4.000 ;
    END
  END wbs_addr_i[18]
  PIN wbs_addr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2366.330 0.000 2366.610 4.000 ;
    END
  END wbs_addr_i[19]
  PIN wbs_addr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1150.600 4.000 1151.200 ;
    END
  END wbs_addr_i[1]
  PIN wbs_addr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1918.320 2850.000 1918.920 ;
    END
  END wbs_addr_i[20]
  PIN wbs_addr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2417.390 0.000 2417.670 4.000 ;
    END
  END wbs_addr_i[21]
  PIN wbs_addr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2028.480 2850.000 2029.080 ;
    END
  END wbs_addr_i[22]
  PIN wbs_addr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2137.960 2850.000 2138.560 ;
    END
  END wbs_addr_i[23]
  PIN wbs_addr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2467.990 0.000 2468.270 4.000 ;
    END
  END wbs_addr_i[24]
  PIN wbs_addr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2247.440 2850.000 2248.040 ;
    END
  END wbs_addr_i[25]
  PIN wbs_addr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1589.390 3396.000 1589.670 3400.000 ;
    END
  END wbs_addr_i[26]
  PIN wbs_addr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1699.360 4.000 1699.960 ;
    END
  END wbs_addr_i[27]
  PIN wbs_addr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1698.870 3396.000 1699.150 3400.000 ;
    END
  END wbs_addr_i[28]
  PIN wbs_addr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1808.840 4.000 1809.440 ;
    END
  END wbs_addr_i[29]
  PIN wbs_addr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1369.970 3396.000 1370.250 3400.000 ;
    END
  END wbs_addr_i[2]
  PIN wbs_addr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2357.600 2850.000 2358.200 ;
    END
  END wbs_addr_i[30]
  PIN wbs_addr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1808.350 3396.000 1808.630 3400.000 ;
    END
  END wbs_addr_i[31]
  PIN wbs_addr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1370.240 2850.000 1370.840 ;
    END
  END wbs_addr_i[3]
  PIN wbs_addr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1260.760 4.000 1261.360 ;
    END
  END wbs_addr_i[4]
  PIN wbs_addr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1479.720 2850.000 1480.320 ;
    END
  END wbs_addr_i[5]
  PIN wbs_addr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1370.240 4.000 1370.840 ;
    END
  END wbs_addr_i[6]
  PIN wbs_addr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2060.890 0.000 2061.170 4.000 ;
    END
  END wbs_addr_i[7]
  PIN wbs_addr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1479.720 4.000 1480.320 ;
    END
  END wbs_addr_i[8]
  PIN wbs_addr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2111.950 0.000 2112.230 4.000 ;
    END
  END wbs_addr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1918.290 3396.000 1918.570 3400.000 ;
    END
  END wbs_cyc_i
  PIN wbs_data_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2519.050 0.000 2519.330 4.000 ;
    END
  END wbs_data_i[0]
  PIN wbs_data_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2027.770 3396.000 2028.050 3400.000 ;
    END
  END wbs_data_i[10]
  PIN wbs_data_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2722.830 0.000 2723.110 4.000 ;
    END
  END wbs_data_i[11]
  PIN wbs_data_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2137.250 3396.000 2137.530 3400.000 ;
    END
  END wbs_data_i[12]
  PIN wbs_data_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2247.190 3396.000 2247.470 3400.000 ;
    END
  END wbs_data_i[13]
  PIN wbs_data_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2686.040 2850.000 2686.640 ;
    END
  END wbs_data_i[14]
  PIN wbs_data_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2357.600 4.000 2358.200 ;
    END
  END wbs_data_i[15]
  PIN wbs_data_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2467.080 4.000 2467.680 ;
    END
  END wbs_data_i[16]
  PIN wbs_data_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2576.560 4.000 2577.160 ;
    END
  END wbs_data_i[17]
  PIN wbs_data_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2796.200 2850.000 2796.800 ;
    END
  END wbs_data_i[18]
  PIN wbs_data_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2686.040 4.000 2686.640 ;
    END
  END wbs_data_i[19]
  PIN wbs_data_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2570.110 0.000 2570.390 4.000 ;
    END
  END wbs_data_i[1]
  PIN wbs_data_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2356.670 3396.000 2356.950 3400.000 ;
    END
  END wbs_data_i[20]
  PIN wbs_data_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2796.200 4.000 2796.800 ;
    END
  END wbs_data_i[21]
  PIN wbs_data_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2905.680 4.000 2906.280 ;
    END
  END wbs_data_i[22]
  PIN wbs_data_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3015.160 4.000 3015.760 ;
    END
  END wbs_data_i[23]
  PIN wbs_data_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3125.320 4.000 3125.920 ;
    END
  END wbs_data_i[24]
  PIN wbs_data_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2466.150 3396.000 2466.430 3400.000 ;
    END
  END wbs_data_i[25]
  PIN wbs_data_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2905.680 2850.000 2906.280 ;
    END
  END wbs_data_i[26]
  PIN wbs_data_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2576.090 3396.000 2576.370 3400.000 ;
    END
  END wbs_data_i[27]
  PIN wbs_data_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2685.570 3396.000 2685.850 3400.000 ;
    END
  END wbs_data_i[28]
  PIN wbs_data_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2795.050 3396.000 2795.330 3400.000 ;
    END
  END wbs_data_i[29]
  PIN wbs_data_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1918.320 4.000 1918.920 ;
    END
  END wbs_data_i[2]
  PIN wbs_data_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 3015.160 2850.000 3015.760 ;
    END
  END wbs_data_i[30]
  PIN wbs_data_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 3125.320 2850.000 3125.920 ;
    END
  END wbs_data_i[31]
  PIN wbs_data_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2467.080 2850.000 2467.680 ;
    END
  END wbs_data_i[3]
  PIN wbs_data_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2028.480 4.000 2029.080 ;
    END
  END wbs_data_i[4]
  PIN wbs_data_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2620.710 0.000 2620.990 4.000 ;
    END
  END wbs_data_i[5]
  PIN wbs_data_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2576.560 2850.000 2577.160 ;
    END
  END wbs_data_i[6]
  PIN wbs_data_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2137.960 4.000 2138.560 ;
    END
  END wbs_data_i[7]
  PIN wbs_data_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2671.770 0.000 2672.050 4.000 ;
    END
  END wbs_data_i[8]
  PIN wbs_data_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2247.440 4.000 2248.040 ;
    END
  END wbs_data_i[9]
  PIN wbs_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 432.490 0.000 432.770 4.000 ;
    END
  END wbs_data_o[0]
  PIN wbs_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 941.250 0.000 941.530 4.000 ;
    END
  END wbs_data_o[10]
  PIN wbs_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 992.310 0.000 992.590 4.000 ;
    END
  END wbs_data_o[11]
  PIN wbs_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1042.910 0.000 1043.190 4.000 ;
    END
  END wbs_data_o[12]
  PIN wbs_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1093.970 0.000 1094.250 4.000 ;
    END
  END wbs_data_o[13]
  PIN wbs_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1145.030 0.000 1145.310 4.000 ;
    END
  END wbs_data_o[14]
  PIN wbs_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1195.630 0.000 1195.910 4.000 ;
    END
  END wbs_data_o[15]
  PIN wbs_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1246.690 0.000 1246.970 4.000 ;
    END
  END wbs_data_o[16]
  PIN wbs_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1297.750 0.000 1298.030 4.000 ;
    END
  END wbs_data_o[17]
  PIN wbs_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1348.350 0.000 1348.630 4.000 ;
    END
  END wbs_data_o[18]
  PIN wbs_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1399.410 0.000 1399.690 4.000 ;
    END
  END wbs_data_o[19]
  PIN wbs_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END wbs_data_o[1]
  PIN wbs_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1450.470 0.000 1450.750 4.000 ;
    END
  END wbs_data_o[20]
  PIN wbs_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1501.070 0.000 1501.350 4.000 ;
    END
  END wbs_data_o[21]
  PIN wbs_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1552.130 0.000 1552.410 4.000 ;
    END
  END wbs_data_o[22]
  PIN wbs_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1602.730 0.000 1603.010 4.000 ;
    END
  END wbs_data_o[23]
  PIN wbs_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1653.790 0.000 1654.070 4.000 ;
    END
  END wbs_data_o[24]
  PIN wbs_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1704.850 0.000 1705.130 4.000 ;
    END
  END wbs_data_o[25]
  PIN wbs_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1755.450 0.000 1755.730 4.000 ;
    END
  END wbs_data_o[26]
  PIN wbs_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1806.510 0.000 1806.790 4.000 ;
    END
  END wbs_data_o[27]
  PIN wbs_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1857.570 0.000 1857.850 4.000 ;
    END
  END wbs_data_o[28]
  PIN wbs_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1908.170 0.000 1908.450 4.000 ;
    END
  END wbs_data_o[29]
  PIN wbs_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 534.150 0.000 534.430 4.000 ;
    END
  END wbs_data_o[2]
  PIN wbs_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1959.230 0.000 1959.510 4.000 ;
    END
  END wbs_data_o[30]
  PIN wbs_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2010.290 0.000 2010.570 4.000 ;
    END
  END wbs_data_o[31]
  PIN wbs_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 585.210 0.000 585.490 4.000 ;
    END
  END wbs_data_o[3]
  PIN wbs_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 635.810 0.000 636.090 4.000 ;
    END
  END wbs_data_o[4]
  PIN wbs_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 686.870 0.000 687.150 4.000 ;
    END
  END wbs_data_o[5]
  PIN wbs_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 737.930 0.000 738.210 4.000 ;
    END
  END wbs_data_o[6]
  PIN wbs_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 788.530 0.000 788.810 4.000 ;
    END
  END wbs_data_o[7]
  PIN wbs_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 839.590 0.000 839.870 4.000 ;
    END
  END wbs_data_o[8]
  PIN wbs_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 890.190 0.000 890.470 4.000 ;
    END
  END wbs_data_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 3234.800 2850.000 3235.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3234.800 4.000 3235.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 3344.280 2850.000 3344.880 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2773.430 0.000 2773.710 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2824.490 0.000 2824.770 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3344.280 4.000 3344.880 ;
    END
  END wbs_we_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 2844.180 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 64.785 2844.180 66.385 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2844.180 3389.205 ;
      LAYER met1 ;
        RECT 5.520 4.460 2844.180 3389.360 ;
      LAYER met2 ;
        RECT 14.350 3395.720 54.550 3396.000 ;
        RECT 55.390 3395.720 164.030 3396.000 ;
        RECT 164.870 3395.720 273.510 3396.000 ;
        RECT 274.350 3395.720 382.990 3396.000 ;
        RECT 383.830 3395.720 492.930 3396.000 ;
        RECT 493.770 3395.720 602.410 3396.000 ;
        RECT 603.250 3395.720 711.890 3396.000 ;
        RECT 712.730 3395.720 821.830 3396.000 ;
        RECT 822.670 3395.720 931.310 3396.000 ;
        RECT 932.150 3395.720 1040.790 3396.000 ;
        RECT 1041.630 3395.720 1150.730 3396.000 ;
        RECT 1151.570 3395.720 1260.210 3396.000 ;
        RECT 1261.050 3395.720 1369.690 3396.000 ;
        RECT 1370.530 3395.720 1479.630 3396.000 ;
        RECT 1480.470 3395.720 1589.110 3396.000 ;
        RECT 1589.950 3395.720 1698.590 3396.000 ;
        RECT 1699.430 3395.720 1808.070 3396.000 ;
        RECT 1808.910 3395.720 1918.010 3396.000 ;
        RECT 1918.850 3395.720 2027.490 3396.000 ;
        RECT 2028.330 3395.720 2136.970 3396.000 ;
        RECT 2137.810 3395.720 2246.910 3396.000 ;
        RECT 2247.750 3395.720 2356.390 3396.000 ;
        RECT 2357.230 3395.720 2465.870 3396.000 ;
        RECT 2466.710 3395.720 2575.810 3396.000 ;
        RECT 2576.650 3395.720 2685.290 3396.000 ;
        RECT 2686.130 3395.720 2794.770 3396.000 ;
        RECT 2795.610 3395.720 2835.810 3396.000 ;
        RECT 14.350 4.280 2835.810 3395.720 ;
        RECT 14.350 4.000 25.110 4.280 ;
        RECT 25.950 4.000 75.710 4.280 ;
        RECT 76.550 4.000 126.770 4.280 ;
        RECT 127.610 4.000 177.370 4.280 ;
        RECT 178.210 4.000 228.430 4.280 ;
        RECT 229.270 4.000 279.490 4.280 ;
        RECT 280.330 4.000 330.090 4.280 ;
        RECT 330.930 4.000 381.150 4.280 ;
        RECT 381.990 4.000 432.210 4.280 ;
        RECT 433.050 4.000 482.810 4.280 ;
        RECT 483.650 4.000 533.870 4.280 ;
        RECT 534.710 4.000 584.930 4.280 ;
        RECT 585.770 4.000 635.530 4.280 ;
        RECT 636.370 4.000 686.590 4.280 ;
        RECT 687.430 4.000 737.650 4.280 ;
        RECT 738.490 4.000 788.250 4.280 ;
        RECT 789.090 4.000 839.310 4.280 ;
        RECT 840.150 4.000 889.910 4.280 ;
        RECT 890.750 4.000 940.970 4.280 ;
        RECT 941.810 4.000 992.030 4.280 ;
        RECT 992.870 4.000 1042.630 4.280 ;
        RECT 1043.470 4.000 1093.690 4.280 ;
        RECT 1094.530 4.000 1144.750 4.280 ;
        RECT 1145.590 4.000 1195.350 4.280 ;
        RECT 1196.190 4.000 1246.410 4.280 ;
        RECT 1247.250 4.000 1297.470 4.280 ;
        RECT 1298.310 4.000 1348.070 4.280 ;
        RECT 1348.910 4.000 1399.130 4.280 ;
        RECT 1399.970 4.000 1450.190 4.280 ;
        RECT 1451.030 4.000 1500.790 4.280 ;
        RECT 1501.630 4.000 1551.850 4.280 ;
        RECT 1552.690 4.000 1602.450 4.280 ;
        RECT 1603.290 4.000 1653.510 4.280 ;
        RECT 1654.350 4.000 1704.570 4.280 ;
        RECT 1705.410 4.000 1755.170 4.280 ;
        RECT 1756.010 4.000 1806.230 4.280 ;
        RECT 1807.070 4.000 1857.290 4.280 ;
        RECT 1858.130 4.000 1907.890 4.280 ;
        RECT 1908.730 4.000 1958.950 4.280 ;
        RECT 1959.790 4.000 2010.010 4.280 ;
        RECT 2010.850 4.000 2060.610 4.280 ;
        RECT 2061.450 4.000 2111.670 4.280 ;
        RECT 2112.510 4.000 2162.730 4.280 ;
        RECT 2163.570 4.000 2213.330 4.280 ;
        RECT 2214.170 4.000 2264.390 4.280 ;
        RECT 2265.230 4.000 2314.990 4.280 ;
        RECT 2315.830 4.000 2366.050 4.280 ;
        RECT 2366.890 4.000 2417.110 4.280 ;
        RECT 2417.950 4.000 2467.710 4.280 ;
        RECT 2468.550 4.000 2518.770 4.280 ;
        RECT 2519.610 4.000 2569.830 4.280 ;
        RECT 2570.670 4.000 2620.430 4.280 ;
        RECT 2621.270 4.000 2671.490 4.280 ;
        RECT 2672.330 4.000 2722.550 4.280 ;
        RECT 2723.390 4.000 2773.150 4.280 ;
        RECT 2773.990 4.000 2824.210 4.280 ;
        RECT 2825.050 4.000 2835.810 4.280 ;
      LAYER met3 ;
        RECT 4.000 3345.280 2846.000 3395.745 ;
        RECT 4.400 3343.880 2845.600 3345.280 ;
        RECT 4.000 3235.800 2846.000 3343.880 ;
        RECT 4.400 3234.400 2845.600 3235.800 ;
        RECT 4.000 3126.320 2846.000 3234.400 ;
        RECT 4.400 3124.920 2845.600 3126.320 ;
        RECT 4.000 3016.160 2846.000 3124.920 ;
        RECT 4.400 3014.760 2845.600 3016.160 ;
        RECT 4.000 2906.680 2846.000 3014.760 ;
        RECT 4.400 2905.280 2845.600 2906.680 ;
        RECT 4.000 2797.200 2846.000 2905.280 ;
        RECT 4.400 2795.800 2845.600 2797.200 ;
        RECT 4.000 2687.040 2846.000 2795.800 ;
        RECT 4.400 2685.640 2845.600 2687.040 ;
        RECT 4.000 2577.560 2846.000 2685.640 ;
        RECT 4.400 2576.160 2845.600 2577.560 ;
        RECT 4.000 2468.080 2846.000 2576.160 ;
        RECT 4.400 2466.680 2845.600 2468.080 ;
        RECT 4.000 2358.600 2846.000 2466.680 ;
        RECT 4.400 2357.200 2845.600 2358.600 ;
        RECT 4.000 2248.440 2846.000 2357.200 ;
        RECT 4.400 2247.040 2845.600 2248.440 ;
        RECT 4.000 2138.960 2846.000 2247.040 ;
        RECT 4.400 2137.560 2845.600 2138.960 ;
        RECT 4.000 2029.480 2846.000 2137.560 ;
        RECT 4.400 2028.080 2845.600 2029.480 ;
        RECT 4.000 1919.320 2846.000 2028.080 ;
        RECT 4.400 1917.920 2845.600 1919.320 ;
        RECT 4.000 1809.840 2846.000 1917.920 ;
        RECT 4.400 1808.440 2845.600 1809.840 ;
        RECT 4.000 1700.360 2846.000 1808.440 ;
        RECT 4.400 1698.960 2845.600 1700.360 ;
        RECT 4.000 1590.880 2846.000 1698.960 ;
        RECT 4.400 1589.480 2845.600 1590.880 ;
        RECT 4.000 1480.720 2846.000 1589.480 ;
        RECT 4.400 1479.320 2845.600 1480.720 ;
        RECT 4.000 1371.240 2846.000 1479.320 ;
        RECT 4.400 1369.840 2845.600 1371.240 ;
        RECT 4.000 1261.760 2846.000 1369.840 ;
        RECT 4.400 1260.360 2845.600 1261.760 ;
        RECT 4.000 1151.600 2846.000 1260.360 ;
        RECT 4.400 1150.200 2845.600 1151.600 ;
        RECT 4.000 1042.120 2846.000 1150.200 ;
        RECT 4.400 1040.720 2845.600 1042.120 ;
        RECT 4.000 932.640 2846.000 1040.720 ;
        RECT 4.400 931.240 2845.600 932.640 ;
        RECT 4.000 823.160 2846.000 931.240 ;
        RECT 4.400 821.760 2845.600 823.160 ;
        RECT 4.000 713.000 2846.000 821.760 ;
        RECT 4.400 711.600 2845.600 713.000 ;
        RECT 4.000 603.520 2846.000 711.600 ;
        RECT 4.400 602.120 2845.600 603.520 ;
        RECT 4.000 494.040 2846.000 602.120 ;
        RECT 4.400 492.640 2845.600 494.040 ;
        RECT 4.000 383.880 2846.000 492.640 ;
        RECT 4.400 382.480 2845.600 383.880 ;
        RECT 4.000 274.400 2846.000 382.480 ;
        RECT 4.400 273.000 2845.600 274.400 ;
        RECT 4.000 164.920 2846.000 273.000 ;
        RECT 4.400 163.520 2845.600 164.920 ;
        RECT 4.000 55.440 2846.000 163.520 ;
        RECT 4.400 54.040 2845.600 55.440 ;
        RECT 4.000 10.715 2846.000 54.040 ;
      LAYER met4 ;
        RECT 21.040 10.640 2787.440 3389.360 ;
      LAYER met5 ;
        RECT 5.520 103.080 2844.180 3359.755 ;
  END
END fpga
END LIBRARY


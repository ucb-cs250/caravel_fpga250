magic
tech sky130A
magscale 1 2
timestamp 1608086250
<< locali >>
rect 6193 599063 6227 608549
rect 6193 591787 6227 598893
rect 6193 579751 6227 589237
rect 6101 569959 6135 579581
rect 6101 560303 6135 565097
rect 6101 550647 6135 553401
rect 6101 540991 6135 550477
rect 6009 531335 6043 534089
rect 6101 483123 6135 487781
rect 5917 473467 5951 476153
rect 6101 456739 6135 471937
rect 6101 444499 6135 452149
rect 6101 434775 6135 444329
rect 6101 425119 6135 431613
rect 6193 415463 6227 425017
rect 6101 405739 6135 410533
rect 6193 376771 6227 386325
rect 6193 347871 6227 357221
rect 6377 327811 6411 336685
rect 6193 309247 6227 318733
rect 6193 301971 6227 309077
rect 6193 289935 6227 299421
rect 6193 282795 6227 289765
rect 6193 270623 6227 280109
rect 6193 263347 6227 270453
rect 6193 251311 6227 260797
rect 6101 241519 6135 251141
rect 6101 231863 6135 236657
rect 6101 222207 6135 224961
rect 6101 212551 6135 222037
rect 6101 154683 6135 159341
rect 6101 106335 6135 115889
rect 6101 96679 6135 101405
rect 6193 87023 6227 96577
rect 6101 77299 6135 82093
rect 6193 48331 6227 57885
rect 6193 38675 6227 47413
rect 6285 19363 6319 28917
rect 11529 7735 11563 7837
rect 45569 7463 45603 7633
rect 13737 3791 13771 3961
<< viali >>
rect 6193 608549 6227 608583
rect 6193 599029 6227 599063
rect 6193 598893 6227 598927
rect 6193 591753 6227 591787
rect 6193 589237 6227 589271
rect 6193 579717 6227 579751
rect 6101 579581 6135 579615
rect 6101 569925 6135 569959
rect 6101 565097 6135 565131
rect 6101 560269 6135 560303
rect 6101 553401 6135 553435
rect 6101 550613 6135 550647
rect 6101 550477 6135 550511
rect 6101 540957 6135 540991
rect 6009 534089 6043 534123
rect 6009 531301 6043 531335
rect 6101 487781 6135 487815
rect 6101 483089 6135 483123
rect 5917 476153 5951 476187
rect 5917 473433 5951 473467
rect 6101 471937 6135 471971
rect 6101 456705 6135 456739
rect 6101 452149 6135 452183
rect 6101 444465 6135 444499
rect 6101 444329 6135 444363
rect 6101 434741 6135 434775
rect 6101 431613 6135 431647
rect 6101 425085 6135 425119
rect 6193 425017 6227 425051
rect 6193 415429 6227 415463
rect 6101 410533 6135 410567
rect 6101 405705 6135 405739
rect 6193 386325 6227 386359
rect 6193 376737 6227 376771
rect 6193 357221 6227 357255
rect 6193 347837 6227 347871
rect 6377 336685 6411 336719
rect 6377 327777 6411 327811
rect 6193 318733 6227 318767
rect 6193 309213 6227 309247
rect 6193 309077 6227 309111
rect 6193 301937 6227 301971
rect 6193 299421 6227 299455
rect 6193 289901 6227 289935
rect 6193 289765 6227 289799
rect 6193 282761 6227 282795
rect 6193 280109 6227 280143
rect 6193 270589 6227 270623
rect 6193 270453 6227 270487
rect 6193 263313 6227 263347
rect 6193 260797 6227 260831
rect 6193 251277 6227 251311
rect 6101 251141 6135 251175
rect 6101 241485 6135 241519
rect 6101 236657 6135 236691
rect 6101 231829 6135 231863
rect 6101 224961 6135 224995
rect 6101 222173 6135 222207
rect 6101 222037 6135 222071
rect 6101 212517 6135 212551
rect 6101 159341 6135 159375
rect 6101 154649 6135 154683
rect 6101 115889 6135 115923
rect 6101 106301 6135 106335
rect 6101 101405 6135 101439
rect 6101 96645 6135 96679
rect 6193 96577 6227 96611
rect 6193 86989 6227 87023
rect 6101 82093 6135 82127
rect 6101 77265 6135 77299
rect 6193 57885 6227 57919
rect 6193 48297 6227 48331
rect 6193 47413 6227 47447
rect 6193 38641 6227 38675
rect 6285 28917 6319 28951
rect 6285 19329 6319 19363
rect 11529 7837 11563 7871
rect 11529 7701 11563 7735
rect 45569 7633 45603 7667
rect 45569 7429 45603 7463
rect 13737 3961 13771 3995
rect 13737 3757 13771 3791
<< metal1 >>
rect 164142 700612 164148 700664
rect 164200 700652 164206 700664
rect 235166 700652 235172 700664
rect 164200 700624 235172 700652
rect 164200 700612 164206 700624
rect 235166 700612 235172 700624
rect 235224 700612 235230 700664
rect 135162 700544 135168 700596
rect 135220 700584 135226 700596
rect 300118 700584 300124 700596
rect 135220 700556 300124 700584
rect 135220 700544 135226 700556
rect 300118 700544 300124 700556
rect 300176 700544 300182 700596
rect 105446 700476 105452 700528
rect 105504 700516 105510 700528
rect 106182 700516 106188 700528
rect 105504 700488 106188 700516
rect 105504 700476 105510 700488
rect 106182 700476 106188 700488
rect 106240 700476 106246 700528
rect 107562 700476 107568 700528
rect 107620 700516 107626 700528
rect 364978 700516 364984 700528
rect 107620 700488 364984 700516
rect 107620 700476 107626 700488
rect 364978 700476 364984 700488
rect 365036 700476 365042 700528
rect 40494 700408 40500 700460
rect 40552 700448 40558 700460
rect 41322 700448 41328 700460
rect 40552 700420 41328 700448
rect 40552 700408 40558 700420
rect 41322 700408 41328 700420
rect 41380 700408 41386 700460
rect 78582 700408 78588 700460
rect 78640 700448 78646 700460
rect 429838 700448 429844 700460
rect 78640 700420 429844 700448
rect 78640 700408 78646 700420
rect 429838 700408 429844 700420
rect 429896 700408 429902 700460
rect 49602 700340 49608 700392
rect 49660 700380 49666 700392
rect 494790 700380 494796 700392
rect 49660 700352 494796 700380
rect 49660 700340 49666 700352
rect 494790 700340 494796 700352
rect 494848 700340 494854 700392
rect 22002 700272 22008 700324
rect 22060 700312 22066 700324
rect 559650 700312 559656 700324
rect 22060 700284 559656 700312
rect 22060 700272 22066 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 170306 699660 170312 699712
rect 170364 699700 170370 699712
rect 171042 699700 171048 699712
rect 170364 699672 171048 699700
rect 170364 699660 170370 699672
rect 171042 699660 171048 699672
rect 171100 699660 171106 699712
rect 21174 689528 21180 689580
rect 21232 689568 21238 689580
rect 22002 689568 22008 689580
rect 21232 689540 22008 689568
rect 21232 689528 21238 689540
rect 22002 689528 22008 689540
rect 22060 689528 22066 689580
rect 106642 689528 106648 689580
rect 106700 689568 106706 689580
rect 107562 689568 107568 689580
rect 106700 689540 107568 689568
rect 106700 689528 106706 689540
rect 107562 689528 107568 689540
rect 107620 689528 107626 689580
rect 171042 689392 171048 689444
rect 171100 689432 171106 689444
rect 192110 689432 192116 689444
rect 171100 689404 192116 689432
rect 171100 689392 171106 689404
rect 192110 689392 192116 689404
rect 192168 689392 192174 689444
rect 106182 689324 106188 689376
rect 106240 689364 106246 689376
rect 220630 689364 220636 689376
rect 106240 689336 220636 689364
rect 106240 689324 106246 689336
rect 220630 689324 220636 689336
rect 220688 689324 220694 689376
rect 41322 689256 41328 689308
rect 41380 689296 41386 689308
rect 249150 689296 249156 689308
rect 41380 689268 249156 689296
rect 41380 689256 41386 689268
rect 249150 689256 249156 689268
rect 249208 689256 249214 689308
rect 9306 689120 9312 689172
rect 9364 689160 9370 689172
rect 306190 689160 306196 689172
rect 9364 689132 306196 689160
rect 9364 689120 9370 689132
rect 306190 689120 306196 689132
rect 306248 689120 306254 689172
rect 277670 689052 277676 689104
rect 277728 689092 277734 689104
rect 576118 689092 576124 689104
rect 277728 689064 576124 689092
rect 277728 689052 277734 689064
rect 576118 689052 576124 689064
rect 576176 689052 576182 689104
rect 9582 688984 9588 689036
rect 9640 689024 9646 689036
rect 334618 689024 334624 689036
rect 9640 688996 334624 689024
rect 9640 688984 9646 688996
rect 334618 688984 334624 688996
rect 334676 688984 334682 689036
rect 9030 688916 9036 688968
rect 9088 688956 9094 688968
rect 363138 688956 363144 688968
rect 9088 688928 363144 688956
rect 9088 688916 9094 688928
rect 363138 688916 363144 688928
rect 363196 688916 363202 688968
rect 9490 688848 9496 688900
rect 9548 688888 9554 688900
rect 448698 688888 448704 688900
rect 9548 688860 448704 688888
rect 9548 688848 9554 688860
rect 448698 688848 448704 688860
rect 448756 688848 448762 688900
rect 9122 688780 9128 688832
rect 9180 688820 9186 688832
rect 477126 688820 477132 688832
rect 9180 688792 477132 688820
rect 9180 688780 9186 688792
rect 477126 688780 477132 688792
rect 477184 688780 477190 688832
rect 9214 688712 9220 688764
rect 9272 688752 9278 688764
rect 505646 688752 505652 688764
rect 9272 688724 505652 688752
rect 9272 688712 9278 688724
rect 505646 688712 505652 688724
rect 505704 688712 505710 688764
rect 9398 688644 9404 688696
rect 9456 688684 9462 688696
rect 562686 688684 562692 688696
rect 9456 688656 562692 688684
rect 9456 688644 9462 688656
rect 562686 688644 562692 688656
rect 562744 688644 562750 688696
rect 3510 681708 3516 681760
rect 3568 681748 3574 681760
rect 7558 681748 7564 681760
rect 3568 681720 7564 681748
rect 3568 681708 3574 681720
rect 7558 681708 7564 681720
rect 7616 681708 7622 681760
rect 3142 616836 3148 616888
rect 3200 616876 3206 616888
rect 6362 616876 6368 616888
rect 3200 616848 6368 616876
rect 3200 616836 3206 616848
rect 6362 616836 6368 616848
rect 6420 616836 6426 616888
rect 6178 608580 6184 608592
rect 6139 608552 6184 608580
rect 6178 608540 6184 608552
rect 6236 608540 6242 608592
rect 6178 599060 6184 599072
rect 6139 599032 6184 599060
rect 6178 599020 6184 599032
rect 6236 599020 6242 599072
rect 6178 598924 6184 598936
rect 6139 598896 6184 598924
rect 6178 598884 6184 598896
rect 6236 598884 6242 598936
rect 6178 591784 6184 591796
rect 6139 591756 6184 591784
rect 6178 591744 6184 591756
rect 6236 591744 6242 591796
rect 6178 589268 6184 589280
rect 6139 589240 6184 589268
rect 6178 589228 6184 589240
rect 6236 589228 6242 589280
rect 6178 579748 6184 579760
rect 6139 579720 6184 579748
rect 6178 579708 6184 579720
rect 6236 579708 6242 579760
rect 6089 579615 6147 579621
rect 6089 579581 6101 579615
rect 6135 579612 6147 579615
rect 6178 579612 6184 579624
rect 6135 579584 6184 579612
rect 6135 579581 6147 579584
rect 6089 579575 6147 579581
rect 6178 579572 6184 579584
rect 6236 579572 6242 579624
rect 6086 569956 6092 569968
rect 6047 569928 6092 569956
rect 6086 569916 6092 569928
rect 6144 569916 6150 569968
rect 3326 567264 3332 567316
rect 3384 567304 3390 567316
rect 7650 567304 7656 567316
rect 3384 567276 7656 567304
rect 3384 567264 3390 567276
rect 7650 567264 7656 567276
rect 7708 567264 7714 567316
rect 6086 565128 6092 565140
rect 6047 565100 6092 565128
rect 6086 565088 6092 565100
rect 6144 565088 6150 565140
rect 6086 560300 6092 560312
rect 6047 560272 6092 560300
rect 6086 560260 6092 560272
rect 6144 560260 6150 560312
rect 6086 553432 6092 553444
rect 6047 553404 6092 553432
rect 6086 553392 6092 553404
rect 6144 553392 6150 553444
rect 6086 550644 6092 550656
rect 6047 550616 6092 550644
rect 6086 550604 6092 550616
rect 6144 550604 6150 550656
rect 6086 550508 6092 550520
rect 6047 550480 6092 550508
rect 6086 550468 6092 550480
rect 6144 550468 6150 550520
rect 6086 540988 6092 541000
rect 6047 540960 6092 540988
rect 6086 540948 6092 540960
rect 6144 540948 6150 541000
rect 5997 534123 6055 534129
rect 5997 534089 6009 534123
rect 6043 534120 6055 534123
rect 6086 534120 6092 534132
rect 6043 534092 6092 534120
rect 6043 534089 6055 534092
rect 5997 534083 6055 534089
rect 6086 534080 6092 534092
rect 6144 534080 6150 534132
rect 5994 531332 6000 531344
rect 5955 531304 6000 531332
rect 5994 531292 6000 531304
rect 6052 531292 6058 531344
rect 5810 521636 5816 521688
rect 5868 521676 5874 521688
rect 6086 521676 6092 521688
rect 5868 521648 6092 521676
rect 5868 521636 5874 521648
rect 6086 521636 6092 521648
rect 6144 521636 6150 521688
rect 6086 514768 6092 514820
rect 6144 514768 6150 514820
rect 6104 514740 6132 514768
rect 6178 514740 6184 514752
rect 6104 514712 6184 514740
rect 6178 514700 6184 514712
rect 6236 514700 6242 514752
rect 3142 509260 3148 509312
rect 3200 509300 3206 509312
rect 7742 509300 7748 509312
rect 3200 509272 7748 509300
rect 3200 509260 3206 509272
rect 7742 509260 7748 509272
rect 7800 509260 7806 509312
rect 6270 502324 6276 502376
rect 6328 502364 6334 502376
rect 6454 502364 6460 502376
rect 6328 502336 6460 502364
rect 6328 502324 6334 502336
rect 6454 502324 6460 502336
rect 6512 502324 6518 502376
rect 6086 487812 6092 487824
rect 6047 487784 6092 487812
rect 6086 487772 6092 487784
rect 6144 487772 6150 487824
rect 576118 487092 576124 487144
rect 576176 487132 576182 487144
rect 579706 487132 579712 487144
rect 576176 487104 579712 487132
rect 576176 487092 576182 487104
rect 579706 487092 579712 487104
rect 579764 487092 579770 487144
rect 6089 483123 6147 483129
rect 6089 483089 6101 483123
rect 6135 483120 6147 483123
rect 6178 483120 6184 483132
rect 6135 483092 6184 483120
rect 6135 483089 6147 483092
rect 6089 483083 6147 483089
rect 6178 483080 6184 483092
rect 6236 483080 6242 483132
rect 5905 476187 5963 476193
rect 5905 476153 5917 476187
rect 5951 476184 5963 476187
rect 6178 476184 6184 476196
rect 5951 476156 6184 476184
rect 5951 476153 5963 476156
rect 5905 476147 5963 476153
rect 6178 476144 6184 476156
rect 6236 476144 6242 476196
rect 5902 473464 5908 473476
rect 5863 473436 5908 473464
rect 5902 473424 5908 473436
rect 5960 473424 5966 473476
rect 5902 471928 5908 471980
rect 5960 471968 5966 471980
rect 6089 471971 6147 471977
rect 6089 471968 6101 471971
rect 5960 471940 6101 471968
rect 5960 471928 5966 471940
rect 6089 471937 6101 471940
rect 6135 471937 6147 471971
rect 6089 471931 6147 471937
rect 6086 456736 6092 456748
rect 6047 456708 6092 456736
rect 6086 456696 6092 456708
rect 6144 456696 6150 456748
rect 6086 452180 6092 452192
rect 6047 452152 6092 452180
rect 6086 452140 6092 452152
rect 6144 452140 6150 452192
rect 6089 444499 6147 444505
rect 6089 444465 6101 444499
rect 6135 444496 6147 444499
rect 6178 444496 6184 444508
rect 6135 444468 6184 444496
rect 6135 444465 6147 444468
rect 6089 444459 6147 444465
rect 6178 444456 6184 444468
rect 6236 444456 6242 444508
rect 6089 444363 6147 444369
rect 6089 444329 6101 444363
rect 6135 444360 6147 444363
rect 6178 444360 6184 444372
rect 6135 444332 6184 444360
rect 6135 444329 6147 444332
rect 6089 444323 6147 444329
rect 6178 444320 6184 444332
rect 6236 444320 6242 444372
rect 6086 434772 6092 434784
rect 6047 434744 6092 434772
rect 6086 434732 6092 434744
rect 6144 434732 6150 434784
rect 6086 431644 6092 431656
rect 6047 431616 6092 431644
rect 6086 431604 6092 431616
rect 6144 431604 6150 431656
rect 6086 425116 6092 425128
rect 6047 425088 6092 425116
rect 6086 425076 6092 425088
rect 6144 425076 6150 425128
rect 6178 425048 6184 425060
rect 6139 425020 6184 425048
rect 6178 425008 6184 425020
rect 6236 425008 6242 425060
rect 6086 415420 6092 415472
rect 6144 415460 6150 415472
rect 6181 415463 6239 415469
rect 6181 415460 6193 415463
rect 6144 415432 6193 415460
rect 6144 415420 6150 415432
rect 6181 415429 6193 415432
rect 6227 415429 6239 415463
rect 6181 415423 6239 415429
rect 6086 410564 6092 410576
rect 6047 410536 6092 410564
rect 6086 410524 6092 410536
rect 6144 410524 6150 410576
rect 6086 405736 6092 405748
rect 6047 405708 6092 405736
rect 6086 405696 6092 405708
rect 6144 405696 6150 405748
rect 6086 398828 6092 398880
rect 6144 398828 6150 398880
rect 6104 398800 6132 398828
rect 6178 398800 6184 398812
rect 6104 398772 6184 398800
rect 6178 398760 6184 398772
rect 6236 398760 6242 398812
rect 6178 389172 6184 389224
rect 6236 389172 6242 389224
rect 6086 389104 6092 389156
rect 6144 389144 6150 389156
rect 6196 389144 6224 389172
rect 6144 389116 6224 389144
rect 6144 389104 6150 389116
rect 6178 386356 6184 386368
rect 6139 386328 6184 386356
rect 6178 386316 6184 386328
rect 6236 386316 6242 386368
rect 6178 376768 6184 376780
rect 6139 376740 6184 376768
rect 6178 376728 6184 376740
rect 6236 376728 6242 376780
rect 6178 369900 6184 369912
rect 6104 369872 6184 369900
rect 6104 369844 6132 369872
rect 6178 369860 6184 369872
rect 6236 369860 6242 369912
rect 6086 369792 6092 369844
rect 6144 369792 6150 369844
rect 6086 360204 6092 360256
rect 6144 360204 6150 360256
rect 6104 360176 6132 360204
rect 6178 360176 6184 360188
rect 6104 360148 6184 360176
rect 6178 360136 6184 360148
rect 6236 360136 6242 360188
rect 6178 357252 6184 357264
rect 6139 357224 6184 357252
rect 6178 357212 6184 357224
rect 6236 357212 6242 357264
rect 6178 347868 6184 347880
rect 6139 347840 6184 347868
rect 6178 347828 6184 347840
rect 6236 347828 6242 347880
rect 6178 340892 6184 340944
rect 6236 340892 6242 340944
rect 6196 340740 6224 340892
rect 6178 340688 6184 340740
rect 6236 340688 6242 340740
rect 6178 338036 6184 338088
rect 6236 338076 6242 338088
rect 6362 338076 6368 338088
rect 6236 338048 6368 338076
rect 6236 338036 6242 338048
rect 6362 338036 6368 338048
rect 6420 338036 6426 338088
rect 6362 336716 6368 336728
rect 6323 336688 6368 336716
rect 6362 336676 6368 336688
rect 6420 336676 6426 336728
rect 6362 327808 6368 327820
rect 6323 327780 6368 327808
rect 6362 327768 6368 327780
rect 6420 327768 6426 327820
rect 6178 318764 6184 318776
rect 6139 318736 6184 318764
rect 6178 318724 6184 318736
rect 6236 318724 6242 318776
rect 6178 309244 6184 309256
rect 6139 309216 6184 309244
rect 6178 309204 6184 309216
rect 6236 309204 6242 309256
rect 6178 309108 6184 309120
rect 6139 309080 6184 309108
rect 6178 309068 6184 309080
rect 6236 309068 6242 309120
rect 6178 301968 6184 301980
rect 6139 301940 6184 301968
rect 6178 301928 6184 301940
rect 6236 301928 6242 301980
rect 6178 299452 6184 299464
rect 6139 299424 6184 299452
rect 6178 299412 6184 299424
rect 6236 299412 6242 299464
rect 6178 289932 6184 289944
rect 6139 289904 6184 289932
rect 6178 289892 6184 289904
rect 6236 289892 6242 289944
rect 6178 289796 6184 289808
rect 6139 289768 6184 289796
rect 6178 289756 6184 289768
rect 6236 289756 6242 289808
rect 6178 282792 6184 282804
rect 6139 282764 6184 282792
rect 6178 282752 6184 282764
rect 6236 282752 6242 282804
rect 6178 280140 6184 280152
rect 6139 280112 6184 280140
rect 6178 280100 6184 280112
rect 6236 280100 6242 280152
rect 6178 270620 6184 270632
rect 6139 270592 6184 270620
rect 6178 270580 6184 270592
rect 6236 270580 6242 270632
rect 6178 270484 6184 270496
rect 6139 270456 6184 270484
rect 6178 270444 6184 270456
rect 6236 270444 6242 270496
rect 6178 263344 6184 263356
rect 6139 263316 6184 263344
rect 6178 263304 6184 263316
rect 6236 263304 6242 263356
rect 6178 260828 6184 260840
rect 6139 260800 6184 260828
rect 6178 260788 6184 260800
rect 6236 260788 6242 260840
rect 6178 251308 6184 251320
rect 6139 251280 6184 251308
rect 6178 251268 6184 251280
rect 6236 251268 6242 251320
rect 6089 251175 6147 251181
rect 6089 251141 6101 251175
rect 6135 251172 6147 251175
rect 6178 251172 6184 251184
rect 6135 251144 6184 251172
rect 6135 251141 6147 251144
rect 6089 251135 6147 251141
rect 6178 251132 6184 251144
rect 6236 251132 6242 251184
rect 6086 241516 6092 241528
rect 6047 241488 6092 241516
rect 6086 241476 6092 241488
rect 6144 241476 6150 241528
rect 6086 236688 6092 236700
rect 6047 236660 6092 236688
rect 6086 236648 6092 236660
rect 6144 236648 6150 236700
rect 6086 231860 6092 231872
rect 6047 231832 6092 231860
rect 6086 231820 6092 231832
rect 6144 231820 6150 231872
rect 6086 224992 6092 225004
rect 6047 224964 6092 224992
rect 6086 224952 6092 224964
rect 6144 224952 6150 225004
rect 6086 222204 6092 222216
rect 6047 222176 6092 222204
rect 6086 222164 6092 222176
rect 6144 222164 6150 222216
rect 6086 222068 6092 222080
rect 6047 222040 6092 222068
rect 6086 222028 6092 222040
rect 6144 222028 6150 222080
rect 6086 212548 6092 212560
rect 6047 212520 6092 212548
rect 6086 212508 6092 212520
rect 6144 212508 6150 212560
rect 578142 209380 578148 209432
rect 578200 209420 578206 209432
rect 580626 209420 580632 209432
rect 578200 209392 580632 209420
rect 578200 209380 578206 209392
rect 580626 209380 580632 209392
rect 580684 209380 580690 209432
rect 6086 205640 6092 205692
rect 6144 205640 6150 205692
rect 6104 205612 6132 205640
rect 6178 205612 6184 205624
rect 6104 205584 6184 205612
rect 6178 205572 6184 205584
rect 6236 205572 6242 205624
rect 6270 193196 6276 193248
rect 6328 193236 6334 193248
rect 6454 193236 6460 193248
rect 6328 193208 6460 193236
rect 6328 193196 6334 193208
rect 6454 193196 6460 193208
rect 6512 193196 6518 193248
rect 578142 187620 578148 187672
rect 578200 187660 578206 187672
rect 580718 187660 580724 187672
rect 578200 187632 580724 187660
rect 578200 187620 578206 187632
rect 580718 187620 580724 187632
rect 580776 187620 580782 187672
rect 6086 183540 6092 183592
rect 6144 183580 6150 183592
rect 6270 183580 6276 183592
rect 6144 183552 6276 183580
rect 6144 183540 6150 183552
rect 6270 183540 6276 183552
rect 6328 183540 6334 183592
rect 6270 173884 6276 173936
rect 6328 173924 6334 173936
rect 6454 173924 6460 173936
rect 6328 173896 6460 173924
rect 6328 173884 6334 173896
rect 6454 173884 6460 173896
rect 6512 173884 6518 173936
rect 578142 166948 578148 167000
rect 578200 166988 578206 167000
rect 580810 166988 580816 167000
rect 578200 166960 580816 166988
rect 578200 166948 578206 166960
rect 580810 166948 580816 166960
rect 580868 166948 580874 167000
rect 6086 159372 6092 159384
rect 6047 159344 6092 159372
rect 6086 159332 6092 159344
rect 6144 159332 6150 159384
rect 6089 154683 6147 154689
rect 6089 154649 6101 154683
rect 6135 154680 6147 154683
rect 6178 154680 6184 154692
rect 6135 154652 6184 154680
rect 6135 154649 6147 154652
rect 6089 154643 6147 154649
rect 6178 154640 6184 154652
rect 6236 154640 6242 154692
rect 5902 154504 5908 154556
rect 5960 154544 5966 154556
rect 6178 154544 6184 154556
rect 5960 154516 6184 154544
rect 5960 154504 5966 154516
rect 6178 154504 6184 154516
rect 6236 154504 6242 154556
rect 578142 145732 578148 145784
rect 578200 145772 578206 145784
rect 580902 145772 580908 145784
rect 578200 145744 580908 145772
rect 578200 145732 578206 145744
rect 580902 145732 580908 145744
rect 580960 145732 580966 145784
rect 6086 138048 6092 138100
rect 6144 138048 6150 138100
rect 6104 137964 6132 138048
rect 6086 137912 6092 137964
rect 6144 137912 6150 137964
rect 5902 135192 5908 135244
rect 5960 135232 5966 135244
rect 6178 135232 6184 135244
rect 5960 135204 6184 135232
rect 5960 135192 5966 135204
rect 6178 135192 6184 135204
rect 6236 135192 6242 135244
rect 6086 118668 6092 118720
rect 6144 118668 6150 118720
rect 6104 118640 6132 118668
rect 6178 118640 6184 118652
rect 6104 118612 6184 118640
rect 6178 118600 6184 118612
rect 6236 118600 6242 118652
rect 6089 115923 6147 115929
rect 6089 115889 6101 115923
rect 6135 115920 6147 115923
rect 6178 115920 6184 115932
rect 6135 115892 6184 115920
rect 6135 115889 6147 115892
rect 6089 115883 6147 115889
rect 6178 115880 6184 115892
rect 6236 115880 6242 115932
rect 6086 106332 6092 106344
rect 6047 106304 6092 106332
rect 6086 106292 6092 106304
rect 6144 106292 6150 106344
rect 578142 103164 578148 103216
rect 578200 103204 578206 103216
rect 580626 103204 580632 103216
rect 578200 103176 580632 103204
rect 578200 103164 578206 103176
rect 580626 103164 580632 103176
rect 580684 103164 580690 103216
rect 6086 101436 6092 101448
rect 6047 101408 6092 101436
rect 6086 101396 6092 101408
rect 6144 101396 6150 101448
rect 6086 96676 6092 96688
rect 6047 96648 6092 96676
rect 6086 96636 6092 96648
rect 6144 96636 6150 96688
rect 6178 96608 6184 96620
rect 6139 96580 6184 96608
rect 6178 96568 6184 96580
rect 6236 96568 6242 96620
rect 6086 86980 6092 87032
rect 6144 87020 6150 87032
rect 6181 87023 6239 87029
rect 6181 87020 6193 87023
rect 6144 86992 6193 87020
rect 6144 86980 6150 86992
rect 6181 86989 6193 86992
rect 6227 86989 6239 87023
rect 6181 86983 6239 86989
rect 6086 82124 6092 82136
rect 6047 82096 6092 82124
rect 6086 82084 6092 82096
rect 6144 82084 6150 82136
rect 578142 81336 578148 81388
rect 578200 81376 578206 81388
rect 580718 81376 580724 81388
rect 578200 81348 580724 81376
rect 578200 81336 578206 81348
rect 580718 81336 580724 81348
rect 580776 81336 580782 81388
rect 6086 77296 6092 77308
rect 6047 77268 6092 77296
rect 6086 77256 6092 77268
rect 6144 77256 6150 77308
rect 6086 70388 6092 70440
rect 6144 70388 6150 70440
rect 6104 70360 6132 70388
rect 6178 70360 6184 70372
rect 6104 70332 6184 70360
rect 6178 70320 6184 70332
rect 6236 70320 6242 70372
rect 6178 60732 6184 60784
rect 6236 60732 6242 60784
rect 6086 60664 6092 60716
rect 6144 60704 6150 60716
rect 6196 60704 6224 60732
rect 6144 60676 6224 60704
rect 6144 60664 6150 60676
rect 578142 60596 578148 60648
rect 578200 60636 578206 60648
rect 580810 60636 580816 60648
rect 578200 60608 580816 60636
rect 578200 60596 578206 60608
rect 580810 60596 580816 60608
rect 580868 60596 580874 60648
rect 6178 57916 6184 57928
rect 6139 57888 6184 57916
rect 6178 57876 6184 57888
rect 6236 57876 6242 57928
rect 6178 48328 6184 48340
rect 6139 48300 6184 48328
rect 6178 48288 6184 48300
rect 6236 48288 6242 48340
rect 6178 47444 6184 47456
rect 6139 47416 6184 47444
rect 6178 47404 6184 47416
rect 6236 47404 6242 47456
rect 578142 39516 578148 39568
rect 578200 39556 578206 39568
rect 580626 39556 580632 39568
rect 578200 39528 580632 39556
rect 578200 39516 578206 39528
rect 580626 39516 580632 39528
rect 580684 39516 580690 39568
rect 6178 38672 6184 38684
rect 6139 38644 6184 38672
rect 6178 38632 6184 38644
rect 6236 38632 6242 38684
rect 6178 31696 6184 31748
rect 6236 31736 6242 31748
rect 6362 31736 6368 31748
rect 6236 31708 6368 31736
rect 6236 31696 6242 31708
rect 6362 31696 6368 31708
rect 6420 31696 6426 31748
rect 6273 28951 6331 28957
rect 6273 28917 6285 28951
rect 6319 28948 6331 28951
rect 6362 28948 6368 28960
rect 6319 28920 6368 28948
rect 6319 28917 6331 28920
rect 6273 28911 6331 28917
rect 6362 28908 6368 28920
rect 6420 28908 6426 28960
rect 6270 19360 6276 19372
rect 6231 19332 6276 19360
rect 6270 19320 6276 19332
rect 6328 19320 6334 19372
rect 9122 7828 9128 7880
rect 9180 7868 9186 7880
rect 11517 7871 11575 7877
rect 11517 7868 11529 7871
rect 9180 7840 11529 7868
rect 9180 7828 9186 7840
rect 11517 7837 11529 7840
rect 11563 7837 11575 7871
rect 11517 7831 11575 7837
rect 9490 7760 9496 7812
rect 9548 7800 9554 7812
rect 9548 7772 45784 7800
rect 9548 7760 9554 7772
rect 45756 7744 45784 7772
rect 9214 7692 9220 7744
rect 9272 7732 9278 7744
rect 11517 7735 11575 7741
rect 9272 7704 11468 7732
rect 9272 7692 9278 7704
rect 9306 7624 9312 7676
rect 9364 7664 9370 7676
rect 11440 7664 11468 7704
rect 11517 7701 11529 7735
rect 11563 7732 11575 7735
rect 11563 7704 45692 7732
rect 11563 7701 11575 7704
rect 11517 7695 11575 7701
rect 45557 7667 45615 7673
rect 45557 7664 45569 7667
rect 9364 7636 11376 7664
rect 11440 7636 45569 7664
rect 9364 7624 9370 7636
rect 9398 7556 9404 7608
rect 9456 7596 9462 7608
rect 11238 7596 11244 7608
rect 9456 7568 11244 7596
rect 9456 7556 9462 7568
rect 11238 7556 11244 7568
rect 11296 7556 11302 7608
rect 11348 7596 11376 7636
rect 45557 7633 45569 7636
rect 45603 7633 45615 7667
rect 45664 7664 45692 7704
rect 45738 7692 45744 7744
rect 45796 7692 45802 7744
rect 49326 7664 49332 7676
rect 45664 7636 49332 7664
rect 45557 7627 45615 7633
rect 49326 7624 49332 7636
rect 49384 7624 49390 7676
rect 12434 7596 12440 7608
rect 11348 7568 12440 7596
rect 12434 7556 12440 7568
rect 12492 7556 12498 7608
rect 62390 7596 62396 7608
rect 12544 7568 62396 7596
rect 9030 7352 9036 7404
rect 9088 7392 9094 7404
rect 12544 7392 12572 7568
rect 62390 7556 62396 7568
rect 62448 7556 62454 7608
rect 45557 7463 45615 7469
rect 45557 7429 45569 7463
rect 45603 7460 45615 7463
rect 52822 7460 52828 7472
rect 45603 7432 52828 7460
rect 45603 7429 45615 7432
rect 45557 7423 45615 7429
rect 52822 7420 52828 7432
rect 52880 7420 52886 7472
rect 9088 7364 12572 7392
rect 9088 7352 9094 7364
rect 8846 6876 8852 6928
rect 8904 6916 8910 6928
rect 8904 6888 9720 6916
rect 8904 6876 8910 6888
rect 9692 6848 9720 6888
rect 11054 6848 11060 6860
rect 9692 6820 11060 6848
rect 11054 6808 11060 6820
rect 11112 6808 11118 6860
rect 50430 6808 50436 6860
rect 50488 6848 50494 6860
rect 580534 6848 580540 6860
rect 50488 6820 580540 6848
rect 50488 6808 50494 6820
rect 580534 6808 580540 6820
rect 580592 6808 580598 6860
rect 60090 6740 60096 6792
rect 60148 6780 60154 6792
rect 580442 6780 580448 6792
rect 60148 6752 580448 6780
rect 60148 6740 60154 6752
rect 580442 6740 580448 6752
rect 580500 6740 580506 6792
rect 69750 6672 69756 6724
rect 69808 6712 69814 6724
rect 580350 6712 580356 6724
rect 69808 6684 580356 6712
rect 69808 6672 69814 6684
rect 580350 6672 580356 6684
rect 580408 6672 580414 6724
rect 79410 6604 79416 6656
rect 79468 6644 79474 6656
rect 580258 6644 580264 6656
rect 79468 6616 580264 6644
rect 79468 6604 79474 6616
rect 580258 6604 580264 6616
rect 580316 6604 580322 6656
rect 87322 6536 87328 6588
rect 87380 6576 87386 6588
rect 578786 6576 578792 6588
rect 87380 6548 578792 6576
rect 87380 6536 87386 6548
rect 578786 6536 578792 6548
rect 578844 6536 578850 6588
rect 76650 6468 76656 6520
rect 76708 6508 76714 6520
rect 578878 6508 578884 6520
rect 76708 6480 578884 6508
rect 76708 6468 76714 6480
rect 578878 6468 578884 6480
rect 578936 6468 578942 6520
rect 65978 6400 65984 6452
rect 66036 6440 66042 6452
rect 578970 6440 578976 6452
rect 66036 6412 578976 6440
rect 66036 6400 66042 6412
rect 578970 6400 578976 6412
rect 579028 6400 579034 6452
rect 55214 6332 55220 6384
rect 55272 6372 55278 6384
rect 579062 6372 579068 6384
rect 55272 6344 579068 6372
rect 55272 6332 55278 6344
rect 579062 6332 579068 6344
rect 579120 6332 579126 6384
rect 48130 6264 48136 6316
rect 48188 6304 48194 6316
rect 579154 6304 579160 6316
rect 48188 6276 579160 6304
rect 48188 6264 48194 6276
rect 579154 6264 579160 6276
rect 579212 6264 579218 6316
rect 7466 6196 7472 6248
rect 7524 6236 7530 6248
rect 579430 6236 579436 6248
rect 7524 6208 579436 6236
rect 7524 6196 7530 6208
rect 579430 6196 579436 6208
rect 579488 6196 579494 6248
rect 566 6128 572 6180
rect 624 6168 630 6180
rect 579522 6168 579528 6180
rect 624 6140 579528 6168
rect 624 6128 630 6140
rect 579522 6128 579528 6140
rect 579580 6128 579586 6180
rect 105170 6060 105176 6112
rect 105228 6100 105234 6112
rect 578694 6100 578700 6112
rect 105228 6072 578700 6100
rect 105228 6060 105234 6072
rect 578694 6060 578700 6072
rect 578752 6060 578758 6112
rect 108758 5992 108764 6044
rect 108816 6032 108822 6044
rect 578602 6032 578608 6044
rect 108816 6004 578608 6032
rect 108816 5992 108822 6004
rect 578602 5992 578608 6004
rect 578660 5992 578666 6044
rect 115934 5924 115940 5976
rect 115992 5964 115998 5976
rect 578510 5964 578516 5976
rect 115992 5936 578516 5964
rect 115992 5924 115998 5936
rect 578510 5924 578516 5936
rect 578568 5924 578574 5976
rect 119430 5856 119436 5908
rect 119488 5896 119494 5908
rect 578418 5896 578424 5908
rect 119488 5868 578424 5896
rect 119488 5856 119494 5868
rect 578418 5856 578424 5868
rect 578476 5856 578482 5908
rect 7558 5448 7564 5500
rect 7616 5488 7622 5500
rect 11790 5488 11796 5500
rect 7616 5460 11796 5488
rect 7616 5448 7622 5460
rect 11790 5448 11796 5460
rect 11848 5448 11854 5500
rect 93302 5448 93308 5500
rect 93360 5488 93366 5500
rect 301590 5488 301596 5500
rect 93360 5460 301596 5488
rect 93360 5448 93366 5460
rect 301590 5448 301596 5460
rect 301648 5448 301654 5500
rect 5258 5380 5264 5432
rect 5316 5420 5322 5432
rect 70670 5420 70676 5432
rect 5316 5392 70676 5420
rect 5316 5380 5322 5392
rect 70670 5380 70676 5392
rect 70728 5380 70734 5432
rect 100478 5380 100484 5432
rect 100536 5420 100542 5432
rect 320910 5420 320916 5432
rect 100536 5392 320916 5420
rect 100536 5380 100542 5392
rect 320910 5380 320916 5392
rect 320968 5380 320974 5432
rect 11054 5312 11060 5364
rect 11112 5352 11118 5364
rect 83826 5352 83832 5364
rect 11112 5324 83832 5352
rect 11112 5312 11118 5324
rect 83826 5312 83832 5324
rect 83884 5312 83890 5364
rect 107562 5312 107568 5364
rect 107620 5352 107626 5364
rect 340230 5352 340236 5364
rect 107620 5324 340236 5352
rect 107620 5312 107626 5324
rect 340230 5312 340236 5324
rect 340288 5312 340294 5364
rect 8938 5244 8944 5296
rect 8996 5284 9002 5296
rect 90910 5284 90916 5296
rect 8996 5256 90916 5284
rect 8996 5244 9002 5256
rect 90910 5244 90916 5256
rect 90968 5244 90974 5296
rect 114738 5244 114744 5296
rect 114796 5284 114802 5296
rect 359550 5284 359556 5296
rect 114796 5256 359556 5284
rect 114796 5244 114802 5256
rect 359550 5244 359556 5256
rect 359608 5244 359614 5296
rect 19518 5176 19524 5228
rect 19576 5216 19582 5228
rect 108390 5216 108396 5228
rect 19576 5188 108396 5216
rect 19576 5176 19582 5188
rect 108390 5176 108396 5188
rect 108448 5176 108454 5228
rect 121822 5176 121828 5228
rect 121880 5216 121886 5228
rect 378870 5216 378876 5228
rect 121880 5188 378876 5216
rect 121880 5176 121886 5188
rect 378870 5176 378876 5188
rect 378928 5176 378934 5228
rect 7650 5108 7656 5160
rect 7708 5148 7714 5160
rect 31110 5148 31116 5160
rect 7708 5120 31116 5148
rect 7708 5108 7714 5120
rect 31110 5108 31116 5120
rect 31168 5108 31174 5160
rect 57606 5108 57612 5160
rect 57664 5148 57670 5160
rect 204990 5148 204996 5160
rect 57664 5120 204996 5148
rect 57664 5108 57670 5120
rect 204990 5108 204996 5120
rect 205048 5108 205054 5160
rect 220722 5108 220728 5160
rect 220780 5148 220786 5160
rect 572070 5148 572076 5160
rect 220780 5120 572076 5148
rect 220780 5108 220786 5120
rect 572070 5108 572076 5120
rect 572128 5108 572134 5160
rect 7742 5040 7748 5092
rect 7800 5080 7806 5092
rect 40770 5080 40776 5092
rect 7800 5052 40776 5080
rect 7800 5040 7806 5052
rect 40770 5040 40776 5052
rect 40828 5040 40834 5092
rect 58802 5040 58808 5092
rect 58860 5080 58866 5092
rect 436830 5080 436836 5092
rect 58860 5052 436836 5080
rect 58860 5040 58866 5052
rect 436830 5040 436836 5052
rect 436888 5040 436894 5092
rect 2866 4972 2872 5024
rect 2924 5012 2930 5024
rect 407850 5012 407856 5024
rect 2924 4984 407856 5012
rect 2924 4972 2930 4984
rect 407850 4972 407856 4984
rect 407908 4972 407914 5024
rect 4614 4904 4620 4956
rect 4672 4944 4678 4956
rect 94498 4944 94504 4956
rect 4672 4916 94504 4944
rect 4672 4904 4678 4916
rect 94498 4904 94504 4916
rect 94556 4904 94562 4956
rect 117130 4904 117136 4956
rect 117188 4944 117194 4956
rect 533430 4944 533436 4956
rect 117188 4916 533436 4944
rect 117188 4904 117194 4916
rect 533430 4904 533436 4916
rect 533488 4904 533494 4956
rect 5442 4836 5448 4888
rect 5500 4876 5506 4888
rect 95694 4876 95700 4888
rect 5500 4848 95700 4876
rect 5500 4836 5506 4848
rect 95694 4836 95700 4848
rect 95752 4836 95758 4888
rect 120626 4836 120632 4888
rect 120684 4876 120690 4888
rect 543090 4876 543096 4888
rect 120684 4848 543096 4876
rect 120684 4836 120690 4848
rect 543090 4836 543096 4848
rect 543148 4836 543154 4888
rect 6638 4768 6644 4820
rect 6696 4808 6702 4820
rect 21450 4808 21456 4820
rect 6696 4780 21456 4808
rect 6696 4768 6702 4780
rect 21450 4768 21456 4780
rect 21508 4768 21514 4820
rect 24302 4768 24308 4820
rect 24360 4808 24366 4820
rect 118050 4808 118056 4820
rect 24360 4780 118056 4808
rect 24360 4768 24366 4780
rect 118050 4768 118056 4780
rect 118108 4768 118114 4820
rect 124214 4768 124220 4820
rect 124272 4808 124278 4820
rect 552750 4808 552756 4820
rect 124272 4780 552756 4808
rect 124272 4768 124278 4780
rect 552750 4768 552756 4780
rect 552808 4768 552814 4820
rect 86126 4700 86132 4752
rect 86184 4740 86190 4752
rect 282270 4740 282276 4752
rect 86184 4712 282276 4740
rect 86184 4700 86190 4712
rect 282270 4700 282276 4712
rect 282328 4700 282334 4752
rect 79042 4632 79048 4684
rect 79100 4672 79106 4684
rect 262950 4672 262956 4684
rect 79100 4644 262956 4672
rect 79100 4632 79106 4644
rect 262950 4632 262956 4644
rect 263008 4632 263014 4684
rect 71866 4564 71872 4616
rect 71924 4604 71930 4616
rect 243630 4604 243636 4616
rect 71924 4576 243636 4604
rect 71924 4564 71930 4576
rect 243630 4564 243636 4576
rect 243688 4564 243694 4616
rect 64782 4496 64788 4548
rect 64840 4536 64846 4548
rect 224310 4536 224316 4548
rect 64840 4508 224316 4536
rect 64840 4496 64846 4508
rect 224310 4496 224316 4508
rect 224368 4496 224374 4548
rect 54018 4428 54024 4480
rect 54076 4468 54082 4480
rect 195330 4468 195336 4480
rect 54076 4440 195336 4468
rect 54076 4428 54082 4440
rect 195330 4428 195336 4440
rect 195388 4428 195394 4480
rect 50522 4360 50528 4412
rect 50580 4400 50586 4412
rect 185670 4400 185676 4412
rect 50580 4372 185676 4400
rect 50580 4360 50586 4372
rect 185670 4360 185676 4372
rect 185728 4360 185734 4412
rect 46934 4292 46940 4344
rect 46992 4332 46998 4344
rect 176010 4332 176016 4344
rect 46992 4304 176016 4332
rect 46992 4292 46998 4304
rect 176010 4292 176016 4304
rect 176068 4292 176074 4344
rect 39758 4224 39764 4276
rect 39816 4264 39822 4276
rect 156690 4264 156696 4276
rect 39816 4236 156696 4264
rect 39816 4224 39822 4236
rect 156690 4224 156696 4236
rect 156748 4224 156754 4276
rect 156782 4224 156788 4276
rect 156840 4264 156846 4276
rect 253290 4264 253296 4276
rect 156840 4236 253296 4264
rect 156840 4224 156846 4236
rect 253290 4224 253296 4236
rect 253348 4224 253354 4276
rect 32674 4156 32680 4208
rect 32732 4196 32738 4208
rect 137370 4196 137376 4208
rect 32732 4168 137376 4196
rect 32732 4156 32738 4168
rect 137370 4156 137376 4168
rect 137428 4156 137434 4208
rect 5258 4088 5264 4140
rect 5316 4128 5322 4140
rect 220722 4128 220728 4140
rect 5316 4100 220728 4128
rect 5316 4088 5322 4100
rect 220722 4088 220728 4100
rect 220780 4088 220786 4140
rect 10042 4020 10048 4072
rect 10100 4060 10106 4072
rect 89070 4060 89076 4072
rect 10100 4032 89076 4060
rect 10100 4020 10106 4032
rect 89070 4020 89076 4032
rect 89128 4020 89134 4072
rect 103974 4020 103980 4072
rect 104032 4060 104038 4072
rect 330570 4060 330576 4072
rect 104032 4032 330576 4060
rect 104032 4020 104038 4032
rect 330570 4020 330576 4032
rect 330628 4020 330634 4072
rect 7006 3952 7012 4004
rect 7064 3992 7070 4004
rect 13725 3995 13783 4001
rect 13725 3992 13737 3995
rect 7064 3964 13737 3992
rect 7064 3952 7070 3964
rect 13725 3961 13737 3964
rect 13771 3961 13783 3995
rect 13725 3955 13783 3961
rect 14826 3952 14832 4004
rect 14884 3992 14890 4004
rect 98730 3992 98736 4004
rect 14884 3964 98736 3992
rect 14884 3952 14890 3964
rect 98730 3952 98736 3964
rect 98788 3952 98794 4004
rect 111150 3952 111156 4004
rect 111208 3992 111214 4004
rect 349890 3992 349896 4004
rect 111208 3964 349896 3992
rect 111208 3952 111214 3964
rect 349890 3952 349896 3964
rect 349948 3952 349954 4004
rect 4798 3884 4804 3936
rect 4856 3924 4862 3936
rect 101582 3924 101588 3936
rect 4856 3896 101588 3924
rect 4856 3884 4862 3896
rect 101582 3884 101588 3896
rect 101640 3884 101646 3936
rect 118234 3884 118240 3936
rect 118292 3924 118298 3936
rect 369210 3924 369216 3936
rect 118292 3896 369216 3924
rect 118292 3884 118298 3896
rect 369210 3884 369216 3896
rect 369268 3884 369274 3936
rect 4890 3816 4896 3868
rect 4948 3856 4954 3868
rect 112346 3856 112352 3868
rect 4948 3828 112352 3856
rect 4948 3816 4954 3828
rect 112346 3816 112352 3828
rect 112404 3816 112410 3868
rect 125410 3816 125416 3868
rect 125468 3856 125474 3868
rect 388530 3856 388536 3868
rect 125468 3828 388536 3856
rect 125468 3816 125474 3828
rect 388530 3816 388536 3828
rect 388588 3816 388594 3868
rect 6914 3748 6920 3800
rect 6972 3788 6978 3800
rect 13630 3788 13636 3800
rect 6972 3760 13636 3788
rect 6972 3748 6978 3760
rect 13630 3748 13636 3760
rect 13688 3748 13694 3800
rect 13725 3791 13783 3797
rect 13725 3757 13737 3791
rect 13771 3788 13783 3791
rect 30282 3788 30288 3800
rect 13771 3760 30288 3788
rect 13771 3757 13783 3760
rect 13725 3751 13783 3757
rect 30282 3748 30288 3760
rect 30340 3748 30346 3800
rect 37366 3748 37372 3800
rect 37424 3788 37430 3800
rect 417510 3788 417516 3800
rect 37424 3760 417516 3788
rect 37424 3748 37430 3760
rect 417510 3748 417516 3760
rect 417568 3748 417574 3800
rect 4154 3680 4160 3732
rect 4212 3720 4218 3732
rect 40954 3720 40960 3732
rect 4212 3692 40960 3720
rect 4212 3680 4218 3692
rect 40954 3680 40960 3692
rect 41012 3680 41018 3732
rect 44542 3680 44548 3732
rect 44600 3720 44606 3732
rect 427170 3720 427176 3732
rect 44600 3692 427176 3720
rect 44600 3680 44606 3692
rect 427170 3680 427176 3692
rect 427228 3680 427234 3732
rect 5350 3612 5356 3664
rect 5408 3652 5414 3664
rect 88518 3652 88524 3664
rect 5408 3624 88524 3652
rect 5408 3612 5414 3624
rect 88518 3612 88524 3624
rect 88576 3612 88582 3664
rect 92106 3612 92112 3664
rect 92164 3652 92170 3664
rect 514110 3652 514116 3664
rect 92164 3624 514116 3652
rect 92164 3612 92170 3624
rect 514110 3612 514116 3624
rect 514168 3612 514174 3664
rect 4706 3544 4712 3596
rect 4764 3584 4770 3596
rect 98086 3584 98092 3596
rect 4764 3556 98092 3584
rect 4764 3544 4770 3556
rect 98086 3544 98092 3556
rect 98144 3544 98150 3596
rect 99282 3544 99288 3596
rect 99340 3584 99346 3596
rect 523770 3584 523776 3596
rect 99340 3556 523776 3584
rect 99340 3544 99346 3556
rect 523770 3544 523776 3556
rect 523828 3544 523834 3596
rect 5166 3476 5172 3528
rect 5224 3516 5230 3528
rect 56410 3516 56416 3528
rect 5224 3488 56416 3516
rect 5224 3476 5230 3488
rect 56410 3476 56416 3488
rect 56468 3476 56474 3528
rect 59998 3476 60004 3528
rect 60056 3516 60062 3528
rect 494790 3516 494796 3528
rect 60056 3488 494796 3516
rect 60056 3476 60062 3488
rect 494790 3476 494796 3488
rect 494848 3476 494854 3528
rect 4062 3408 4068 3460
rect 4120 3448 4126 3460
rect 446490 3448 446496 3460
rect 4120 3420 446496 3448
rect 4120 3408 4126 3420
rect 446490 3408 446496 3420
rect 446548 3408 446554 3460
rect 4522 3340 4528 3392
rect 4580 3380 4586 3392
rect 80238 3380 80244 3392
rect 4580 3352 80244 3380
rect 4580 3340 4586 3352
rect 80238 3340 80244 3352
rect 80296 3340 80302 3392
rect 96890 3340 96896 3392
rect 96948 3380 96954 3392
rect 311250 3380 311256 3392
rect 96948 3352 311256 3380
rect 96948 3340 96954 3352
rect 311250 3340 311256 3352
rect 311308 3340 311314 3392
rect 4430 3272 4436 3324
rect 4488 3312 4494 3324
rect 73062 3312 73068 3324
rect 4488 3284 73068 3312
rect 4488 3272 4494 3284
rect 73062 3272 73068 3284
rect 73120 3272 73126 3324
rect 89714 3272 89720 3324
rect 89772 3312 89778 3324
rect 291930 3312 291936 3324
rect 89772 3284 291936 3312
rect 89772 3272 89778 3284
rect 291930 3272 291936 3284
rect 291988 3272 291994 3324
rect 4338 3204 4344 3256
rect 4396 3244 4402 3256
rect 69474 3244 69480 3256
rect 4396 3216 69480 3244
rect 4396 3204 4402 3216
rect 69474 3204 69480 3216
rect 69532 3204 69538 3256
rect 82630 3204 82636 3256
rect 82688 3244 82694 3256
rect 272610 3244 272616 3256
rect 82688 3216 272616 3244
rect 82688 3204 82694 3216
rect 272610 3204 272616 3216
rect 272668 3204 272674 3256
rect 4246 3136 4252 3188
rect 4304 3176 4310 3188
rect 51626 3176 51632 3188
rect 4304 3148 51632 3176
rect 4304 3136 4310 3148
rect 51626 3136 51632 3148
rect 51684 3136 51690 3188
rect 68278 3136 68284 3188
rect 68336 3176 68342 3188
rect 233970 3176 233976 3188
rect 68336 3148 233976 3176
rect 68336 3136 68342 3148
rect 233970 3136 233976 3148
rect 234028 3136 234034 3188
rect 5074 3068 5080 3120
rect 5132 3108 5138 3120
rect 23106 3108 23112 3120
rect 5132 3080 23112 3108
rect 5132 3068 5138 3080
rect 23106 3068 23112 3080
rect 23164 3068 23170 3120
rect 61194 3068 61200 3120
rect 61252 3108 61258 3120
rect 214650 3108 214656 3120
rect 61252 3080 214656 3108
rect 61252 3068 61258 3080
rect 214650 3068 214656 3080
rect 214708 3068 214714 3120
rect 9582 3000 9588 3052
rect 9640 3040 9646 3052
rect 26694 3040 26700 3052
rect 9640 3012 26700 3040
rect 9640 3000 9646 3012
rect 26694 3000 26700 3012
rect 26752 3000 26758 3052
rect 43346 3000 43352 3052
rect 43404 3040 43410 3052
rect 166350 3040 166356 3052
rect 43404 3012 166356 3040
rect 43404 3000 43410 3012
rect 166350 3000 166356 3012
rect 166408 3000 166414 3052
rect 6822 2932 6828 2984
rect 6880 2972 6886 2984
rect 20714 2972 20720 2984
rect 6880 2944 20720 2972
rect 6880 2932 6886 2944
rect 20714 2932 20720 2944
rect 20772 2932 20778 2984
rect 36170 2932 36176 2984
rect 36228 2972 36234 2984
rect 147030 2972 147036 2984
rect 36228 2944 147036 2972
rect 36228 2932 36234 2944
rect 147030 2932 147036 2944
rect 147088 2932 147094 2984
rect 4982 2864 4988 2916
rect 5040 2904 5046 2916
rect 18322 2904 18328 2916
rect 5040 2876 18328 2904
rect 5040 2864 5046 2876
rect 18322 2864 18328 2876
rect 18380 2864 18386 2916
rect 29086 2864 29092 2916
rect 29144 2904 29150 2916
rect 127710 2904 127716 2916
rect 29144 2876 127716 2904
rect 29144 2864 29150 2876
rect 127710 2864 127716 2876
rect 127768 2864 127774 2916
rect 7098 2796 7104 2848
rect 7156 2836 7162 2848
rect 21910 2836 21916 2848
rect 7156 2808 21916 2836
rect 7156 2796 7162 2808
rect 21910 2796 21916 2808
rect 21968 2796 21974 2848
rect 75454 2796 75460 2848
rect 75512 2836 75518 2848
rect 156782 2836 156788 2848
rect 75512 2808 156788 2836
rect 75512 2796 75518 2808
rect 156782 2796 156788 2808
rect 156840 2796 156846 2848
rect 1670 2048 1676 2100
rect 1728 2088 1734 2100
rect 398190 2088 398196 2100
rect 1728 2060 398196 2088
rect 1728 2048 1734 2060
rect 398190 2048 398196 2060
rect 398248 2048 398254 2100
rect 5534 552 5540 604
rect 5592 592 5598 604
rect 6454 592 6460 604
rect 5592 564 6460 592
rect 5592 552 5598 564
rect 6454 552 6460 564
rect 6512 552 6518 604
<< via1 >>
rect 164148 700612 164200 700664
rect 235172 700612 235224 700664
rect 135168 700544 135220 700596
rect 300124 700544 300176 700596
rect 105452 700476 105504 700528
rect 106188 700476 106240 700528
rect 107568 700476 107620 700528
rect 364984 700476 365036 700528
rect 40500 700408 40552 700460
rect 41328 700408 41380 700460
rect 78588 700408 78640 700460
rect 429844 700408 429896 700460
rect 49608 700340 49660 700392
rect 494796 700340 494848 700392
rect 22008 700272 22060 700324
rect 559656 700272 559708 700324
rect 170312 699660 170364 699712
rect 171048 699660 171100 699712
rect 21180 689528 21232 689580
rect 22008 689528 22060 689580
rect 106648 689528 106700 689580
rect 107568 689528 107620 689580
rect 171048 689392 171100 689444
rect 192116 689392 192168 689444
rect 106188 689324 106240 689376
rect 220636 689324 220688 689376
rect 41328 689256 41380 689308
rect 249156 689256 249208 689308
rect 9312 689120 9364 689172
rect 306196 689120 306248 689172
rect 277676 689052 277728 689104
rect 576124 689052 576176 689104
rect 9588 688984 9640 689036
rect 334624 688984 334676 689036
rect 9036 688916 9088 688968
rect 363144 688916 363196 688968
rect 9496 688848 9548 688900
rect 448704 688848 448756 688900
rect 9128 688780 9180 688832
rect 477132 688780 477184 688832
rect 9220 688712 9272 688764
rect 505652 688712 505704 688764
rect 9404 688644 9456 688696
rect 562692 688644 562744 688696
rect 3516 681708 3568 681760
rect 7564 681708 7616 681760
rect 3148 616836 3200 616888
rect 6368 616836 6420 616888
rect 6184 608583 6236 608592
rect 6184 608549 6193 608583
rect 6193 608549 6227 608583
rect 6227 608549 6236 608583
rect 6184 608540 6236 608549
rect 6184 599063 6236 599072
rect 6184 599029 6193 599063
rect 6193 599029 6227 599063
rect 6227 599029 6236 599063
rect 6184 599020 6236 599029
rect 6184 598927 6236 598936
rect 6184 598893 6193 598927
rect 6193 598893 6227 598927
rect 6227 598893 6236 598927
rect 6184 598884 6236 598893
rect 6184 591787 6236 591796
rect 6184 591753 6193 591787
rect 6193 591753 6227 591787
rect 6227 591753 6236 591787
rect 6184 591744 6236 591753
rect 6184 589271 6236 589280
rect 6184 589237 6193 589271
rect 6193 589237 6227 589271
rect 6227 589237 6236 589271
rect 6184 589228 6236 589237
rect 6184 579751 6236 579760
rect 6184 579717 6193 579751
rect 6193 579717 6227 579751
rect 6227 579717 6236 579751
rect 6184 579708 6236 579717
rect 6184 579572 6236 579624
rect 6092 569959 6144 569968
rect 6092 569925 6101 569959
rect 6101 569925 6135 569959
rect 6135 569925 6144 569959
rect 6092 569916 6144 569925
rect 3332 567264 3384 567316
rect 7656 567264 7708 567316
rect 6092 565131 6144 565140
rect 6092 565097 6101 565131
rect 6101 565097 6135 565131
rect 6135 565097 6144 565131
rect 6092 565088 6144 565097
rect 6092 560303 6144 560312
rect 6092 560269 6101 560303
rect 6101 560269 6135 560303
rect 6135 560269 6144 560303
rect 6092 560260 6144 560269
rect 6092 553435 6144 553444
rect 6092 553401 6101 553435
rect 6101 553401 6135 553435
rect 6135 553401 6144 553435
rect 6092 553392 6144 553401
rect 6092 550647 6144 550656
rect 6092 550613 6101 550647
rect 6101 550613 6135 550647
rect 6135 550613 6144 550647
rect 6092 550604 6144 550613
rect 6092 550511 6144 550520
rect 6092 550477 6101 550511
rect 6101 550477 6135 550511
rect 6135 550477 6144 550511
rect 6092 550468 6144 550477
rect 6092 540991 6144 541000
rect 6092 540957 6101 540991
rect 6101 540957 6135 540991
rect 6135 540957 6144 540991
rect 6092 540948 6144 540957
rect 6092 534080 6144 534132
rect 6000 531335 6052 531344
rect 6000 531301 6009 531335
rect 6009 531301 6043 531335
rect 6043 531301 6052 531335
rect 6000 531292 6052 531301
rect 5816 521636 5868 521688
rect 6092 521636 6144 521688
rect 6092 514768 6144 514820
rect 6184 514700 6236 514752
rect 3148 509260 3200 509312
rect 7748 509260 7800 509312
rect 6276 502324 6328 502376
rect 6460 502324 6512 502376
rect 6092 487815 6144 487824
rect 6092 487781 6101 487815
rect 6101 487781 6135 487815
rect 6135 487781 6144 487815
rect 6092 487772 6144 487781
rect 576124 487092 576176 487144
rect 579712 487092 579764 487144
rect 6184 483080 6236 483132
rect 6184 476144 6236 476196
rect 5908 473467 5960 473476
rect 5908 473433 5917 473467
rect 5917 473433 5951 473467
rect 5951 473433 5960 473467
rect 5908 473424 5960 473433
rect 5908 471928 5960 471980
rect 6092 456739 6144 456748
rect 6092 456705 6101 456739
rect 6101 456705 6135 456739
rect 6135 456705 6144 456739
rect 6092 456696 6144 456705
rect 6092 452183 6144 452192
rect 6092 452149 6101 452183
rect 6101 452149 6135 452183
rect 6135 452149 6144 452183
rect 6092 452140 6144 452149
rect 6184 444456 6236 444508
rect 6184 444320 6236 444372
rect 6092 434775 6144 434784
rect 6092 434741 6101 434775
rect 6101 434741 6135 434775
rect 6135 434741 6144 434775
rect 6092 434732 6144 434741
rect 6092 431647 6144 431656
rect 6092 431613 6101 431647
rect 6101 431613 6135 431647
rect 6135 431613 6144 431647
rect 6092 431604 6144 431613
rect 6092 425119 6144 425128
rect 6092 425085 6101 425119
rect 6101 425085 6135 425119
rect 6135 425085 6144 425119
rect 6092 425076 6144 425085
rect 6184 425051 6236 425060
rect 6184 425017 6193 425051
rect 6193 425017 6227 425051
rect 6227 425017 6236 425051
rect 6184 425008 6236 425017
rect 6092 415420 6144 415472
rect 6092 410567 6144 410576
rect 6092 410533 6101 410567
rect 6101 410533 6135 410567
rect 6135 410533 6144 410567
rect 6092 410524 6144 410533
rect 6092 405739 6144 405748
rect 6092 405705 6101 405739
rect 6101 405705 6135 405739
rect 6135 405705 6144 405739
rect 6092 405696 6144 405705
rect 6092 398828 6144 398880
rect 6184 398760 6236 398812
rect 6184 389172 6236 389224
rect 6092 389104 6144 389156
rect 6184 386359 6236 386368
rect 6184 386325 6193 386359
rect 6193 386325 6227 386359
rect 6227 386325 6236 386359
rect 6184 386316 6236 386325
rect 6184 376771 6236 376780
rect 6184 376737 6193 376771
rect 6193 376737 6227 376771
rect 6227 376737 6236 376771
rect 6184 376728 6236 376737
rect 6184 369860 6236 369912
rect 6092 369792 6144 369844
rect 6092 360204 6144 360256
rect 6184 360136 6236 360188
rect 6184 357255 6236 357264
rect 6184 357221 6193 357255
rect 6193 357221 6227 357255
rect 6227 357221 6236 357255
rect 6184 357212 6236 357221
rect 6184 347871 6236 347880
rect 6184 347837 6193 347871
rect 6193 347837 6227 347871
rect 6227 347837 6236 347871
rect 6184 347828 6236 347837
rect 6184 340892 6236 340944
rect 6184 340688 6236 340740
rect 6184 338036 6236 338088
rect 6368 338036 6420 338088
rect 6368 336719 6420 336728
rect 6368 336685 6377 336719
rect 6377 336685 6411 336719
rect 6411 336685 6420 336719
rect 6368 336676 6420 336685
rect 6368 327811 6420 327820
rect 6368 327777 6377 327811
rect 6377 327777 6411 327811
rect 6411 327777 6420 327811
rect 6368 327768 6420 327777
rect 6184 318767 6236 318776
rect 6184 318733 6193 318767
rect 6193 318733 6227 318767
rect 6227 318733 6236 318767
rect 6184 318724 6236 318733
rect 6184 309247 6236 309256
rect 6184 309213 6193 309247
rect 6193 309213 6227 309247
rect 6227 309213 6236 309247
rect 6184 309204 6236 309213
rect 6184 309111 6236 309120
rect 6184 309077 6193 309111
rect 6193 309077 6227 309111
rect 6227 309077 6236 309111
rect 6184 309068 6236 309077
rect 6184 301971 6236 301980
rect 6184 301937 6193 301971
rect 6193 301937 6227 301971
rect 6227 301937 6236 301971
rect 6184 301928 6236 301937
rect 6184 299455 6236 299464
rect 6184 299421 6193 299455
rect 6193 299421 6227 299455
rect 6227 299421 6236 299455
rect 6184 299412 6236 299421
rect 6184 289935 6236 289944
rect 6184 289901 6193 289935
rect 6193 289901 6227 289935
rect 6227 289901 6236 289935
rect 6184 289892 6236 289901
rect 6184 289799 6236 289808
rect 6184 289765 6193 289799
rect 6193 289765 6227 289799
rect 6227 289765 6236 289799
rect 6184 289756 6236 289765
rect 6184 282795 6236 282804
rect 6184 282761 6193 282795
rect 6193 282761 6227 282795
rect 6227 282761 6236 282795
rect 6184 282752 6236 282761
rect 6184 280143 6236 280152
rect 6184 280109 6193 280143
rect 6193 280109 6227 280143
rect 6227 280109 6236 280143
rect 6184 280100 6236 280109
rect 6184 270623 6236 270632
rect 6184 270589 6193 270623
rect 6193 270589 6227 270623
rect 6227 270589 6236 270623
rect 6184 270580 6236 270589
rect 6184 270487 6236 270496
rect 6184 270453 6193 270487
rect 6193 270453 6227 270487
rect 6227 270453 6236 270487
rect 6184 270444 6236 270453
rect 6184 263347 6236 263356
rect 6184 263313 6193 263347
rect 6193 263313 6227 263347
rect 6227 263313 6236 263347
rect 6184 263304 6236 263313
rect 6184 260831 6236 260840
rect 6184 260797 6193 260831
rect 6193 260797 6227 260831
rect 6227 260797 6236 260831
rect 6184 260788 6236 260797
rect 6184 251311 6236 251320
rect 6184 251277 6193 251311
rect 6193 251277 6227 251311
rect 6227 251277 6236 251311
rect 6184 251268 6236 251277
rect 6184 251132 6236 251184
rect 6092 241519 6144 241528
rect 6092 241485 6101 241519
rect 6101 241485 6135 241519
rect 6135 241485 6144 241519
rect 6092 241476 6144 241485
rect 6092 236691 6144 236700
rect 6092 236657 6101 236691
rect 6101 236657 6135 236691
rect 6135 236657 6144 236691
rect 6092 236648 6144 236657
rect 6092 231863 6144 231872
rect 6092 231829 6101 231863
rect 6101 231829 6135 231863
rect 6135 231829 6144 231863
rect 6092 231820 6144 231829
rect 6092 224995 6144 225004
rect 6092 224961 6101 224995
rect 6101 224961 6135 224995
rect 6135 224961 6144 224995
rect 6092 224952 6144 224961
rect 6092 222207 6144 222216
rect 6092 222173 6101 222207
rect 6101 222173 6135 222207
rect 6135 222173 6144 222207
rect 6092 222164 6144 222173
rect 6092 222071 6144 222080
rect 6092 222037 6101 222071
rect 6101 222037 6135 222071
rect 6135 222037 6144 222071
rect 6092 222028 6144 222037
rect 6092 212551 6144 212560
rect 6092 212517 6101 212551
rect 6101 212517 6135 212551
rect 6135 212517 6144 212551
rect 6092 212508 6144 212517
rect 578148 209380 578200 209432
rect 580632 209380 580684 209432
rect 6092 205640 6144 205692
rect 6184 205572 6236 205624
rect 6276 193196 6328 193248
rect 6460 193196 6512 193248
rect 578148 187620 578200 187672
rect 580724 187620 580776 187672
rect 6092 183540 6144 183592
rect 6276 183540 6328 183592
rect 6276 173884 6328 173936
rect 6460 173884 6512 173936
rect 578148 166948 578200 167000
rect 580816 166948 580868 167000
rect 6092 159375 6144 159384
rect 6092 159341 6101 159375
rect 6101 159341 6135 159375
rect 6135 159341 6144 159375
rect 6092 159332 6144 159341
rect 6184 154640 6236 154692
rect 5908 154504 5960 154556
rect 6184 154504 6236 154556
rect 578148 145732 578200 145784
rect 580908 145732 580960 145784
rect 6092 138048 6144 138100
rect 6092 137912 6144 137964
rect 5908 135192 5960 135244
rect 6184 135192 6236 135244
rect 6092 118668 6144 118720
rect 6184 118600 6236 118652
rect 6184 115880 6236 115932
rect 6092 106335 6144 106344
rect 6092 106301 6101 106335
rect 6101 106301 6135 106335
rect 6135 106301 6144 106335
rect 6092 106292 6144 106301
rect 578148 103164 578200 103216
rect 580632 103164 580684 103216
rect 6092 101439 6144 101448
rect 6092 101405 6101 101439
rect 6101 101405 6135 101439
rect 6135 101405 6144 101439
rect 6092 101396 6144 101405
rect 6092 96679 6144 96688
rect 6092 96645 6101 96679
rect 6101 96645 6135 96679
rect 6135 96645 6144 96679
rect 6092 96636 6144 96645
rect 6184 96611 6236 96620
rect 6184 96577 6193 96611
rect 6193 96577 6227 96611
rect 6227 96577 6236 96611
rect 6184 96568 6236 96577
rect 6092 86980 6144 87032
rect 6092 82127 6144 82136
rect 6092 82093 6101 82127
rect 6101 82093 6135 82127
rect 6135 82093 6144 82127
rect 6092 82084 6144 82093
rect 578148 81336 578200 81388
rect 580724 81336 580776 81388
rect 6092 77299 6144 77308
rect 6092 77265 6101 77299
rect 6101 77265 6135 77299
rect 6135 77265 6144 77299
rect 6092 77256 6144 77265
rect 6092 70388 6144 70440
rect 6184 70320 6236 70372
rect 6184 60732 6236 60784
rect 6092 60664 6144 60716
rect 578148 60596 578200 60648
rect 580816 60596 580868 60648
rect 6184 57919 6236 57928
rect 6184 57885 6193 57919
rect 6193 57885 6227 57919
rect 6227 57885 6236 57919
rect 6184 57876 6236 57885
rect 6184 48331 6236 48340
rect 6184 48297 6193 48331
rect 6193 48297 6227 48331
rect 6227 48297 6236 48331
rect 6184 48288 6236 48297
rect 6184 47447 6236 47456
rect 6184 47413 6193 47447
rect 6193 47413 6227 47447
rect 6227 47413 6236 47447
rect 6184 47404 6236 47413
rect 578148 39516 578200 39568
rect 580632 39516 580684 39568
rect 6184 38675 6236 38684
rect 6184 38641 6193 38675
rect 6193 38641 6227 38675
rect 6227 38641 6236 38675
rect 6184 38632 6236 38641
rect 6184 31696 6236 31748
rect 6368 31696 6420 31748
rect 6368 28908 6420 28960
rect 6276 19363 6328 19372
rect 6276 19329 6285 19363
rect 6285 19329 6319 19363
rect 6319 19329 6328 19363
rect 6276 19320 6328 19329
rect 9128 7828 9180 7880
rect 9496 7760 9548 7812
rect 9220 7692 9272 7744
rect 9312 7624 9364 7676
rect 9404 7556 9456 7608
rect 11244 7556 11296 7608
rect 45744 7692 45796 7744
rect 49332 7624 49384 7676
rect 12440 7556 12492 7608
rect 9036 7352 9088 7404
rect 62396 7556 62448 7608
rect 52828 7420 52880 7472
rect 8852 6876 8904 6928
rect 11060 6808 11112 6860
rect 50436 6808 50488 6860
rect 580540 6808 580592 6860
rect 60096 6740 60148 6792
rect 580448 6740 580500 6792
rect 69756 6672 69808 6724
rect 580356 6672 580408 6724
rect 79416 6604 79468 6656
rect 580264 6604 580316 6656
rect 87328 6536 87380 6588
rect 578792 6536 578844 6588
rect 76656 6468 76708 6520
rect 578884 6468 578936 6520
rect 65984 6400 66036 6452
rect 578976 6400 579028 6452
rect 55220 6332 55272 6384
rect 579068 6332 579120 6384
rect 48136 6264 48188 6316
rect 579160 6264 579212 6316
rect 7472 6196 7524 6248
rect 579436 6196 579488 6248
rect 572 6128 624 6180
rect 579528 6128 579580 6180
rect 105176 6060 105228 6112
rect 578700 6060 578752 6112
rect 108764 5992 108816 6044
rect 578608 5992 578660 6044
rect 115940 5924 115992 5976
rect 578516 5924 578568 5976
rect 119436 5856 119488 5908
rect 578424 5856 578476 5908
rect 7564 5448 7616 5500
rect 11796 5448 11848 5500
rect 93308 5448 93360 5500
rect 301596 5448 301648 5500
rect 5264 5380 5316 5432
rect 70676 5380 70728 5432
rect 100484 5380 100536 5432
rect 320916 5380 320968 5432
rect 11060 5312 11112 5364
rect 83832 5312 83884 5364
rect 107568 5312 107620 5364
rect 340236 5312 340288 5364
rect 8944 5244 8996 5296
rect 90916 5244 90968 5296
rect 114744 5244 114796 5296
rect 359556 5244 359608 5296
rect 19524 5176 19576 5228
rect 108396 5176 108448 5228
rect 121828 5176 121880 5228
rect 378876 5176 378928 5228
rect 7656 5108 7708 5160
rect 31116 5108 31168 5160
rect 57612 5108 57664 5160
rect 204996 5108 205048 5160
rect 220728 5108 220780 5160
rect 572076 5108 572128 5160
rect 7748 5040 7800 5092
rect 40776 5040 40828 5092
rect 58808 5040 58860 5092
rect 436836 5040 436888 5092
rect 2872 4972 2924 5024
rect 407856 4972 407908 5024
rect 4620 4904 4672 4956
rect 94504 4904 94556 4956
rect 117136 4904 117188 4956
rect 533436 4904 533488 4956
rect 5448 4836 5500 4888
rect 95700 4836 95752 4888
rect 120632 4836 120684 4888
rect 543096 4836 543148 4888
rect 6644 4768 6696 4820
rect 21456 4768 21508 4820
rect 24308 4768 24360 4820
rect 118056 4768 118108 4820
rect 124220 4768 124272 4820
rect 552756 4768 552808 4820
rect 86132 4700 86184 4752
rect 282276 4700 282328 4752
rect 79048 4632 79100 4684
rect 262956 4632 263008 4684
rect 71872 4564 71924 4616
rect 243636 4564 243688 4616
rect 64788 4496 64840 4548
rect 224316 4496 224368 4548
rect 54024 4428 54076 4480
rect 195336 4428 195388 4480
rect 50528 4360 50580 4412
rect 185676 4360 185728 4412
rect 46940 4292 46992 4344
rect 176016 4292 176068 4344
rect 39764 4224 39816 4276
rect 156696 4224 156748 4276
rect 156788 4224 156840 4276
rect 253296 4224 253348 4276
rect 32680 4156 32732 4208
rect 137376 4156 137428 4208
rect 5264 4088 5316 4140
rect 220728 4088 220780 4140
rect 10048 4020 10100 4072
rect 89076 4020 89128 4072
rect 103980 4020 104032 4072
rect 330576 4020 330628 4072
rect 7012 3952 7064 4004
rect 14832 3952 14884 4004
rect 98736 3952 98788 4004
rect 111156 3952 111208 4004
rect 349896 3952 349948 4004
rect 4804 3884 4856 3936
rect 101588 3884 101640 3936
rect 118240 3884 118292 3936
rect 369216 3884 369268 3936
rect 4896 3816 4948 3868
rect 112352 3816 112404 3868
rect 125416 3816 125468 3868
rect 388536 3816 388588 3868
rect 6920 3748 6972 3800
rect 13636 3748 13688 3800
rect 30288 3748 30340 3800
rect 37372 3748 37424 3800
rect 417516 3748 417568 3800
rect 4160 3680 4212 3732
rect 40960 3680 41012 3732
rect 44548 3680 44600 3732
rect 427176 3680 427228 3732
rect 5356 3612 5408 3664
rect 88524 3612 88576 3664
rect 92112 3612 92164 3664
rect 514116 3612 514168 3664
rect 4712 3544 4764 3596
rect 98092 3544 98144 3596
rect 99288 3544 99340 3596
rect 523776 3544 523828 3596
rect 5172 3476 5224 3528
rect 56416 3476 56468 3528
rect 60004 3476 60056 3528
rect 494796 3476 494848 3528
rect 4068 3408 4120 3460
rect 446496 3408 446548 3460
rect 4528 3340 4580 3392
rect 80244 3340 80296 3392
rect 96896 3340 96948 3392
rect 311256 3340 311308 3392
rect 4436 3272 4488 3324
rect 73068 3272 73120 3324
rect 89720 3272 89772 3324
rect 291936 3272 291988 3324
rect 4344 3204 4396 3256
rect 69480 3204 69532 3256
rect 82636 3204 82688 3256
rect 272616 3204 272668 3256
rect 4252 3136 4304 3188
rect 51632 3136 51684 3188
rect 68284 3136 68336 3188
rect 233976 3136 234028 3188
rect 5080 3068 5132 3120
rect 23112 3068 23164 3120
rect 61200 3068 61252 3120
rect 214656 3068 214708 3120
rect 9588 3000 9640 3052
rect 26700 3000 26752 3052
rect 43352 3000 43404 3052
rect 166356 3000 166408 3052
rect 6828 2932 6880 2984
rect 20720 2932 20772 2984
rect 36176 2932 36228 2984
rect 147036 2932 147088 2984
rect 4988 2864 5040 2916
rect 18328 2864 18380 2916
rect 29092 2864 29144 2916
rect 127716 2864 127768 2916
rect 7104 2796 7156 2848
rect 21916 2796 21968 2848
rect 75460 2796 75512 2848
rect 156788 2796 156840 2848
rect 1676 2048 1728 2100
rect 398196 2048 398248 2100
rect 5540 552 5592 604
rect 6460 552 6512 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 40512 700466 40540 703520
rect 105464 700534 105492 703520
rect 164148 700664 164200 700670
rect 164148 700606 164200 700612
rect 135168 700596 135220 700602
rect 135168 700538 135220 700544
rect 105452 700528 105504 700534
rect 105452 700470 105504 700476
rect 106188 700528 106240 700534
rect 106188 700470 106240 700476
rect 107568 700528 107620 700534
rect 107568 700470 107620 700476
rect 40500 700460 40552 700466
rect 40500 700402 40552 700408
rect 41328 700460 41380 700466
rect 41328 700402 41380 700408
rect 78588 700460 78640 700466
rect 78588 700402 78640 700408
rect 22008 700324 22060 700330
rect 22008 700266 22060 700272
rect 22020 689586 22048 700266
rect 21180 689580 21232 689586
rect 21180 689522 21232 689528
rect 22008 689580 22060 689586
rect 22008 689522 22060 689528
rect 9312 689172 9364 689178
rect 9312 689114 9364 689120
rect 9036 688968 9088 688974
rect 9036 688910 9088 688916
rect 8850 685264 8906 685273
rect 8850 685199 8906 685208
rect 3514 682272 3570 682281
rect 3514 682207 3570 682216
rect 3528 681766 3556 682207
rect 3516 681760 3568 681766
rect 3516 681702 3568 681708
rect 7564 681760 7616 681766
rect 7564 681702 7616 681708
rect 5538 676424 5594 676433
rect 5538 676359 5594 676368
rect 3146 624880 3202 624889
rect 3146 624815 3202 624824
rect 3160 616894 3188 624815
rect 3148 616888 3200 616894
rect 3148 616830 3200 616836
rect 5446 572928 5502 572937
rect 5446 572863 5502 572872
rect 3330 567352 3386 567361
rect 3330 567287 3332 567296
rect 3384 567287 3386 567296
rect 3332 567258 3384 567264
rect 5354 552392 5410 552401
rect 5354 552327 5410 552336
rect 5262 531720 5318 531729
rect 5262 531655 5318 531664
rect 5170 511184 5226 511193
rect 5170 511119 5226 511128
rect 3146 509960 3202 509969
rect 3146 509895 3202 509904
rect 3160 509318 3188 509895
rect 3148 509312 3200 509318
rect 3148 509254 3200 509260
rect 5078 490512 5134 490521
rect 5078 490447 5134 490456
rect 4986 469976 5042 469985
rect 4986 469911 5042 469920
rect 3422 452432 3478 452441
rect 3422 452367 3478 452376
rect 3238 165064 3294 165073
rect 3238 164999 3294 165008
rect 3252 141545 3280 164999
rect 3330 160848 3386 160857
rect 3330 160783 3386 160792
rect 3238 141536 3294 141545
rect 3238 141471 3294 141480
rect 3344 122097 3372 160783
rect 3330 122088 3386 122097
rect 3330 122023 3386 122032
rect 3436 17921 3464 452367
rect 4894 429312 4950 429321
rect 4894 429247 4950 429256
rect 4802 408640 4858 408649
rect 4802 408575 4858 408584
rect 3514 395040 3570 395049
rect 3514 394975 3570 394984
rect 3528 38321 3556 394975
rect 4710 387832 4766 387841
rect 4710 387767 4766 387776
rect 4618 367296 4674 367305
rect 4618 367231 4674 367240
rect 4526 346488 4582 346497
rect 4526 346423 4582 346432
rect 3606 337512 3662 337521
rect 3606 337447 3662 337456
rect 3620 59129 3648 337447
rect 4434 325816 4490 325825
rect 4434 325751 4490 325760
rect 4342 305144 4398 305153
rect 4342 305079 4398 305088
rect 3698 294400 3754 294409
rect 3698 294335 3754 294344
rect 3712 79665 3740 294335
rect 4250 284472 4306 284481
rect 4250 284407 4306 284416
rect 4158 263936 4214 263945
rect 4158 263871 4214 263880
rect 3882 251288 3938 251297
rect 3882 251223 3938 251232
rect 3790 202056 3846 202065
rect 3790 201991 3846 202000
rect 3698 79656 3754 79665
rect 3698 79591 3754 79600
rect 3606 59120 3662 59129
rect 3606 59055 3662 59064
rect 3514 38312 3570 38321
rect 3514 38247 3570 38256
rect 3804 35873 3832 201991
rect 3896 100337 3924 251223
rect 4066 208176 4122 208185
rect 4066 208111 4122 208120
rect 3974 181520 4030 181529
rect 3974 181455 4030 181464
rect 3882 100328 3938 100337
rect 3882 100263 3938 100272
rect 3988 78985 4016 181455
rect 4080 120873 4108 208111
rect 4066 120864 4122 120873
rect 4066 120799 4122 120808
rect 3974 78976 4030 78985
rect 3974 78911 4030 78920
rect 3790 35864 3846 35873
rect 3790 35799 3846 35808
rect 3422 17912 3478 17921
rect 3422 17847 3478 17856
rect 572 6180 624 6186
rect 572 6122 624 6128
rect 584 480 612 6122
rect 2872 5024 2924 5030
rect 2872 4966 2924 4972
rect 1676 2100 1728 2106
rect 1676 2042 1728 2048
rect 1688 480 1716 2042
rect 2884 480 2912 4966
rect 4172 3738 4200 263871
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 4068 3460 4120 3466
rect 4068 3402 4120 3408
rect 4080 480 4108 3402
rect 4264 3194 4292 284407
rect 4356 3262 4384 305079
rect 4448 3330 4476 325751
rect 4540 3398 4568 346423
rect 4632 4962 4660 367231
rect 4620 4956 4672 4962
rect 4620 4898 4672 4904
rect 4724 3602 4752 387767
rect 4816 3942 4844 408575
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4908 3874 4936 429247
rect 4896 3868 4948 3874
rect 4896 3810 4948 3816
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4528 3392 4580 3398
rect 4528 3334 4580 3340
rect 4436 3324 4488 3330
rect 4436 3266 4488 3272
rect 4344 3256 4396 3262
rect 4344 3198 4396 3204
rect 4252 3188 4304 3194
rect 4252 3130 4304 3136
rect 5000 2922 5028 469911
rect 5092 3126 5120 490447
rect 5184 3534 5212 511119
rect 5276 5438 5304 531655
rect 5264 5432 5316 5438
rect 5264 5374 5316 5380
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 5172 3528 5224 3534
rect 5172 3470 5224 3476
rect 5080 3120 5132 3126
rect 5080 3062 5132 3068
rect 4988 2916 5040 2922
rect 4988 2858 5040 2864
rect 5276 480 5304 4082
rect 5368 3670 5396 552327
rect 5460 4894 5488 572863
rect 5448 4888 5500 4894
rect 5448 4830 5500 4836
rect 5356 3664 5408 3670
rect 5356 3606 5408 3612
rect 5552 610 5580 676359
rect 6826 655752 6882 655761
rect 6826 655687 6882 655696
rect 6368 616888 6420 616894
rect 6368 616830 6420 616836
rect 6380 608682 6408 616830
rect 6196 608654 6408 608682
rect 6196 608598 6224 608654
rect 6184 608592 6236 608598
rect 6184 608534 6236 608540
rect 6184 599072 6236 599078
rect 6184 599014 6236 599020
rect 6196 598942 6224 599014
rect 6184 598936 6236 598942
rect 6184 598878 6236 598884
rect 6184 591796 6236 591802
rect 6184 591738 6236 591744
rect 6196 589286 6224 591738
rect 6184 589280 6236 589286
rect 6184 589222 6236 589228
rect 6184 579760 6236 579766
rect 6184 579702 6236 579708
rect 6196 579630 6224 579702
rect 6184 579624 6236 579630
rect 6184 579566 6236 579572
rect 6092 569968 6144 569974
rect 6092 569910 6144 569916
rect 6104 565146 6132 569910
rect 6092 565140 6144 565146
rect 6092 565082 6144 565088
rect 6092 560312 6144 560318
rect 6092 560254 6144 560260
rect 6104 553450 6132 560254
rect 6092 553444 6144 553450
rect 6092 553386 6144 553392
rect 6092 550656 6144 550662
rect 6092 550598 6144 550604
rect 6104 550526 6132 550598
rect 6092 550520 6144 550526
rect 6092 550462 6144 550468
rect 6092 541000 6144 541006
rect 6092 540942 6144 540948
rect 6104 534138 6132 540942
rect 6092 534132 6144 534138
rect 6092 534074 6144 534080
rect 6000 531344 6052 531350
rect 5814 531312 5870 531321
rect 5814 531247 5870 531256
rect 5998 531312 6000 531321
rect 6052 531312 6054 531321
rect 5998 531247 6054 531256
rect 5828 521694 5856 531247
rect 5816 521688 5868 521694
rect 5816 521630 5868 521636
rect 6092 521688 6144 521694
rect 6092 521630 6144 521636
rect 6104 514826 6132 521630
rect 6092 514820 6144 514826
rect 6092 514762 6144 514768
rect 6184 514752 6236 514758
rect 6184 514694 6236 514700
rect 6196 512009 6224 514694
rect 6182 512000 6238 512009
rect 6182 511935 6238 511944
rect 6458 512000 6514 512009
rect 6458 511935 6514 511944
rect 6472 502382 6500 511935
rect 6276 502376 6328 502382
rect 6276 502318 6328 502324
rect 6460 502376 6512 502382
rect 6460 502318 6512 502324
rect 6288 492697 6316 502318
rect 6090 492688 6146 492697
rect 6090 492623 6146 492632
rect 6274 492688 6330 492697
rect 6274 492623 6330 492632
rect 6104 487830 6132 492623
rect 6092 487824 6144 487830
rect 6092 487766 6144 487772
rect 6184 483132 6236 483138
rect 6184 483074 6236 483080
rect 6196 476202 6224 483074
rect 6184 476196 6236 476202
rect 6184 476138 6236 476144
rect 5908 473476 5960 473482
rect 5908 473418 5960 473424
rect 5920 471986 5948 473418
rect 5908 471980 5960 471986
rect 5908 471922 5960 471928
rect 6092 456748 6144 456754
rect 6092 456690 6144 456696
rect 6104 452198 6132 456690
rect 6092 452192 6144 452198
rect 6092 452134 6144 452140
rect 6184 444508 6236 444514
rect 6184 444450 6236 444456
rect 6196 444378 6224 444450
rect 6184 444372 6236 444378
rect 6184 444314 6236 444320
rect 6092 434784 6144 434790
rect 6092 434726 6144 434732
rect 6104 431662 6132 434726
rect 6092 431656 6144 431662
rect 6092 431598 6144 431604
rect 6092 425128 6144 425134
rect 6144 425076 6224 425082
rect 6092 425070 6224 425076
rect 6104 425066 6224 425070
rect 6104 425060 6236 425066
rect 6104 425054 6184 425060
rect 6184 425002 6236 425008
rect 6196 424971 6224 425002
rect 6092 415472 6144 415478
rect 6092 415414 6144 415420
rect 6104 410582 6132 415414
rect 6092 410576 6144 410582
rect 6092 410518 6144 410524
rect 6092 405748 6144 405754
rect 6092 405690 6144 405696
rect 6104 398886 6132 405690
rect 6092 398880 6144 398886
rect 6092 398822 6144 398828
rect 6184 398812 6236 398818
rect 6184 398754 6236 398760
rect 6196 389230 6224 398754
rect 6184 389224 6236 389230
rect 6184 389166 6236 389172
rect 6092 389156 6144 389162
rect 6092 389098 6144 389104
rect 6104 386458 6132 389098
rect 6104 386430 6224 386458
rect 6196 386374 6224 386430
rect 6184 386368 6236 386374
rect 6184 386310 6236 386316
rect 6184 376780 6236 376786
rect 6184 376722 6236 376728
rect 6196 369918 6224 376722
rect 6184 369912 6236 369918
rect 6184 369854 6236 369860
rect 6092 369844 6144 369850
rect 6092 369786 6144 369792
rect 6104 360262 6132 369786
rect 6092 360256 6144 360262
rect 6092 360198 6144 360204
rect 6184 360188 6236 360194
rect 6184 360130 6236 360136
rect 6196 357270 6224 360130
rect 6184 357264 6236 357270
rect 6184 357206 6236 357212
rect 6184 347880 6236 347886
rect 6184 347822 6236 347828
rect 6196 340950 6224 347822
rect 6184 340944 6236 340950
rect 6184 340886 6236 340892
rect 6184 340740 6236 340746
rect 6184 340682 6236 340688
rect 6196 338094 6224 340682
rect 6184 338088 6236 338094
rect 6184 338030 6236 338036
rect 6368 338088 6420 338094
rect 6368 338030 6420 338036
rect 6380 336734 6408 338030
rect 6368 336728 6420 336734
rect 6368 336670 6420 336676
rect 6368 327820 6420 327826
rect 6368 327762 6420 327768
rect 6380 321450 6408 327762
rect 6196 321422 6408 321450
rect 6196 318782 6224 321422
rect 6184 318776 6236 318782
rect 6184 318718 6236 318724
rect 6184 309256 6236 309262
rect 6184 309198 6236 309204
rect 6196 309126 6224 309198
rect 6184 309120 6236 309126
rect 6184 309062 6236 309068
rect 6184 301980 6236 301986
rect 6184 301922 6236 301928
rect 6196 299470 6224 301922
rect 6184 299464 6236 299470
rect 6184 299406 6236 299412
rect 6184 289944 6236 289950
rect 6184 289886 6236 289892
rect 6196 289814 6224 289886
rect 6184 289808 6236 289814
rect 6184 289750 6236 289756
rect 6184 282804 6236 282810
rect 6184 282746 6236 282752
rect 6196 280158 6224 282746
rect 6184 280152 6236 280158
rect 6184 280094 6236 280100
rect 6184 270632 6236 270638
rect 6184 270574 6236 270580
rect 6196 270502 6224 270574
rect 6184 270496 6236 270502
rect 6184 270438 6236 270444
rect 6184 263356 6236 263362
rect 6184 263298 6236 263304
rect 6196 260846 6224 263298
rect 6184 260840 6236 260846
rect 6184 260782 6236 260788
rect 6184 251320 6236 251326
rect 6184 251262 6236 251268
rect 6196 251190 6224 251262
rect 6184 251184 6236 251190
rect 6184 251126 6236 251132
rect 6092 241528 6144 241534
rect 6092 241470 6144 241476
rect 6104 236706 6132 241470
rect 6092 236700 6144 236706
rect 6092 236642 6144 236648
rect 6092 231872 6144 231878
rect 6092 231814 6144 231820
rect 6104 225010 6132 231814
rect 6092 225004 6144 225010
rect 6092 224946 6144 224952
rect 6092 222216 6144 222222
rect 6092 222158 6144 222164
rect 6104 222086 6132 222158
rect 6092 222080 6144 222086
rect 6092 222022 6144 222028
rect 6092 212560 6144 212566
rect 6092 212502 6144 212508
rect 6104 205698 6132 212502
rect 6092 205692 6144 205698
rect 6092 205634 6144 205640
rect 6184 205624 6236 205630
rect 6184 205566 6236 205572
rect 6196 202881 6224 205566
rect 6182 202872 6238 202881
rect 6182 202807 6238 202816
rect 6458 202872 6514 202881
rect 6458 202807 6514 202816
rect 6472 193254 6500 202807
rect 6276 193248 6328 193254
rect 6276 193190 6328 193196
rect 6460 193248 6512 193254
rect 6460 193190 6512 193196
rect 6104 183598 6132 183629
rect 6288 183598 6316 193190
rect 6092 183592 6144 183598
rect 6276 183592 6328 183598
rect 6182 183560 6238 183569
rect 6144 183540 6182 183546
rect 6092 183534 6182 183540
rect 6104 183518 6182 183534
rect 6276 183534 6328 183540
rect 6458 183560 6514 183569
rect 6182 183495 6238 183504
rect 6458 183495 6514 183504
rect 6472 173942 6500 183495
rect 6276 173936 6328 173942
rect 6276 173878 6328 173884
rect 6460 173936 6512 173942
rect 6460 173878 6512 173884
rect 6288 164257 6316 173878
rect 6090 164248 6146 164257
rect 6090 164183 6146 164192
rect 6274 164248 6330 164257
rect 6274 164183 6330 164192
rect 6104 159390 6132 164183
rect 6092 159384 6144 159390
rect 6092 159326 6144 159332
rect 6184 154692 6236 154698
rect 6184 154634 6236 154640
rect 6196 154562 6224 154634
rect 5908 154556 5960 154562
rect 5908 154498 5960 154504
rect 6184 154556 6236 154562
rect 6184 154498 6236 154504
rect 5920 144945 5948 154498
rect 5906 144936 5962 144945
rect 5906 144871 5962 144880
rect 6090 144936 6146 144945
rect 6090 144871 6146 144880
rect 6104 138106 6132 144871
rect 6092 138100 6144 138106
rect 6092 138042 6144 138048
rect 6092 137964 6144 137970
rect 6092 137906 6144 137912
rect 6104 135266 6132 137906
rect 6104 135250 6224 135266
rect 5908 135244 5960 135250
rect 6104 135244 6236 135250
rect 6104 135238 6184 135244
rect 5908 135186 5960 135192
rect 6184 135186 6236 135192
rect 5920 125633 5948 135186
rect 6196 135155 6224 135186
rect 5906 125624 5962 125633
rect 5906 125559 5962 125568
rect 6090 125624 6146 125633
rect 6090 125559 6146 125568
rect 6104 118726 6132 125559
rect 6092 118720 6144 118726
rect 6092 118662 6144 118668
rect 6184 118652 6236 118658
rect 6184 118594 6236 118600
rect 6196 115938 6224 118594
rect 6184 115932 6236 115938
rect 6184 115874 6236 115880
rect 6092 106344 6144 106350
rect 6092 106286 6144 106292
rect 6104 101454 6132 106286
rect 6092 101448 6144 101454
rect 6092 101390 6144 101396
rect 6092 96688 6144 96694
rect 6144 96636 6224 96642
rect 6092 96630 6224 96636
rect 6104 96626 6224 96630
rect 6104 96620 6236 96626
rect 6104 96614 6184 96620
rect 6184 96562 6236 96568
rect 6196 96531 6224 96562
rect 6092 87032 6144 87038
rect 6092 86974 6144 86980
rect 6104 82142 6132 86974
rect 6092 82136 6144 82142
rect 6092 82078 6144 82084
rect 6092 77308 6144 77314
rect 6092 77250 6144 77256
rect 6104 70446 6132 77250
rect 6092 70440 6144 70446
rect 6092 70382 6144 70388
rect 6184 70372 6236 70378
rect 6184 70314 6236 70320
rect 6196 60790 6224 70314
rect 6184 60784 6236 60790
rect 6184 60726 6236 60732
rect 6092 60716 6144 60722
rect 6092 60658 6144 60664
rect 6104 58018 6132 60658
rect 6104 57990 6224 58018
rect 6196 57934 6224 57990
rect 6184 57928 6236 57934
rect 6184 57870 6236 57876
rect 6184 48340 6236 48346
rect 6184 48282 6236 48288
rect 6196 47462 6224 48282
rect 6184 47456 6236 47462
rect 6184 47398 6236 47404
rect 6184 38684 6236 38690
rect 6184 38626 6236 38632
rect 6196 31754 6224 38626
rect 6184 31748 6236 31754
rect 6184 31690 6236 31696
rect 6368 31748 6420 31754
rect 6368 31690 6420 31696
rect 6380 28966 6408 31690
rect 6368 28960 6420 28966
rect 6368 28902 6420 28908
rect 6276 19372 6328 19378
rect 6276 19314 6328 19320
rect 6288 12458 6316 19314
rect 6288 12430 6684 12458
rect 6656 4826 6684 12430
rect 6644 4820 6696 4826
rect 6644 4762 6696 4768
rect 6840 2990 6868 655687
rect 6918 449712 6974 449721
rect 6918 449647 6974 449656
rect 6932 3806 6960 449647
rect 7010 243264 7066 243273
rect 7010 243199 7066 243208
rect 7024 4010 7052 243199
rect 7102 222728 7158 222737
rect 7102 222663 7158 222672
rect 7012 4004 7064 4010
rect 7012 3946 7064 3952
rect 6920 3800 6972 3806
rect 6920 3742 6972 3748
rect 6828 2984 6880 2990
rect 6828 2926 6880 2932
rect 7116 2854 7144 222663
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 7104 2848 7156 2854
rect 7104 2790 7156 2796
rect 7484 2802 7512 6190
rect 7576 5506 7604 681702
rect 7656 567316 7708 567322
rect 7656 567258 7708 567264
rect 7564 5500 7616 5506
rect 7564 5442 7616 5448
rect 7668 5166 7696 567258
rect 7748 509312 7800 509318
rect 7748 509254 7800 509260
rect 7656 5160 7708 5166
rect 7656 5102 7708 5108
rect 7760 5098 7788 509254
rect 8864 6934 8892 685199
rect 8942 685128 8998 685137
rect 8942 685063 8998 685072
rect 8852 6928 8904 6934
rect 8852 6870 8904 6876
rect 8956 5302 8984 685063
rect 9048 7410 9076 688910
rect 9128 688832 9180 688838
rect 9128 688774 9180 688780
rect 9140 7886 9168 688774
rect 9220 688764 9272 688770
rect 9220 688706 9272 688712
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9232 7750 9260 688706
rect 9220 7744 9272 7750
rect 9220 7686 9272 7692
rect 9324 7682 9352 689114
rect 9588 689036 9640 689042
rect 9588 688978 9640 688984
rect 9496 688900 9548 688906
rect 9496 688842 9548 688848
rect 9404 688696 9456 688702
rect 9404 688638 9456 688644
rect 9312 7676 9364 7682
rect 9312 7618 9364 7624
rect 9416 7614 9444 688638
rect 9508 7818 9536 688842
rect 9496 7812 9548 7818
rect 9496 7754 9548 7760
rect 9404 7608 9456 7614
rect 9404 7550 9456 7556
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 8944 5296 8996 5302
rect 8944 5238 8996 5244
rect 7748 5092 7800 5098
rect 7748 5034 7800 5040
rect 8850 4992 8906 5001
rect 8850 4927 8906 4936
rect 7484 2774 7696 2802
rect 5540 604 5592 610
rect 5540 546 5592 552
rect 6460 604 6512 610
rect 6460 546 6512 552
rect 6472 480 6500 546
rect 7668 480 7696 2774
rect 8864 480 8892 4927
rect 9600 3058 9628 688978
rect 21192 686868 21220 689522
rect 41340 689314 41368 700402
rect 49608 700392 49660 700398
rect 49608 700334 49660 700340
rect 41328 689308 41380 689314
rect 41328 689250 41380 689256
rect 49620 686868 49648 700334
rect 78600 686882 78628 700402
rect 106200 689382 106228 700470
rect 107580 689586 107608 700470
rect 106648 689580 106700 689586
rect 106648 689522 106700 689528
rect 107568 689580 107620 689586
rect 107568 689522 107620 689528
rect 106188 689376 106240 689382
rect 106188 689318 106240 689324
rect 78154 686854 78628 686882
rect 106660 686868 106688 689522
rect 135180 686868 135208 700538
rect 164160 686882 164188 700606
rect 170324 699718 170352 703520
rect 235184 700670 235212 703520
rect 235172 700664 235224 700670
rect 235172 700606 235224 700612
rect 300136 700602 300164 703520
rect 300124 700596 300176 700602
rect 300124 700538 300176 700544
rect 364996 700534 365024 703520
rect 364984 700528 365036 700534
rect 364984 700470 365036 700476
rect 429856 700466 429884 703520
rect 429844 700460 429896 700466
rect 429844 700402 429896 700408
rect 494808 700398 494836 703520
rect 494796 700392 494848 700398
rect 494796 700334 494848 700340
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 170312 699712 170364 699718
rect 170312 699654 170364 699660
rect 171048 699712 171100 699718
rect 171048 699654 171100 699660
rect 171060 689450 171088 699654
rect 171048 689444 171100 689450
rect 171048 689386 171100 689392
rect 192116 689444 192168 689450
rect 192116 689386 192168 689392
rect 163714 686854 164188 686882
rect 192128 686868 192156 689386
rect 220636 689376 220688 689382
rect 220636 689318 220688 689324
rect 220648 686868 220676 689318
rect 249156 689308 249208 689314
rect 249156 689250 249208 689256
rect 249168 686868 249196 689250
rect 306196 689172 306248 689178
rect 306196 689114 306248 689120
rect 277676 689104 277728 689110
rect 277676 689046 277728 689052
rect 277688 686868 277716 689046
rect 306208 686868 306236 689114
rect 576124 689104 576176 689110
rect 576124 689046 576176 689052
rect 334624 689036 334676 689042
rect 334624 688978 334676 688984
rect 334636 686868 334664 688978
rect 363144 688968 363196 688974
rect 363144 688910 363196 688916
rect 363156 686868 363184 688910
rect 448704 688900 448756 688906
rect 448704 688842 448756 688848
rect 448716 686868 448744 688842
rect 477132 688832 477184 688838
rect 477132 688774 477184 688780
rect 477144 686868 477172 688774
rect 505652 688764 505704 688770
rect 505652 688706 505704 688712
rect 505664 686868 505692 688706
rect 562692 688696 562744 688702
rect 534170 688664 534226 688673
rect 562692 688638 562744 688644
rect 534170 688599 534226 688608
rect 534184 686868 534212 688599
rect 562704 686868 562732 688638
rect 391478 686352 391534 686361
rect 419998 686352 420054 686361
rect 391534 686310 391690 686338
rect 391478 686287 391534 686296
rect 420054 686310 420210 686338
rect 419998 686287 420054 686296
rect 576136 487150 576164 689046
rect 580262 674656 580318 674665
rect 580262 674591 580318 674600
rect 578238 527232 578294 527241
rect 578238 527167 578294 527176
rect 576124 487144 576176 487150
rect 576124 487086 576176 487092
rect 578148 209432 578200 209438
rect 578146 209400 578148 209409
rect 578200 209400 578202 209409
rect 578146 209335 578202 209344
rect 578148 187672 578200 187678
rect 578146 187640 578148 187649
rect 578200 187640 578202 187649
rect 578146 187575 578202 187584
rect 578148 167000 578200 167006
rect 578146 166968 578148 166977
rect 578200 166968 578202 166977
rect 578146 166903 578202 166912
rect 578148 145784 578200 145790
rect 578146 145752 578148 145761
rect 578200 145752 578202 145761
rect 578146 145687 578202 145696
rect 578148 103216 578200 103222
rect 578146 103184 578148 103193
rect 578200 103184 578202 103193
rect 578146 103119 578202 103128
rect 578146 81424 578202 81433
rect 578146 81359 578148 81368
rect 578200 81359 578202 81368
rect 578148 81330 578200 81336
rect 578148 60648 578200 60654
rect 578146 60616 578148 60625
rect 578200 60616 578202 60625
rect 578146 60551 578202 60560
rect 578148 39568 578200 39574
rect 578146 39536 578148 39545
rect 578200 39536 578202 39545
rect 578146 39471 578202 39480
rect 45744 7744 45796 7750
rect 45744 7686 45796 7692
rect 11244 7608 11296 7614
rect 11244 7550 11296 7556
rect 12440 7608 12492 7614
rect 12440 7550 12492 7556
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 11072 5370 11100 6802
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 10048 4072 10100 4078
rect 10048 4014 10100 4020
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 10060 480 10088 4014
rect 11256 480 11284 7550
rect 11808 5506 11836 7004
rect 11796 5500 11848 5506
rect 11796 5442 11848 5448
rect 12452 480 12480 7550
rect 19524 5228 19576 5234
rect 19524 5170 19576 5176
rect 14832 4004 14884 4010
rect 14832 3946 14884 3952
rect 13636 3800 13688 3806
rect 13636 3742 13688 3748
rect 13648 480 13676 3742
rect 14844 480 14872 3946
rect 17222 3496 17278 3505
rect 17222 3431 17278 3440
rect 16026 3360 16082 3369
rect 16026 3295 16082 3304
rect 16040 480 16068 3295
rect 17236 480 17264 3431
rect 18328 2916 18380 2922
rect 18328 2858 18380 2864
rect 18340 480 18368 2858
rect 19536 480 19564 5170
rect 21468 4826 21496 7004
rect 31128 5166 31156 7004
rect 31482 5536 31538 5545
rect 31482 5471 31538 5480
rect 31116 5160 31168 5166
rect 31116 5102 31168 5108
rect 25502 4856 25558 4865
rect 21456 4820 21508 4826
rect 21456 4762 21508 4768
rect 24308 4820 24360 4826
rect 25502 4791 25558 4800
rect 24308 4762 24360 4768
rect 23112 3120 23164 3126
rect 23112 3062 23164 3068
rect 20720 2984 20772 2990
rect 20720 2926 20772 2932
rect 20732 480 20760 2926
rect 21916 2848 21968 2854
rect 21916 2790 21968 2796
rect 21928 480 21956 2790
rect 23124 480 23152 3062
rect 24320 480 24348 4762
rect 25516 480 25544 4791
rect 30288 3800 30340 3806
rect 30288 3742 30340 3748
rect 27894 3632 27950 3641
rect 27894 3567 27950 3576
rect 26700 3052 26752 3058
rect 26700 2994 26752 3000
rect 26712 480 26740 2994
rect 27908 480 27936 3567
rect 29092 2916 29144 2922
rect 29092 2858 29144 2864
rect 29104 480 29132 2858
rect 30300 480 30328 3742
rect 31496 480 31524 5471
rect 38566 5400 38622 5409
rect 38566 5335 38622 5344
rect 32680 4208 32732 4214
rect 32680 4150 32732 4156
rect 32692 480 32720 4150
rect 34978 3904 35034 3913
rect 34978 3839 35034 3848
rect 33874 3768 33930 3777
rect 33874 3703 33930 3712
rect 33888 480 33916 3703
rect 34992 480 35020 3839
rect 37372 3800 37424 3806
rect 37372 3742 37424 3748
rect 36176 2984 36228 2990
rect 36176 2926 36228 2932
rect 36188 480 36216 2926
rect 37384 480 37412 3742
rect 38580 480 38608 5335
rect 40788 5098 40816 7004
rect 42154 5128 42210 5137
rect 40776 5092 40828 5098
rect 42154 5063 42210 5072
rect 40776 5034 40828 5040
rect 39764 4276 39816 4282
rect 39764 4218 39816 4224
rect 39776 480 39804 4218
rect 40960 3732 41012 3738
rect 40960 3674 41012 3680
rect 40972 480 41000 3674
rect 42168 480 42196 5063
rect 44548 3732 44600 3738
rect 44548 3674 44600 3680
rect 43352 3052 43404 3058
rect 43352 2994 43404 3000
rect 43364 480 43392 2994
rect 44560 480 44588 3674
rect 45756 480 45784 7686
rect 49332 7676 49384 7682
rect 49332 7618 49384 7624
rect 48136 6316 48188 6322
rect 48136 6258 48188 6264
rect 46940 4344 46992 4350
rect 46940 4286 46992 4292
rect 46952 480 46980 4286
rect 48148 480 48176 6258
rect 49344 480 49372 7618
rect 62396 7608 62448 7614
rect 62396 7550 62448 7556
rect 77850 7576 77906 7585
rect 52828 7472 52880 7478
rect 52828 7414 52880 7420
rect 50448 6866 50476 7004
rect 50436 6860 50488 6866
rect 50436 6802 50488 6808
rect 50528 4412 50580 4418
rect 50528 4354 50580 4360
rect 50540 480 50568 4354
rect 51632 3188 51684 3194
rect 51632 3130 51684 3136
rect 51644 480 51672 3130
rect 52840 480 52868 7414
rect 60108 6798 60136 7004
rect 60096 6792 60148 6798
rect 60096 6734 60148 6740
rect 55220 6384 55272 6390
rect 55220 6326 55272 6332
rect 54024 4480 54076 4486
rect 54024 4422 54076 4428
rect 54036 480 54064 4422
rect 55232 480 55260 6326
rect 57612 5160 57664 5166
rect 57612 5102 57664 5108
rect 56416 3528 56468 3534
rect 56416 3470 56468 3476
rect 56428 480 56456 3470
rect 57624 480 57652 5102
rect 58808 5092 58860 5098
rect 58808 5034 58860 5040
rect 58820 480 58848 5034
rect 60004 3528 60056 3534
rect 60004 3470 60056 3476
rect 60016 480 60044 3470
rect 61200 3120 61252 3126
rect 61200 3062 61252 3068
rect 61212 480 61240 3062
rect 62408 480 62436 7550
rect 77850 7511 77906 7520
rect 69768 6730 69796 7004
rect 69756 6724 69808 6730
rect 69756 6666 69808 6672
rect 76656 6520 76708 6526
rect 76656 6462 76708 6468
rect 65984 6452 66036 6458
rect 65984 6394 66036 6400
rect 63590 6216 63646 6225
rect 63590 6151 63646 6160
rect 63604 480 63632 6151
rect 64788 4548 64840 4554
rect 64788 4490 64840 4496
rect 64800 480 64828 4490
rect 65996 480 66024 6394
rect 74262 6352 74318 6361
rect 74262 6287 74318 6296
rect 70676 5432 70728 5438
rect 70676 5374 70728 5380
rect 67178 5264 67234 5273
rect 67178 5199 67234 5208
rect 67192 480 67220 5199
rect 69480 3256 69532 3262
rect 69480 3198 69532 3204
rect 68284 3188 68336 3194
rect 68284 3130 68336 3136
rect 68296 480 68324 3130
rect 69492 480 69520 3198
rect 70688 480 70716 5374
rect 71872 4616 71924 4622
rect 71872 4558 71924 4564
rect 71884 480 71912 4558
rect 73068 3324 73120 3330
rect 73068 3266 73120 3272
rect 73080 480 73108 3266
rect 74276 480 74304 6287
rect 75460 2848 75512 2854
rect 75460 2790 75512 2796
rect 75472 480 75500 2790
rect 76668 480 76696 6462
rect 77864 480 77892 7511
rect 79428 6662 79456 7004
rect 79416 6656 79468 6662
rect 79416 6598 79468 6604
rect 84934 6624 84990 6633
rect 84934 6559 84990 6568
rect 87328 6588 87380 6594
rect 81438 6488 81494 6497
rect 81438 6423 81494 6432
rect 79048 4684 79100 4690
rect 79048 4626 79100 4632
rect 79060 480 79088 4626
rect 80244 3392 80296 3398
rect 80244 3334 80296 3340
rect 80256 480 80284 3334
rect 81452 480 81480 6423
rect 83832 5364 83884 5370
rect 83832 5306 83884 5312
rect 82636 3256 82688 3262
rect 82636 3198 82688 3204
rect 82648 480 82676 3198
rect 83844 480 83872 5306
rect 84948 480 84976 6559
rect 87328 6530 87380 6536
rect 86132 4752 86184 4758
rect 86132 4694 86184 4700
rect 86144 480 86172 4694
rect 87340 480 87368 6530
rect 89088 4078 89116 7004
rect 93308 5500 93360 5506
rect 93308 5442 93360 5448
rect 90916 5296 90968 5302
rect 90916 5238 90968 5244
rect 89076 4072 89128 4078
rect 89076 4014 89128 4020
rect 88524 3664 88576 3670
rect 88524 3606 88576 3612
rect 88536 480 88564 3606
rect 89720 3324 89772 3330
rect 89720 3266 89772 3272
rect 89732 480 89760 3266
rect 90928 480 90956 5238
rect 92112 3664 92164 3670
rect 92112 3606 92164 3612
rect 92124 480 92152 3606
rect 93320 480 93348 5442
rect 94504 4956 94556 4962
rect 94504 4898 94556 4904
rect 94516 480 94544 4898
rect 95700 4888 95752 4894
rect 95700 4830 95752 4836
rect 95712 480 95740 4830
rect 98748 4010 98776 7004
rect 102782 6760 102838 6769
rect 102782 6695 102838 6704
rect 100484 5432 100536 5438
rect 100484 5374 100536 5380
rect 98736 4004 98788 4010
rect 98736 3946 98788 3952
rect 98092 3596 98144 3602
rect 98092 3538 98144 3544
rect 99288 3596 99340 3602
rect 99288 3538 99340 3544
rect 96896 3392 96948 3398
rect 96896 3334 96948 3340
rect 96908 480 96936 3334
rect 98104 480 98132 3538
rect 99300 480 99328 3538
rect 100496 480 100524 5374
rect 101588 3936 101640 3942
rect 101588 3878 101640 3884
rect 101600 480 101628 3878
rect 102796 480 102824 6695
rect 105176 6112 105228 6118
rect 105176 6054 105228 6060
rect 103980 4072 104032 4078
rect 103980 4014 104032 4020
rect 103992 480 104020 4014
rect 105188 480 105216 6054
rect 107568 5364 107620 5370
rect 107568 5306 107620 5312
rect 106370 4720 106426 4729
rect 106370 4655 106426 4664
rect 106384 480 106412 4655
rect 107580 480 107608 5306
rect 108408 5234 108436 7004
rect 108764 6044 108816 6050
rect 108764 5986 108816 5992
rect 108396 5228 108448 5234
rect 108396 5170 108448 5176
rect 108776 480 108804 5986
rect 115940 5976 115992 5982
rect 115940 5918 115992 5924
rect 114744 5296 114796 5302
rect 114744 5238 114796 5244
rect 113546 4040 113602 4049
rect 111156 4004 111208 4010
rect 113546 3975 113602 3984
rect 111156 3946 111208 3952
rect 109958 3224 110014 3233
rect 109958 3159 110014 3168
rect 109972 480 110000 3159
rect 111168 480 111196 3946
rect 112352 3868 112404 3874
rect 112352 3810 112404 3816
rect 112364 480 112392 3810
rect 113560 480 113588 3975
rect 114756 480 114784 5238
rect 115952 480 115980 5918
rect 117136 4956 117188 4962
rect 117136 4898 117188 4904
rect 117148 480 117176 4898
rect 118068 4826 118096 7004
rect 119436 5908 119488 5914
rect 119436 5850 119488 5856
rect 118056 4820 118108 4826
rect 118056 4762 118108 4768
rect 118240 3936 118292 3942
rect 118240 3878 118292 3884
rect 118252 480 118280 3878
rect 119448 480 119476 5850
rect 121828 5228 121880 5234
rect 121828 5170 121880 5176
rect 120632 4888 120684 4894
rect 120632 4830 120684 4836
rect 120644 480 120672 4830
rect 121840 480 121868 5170
rect 124220 4820 124272 4826
rect 124220 4762 124272 4768
rect 123022 4040 123078 4049
rect 123022 3975 123078 3984
rect 123036 480 123064 3975
rect 124232 480 124260 4762
rect 125416 3868 125468 3874
rect 125416 3810 125468 3816
rect 125428 480 125456 3810
rect 127728 2922 127756 7004
rect 137388 4214 137416 7004
rect 137376 4208 137428 4214
rect 137376 4150 137428 4156
rect 147048 2990 147076 7004
rect 156708 4282 156736 7004
rect 156696 4276 156748 4282
rect 156696 4218 156748 4224
rect 156788 4276 156840 4282
rect 156788 4218 156840 4224
rect 147036 2984 147088 2990
rect 147036 2926 147088 2932
rect 127716 2916 127768 2922
rect 127716 2858 127768 2864
rect 156800 2854 156828 4218
rect 166368 3058 166396 7004
rect 176028 4350 176056 7004
rect 185688 4418 185716 7004
rect 195348 4486 195376 7004
rect 205008 5166 205036 7004
rect 204996 5160 205048 5166
rect 204996 5102 205048 5108
rect 195336 4480 195388 4486
rect 195336 4422 195388 4428
rect 185676 4412 185728 4418
rect 185676 4354 185728 4360
rect 176016 4344 176068 4350
rect 176016 4286 176068 4292
rect 214668 3126 214696 7004
rect 220728 5160 220780 5166
rect 220728 5102 220780 5108
rect 220740 4146 220768 5102
rect 224328 4554 224356 7004
rect 224316 4548 224368 4554
rect 224316 4490 224368 4496
rect 220728 4140 220780 4146
rect 220728 4082 220780 4088
rect 233988 3194 234016 7004
rect 243648 4622 243676 7004
rect 243636 4616 243688 4622
rect 243636 4558 243688 4564
rect 253308 4282 253336 7004
rect 262968 4690 262996 7004
rect 262956 4684 263008 4690
rect 262956 4626 263008 4632
rect 253296 4276 253348 4282
rect 253296 4218 253348 4224
rect 272628 3262 272656 7004
rect 282288 4758 282316 7004
rect 282276 4752 282328 4758
rect 282276 4694 282328 4700
rect 291948 3330 291976 7004
rect 301608 5506 301636 7004
rect 301596 5500 301648 5506
rect 301596 5442 301648 5448
rect 311268 3398 311296 7004
rect 320928 5438 320956 7004
rect 320916 5432 320968 5438
rect 320916 5374 320968 5380
rect 330588 4078 330616 7004
rect 340248 5370 340276 7004
rect 340236 5364 340288 5370
rect 340236 5306 340288 5312
rect 330576 4072 330628 4078
rect 330576 4014 330628 4020
rect 349908 4010 349936 7004
rect 359568 5302 359596 7004
rect 359556 5296 359608 5302
rect 359556 5238 359608 5244
rect 349896 4004 349948 4010
rect 349896 3946 349948 3952
rect 369228 3942 369256 7004
rect 378888 5234 378916 7004
rect 378876 5228 378928 5234
rect 378876 5170 378928 5176
rect 369216 3936 369268 3942
rect 369216 3878 369268 3884
rect 388548 3874 388576 7004
rect 388536 3868 388588 3874
rect 388536 3810 388588 3816
rect 311256 3392 311308 3398
rect 311256 3334 311308 3340
rect 291936 3324 291988 3330
rect 291936 3266 291988 3272
rect 272616 3256 272668 3262
rect 272616 3198 272668 3204
rect 233976 3188 234028 3194
rect 233976 3130 234028 3136
rect 214656 3120 214708 3126
rect 214656 3062 214708 3068
rect 166356 3052 166408 3058
rect 166356 2994 166408 3000
rect 156788 2848 156840 2854
rect 156788 2790 156840 2796
rect 398208 2106 398236 7004
rect 407868 5030 407896 7004
rect 407856 5024 407908 5030
rect 407856 4966 407908 4972
rect 417528 3806 417556 7004
rect 417516 3800 417568 3806
rect 417516 3742 417568 3748
rect 427188 3738 427216 7004
rect 436848 5098 436876 7004
rect 436836 5092 436888 5098
rect 436836 5034 436888 5040
rect 427176 3732 427228 3738
rect 427176 3674 427228 3680
rect 446508 3466 446536 7004
rect 456168 5001 456196 7004
rect 465828 5545 465856 7004
rect 465814 5536 465870 5545
rect 465814 5471 465870 5480
rect 475488 5409 475516 7004
rect 475474 5400 475530 5409
rect 475474 5335 475530 5344
rect 485148 5137 485176 7004
rect 485134 5128 485190 5137
rect 485134 5063 485190 5072
rect 456154 4992 456210 5001
rect 456154 4927 456210 4936
rect 494808 3534 494836 7004
rect 504468 5273 504496 7004
rect 504454 5264 504510 5273
rect 504454 5199 504510 5208
rect 514128 3670 514156 7004
rect 514116 3664 514168 3670
rect 514116 3606 514168 3612
rect 523788 3602 523816 7004
rect 533448 4962 533476 7004
rect 533436 4956 533488 4962
rect 533436 4898 533488 4904
rect 543108 4894 543136 7004
rect 543096 4888 543148 4894
rect 543096 4830 543148 4836
rect 552768 4826 552796 7004
rect 562428 4865 562456 7004
rect 572088 5166 572116 7004
rect 572076 5160 572128 5166
rect 572076 5102 572128 5108
rect 562414 4856 562470 4865
rect 552756 4820 552808 4826
rect 562414 4791 562470 4800
rect 552756 4762 552808 4768
rect 578252 3641 578280 527167
rect 578330 505744 578386 505753
rect 578330 505679 578386 505688
rect 578344 4049 578372 505679
rect 579712 487144 579764 487150
rect 579712 487086 579764 487092
rect 579724 486849 579752 487086
rect 579710 486840 579766 486849
rect 579710 486775 579766 486784
rect 578422 484528 578478 484537
rect 578422 484463 578478 484472
rect 578436 5914 578464 484463
rect 578514 463720 578570 463729
rect 578514 463655 578570 463664
rect 578528 5982 578556 463655
rect 578606 442232 578662 442241
rect 578606 442167 578662 442176
rect 578620 6050 578648 442167
rect 578698 421016 578754 421025
rect 578698 420951 578754 420960
rect 578712 6118 578740 420951
rect 578790 399528 578846 399537
rect 578790 399463 578846 399472
rect 578804 6594 578832 399463
rect 578882 378312 578938 378321
rect 578882 378247 578938 378256
rect 578792 6588 578844 6594
rect 578792 6530 578844 6536
rect 578896 6526 578924 378247
rect 578974 357504 579030 357513
rect 578974 357439 579030 357448
rect 578884 6520 578936 6526
rect 578884 6462 578936 6468
rect 578988 6458 579016 357439
rect 579066 335880 579122 335889
rect 579066 335815 579122 335824
rect 578976 6452 579028 6458
rect 578976 6394 579028 6400
rect 579080 6390 579108 335815
rect 579158 314800 579214 314809
rect 579158 314735 579214 314744
rect 579068 6384 579120 6390
rect 579068 6326 579120 6332
rect 579172 6322 579200 314735
rect 579250 293312 579306 293321
rect 579250 293247 579306 293256
rect 579160 6316 579212 6322
rect 579160 6258 579212 6264
rect 578700 6112 578752 6118
rect 578700 6054 578752 6060
rect 578608 6044 578660 6050
rect 578608 5986 578660 5992
rect 578516 5976 578568 5982
rect 578516 5918 578568 5924
rect 578424 5908 578476 5914
rect 578424 5850 578476 5856
rect 578330 4040 578386 4049
rect 578330 3975 578386 3984
rect 579264 3777 579292 293247
rect 579342 272096 579398 272105
rect 579342 272031 579398 272040
rect 579250 3768 579306 3777
rect 579250 3703 579306 3712
rect 578238 3632 578294 3641
rect 523776 3596 523828 3602
rect 578238 3567 578294 3576
rect 523776 3538 523828 3544
rect 494796 3528 494848 3534
rect 579356 3505 579384 272031
rect 580170 252240 580226 252249
rect 580170 252175 580226 252184
rect 579434 251288 579490 251297
rect 579434 251223 579490 251232
rect 579448 6254 579476 251223
rect 579526 229664 579582 229673
rect 579526 229599 579582 229608
rect 579436 6248 579488 6254
rect 579436 6190 579488 6196
rect 579540 6186 579568 229599
rect 580184 124137 580212 252175
rect 580170 124128 580226 124137
rect 580170 124063 580226 124072
rect 580276 6662 580304 674591
rect 580354 627736 580410 627745
rect 580354 627671 580410 627680
rect 580368 6730 580396 627671
rect 580446 580816 580502 580825
rect 580446 580751 580502 580760
rect 580460 6798 580488 580751
rect 580538 533896 580594 533905
rect 580538 533831 580594 533840
rect 580552 6866 580580 533831
rect 580630 439920 580686 439929
rect 580630 439855 580686 439864
rect 580644 209438 580672 439855
rect 580722 393000 580778 393009
rect 580722 392935 580778 392944
rect 580632 209432 580684 209438
rect 580632 209374 580684 209380
rect 580630 205320 580686 205329
rect 580630 205255 580686 205264
rect 580644 103222 580672 205255
rect 580736 187678 580764 392935
rect 580814 346080 580870 346089
rect 580814 346015 580870 346024
rect 580724 187672 580776 187678
rect 580724 187614 580776 187620
rect 580828 167006 580856 346015
rect 580906 299160 580962 299169
rect 580906 299095 580962 299104
rect 580816 167000 580868 167006
rect 580816 166942 580868 166948
rect 580722 158400 580778 158409
rect 580722 158335 580778 158344
rect 580632 103216 580684 103222
rect 580632 103158 580684 103164
rect 580736 81394 580764 158335
rect 580920 145790 580948 299095
rect 580908 145784 580960 145790
rect 580908 145726 580960 145732
rect 580814 111480 580870 111489
rect 580814 111415 580870 111424
rect 580724 81388 580776 81394
rect 580724 81330 580776 81336
rect 580630 64560 580686 64569
rect 580630 64495 580686 64504
rect 580644 39574 580672 64495
rect 580828 60654 580856 111415
rect 580816 60648 580868 60654
rect 580816 60590 580868 60596
rect 580632 39568 580684 39574
rect 580632 39510 580684 39516
rect 580540 6860 580592 6866
rect 580540 6802 580592 6808
rect 580448 6792 580500 6798
rect 580448 6734 580500 6740
rect 580356 6724 580408 6730
rect 580356 6666 580408 6672
rect 580264 6656 580316 6662
rect 580264 6598 580316 6604
rect 579528 6180 579580 6186
rect 579528 6122 579580 6128
rect 494796 3470 494848 3476
rect 579342 3496 579398 3505
rect 446496 3460 446548 3466
rect 579342 3431 579398 3440
rect 446496 3402 446548 3408
rect 398196 2100 398248 2106
rect 398196 2042 398248 2048
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 8850 685208 8906 685264
rect 3514 682216 3570 682272
rect 5538 676368 5594 676424
rect 3146 624824 3202 624880
rect 5446 572872 5502 572928
rect 3330 567316 3386 567352
rect 3330 567296 3332 567316
rect 3332 567296 3384 567316
rect 3384 567296 3386 567316
rect 5354 552336 5410 552392
rect 5262 531664 5318 531720
rect 5170 511128 5226 511184
rect 3146 509904 3202 509960
rect 5078 490456 5134 490512
rect 4986 469920 5042 469976
rect 3422 452376 3478 452432
rect 3238 165008 3294 165064
rect 3330 160792 3386 160848
rect 3238 141480 3294 141536
rect 3330 122032 3386 122088
rect 4894 429256 4950 429312
rect 4802 408584 4858 408640
rect 3514 394984 3570 395040
rect 4710 387776 4766 387832
rect 4618 367240 4674 367296
rect 4526 346432 4582 346488
rect 3606 337456 3662 337512
rect 4434 325760 4490 325816
rect 4342 305088 4398 305144
rect 3698 294344 3754 294400
rect 4250 284416 4306 284472
rect 4158 263880 4214 263936
rect 3882 251232 3938 251288
rect 3790 202000 3846 202056
rect 3698 79600 3754 79656
rect 3606 59064 3662 59120
rect 3514 38256 3570 38312
rect 4066 208120 4122 208176
rect 3974 181464 4030 181520
rect 3882 100272 3938 100328
rect 4066 120808 4122 120864
rect 3974 78920 4030 78976
rect 3790 35808 3846 35864
rect 3422 17856 3478 17912
rect 6826 655696 6882 655752
rect 5814 531256 5870 531312
rect 5998 531292 6000 531312
rect 6000 531292 6052 531312
rect 6052 531292 6054 531312
rect 5998 531256 6054 531292
rect 6182 511944 6238 512000
rect 6458 511944 6514 512000
rect 6090 492632 6146 492688
rect 6274 492632 6330 492688
rect 6182 202816 6238 202872
rect 6458 202816 6514 202872
rect 6182 183504 6238 183560
rect 6458 183504 6514 183560
rect 6090 164192 6146 164248
rect 6274 164192 6330 164248
rect 5906 144880 5962 144936
rect 6090 144880 6146 144936
rect 5906 125568 5962 125624
rect 6090 125568 6146 125624
rect 6918 449656 6974 449712
rect 7010 243208 7066 243264
rect 7102 222672 7158 222728
rect 8942 685072 8998 685128
rect 8850 4936 8906 4992
rect 534170 688608 534226 688664
rect 391478 686296 391534 686352
rect 419998 686296 420054 686352
rect 580262 674600 580318 674656
rect 578238 527176 578294 527232
rect 578146 209380 578148 209400
rect 578148 209380 578200 209400
rect 578200 209380 578202 209400
rect 578146 209344 578202 209380
rect 578146 187620 578148 187640
rect 578148 187620 578200 187640
rect 578200 187620 578202 187640
rect 578146 187584 578202 187620
rect 578146 166948 578148 166968
rect 578148 166948 578200 166968
rect 578200 166948 578202 166968
rect 578146 166912 578202 166948
rect 578146 145732 578148 145752
rect 578148 145732 578200 145752
rect 578200 145732 578202 145752
rect 578146 145696 578202 145732
rect 578146 103164 578148 103184
rect 578148 103164 578200 103184
rect 578200 103164 578202 103184
rect 578146 103128 578202 103164
rect 578146 81388 578202 81424
rect 578146 81368 578148 81388
rect 578148 81368 578200 81388
rect 578200 81368 578202 81388
rect 578146 60596 578148 60616
rect 578148 60596 578200 60616
rect 578200 60596 578202 60616
rect 578146 60560 578202 60596
rect 578146 39516 578148 39536
rect 578148 39516 578200 39536
rect 578200 39516 578202 39536
rect 578146 39480 578202 39516
rect 17222 3440 17278 3496
rect 16026 3304 16082 3360
rect 31482 5480 31538 5536
rect 25502 4800 25558 4856
rect 27894 3576 27950 3632
rect 38566 5344 38622 5400
rect 34978 3848 35034 3904
rect 33874 3712 33930 3768
rect 42154 5072 42210 5128
rect 77850 7520 77906 7576
rect 63590 6160 63646 6216
rect 74262 6296 74318 6352
rect 67178 5208 67234 5264
rect 84934 6568 84990 6624
rect 81438 6432 81494 6488
rect 102782 6704 102838 6760
rect 106370 4664 106426 4720
rect 113546 3984 113602 4040
rect 109958 3168 110014 3224
rect 123022 3984 123078 4040
rect 465814 5480 465870 5536
rect 475474 5344 475530 5400
rect 485134 5072 485190 5128
rect 456154 4936 456210 4992
rect 504454 5208 504510 5264
rect 562414 4800 562470 4856
rect 578330 505688 578386 505744
rect 579710 486784 579766 486840
rect 578422 484472 578478 484528
rect 578514 463664 578570 463720
rect 578606 442176 578662 442232
rect 578698 420960 578754 421016
rect 578790 399472 578846 399528
rect 578882 378256 578938 378312
rect 578974 357448 579030 357504
rect 579066 335824 579122 335880
rect 579158 314744 579214 314800
rect 579250 293256 579306 293312
rect 578330 3984 578386 4040
rect 579342 272040 579398 272096
rect 579250 3712 579306 3768
rect 578238 3576 578294 3632
rect 580170 252184 580226 252240
rect 579434 251232 579490 251288
rect 579526 229608 579582 229664
rect 580170 124072 580226 124128
rect 580354 627680 580410 627736
rect 580446 580760 580502 580816
rect 580538 533840 580594 533896
rect 580630 439864 580686 439920
rect 580722 392944 580778 393000
rect 580630 205264 580686 205320
rect 580814 346024 580870 346080
rect 580906 299104 580962 299160
rect 580722 158344 580778 158400
rect 580814 111424 580870 111480
rect 580630 64504 580686 64560
rect 579342 3440 579398 3496
<< metal3 >>
rect 583520 697900 584960 698140
rect -960 696540 480 696780
rect 534165 688666 534231 688669
rect 569718 688666 569724 688668
rect 534165 688664 569724 688666
rect 534165 688608 534170 688664
rect 534226 688608 569724 688664
rect 534165 688606 569724 688608
rect 534165 688603 534231 688606
rect 569718 688604 569724 688606
rect 569788 688604 569794 688668
rect 391473 686356 391539 686357
rect 419993 686356 420059 686357
rect 391422 686354 391428 686356
rect 391382 686294 391428 686354
rect 391492 686352 391539 686356
rect 419942 686354 419948 686356
rect 391534 686296 391539 686352
rect 391422 686292 391428 686294
rect 391492 686292 391539 686296
rect 419902 686294 419948 686354
rect 420012 686352 420059 686356
rect 420054 686296 420059 686352
rect 419942 686292 419948 686294
rect 420012 686292 420059 686296
rect 391473 686291 391539 686292
rect 419993 686291 420059 686292
rect 583520 686204 584960 686444
rect 8845 685266 8911 685269
rect 391422 685266 391428 685268
rect 8845 685264 391428 685266
rect 8845 685208 8850 685264
rect 8906 685208 391428 685264
rect 8845 685206 391428 685208
rect 8845 685203 8911 685206
rect 391422 685204 391428 685206
rect 391492 685204 391498 685268
rect 8937 685130 9003 685133
rect 419942 685130 419948 685132
rect 8937 685128 419948 685130
rect 8937 685072 8942 685128
rect 8998 685072 419948 685128
rect 8937 685070 419948 685072
rect 8937 685067 9003 685070
rect 419942 685068 419948 685070
rect 420012 685068 420018 685132
rect -960 682274 480 682364
rect 3509 682274 3575 682277
rect -960 682272 3575 682274
rect -960 682216 3514 682272
rect 3570 682216 3575 682272
rect -960 682214 3575 682216
rect -960 682124 480 682214
rect 3509 682211 3575 682214
rect 5533 676426 5599 676429
rect 7054 676426 7114 676600
rect 5533 676424 7114 676426
rect 5533 676368 5538 676424
rect 5594 676368 7114 676424
rect 5533 676366 7114 676368
rect 5533 676363 5599 676366
rect 576902 676290 576962 676328
rect 578182 676290 578188 676292
rect 576902 676230 578188 676290
rect 578182 676228 578188 676230
rect 578252 676228 578258 676292
rect 580257 674658 580323 674661
rect 583520 674658 584960 674748
rect 580257 674656 584960 674658
rect 580257 674600 580262 674656
rect 580318 674600 584960 674656
rect 580257 674598 584960 674600
rect 580257 674595 580323 674598
rect 583520 674508 584960 674598
rect -960 667844 480 668084
rect 583520 662676 584960 662916
rect 6821 655754 6887 655757
rect 7054 655754 7114 655928
rect 6821 655752 7114 655754
rect 6821 655696 6826 655752
rect 6882 655696 7114 655752
rect 6821 655694 7114 655696
rect 6821 655691 6887 655694
rect 576902 654666 576962 655112
rect 578366 654666 578372 654668
rect 576902 654606 578372 654666
rect 578366 654604 578372 654606
rect 578436 654604 578442 654668
rect -960 653428 480 653668
rect 583520 650980 584960 651220
rect 583520 639284 584960 639524
rect -960 639012 480 639252
rect 5390 634884 5396 634948
rect 5460 634946 5466 634948
rect 7054 634946 7114 635392
rect 5460 634886 7114 634946
rect 5460 634884 5466 634886
rect 576902 633450 576962 633896
rect 578550 633450 578556 633452
rect 576902 633390 578556 633450
rect 578550 633388 578556 633390
rect 578620 633388 578626 633452
rect 580349 627738 580415 627741
rect 583520 627738 584960 627828
rect 580349 627736 584960 627738
rect 580349 627680 580354 627736
rect 580410 627680 584960 627736
rect 580349 627678 584960 627680
rect 580349 627675 580415 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 3141 624882 3207 624885
rect -960 624880 3207 624882
rect -960 624824 3146 624880
rect 3202 624824 3207 624880
rect -960 624822 3207 624824
rect -960 624732 480 624822
rect 3141 624819 3207 624822
rect 583520 615756 584960 615996
rect 5206 614076 5212 614140
rect 5276 614138 5282 614140
rect 7054 614138 7114 614720
rect 5276 614078 7114 614138
rect 5276 614076 5282 614078
rect 576902 612098 576962 612680
rect 578734 612098 578740 612100
rect 576902 612038 578740 612098
rect 578734 612036 578740 612038
rect 578804 612036 578810 612100
rect -960 610316 480 610556
rect 583520 604060 584960 604300
rect -960 595900 480 596140
rect 5022 593540 5028 593604
rect 5092 593602 5098 593604
rect 7054 593602 7114 594184
rect 5092 593542 7114 593602
rect 5092 593540 5098 593542
rect 583520 592364 584960 592604
rect 576902 590746 576962 591328
rect 578918 590746 578924 590748
rect 576902 590686 578924 590746
rect 578918 590684 578924 590686
rect 578988 590684 578994 590748
rect -960 581620 480 581860
rect 580441 580818 580507 580821
rect 583520 580818 584960 580908
rect 580441 580816 584960 580818
rect 580441 580760 580446 580816
rect 580502 580760 584960 580816
rect 580441 580758 584960 580760
rect 580441 580755 580507 580758
rect 583520 580668 584960 580758
rect 5441 572930 5507 572933
rect 7054 572930 7114 573512
rect 5441 572928 7114 572930
rect 5441 572872 5446 572928
rect 5502 572872 7114 572928
rect 5441 572870 7114 572872
rect 5441 572867 5507 572870
rect 576902 570074 576962 570112
rect 579102 570074 579108 570076
rect 576902 570014 579108 570074
rect 579102 570012 579108 570014
rect 579172 570012 579178 570076
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 3325 567354 3391 567357
rect -960 567352 3391 567354
rect -960 567296 3330 567352
rect 3386 567296 3391 567352
rect -960 567294 3391 567296
rect -960 567204 480 567294
rect 3325 567291 3391 567294
rect 583520 557140 584960 557380
rect -960 552924 480 553164
rect 5349 552394 5415 552397
rect 7054 552394 7114 552976
rect 5349 552392 7114 552394
rect 5349 552336 5354 552392
rect 5410 552336 7114 552392
rect 5349 552334 7114 552336
rect 5349 552331 5415 552334
rect 576902 548450 576962 548896
rect 579286 548450 579292 548452
rect 576902 548390 579292 548450
rect 579286 548388 579292 548390
rect 579356 548388 579362 548452
rect 583520 545444 584960 545684
rect -960 538508 480 538748
rect 580533 533898 580599 533901
rect 583520 533898 584960 533988
rect 580533 533896 584960 533898
rect 580533 533840 580538 533896
rect 580594 533840 584960 533896
rect 580533 533838 584960 533840
rect 580533 533835 580599 533838
rect 583520 533748 584960 533838
rect 5257 531722 5323 531725
rect 7054 531722 7114 532304
rect 5257 531720 7114 531722
rect 5257 531664 5262 531720
rect 5318 531664 7114 531720
rect 5257 531662 7114 531664
rect 5257 531659 5323 531662
rect 5809 531314 5875 531317
rect 5993 531314 6059 531317
rect 5809 531312 6059 531314
rect 5809 531256 5814 531312
rect 5870 531256 5998 531312
rect 6054 531256 6059 531312
rect 5809 531254 6059 531256
rect 5809 531251 5875 531254
rect 5993 531251 6059 531254
rect 576902 527234 576962 527680
rect 578233 527234 578299 527237
rect 576902 527232 578299 527234
rect 576902 527176 578238 527232
rect 578294 527176 578299 527232
rect 576902 527174 578299 527176
rect 578233 527171 578299 527174
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 6177 512002 6243 512005
rect 6453 512002 6519 512005
rect 6177 512000 6519 512002
rect 6177 511944 6182 512000
rect 6238 511944 6458 512000
rect 6514 511944 6519 512000
rect 6177 511942 6519 511944
rect 6177 511939 6243 511942
rect 6453 511939 6519 511942
rect 5165 511186 5231 511189
rect 7054 511186 7114 511768
rect 5165 511184 7114 511186
rect 5165 511128 5170 511184
rect 5226 511128 7114 511184
rect 5165 511126 7114 511128
rect 5165 511123 5231 511126
rect 583520 510220 584960 510460
rect -960 509962 480 510052
rect 3141 509962 3207 509965
rect -960 509960 3207 509962
rect -960 509904 3146 509960
rect 3202 509904 3207 509960
rect -960 509902 3207 509904
rect -960 509812 480 509902
rect 3141 509899 3207 509902
rect 576902 505746 576962 506328
rect 578325 505746 578391 505749
rect 576902 505744 578391 505746
rect 576902 505688 578330 505744
rect 578386 505688 578391 505744
rect 576902 505686 578391 505688
rect 578325 505683 578391 505686
rect 583520 498524 584960 498764
rect -960 495396 480 495636
rect 6085 492690 6151 492693
rect 6269 492690 6335 492693
rect 6085 492688 6335 492690
rect 6085 492632 6090 492688
rect 6146 492632 6274 492688
rect 6330 492632 6335 492688
rect 6085 492630 6335 492632
rect 6085 492627 6151 492630
rect 6269 492627 6335 492630
rect 5073 490514 5139 490517
rect 7054 490514 7114 491096
rect 5073 490512 7114 490514
rect 5073 490456 5078 490512
rect 5134 490456 7114 490512
rect 5073 490454 7114 490456
rect 5073 490451 5139 490454
rect 579705 486842 579771 486845
rect 583520 486842 584960 486932
rect 579705 486840 584960 486842
rect 579705 486784 579710 486840
rect 579766 486784 584960 486840
rect 579705 486782 584960 486784
rect 579705 486779 579771 486782
rect 583520 486692 584960 486782
rect 576902 484530 576962 485112
rect 578417 484530 578483 484533
rect 576902 484528 578483 484530
rect 576902 484472 578422 484528
rect 578478 484472 578483 484528
rect 576902 484470 578483 484472
rect 578417 484467 578483 484470
rect -960 480980 480 481220
rect 583520 474996 584960 475236
rect 4981 469978 5047 469981
rect 7054 469978 7114 470560
rect 4981 469976 7114 469978
rect 4981 469920 4986 469976
rect 5042 469920 7114 469976
rect 4981 469918 7114 469920
rect 4981 469915 5047 469918
rect -960 466700 480 466940
rect 576902 463722 576962 463896
rect 578509 463722 578575 463725
rect 576902 463720 578575 463722
rect 576902 463664 578514 463720
rect 578570 463664 578575 463720
rect 576902 463662 578575 463664
rect 578509 463659 578575 463662
rect 583520 463300 584960 463540
rect -960 452434 480 452524
rect 3417 452434 3483 452437
rect -960 452432 3483 452434
rect -960 452376 3422 452432
rect 3478 452376 3483 452432
rect -960 452374 3483 452376
rect -960 452284 480 452374
rect 3417 452371 3483 452374
rect 583520 451604 584960 451844
rect 6913 449714 6979 449717
rect 7054 449714 7114 449888
rect 6913 449712 7114 449714
rect 6913 449656 6918 449712
rect 6974 449656 7114 449712
rect 6913 449654 7114 449656
rect 6913 449651 6979 449654
rect 576902 442234 576962 442680
rect 578601 442234 578667 442237
rect 576902 442232 578667 442234
rect 576902 442176 578606 442232
rect 578662 442176 578667 442232
rect 576902 442174 578667 442176
rect 578601 442171 578667 442174
rect 580625 439922 580691 439925
rect 583520 439922 584960 440012
rect 580625 439920 584960 439922
rect 580625 439864 580630 439920
rect 580686 439864 584960 439920
rect 580625 439862 584960 439864
rect 580625 439859 580691 439862
rect 583520 439772 584960 439862
rect -960 437868 480 438108
rect 4889 429314 4955 429317
rect 7054 429314 7114 429352
rect 4889 429312 7114 429314
rect 4889 429256 4894 429312
rect 4950 429256 7114 429312
rect 4889 429254 7114 429256
rect 4889 429251 4955 429254
rect 583520 428076 584960 428316
rect -960 423588 480 423828
rect 576902 421018 576962 421328
rect 578693 421018 578759 421021
rect 576902 421016 578759 421018
rect 576902 420960 578698 421016
rect 578754 420960 578759 421016
rect 576902 420958 578759 420960
rect 578693 420955 578759 420958
rect 583520 416380 584960 416620
rect -960 409172 480 409412
rect 4797 408642 4863 408645
rect 7054 408642 7114 408680
rect 4797 408640 7114 408642
rect 4797 408584 4802 408640
rect 4858 408584 7114 408640
rect 4797 408582 7114 408584
rect 4797 408579 4863 408582
rect 583520 404684 584960 404924
rect 576902 399530 576962 400112
rect 578785 399530 578851 399533
rect 576902 399528 578851 399530
rect 576902 399472 578790 399528
rect 578846 399472 578851 399528
rect 576902 399470 578851 399472
rect 578785 399467 578851 399470
rect -960 395042 480 395132
rect 3509 395042 3575 395045
rect -960 395040 3575 395042
rect -960 394984 3514 395040
rect 3570 394984 3575 395040
rect -960 394982 3575 394984
rect -960 394892 480 394982
rect 3509 394979 3575 394982
rect 580717 393002 580783 393005
rect 583520 393002 584960 393092
rect 580717 393000 584960 393002
rect 580717 392944 580722 393000
rect 580778 392944 584960 393000
rect 580717 392942 584960 392944
rect 580717 392939 580783 392942
rect 583520 392852 584960 392942
rect 4705 387834 4771 387837
rect 7054 387834 7114 388144
rect 4705 387832 7114 387834
rect 4705 387776 4710 387832
rect 4766 387776 7114 387832
rect 4705 387774 7114 387776
rect 4705 387771 4771 387774
rect 583520 381156 584960 381396
rect -960 380476 480 380716
rect 576902 378314 576962 378896
rect 578877 378314 578943 378317
rect 576902 378312 578943 378314
rect 576902 378256 578882 378312
rect 578938 378256 578943 378312
rect 576902 378254 578943 378256
rect 578877 378251 578943 378254
rect 583520 369460 584960 369700
rect 4613 367298 4679 367301
rect 7054 367298 7114 367472
rect 4613 367296 7114 367298
rect 4613 367240 4618 367296
rect 4674 367240 7114 367296
rect 4613 367238 7114 367240
rect 4613 367235 4679 367238
rect -960 366060 480 366300
rect 583520 357764 584960 358004
rect 576902 357506 576962 357680
rect 578969 357506 579035 357509
rect 576902 357504 579035 357506
rect 576902 357448 578974 357504
rect 579030 357448 579035 357504
rect 576902 357446 579035 357448
rect 578969 357443 579035 357446
rect -960 351780 480 352020
rect 4521 346490 4587 346493
rect 7054 346490 7114 346936
rect 4521 346488 7114 346490
rect 4521 346432 4526 346488
rect 4582 346432 7114 346488
rect 4521 346430 7114 346432
rect 4521 346427 4587 346430
rect 580809 346082 580875 346085
rect 583520 346082 584960 346172
rect 580809 346080 584960 346082
rect 580809 346024 580814 346080
rect 580870 346024 584960 346080
rect 580809 346022 584960 346024
rect 580809 346019 580875 346022
rect 583520 345932 584960 346022
rect -960 337514 480 337604
rect 3601 337514 3667 337517
rect -960 337512 3667 337514
rect -960 337456 3606 337512
rect 3662 337456 3667 337512
rect -960 337454 3667 337456
rect -960 337364 480 337454
rect 3601 337451 3667 337454
rect 576902 335882 576962 336328
rect 579061 335882 579127 335885
rect 576902 335880 579127 335882
rect 576902 335824 579066 335880
rect 579122 335824 579127 335880
rect 576902 335822 579127 335824
rect 579061 335819 579127 335822
rect 583520 334236 584960 334476
rect 4429 325818 4495 325821
rect 7054 325818 7114 326264
rect 4429 325816 7114 325818
rect 4429 325760 4434 325816
rect 4490 325760 7114 325816
rect 4429 325758 7114 325760
rect 4429 325755 4495 325758
rect -960 322948 480 323188
rect 583520 322540 584960 322780
rect 576902 314802 576962 315112
rect 579153 314802 579219 314805
rect 576902 314800 579219 314802
rect 576902 314744 579158 314800
rect 579214 314744 579219 314800
rect 576902 314742 579219 314744
rect 579153 314739 579219 314742
rect 583520 310708 584960 310948
rect -960 308668 480 308908
rect 4337 305146 4403 305149
rect 7054 305146 7114 305728
rect 4337 305144 7114 305146
rect 4337 305088 4342 305144
rect 4398 305088 7114 305144
rect 4337 305086 7114 305088
rect 4337 305083 4403 305086
rect 580901 299162 580967 299165
rect 583520 299162 584960 299252
rect 580901 299160 584960 299162
rect 580901 299104 580906 299160
rect 580962 299104 584960 299160
rect 580901 299102 584960 299104
rect 580901 299099 580967 299102
rect 583520 299012 584960 299102
rect -960 294402 480 294492
rect 3693 294402 3759 294405
rect -960 294400 3759 294402
rect -960 294344 3698 294400
rect 3754 294344 3759 294400
rect -960 294342 3759 294344
rect -960 294252 480 294342
rect 3693 294339 3759 294342
rect 576902 293314 576962 293896
rect 579245 293314 579311 293317
rect 576902 293312 579311 293314
rect 576902 293256 579250 293312
rect 579306 293256 579311 293312
rect 576902 293254 579311 293256
rect 579245 293251 579311 293254
rect 583520 287316 584960 287556
rect 4245 284474 4311 284477
rect 7054 284474 7114 285056
rect 4245 284472 7114 284474
rect 4245 284416 4250 284472
rect 4306 284416 7114 284472
rect 4245 284414 7114 284416
rect 4245 284411 4311 284414
rect -960 279972 480 280212
rect 583520 275620 584960 275860
rect 576902 272098 576962 272680
rect 579337 272098 579403 272101
rect 576902 272096 579403 272098
rect 576902 272040 579342 272096
rect 579398 272040 579403 272096
rect 576902 272038 579403 272040
rect 579337 272035 579403 272038
rect -960 265556 480 265796
rect 4153 263938 4219 263941
rect 7054 263938 7114 264520
rect 4153 263936 7114 263938
rect 4153 263880 4158 263936
rect 4214 263880 7114 263936
rect 4153 263878 7114 263880
rect 4153 263875 4219 263878
rect 583520 263788 584960 264028
rect 580165 252242 580231 252245
rect 583520 252242 584960 252332
rect 580165 252240 584960 252242
rect 580165 252184 580170 252240
rect 580226 252184 584960 252240
rect 580165 252182 584960 252184
rect 580165 252179 580231 252182
rect 583520 252092 584960 252182
rect -960 251290 480 251380
rect 3877 251290 3943 251293
rect -960 251288 3943 251290
rect -960 251232 3882 251288
rect 3938 251232 3943 251288
rect -960 251230 3943 251232
rect 576902 251290 576962 251328
rect 579429 251290 579495 251293
rect 576902 251288 579495 251290
rect 576902 251232 579434 251288
rect 579490 251232 579495 251288
rect 576902 251230 579495 251232
rect -960 251140 480 251230
rect 3877 251227 3943 251230
rect 579429 251227 579495 251230
rect 7054 243269 7114 243848
rect 7005 243264 7114 243269
rect 7005 243208 7010 243264
rect 7066 243208 7114 243264
rect 7005 243206 7114 243208
rect 7005 243203 7071 243206
rect 583520 240396 584960 240636
rect -960 236860 480 237100
rect 576902 229666 576962 230112
rect 579521 229666 579587 229669
rect 576902 229664 579587 229666
rect 576902 229608 579526 229664
rect 579582 229608 579587 229664
rect 576902 229606 579587 229608
rect 579521 229603 579587 229606
rect 583520 228700 584960 228940
rect 7054 222733 7114 223312
rect 7054 222728 7163 222733
rect -960 222444 480 222684
rect 7054 222672 7102 222728
rect 7158 222672 7163 222728
rect 7054 222670 7163 222672
rect 7097 222667 7163 222670
rect 583520 216868 584960 217108
rect 578141 209402 578207 209405
rect 576902 209400 578207 209402
rect 576902 209344 578146 209400
rect 578202 209344 578207 209400
rect 576902 209342 578207 209344
rect 576902 208896 576962 209342
rect 578141 209339 578207 209342
rect -960 208178 480 208268
rect 4061 208178 4127 208181
rect -960 208176 4127 208178
rect -960 208120 4066 208176
rect 4122 208120 4127 208176
rect -960 208118 4127 208120
rect -960 208028 480 208118
rect 4061 208115 4127 208118
rect 580625 205322 580691 205325
rect 583520 205322 584960 205412
rect 580625 205320 584960 205322
rect 580625 205264 580630 205320
rect 580686 205264 584960 205320
rect 580625 205262 584960 205264
rect 580625 205259 580691 205262
rect 583520 205172 584960 205262
rect 6177 202874 6243 202877
rect 6453 202874 6519 202877
rect 6177 202872 6519 202874
rect 6177 202816 6182 202872
rect 6238 202816 6458 202872
rect 6514 202816 6519 202872
rect 6177 202814 6519 202816
rect 6177 202811 6243 202814
rect 6453 202811 6519 202814
rect 3785 202058 3851 202061
rect 7054 202058 7114 202640
rect 3785 202056 7114 202058
rect 3785 202000 3790 202056
rect 3846 202000 7114 202056
rect 3785 201998 7114 202000
rect 3785 201995 3851 201998
rect -960 193748 480 193988
rect 583520 193476 584960 193716
rect 576902 187642 576962 187680
rect 578141 187642 578207 187645
rect 576902 187640 578207 187642
rect 576902 187584 578146 187640
rect 578202 187584 578207 187640
rect 576902 187582 578207 187584
rect 578141 187579 578207 187582
rect 6177 183562 6243 183565
rect 6453 183562 6519 183565
rect 6177 183560 6519 183562
rect 6177 183504 6182 183560
rect 6238 183504 6458 183560
rect 6514 183504 6519 183560
rect 6177 183502 6519 183504
rect 6177 183499 6243 183502
rect 6453 183499 6519 183502
rect 3969 181522 4035 181525
rect 7054 181522 7114 182104
rect 583520 181780 584960 182020
rect 3969 181520 7114 181522
rect 3969 181464 3974 181520
rect 4030 181464 7114 181520
rect 3969 181462 7114 181464
rect 3969 181459 4035 181462
rect -960 179332 480 179572
rect 583520 169948 584960 170188
rect 578141 166970 578207 166973
rect 576902 166968 578207 166970
rect 576902 166912 578146 166968
rect 578202 166912 578207 166968
rect 576902 166910 578207 166912
rect 576902 166328 576962 166910
rect 578141 166907 578207 166910
rect -960 165066 480 165156
rect 3233 165066 3299 165069
rect -960 165064 3299 165066
rect -960 165008 3238 165064
rect 3294 165008 3299 165064
rect -960 165006 3299 165008
rect -960 164916 480 165006
rect 3233 165003 3299 165006
rect 6085 164250 6151 164253
rect 6269 164250 6335 164253
rect 6085 164248 6335 164250
rect 6085 164192 6090 164248
rect 6146 164192 6274 164248
rect 6330 164192 6335 164248
rect 6085 164190 6335 164192
rect 6085 164187 6151 164190
rect 6269 164187 6335 164190
rect 3325 160850 3391 160853
rect 7054 160850 7114 161432
rect 3325 160848 7114 160850
rect 3325 160792 3330 160848
rect 3386 160792 7114 160848
rect 3325 160790 7114 160792
rect 3325 160787 3391 160790
rect 580717 158402 580783 158405
rect 583520 158402 584960 158492
rect 580717 158400 584960 158402
rect 580717 158344 580722 158400
rect 580778 158344 584960 158400
rect 580717 158342 584960 158344
rect 580717 158339 580783 158342
rect 583520 158252 584960 158342
rect -960 150636 480 150876
rect 583520 146556 584960 146796
rect 578141 145754 578207 145757
rect 576902 145752 578207 145754
rect 576902 145696 578146 145752
rect 578202 145696 578207 145752
rect 576902 145694 578207 145696
rect 576902 145112 576962 145694
rect 578141 145691 578207 145694
rect 5901 144938 5967 144941
rect 6085 144938 6151 144941
rect 5901 144936 6151 144938
rect 5901 144880 5906 144936
rect 5962 144880 6090 144936
rect 6146 144880 6151 144936
rect 5901 144878 6151 144880
rect 5901 144875 5967 144878
rect 6085 144875 6151 144878
rect 3233 141538 3299 141541
rect 3233 141536 7114 141538
rect 3233 141480 3238 141536
rect 3294 141480 7114 141536
rect 3233 141478 7114 141480
rect 3233 141475 3299 141478
rect 7054 140896 7114 141478
rect -960 136220 480 136460
rect 583520 134724 584960 134964
rect 5901 125626 5967 125629
rect 6085 125626 6151 125629
rect 5901 125624 6151 125626
rect 5901 125568 5906 125624
rect 5962 125568 6090 125624
rect 6146 125568 6151 125624
rect 5901 125566 6151 125568
rect 5901 125563 5967 125566
rect 6085 125563 6151 125566
rect 580165 124130 580231 124133
rect 576902 124128 580231 124130
rect 576902 124072 580170 124128
rect 580226 124072 580231 124128
rect 576902 124070 580231 124072
rect 576902 123896 576962 124070
rect 580165 124067 580231 124070
rect 583520 123028 584960 123268
rect -960 122090 480 122180
rect 3325 122090 3391 122093
rect -960 122088 3391 122090
rect -960 122032 3330 122088
rect 3386 122032 3391 122088
rect -960 122030 3391 122032
rect -960 121940 480 122030
rect 3325 122027 3391 122030
rect 4061 120866 4127 120869
rect 4061 120864 7114 120866
rect 4061 120808 4066 120864
rect 4122 120808 7114 120864
rect 4061 120806 7114 120808
rect 4061 120803 4127 120806
rect 7054 120224 7114 120806
rect 580809 111482 580875 111485
rect 583520 111482 584960 111572
rect 580809 111480 584960 111482
rect 580809 111424 580814 111480
rect 580870 111424 584960 111480
rect 580809 111422 584960 111424
rect 580809 111419 580875 111422
rect 583520 111332 584960 111422
rect -960 107524 480 107764
rect 578141 103186 578207 103189
rect 576902 103184 578207 103186
rect 576902 103128 578146 103184
rect 578202 103128 578207 103184
rect 576902 103126 578207 103128
rect 576902 102680 576962 103126
rect 578141 103123 578207 103126
rect 3877 100330 3943 100333
rect 3877 100328 7114 100330
rect 3877 100272 3882 100328
rect 3938 100272 7114 100328
rect 3877 100270 7114 100272
rect 3877 100267 3943 100270
rect 7054 99688 7114 100270
rect 583520 99636 584960 99876
rect -960 93108 480 93348
rect 583520 87804 584960 88044
rect 578141 81426 578207 81429
rect 576902 81424 578207 81426
rect 576902 81368 578146 81424
rect 578202 81368 578207 81424
rect 576902 81366 578207 81368
rect 576902 81328 576962 81366
rect 578141 81363 578207 81366
rect 3693 79658 3759 79661
rect 3693 79656 7114 79658
rect 3693 79600 3698 79656
rect 3754 79600 7114 79656
rect 3693 79598 7114 79600
rect 3693 79595 3759 79598
rect -960 78978 480 79068
rect 7054 79016 7114 79598
rect 3969 78978 4035 78981
rect -960 78976 4035 78978
rect -960 78920 3974 78976
rect 4030 78920 4035 78976
rect -960 78918 4035 78920
rect -960 78828 480 78918
rect 3969 78915 4035 78918
rect 583520 76108 584960 76348
rect -960 64412 480 64652
rect 580625 64562 580691 64565
rect 583520 64562 584960 64652
rect 580625 64560 584960 64562
rect 580625 64504 580630 64560
rect 580686 64504 584960 64560
rect 580625 64502 584960 64504
rect 580625 64499 580691 64502
rect 583520 64412 584960 64502
rect 578141 60618 578207 60621
rect 576902 60616 578207 60618
rect 576902 60560 578146 60616
rect 578202 60560 578207 60616
rect 576902 60558 578207 60560
rect 576902 60112 576962 60558
rect 578141 60555 578207 60558
rect 3601 59122 3667 59125
rect 3601 59120 7114 59122
rect 3601 59064 3606 59120
rect 3662 59064 7114 59120
rect 3601 59062 7114 59064
rect 3601 59059 3667 59062
rect 7054 58480 7114 59062
rect 583520 52716 584960 52956
rect -960 49996 480 50236
rect 583520 40884 584960 41124
rect 578141 39538 578207 39541
rect 576902 39536 578207 39538
rect 576902 39480 578146 39536
rect 578202 39480 578207 39536
rect 576902 39478 578207 39480
rect 576902 38896 576962 39478
rect 578141 39475 578207 39478
rect 3509 38314 3575 38317
rect 3509 38312 7114 38314
rect 3509 38256 3514 38312
rect 3570 38256 7114 38312
rect 3509 38254 7114 38256
rect 3509 38251 3575 38254
rect 7054 37808 7114 38254
rect -960 35866 480 35956
rect 3785 35866 3851 35869
rect -960 35864 3851 35866
rect -960 35808 3790 35864
rect 3846 35808 3851 35864
rect -960 35806 3851 35808
rect -960 35716 480 35806
rect 3785 35803 3851 35806
rect 583520 29188 584960 29428
rect -960 21300 480 21540
rect 3417 17914 3483 17917
rect 3417 17912 7114 17914
rect 3417 17856 3422 17912
rect 3478 17856 7114 17912
rect 3417 17854 7114 17856
rect 3417 17851 3483 17854
rect 7054 17272 7114 17854
rect 576902 17642 576962 17680
rect 583520 17642 584960 17732
rect 576902 17582 584960 17642
rect 583520 17492 584960 17582
rect 77845 7578 77911 7581
rect 569718 7578 569724 7580
rect 77845 7576 569724 7578
rect 77845 7520 77850 7576
rect 77906 7520 569724 7576
rect 77845 7518 569724 7520
rect 77845 7515 77911 7518
rect 569718 7516 569724 7518
rect 569788 7516 569794 7580
rect -960 7020 480 7260
rect 102777 6762 102843 6765
rect 578366 6762 578372 6764
rect 102777 6760 578372 6762
rect 102777 6704 102782 6760
rect 102838 6704 578372 6760
rect 102777 6702 578372 6704
rect 102777 6699 102843 6702
rect 578366 6700 578372 6702
rect 578436 6700 578442 6764
rect 84929 6626 84995 6629
rect 578550 6626 578556 6628
rect 84929 6624 578556 6626
rect 84929 6568 84934 6624
rect 84990 6568 578556 6624
rect 84929 6566 578556 6568
rect 84929 6563 84995 6566
rect 578550 6564 578556 6566
rect 578620 6564 578626 6628
rect 81433 6490 81499 6493
rect 578734 6490 578740 6492
rect 81433 6488 578740 6490
rect 81433 6432 81438 6488
rect 81494 6432 578740 6488
rect 81433 6430 578740 6432
rect 81433 6427 81499 6430
rect 578734 6428 578740 6430
rect 578804 6428 578810 6492
rect 74257 6354 74323 6357
rect 578918 6354 578924 6356
rect 74257 6352 578924 6354
rect 74257 6296 74262 6352
rect 74318 6296 578924 6352
rect 74257 6294 578924 6296
rect 74257 6291 74323 6294
rect 578918 6292 578924 6294
rect 578988 6292 578994 6356
rect 63585 6218 63651 6221
rect 579102 6218 579108 6220
rect 63585 6216 579108 6218
rect 63585 6160 63590 6216
rect 63646 6160 579108 6216
rect 63585 6158 579108 6160
rect 63585 6155 63651 6158
rect 579102 6156 579108 6158
rect 579172 6156 579178 6220
rect 583520 5796 584960 6036
rect 31477 5538 31543 5541
rect 465809 5538 465875 5541
rect 31477 5536 465875 5538
rect 31477 5480 31482 5536
rect 31538 5480 465814 5536
rect 465870 5480 465875 5536
rect 31477 5478 465875 5480
rect 31477 5475 31543 5478
rect 465809 5475 465875 5478
rect 38561 5402 38627 5405
rect 475469 5402 475535 5405
rect 38561 5400 475535 5402
rect 38561 5344 38566 5400
rect 38622 5344 475474 5400
rect 475530 5344 475535 5400
rect 38561 5342 475535 5344
rect 38561 5339 38627 5342
rect 475469 5339 475535 5342
rect 67173 5266 67239 5269
rect 504449 5266 504515 5269
rect 67173 5264 504515 5266
rect 67173 5208 67178 5264
rect 67234 5208 504454 5264
rect 504510 5208 504515 5264
rect 67173 5206 504515 5208
rect 67173 5203 67239 5206
rect 504449 5203 504515 5206
rect 42149 5130 42215 5133
rect 485129 5130 485195 5133
rect 42149 5128 485195 5130
rect 42149 5072 42154 5128
rect 42210 5072 485134 5128
rect 485190 5072 485195 5128
rect 42149 5070 485195 5072
rect 42149 5067 42215 5070
rect 485129 5067 485195 5070
rect 8845 4994 8911 4997
rect 456149 4994 456215 4997
rect 8845 4992 456215 4994
rect 8845 4936 8850 4992
rect 8906 4936 456154 4992
rect 456210 4936 456215 4992
rect 8845 4934 456215 4936
rect 8845 4931 8911 4934
rect 456149 4931 456215 4934
rect 25497 4858 25563 4861
rect 562409 4858 562475 4861
rect 25497 4856 562475 4858
rect 25497 4800 25502 4856
rect 25558 4800 562414 4856
rect 562470 4800 562475 4856
rect 25497 4798 562475 4800
rect 25497 4795 25563 4798
rect 562409 4795 562475 4798
rect 5022 4660 5028 4724
rect 5092 4722 5098 4724
rect 106365 4722 106431 4725
rect 5092 4720 106431 4722
rect 5092 4664 106370 4720
rect 106426 4664 106431 4720
rect 5092 4662 106431 4664
rect 5092 4660 5098 4662
rect 106365 4659 106431 4662
rect 5390 3980 5396 4044
rect 5460 4042 5466 4044
rect 113541 4042 113607 4045
rect 5460 4040 113607 4042
rect 5460 3984 113546 4040
rect 113602 3984 113607 4040
rect 5460 3982 113607 3984
rect 5460 3980 5466 3982
rect 113541 3979 113607 3982
rect 123017 4042 123083 4045
rect 578325 4042 578391 4045
rect 123017 4040 578391 4042
rect 123017 3984 123022 4040
rect 123078 3984 578330 4040
rect 578386 3984 578391 4040
rect 123017 3982 578391 3984
rect 123017 3979 123083 3982
rect 578325 3979 578391 3982
rect 34973 3906 35039 3909
rect 579286 3906 579292 3908
rect 34973 3904 579292 3906
rect 34973 3848 34978 3904
rect 35034 3848 579292 3904
rect 34973 3846 579292 3848
rect 34973 3843 35039 3846
rect 579286 3844 579292 3846
rect 579356 3844 579362 3908
rect 33869 3770 33935 3773
rect 579245 3770 579311 3773
rect 33869 3768 579311 3770
rect 33869 3712 33874 3768
rect 33930 3712 579250 3768
rect 579306 3712 579311 3768
rect 33869 3710 579311 3712
rect 33869 3707 33935 3710
rect 579245 3707 579311 3710
rect 27889 3634 27955 3637
rect 578233 3634 578299 3637
rect 27889 3632 578299 3634
rect 27889 3576 27894 3632
rect 27950 3576 578238 3632
rect 578294 3576 578299 3632
rect 27889 3574 578299 3576
rect 27889 3571 27955 3574
rect 578233 3571 578299 3574
rect 17217 3498 17283 3501
rect 579337 3498 579403 3501
rect 17217 3496 579403 3498
rect 17217 3440 17222 3496
rect 17278 3440 579342 3496
rect 579398 3440 579403 3496
rect 17217 3438 579403 3440
rect 17217 3435 17283 3438
rect 579337 3435 579403 3438
rect 16021 3362 16087 3365
rect 578182 3362 578188 3364
rect 16021 3360 578188 3362
rect 16021 3304 16026 3360
rect 16082 3304 578188 3360
rect 16021 3302 578188 3304
rect 16021 3299 16087 3302
rect 578182 3300 578188 3302
rect 578252 3300 578258 3364
rect 5206 3164 5212 3228
rect 5276 3226 5282 3228
rect 109953 3226 110019 3229
rect 5276 3224 110019 3226
rect 5276 3168 109958 3224
rect 110014 3168 110019 3224
rect 5276 3166 110019 3168
rect 5276 3164 5282 3166
rect 109953 3163 110019 3166
<< via3 >>
rect 569724 688604 569788 688668
rect 391428 686352 391492 686356
rect 391428 686296 391478 686352
rect 391478 686296 391492 686352
rect 391428 686292 391492 686296
rect 419948 686352 420012 686356
rect 419948 686296 419998 686352
rect 419998 686296 420012 686352
rect 419948 686292 420012 686296
rect 391428 685204 391492 685268
rect 419948 685068 420012 685132
rect 578188 676228 578252 676292
rect 578372 654604 578436 654668
rect 5396 634884 5460 634948
rect 578556 633388 578620 633452
rect 5212 614076 5276 614140
rect 578740 612036 578804 612100
rect 5028 593540 5092 593604
rect 578924 590684 578988 590748
rect 579108 570012 579172 570076
rect 579292 548388 579356 548452
rect 569724 7516 569788 7580
rect 578372 6700 578436 6764
rect 578556 6564 578620 6628
rect 578740 6428 578804 6492
rect 578924 6292 578988 6356
rect 579108 6156 579172 6220
rect 5028 4660 5092 4724
rect 5396 3980 5460 4044
rect 579292 3844 579356 3908
rect 578188 3300 578252 3364
rect 5212 3164 5276 3228
<< metal4 >>
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 -3166 -4216 707102
rect 23424 707658 24024 707680
rect 23424 707422 23606 707658
rect 23842 707422 24024 707658
rect 23424 707338 24024 707422
rect 23424 707102 23606 707338
rect 23842 707102 24024 707338
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 -2226 -3276 706162
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 -1286 -2336 705222
rect 23424 705778 24024 707102
rect 23424 705542 23606 705778
rect 23842 705542 24024 705778
rect 23424 705458 24024 705542
rect 23424 705222 23606 705458
rect 23842 705222 24024 705458
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 -346 -1396 704282
rect 5395 634948 5461 634949
rect 5395 634884 5396 634948
rect 5460 634884 5461 634948
rect 5395 634883 5461 634884
rect 5211 614140 5277 614141
rect 5211 614076 5212 614140
rect 5276 614076 5277 614140
rect 5211 614075 5277 614076
rect 5027 593604 5093 593605
rect 5027 593540 5028 593604
rect 5092 593540 5093 593604
rect 5027 593539 5093 593540
rect 5030 4725 5090 593539
rect 5027 4724 5093 4725
rect 5027 4660 5028 4724
rect 5092 4660 5093 4724
rect 5027 4659 5093 4660
rect 5214 3229 5274 614075
rect 5398 4045 5458 634883
rect 5395 4044 5461 4045
rect 5395 3980 5396 4044
rect 5460 3980 5461 4044
rect 5395 3979 5461 3980
rect 5211 3228 5277 3229
rect 5211 3164 5212 3228
rect 5276 3164 5277 3228
rect 5211 3163 5277 3164
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 23424 -1286 24024 705222
rect 23424 -1522 23606 -1286
rect 23842 -1522 24024 -1286
rect 23424 -1606 24024 -1522
rect 23424 -1842 23606 -1606
rect 23842 -1842 24024 -1606
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 23424 -3166 24024 -1842
rect 23424 -3402 23606 -3166
rect 23842 -3402 24024 -3166
rect 23424 -3486 24024 -3402
rect 23424 -3722 23606 -3486
rect 23842 -3722 24024 -3486
rect 23424 -3744 24024 -3722
rect 99424 706718 100024 707680
rect 99424 706482 99606 706718
rect 99842 706482 100024 706718
rect 99424 706398 100024 706482
rect 99424 706162 99606 706398
rect 99842 706162 100024 706398
rect 99424 704838 100024 706162
rect 99424 704602 99606 704838
rect 99842 704602 100024 704838
rect 99424 704518 100024 704602
rect 99424 704282 99606 704518
rect 99842 704282 100024 704518
rect 99424 -346 100024 704282
rect 99424 -582 99606 -346
rect 99842 -582 100024 -346
rect 99424 -666 100024 -582
rect 99424 -902 99606 -666
rect 99842 -902 100024 -666
rect 99424 -2226 100024 -902
rect 99424 -2462 99606 -2226
rect 99842 -2462 100024 -2226
rect 99424 -2546 100024 -2462
rect 99424 -2782 99606 -2546
rect 99842 -2782 100024 -2546
rect 99424 -3744 100024 -2782
rect 175424 707658 176024 707680
rect 175424 707422 175606 707658
rect 175842 707422 176024 707658
rect 175424 707338 176024 707422
rect 175424 707102 175606 707338
rect 175842 707102 176024 707338
rect 175424 705778 176024 707102
rect 175424 705542 175606 705778
rect 175842 705542 176024 705778
rect 175424 705458 176024 705542
rect 175424 705222 175606 705458
rect 175842 705222 176024 705458
rect 175424 -1286 176024 705222
rect 175424 -1522 175606 -1286
rect 175842 -1522 176024 -1286
rect 175424 -1606 176024 -1522
rect 175424 -1842 175606 -1606
rect 175842 -1842 176024 -1606
rect 175424 -3166 176024 -1842
rect 175424 -3402 175606 -3166
rect 175842 -3402 176024 -3166
rect 175424 -3486 176024 -3402
rect 175424 -3722 175606 -3486
rect 175842 -3722 176024 -3486
rect 175424 -3744 176024 -3722
rect 251424 706718 252024 707680
rect 251424 706482 251606 706718
rect 251842 706482 252024 706718
rect 251424 706398 252024 706482
rect 251424 706162 251606 706398
rect 251842 706162 252024 706398
rect 251424 704838 252024 706162
rect 251424 704602 251606 704838
rect 251842 704602 252024 704838
rect 251424 704518 252024 704602
rect 251424 704282 251606 704518
rect 251842 704282 252024 704518
rect 251424 -346 252024 704282
rect 251424 -582 251606 -346
rect 251842 -582 252024 -346
rect 251424 -666 252024 -582
rect 251424 -902 251606 -666
rect 251842 -902 252024 -666
rect 251424 -2226 252024 -902
rect 251424 -2462 251606 -2226
rect 251842 -2462 252024 -2226
rect 251424 -2546 252024 -2462
rect 251424 -2782 251606 -2546
rect 251842 -2782 252024 -2546
rect 251424 -3744 252024 -2782
rect 327424 707658 328024 707680
rect 327424 707422 327606 707658
rect 327842 707422 328024 707658
rect 327424 707338 328024 707422
rect 327424 707102 327606 707338
rect 327842 707102 328024 707338
rect 327424 705778 328024 707102
rect 327424 705542 327606 705778
rect 327842 705542 328024 705778
rect 327424 705458 328024 705542
rect 327424 705222 327606 705458
rect 327842 705222 328024 705458
rect 327424 -1286 328024 705222
rect 403424 706718 404024 707680
rect 403424 706482 403606 706718
rect 403842 706482 404024 706718
rect 403424 706398 404024 706482
rect 403424 706162 403606 706398
rect 403842 706162 404024 706398
rect 403424 704838 404024 706162
rect 403424 704602 403606 704838
rect 403842 704602 404024 704838
rect 403424 704518 404024 704602
rect 403424 704282 403606 704518
rect 403842 704282 404024 704518
rect 391427 686356 391493 686357
rect 391427 686292 391428 686356
rect 391492 686292 391493 686356
rect 391427 686291 391493 686292
rect 391430 685269 391490 686291
rect 391427 685268 391493 685269
rect 391427 685204 391428 685268
rect 391492 685204 391493 685268
rect 391427 685203 391493 685204
rect 327424 -1522 327606 -1286
rect 327842 -1522 328024 -1286
rect 327424 -1606 328024 -1522
rect 327424 -1842 327606 -1606
rect 327842 -1842 328024 -1606
rect 327424 -3166 328024 -1842
rect 327424 -3402 327606 -3166
rect 327842 -3402 328024 -3166
rect 327424 -3486 328024 -3402
rect 327424 -3722 327606 -3486
rect 327842 -3722 328024 -3486
rect 327424 -3744 328024 -3722
rect 403424 -346 404024 704282
rect 479424 707658 480024 707680
rect 479424 707422 479606 707658
rect 479842 707422 480024 707658
rect 479424 707338 480024 707422
rect 479424 707102 479606 707338
rect 479842 707102 480024 707338
rect 479424 705778 480024 707102
rect 479424 705542 479606 705778
rect 479842 705542 480024 705778
rect 479424 705458 480024 705542
rect 479424 705222 479606 705458
rect 479842 705222 480024 705458
rect 419947 686356 420013 686357
rect 419947 686292 419948 686356
rect 420012 686292 420013 686356
rect 419947 686291 420013 686292
rect 419950 685133 420010 686291
rect 419947 685132 420013 685133
rect 419947 685068 419948 685132
rect 420012 685068 420013 685132
rect 419947 685067 420013 685068
rect 403424 -582 403606 -346
rect 403842 -582 404024 -346
rect 403424 -666 404024 -582
rect 403424 -902 403606 -666
rect 403842 -902 404024 -666
rect 403424 -2226 404024 -902
rect 403424 -2462 403606 -2226
rect 403842 -2462 404024 -2226
rect 403424 -2546 404024 -2462
rect 403424 -2782 403606 -2546
rect 403842 -2782 404024 -2546
rect 403424 -3744 404024 -2782
rect 479424 -1286 480024 705222
rect 479424 -1522 479606 -1286
rect 479842 -1522 480024 -1286
rect 479424 -1606 480024 -1522
rect 479424 -1842 479606 -1606
rect 479842 -1842 480024 -1606
rect 479424 -3166 480024 -1842
rect 479424 -3402 479606 -3166
rect 479842 -3402 480024 -3166
rect 479424 -3486 480024 -3402
rect 479424 -3722 479606 -3486
rect 479842 -3722 480024 -3486
rect 479424 -3744 480024 -3722
rect 555424 706718 556024 707680
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect 555424 706482 555606 706718
rect 555842 706482 556024 706718
rect 555424 706398 556024 706482
rect 555424 706162 555606 706398
rect 555842 706162 556024 706398
rect 555424 704838 556024 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 555424 704602 555606 704838
rect 555842 704602 556024 704838
rect 555424 704518 556024 704602
rect 555424 704282 555606 704518
rect 555842 704282 556024 704518
rect 555424 -346 556024 704282
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 569723 688668 569789 688669
rect 569723 688604 569724 688668
rect 569788 688604 569789 688668
rect 569723 688603 569789 688604
rect 569726 685810 569786 688603
rect 569726 685750 570154 685810
rect 570094 685130 570154 685750
rect 570094 685070 570338 685130
rect 570278 675610 570338 685070
rect 578187 676292 578253 676293
rect 578187 676228 578188 676292
rect 578252 676228 578253 676292
rect 578187 676227 578253 676228
rect 570278 675550 570522 675610
rect 570462 674250 570522 675550
rect 570462 674190 570706 674250
rect 570646 659290 570706 674190
rect 570462 659230 570706 659290
rect 570462 649090 570522 659230
rect 570094 649030 570522 649090
rect 570094 642290 570154 649030
rect 570094 642230 570338 642290
rect 570278 637530 570338 642230
rect 570278 637470 570522 637530
rect 570462 628010 570522 637470
rect 570462 627950 570706 628010
rect 570646 621210 570706 627950
rect 570462 621150 570706 621210
rect 570462 611690 570522 621150
rect 570278 611630 570522 611690
rect 570278 601490 570338 611630
rect 570278 601430 570522 601490
rect 570462 591970 570522 601430
rect 570094 591910 570522 591970
rect 570094 589250 570154 591910
rect 570094 589190 571074 589250
rect 571014 581770 571074 589190
rect 569910 581710 571074 581770
rect 569910 579050 569970 581710
rect 569910 578990 570338 579050
rect 570278 572930 570338 578990
rect 569910 572870 570338 572930
rect 569910 570074 569970 572870
rect 569910 570014 570338 570074
rect 570278 562730 570338 570014
rect 570094 562670 570338 562730
rect 570094 553210 570154 562670
rect 570094 553150 570338 553210
rect 570278 543010 570338 553150
rect 569910 542950 570338 543010
rect 569910 540970 569970 542950
rect 569910 540910 571074 540970
rect 571014 531450 571074 540910
rect 570278 531390 571074 531450
rect 570278 524650 570338 531390
rect 570094 524590 570338 524650
rect 570094 521250 570154 524590
rect 570094 521190 570338 521250
rect 570278 519890 570338 521190
rect 570278 519830 571258 519890
rect 571198 512410 571258 519830
rect 570278 512350 571258 512410
rect 570278 504250 570338 512350
rect 569910 504190 570338 504250
rect 569910 495410 569970 504190
rect 569910 495350 570154 495410
rect 570094 492010 570154 495350
rect 570094 491950 570338 492010
rect 570278 485210 570338 491950
rect 570278 485150 570706 485210
rect 570646 475690 570706 485150
rect 570462 475630 570706 475690
rect 570462 467530 570522 475630
rect 570462 467470 571258 467530
rect 571198 466170 571258 467470
rect 570094 466110 571258 466170
rect 570094 458690 570154 466110
rect 570094 458630 570338 458690
rect 570278 432850 570338 458630
rect 570278 432790 571258 432850
rect 571198 431490 571258 432790
rect 570278 431430 571258 431490
rect 570278 426730 570338 431430
rect 569910 426670 570338 426730
rect 569910 421970 569970 426670
rect 569910 421910 571074 421970
rect 571014 413130 571074 421910
rect 570094 413070 571074 413130
rect 570094 383890 570154 413070
rect 570094 383830 570522 383890
rect 570462 381850 570522 383830
rect 570462 381790 570706 381850
rect 570646 369610 570706 381790
rect 570462 369550 570706 369610
rect 570462 360090 570522 369550
rect 570462 360030 570706 360090
rect 570646 351250 570706 360030
rect 570462 351190 570706 351250
rect 570462 347850 570522 351190
rect 570278 347790 570522 347850
rect 570278 347170 570338 347790
rect 570278 347110 570522 347170
rect 570462 345810 570522 347110
rect 570462 345750 570706 345810
rect 570646 330850 570706 345750
rect 570462 330790 570706 330850
rect 570462 320650 570522 330790
rect 570094 320590 570522 320650
rect 570094 313850 570154 320590
rect 570094 313790 570338 313850
rect 570278 309090 570338 313790
rect 570278 309030 570522 309090
rect 570462 299570 570522 309030
rect 570462 299510 570706 299570
rect 570646 292770 570706 299510
rect 570462 292710 570706 292770
rect 570462 283250 570522 292710
rect 570278 283190 570522 283250
rect 570278 275090 570338 283190
rect 570278 275030 570706 275090
rect 570646 263530 570706 275030
rect 570094 263470 570706 263530
rect 570094 260810 570154 263470
rect 570094 260750 571074 260810
rect 571014 253330 571074 260750
rect 569910 253270 571074 253330
rect 569910 250610 569970 253270
rect 569910 250550 570338 250610
rect 570278 249930 570338 250550
rect 570278 249870 571258 249930
rect 571198 241770 571258 249870
rect 570278 241710 571258 241770
rect 570278 234290 570338 241710
rect 570094 234230 570338 234290
rect 570094 224770 570154 234230
rect 570094 224710 570338 224770
rect 570278 214570 570338 224710
rect 569910 214510 570338 214570
rect 569910 212530 569970 214510
rect 569910 212470 571074 212530
rect 571014 203010 571074 212470
rect 570278 202950 571074 203010
rect 570278 196210 570338 202950
rect 570094 196150 570338 196210
rect 570094 192810 570154 196150
rect 570094 192750 571074 192810
rect 571014 185330 571074 192750
rect 570094 185270 571074 185330
rect 570094 183970 570154 185270
rect 569910 183910 570154 183970
rect 569910 176490 569970 183910
rect 569910 176430 570154 176490
rect 570094 173770 570154 176430
rect 570094 173710 570338 173770
rect 570278 166970 570338 173710
rect 570094 166910 570338 166970
rect 570094 164250 570154 166910
rect 570094 164190 570338 164250
rect 570278 156770 570338 164190
rect 569910 156710 570338 156770
rect 569910 154050 569970 156710
rect 569910 153990 570338 154050
rect 570278 153370 570338 153990
rect 570278 153310 571074 153370
rect 571014 145210 571074 153310
rect 570278 145150 571074 145210
rect 570278 137730 570338 145150
rect 570094 137670 570338 137730
rect 570094 130250 570154 137670
rect 570094 130190 570338 130250
rect 570278 104410 570338 130190
rect 570278 104350 571258 104410
rect 571198 103050 571258 104350
rect 570278 102990 571258 103050
rect 570278 98290 570338 102990
rect 569910 98230 570338 98290
rect 569910 93530 569970 98230
rect 569910 93470 571074 93530
rect 571014 84690 571074 93470
rect 570094 84630 571074 84690
rect 570094 64970 570154 84630
rect 569910 64910 570154 64970
rect 569910 59530 569970 64910
rect 569910 59470 570522 59530
rect 570462 51370 570522 59470
rect 570278 51310 570522 51370
rect 570278 37770 570338 51310
rect 570094 37710 570338 37770
rect 570094 33690 570154 37710
rect 570094 33630 570338 33690
rect 570278 22810 570338 33630
rect 570094 22750 570338 22810
rect 570094 19410 570154 22750
rect 569910 19350 570154 19410
rect 569910 17458 569970 19350
rect 569910 8530 569970 15862
rect 569726 8470 569970 8530
rect 569726 7581 569786 8470
rect 569723 7580 569789 7581
rect 569723 7516 569724 7580
rect 569788 7516 569789 7580
rect 569723 7515 569789 7516
rect 578190 3365 578250 676227
rect 578371 654668 578437 654669
rect 578371 654604 578372 654668
rect 578436 654604 578437 654668
rect 578371 654603 578437 654604
rect 578374 6765 578434 654603
rect 578555 633452 578621 633453
rect 578555 633388 578556 633452
rect 578620 633388 578621 633452
rect 578555 633387 578621 633388
rect 578371 6764 578437 6765
rect 578371 6700 578372 6764
rect 578436 6700 578437 6764
rect 578371 6699 578437 6700
rect 578558 6629 578618 633387
rect 578739 612100 578805 612101
rect 578739 612036 578740 612100
rect 578804 612036 578805 612100
rect 578739 612035 578805 612036
rect 578555 6628 578621 6629
rect 578555 6564 578556 6628
rect 578620 6564 578621 6628
rect 578555 6563 578621 6564
rect 578742 6493 578802 612035
rect 578923 590748 578989 590749
rect 578923 590684 578924 590748
rect 578988 590684 578989 590748
rect 578923 590683 578989 590684
rect 578739 6492 578805 6493
rect 578739 6428 578740 6492
rect 578804 6428 578805 6492
rect 578739 6427 578805 6428
rect 578926 6357 578986 590683
rect 579107 570076 579173 570077
rect 579107 570012 579108 570076
rect 579172 570012 579173 570076
rect 579107 570011 579173 570012
rect 578923 6356 578989 6357
rect 578923 6292 578924 6356
rect 578988 6292 578989 6356
rect 578923 6291 578989 6292
rect 579110 6221 579170 570011
rect 579291 548452 579357 548453
rect 579291 548388 579292 548452
rect 579356 548388 579357 548452
rect 579291 548387 579357 548388
rect 579107 6220 579173 6221
rect 579107 6156 579108 6220
rect 579172 6156 579173 6220
rect 579107 6155 579173 6156
rect 579294 3909 579354 548387
rect 579291 3908 579357 3909
rect 579291 3844 579292 3908
rect 579356 3844 579357 3908
rect 579291 3843 579357 3844
rect 578187 3364 578253 3365
rect 578187 3300 578188 3364
rect 578252 3300 578253 3364
rect 578187 3299 578253 3300
rect 555424 -582 555606 -346
rect 555842 -582 556024 -346
rect 555424 -666 556024 -582
rect 555424 -902 555606 -666
rect 555842 -902 556024 -666
rect 555424 -2226 556024 -902
rect 585320 -346 585920 704282
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 -1286 586860 705222
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect 555424 -2462 555606 -2226
rect 555842 -2462 556024 -2226
rect 555424 -2546 556024 -2462
rect 555424 -2782 555606 -2546
rect 555842 -2782 556024 -2546
rect 555424 -3744 556024 -2782
rect 587200 -2226 587800 706162
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect 588140 -3166 588740 707102
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
<< via4 >>
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect 23606 707422 23842 707658
rect 23606 707102 23842 707338
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect 23606 705542 23842 705778
rect 23606 705222 23842 705458
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 23606 -1522 23842 -1286
rect 23606 -1842 23842 -1606
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect 23606 -3402 23842 -3166
rect 23606 -3722 23842 -3486
rect 99606 706482 99842 706718
rect 99606 706162 99842 706398
rect 99606 704602 99842 704838
rect 99606 704282 99842 704518
rect 99606 -582 99842 -346
rect 99606 -902 99842 -666
rect 99606 -2462 99842 -2226
rect 99606 -2782 99842 -2546
rect 175606 707422 175842 707658
rect 175606 707102 175842 707338
rect 175606 705542 175842 705778
rect 175606 705222 175842 705458
rect 175606 -1522 175842 -1286
rect 175606 -1842 175842 -1606
rect 175606 -3402 175842 -3166
rect 175606 -3722 175842 -3486
rect 251606 706482 251842 706718
rect 251606 706162 251842 706398
rect 251606 704602 251842 704838
rect 251606 704282 251842 704518
rect 251606 -582 251842 -346
rect 251606 -902 251842 -666
rect 251606 -2462 251842 -2226
rect 251606 -2782 251842 -2546
rect 327606 707422 327842 707658
rect 327606 707102 327842 707338
rect 327606 705542 327842 705778
rect 327606 705222 327842 705458
rect 403606 706482 403842 706718
rect 403606 706162 403842 706398
rect 403606 704602 403842 704838
rect 403606 704282 403842 704518
rect 327606 -1522 327842 -1286
rect 327606 -1842 327842 -1606
rect 327606 -3402 327842 -3166
rect 327606 -3722 327842 -3486
rect 479606 707422 479842 707658
rect 479606 707102 479842 707338
rect 479606 705542 479842 705778
rect 479606 705222 479842 705458
rect 403606 -582 403842 -346
rect 403606 -902 403842 -666
rect 403606 -2462 403842 -2226
rect 403606 -2782 403842 -2546
rect 479606 -1522 479842 -1286
rect 479606 -1842 479842 -1606
rect 479606 -3402 479842 -3166
rect 479606 -3722 479842 -3486
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect 555606 706482 555842 706718
rect 555606 706162 555842 706398
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 555606 704602 555842 704838
rect 555606 704282 555842 704518
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 569822 17222 570058 17458
rect 569822 15862 570058 16098
rect 555606 -582 555842 -346
rect 555606 -902 555842 -666
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect 555606 -2462 555842 -2226
rect 555606 -2782 555842 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
<< metal5 >>
rect -4816 707680 -4216 707682
rect 23424 707680 24024 707682
rect 175424 707680 176024 707682
rect 327424 707680 328024 707682
rect 479424 707680 480024 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 23606 707658
rect 23842 707422 175606 707658
rect 175842 707422 327606 707658
rect 327842 707422 479606 707658
rect 479842 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 23606 707338
rect 23842 707102 175606 707338
rect 175842 707102 327606 707338
rect 327842 707102 479606 707338
rect 479842 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 23424 707078 24024 707080
rect 175424 707078 176024 707080
rect 327424 707078 328024 707080
rect 479424 707078 480024 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 99424 706740 100024 706742
rect 251424 706740 252024 706742
rect 403424 706740 404024 706742
rect 555424 706740 556024 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 99606 706718
rect 99842 706482 251606 706718
rect 251842 706482 403606 706718
rect 403842 706482 555606 706718
rect 555842 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 99606 706398
rect 99842 706162 251606 706398
rect 251842 706162 403606 706398
rect 403842 706162 555606 706398
rect 555842 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 99424 706138 100024 706140
rect 251424 706138 252024 706140
rect 403424 706138 404024 706140
rect 555424 706138 556024 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 23424 705800 24024 705802
rect 175424 705800 176024 705802
rect 327424 705800 328024 705802
rect 479424 705800 480024 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 23606 705778
rect 23842 705542 175606 705778
rect 175842 705542 327606 705778
rect 327842 705542 479606 705778
rect 479842 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 23606 705458
rect 23842 705222 175606 705458
rect 175842 705222 327606 705458
rect 327842 705222 479606 705458
rect 479842 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 23424 705198 24024 705200
rect 175424 705198 176024 705200
rect 327424 705198 328024 705200
rect 479424 705198 480024 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 99424 704860 100024 704862
rect 251424 704860 252024 704862
rect 403424 704860 404024 704862
rect 555424 704860 556024 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 99606 704838
rect 99842 704602 251606 704838
rect 251842 704602 403606 704838
rect 403842 704602 555606 704838
rect 555842 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 99606 704518
rect 99842 704282 251606 704518
rect 251842 704282 403606 704518
rect 403842 704282 555606 704518
rect 555842 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 99424 704258 100024 704260
rect 251424 704258 252024 704260
rect 403424 704258 404024 704260
rect 555424 704258 556024 704260
rect 585320 704258 585920 704260
rect 568492 17458 570100 17500
rect 568492 17222 569822 17458
rect 570058 17222 570100 17458
rect 568492 17180 570100 17222
rect 568492 16140 568812 17180
rect 568492 16098 570100 16140
rect 568492 15862 569822 16098
rect 570058 15862 570100 16098
rect 568492 15820 570100 15862
rect -1996 -324 -1396 -322
rect 99424 -324 100024 -322
rect 251424 -324 252024 -322
rect 403424 -324 404024 -322
rect 555424 -324 556024 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 99606 -346
rect 99842 -582 251606 -346
rect 251842 -582 403606 -346
rect 403842 -582 555606 -346
rect 555842 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 99606 -666
rect 99842 -902 251606 -666
rect 251842 -902 403606 -666
rect 403842 -902 555606 -666
rect 555842 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 99424 -926 100024 -924
rect 251424 -926 252024 -924
rect 403424 -926 404024 -924
rect 555424 -926 556024 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 23424 -1264 24024 -1262
rect 175424 -1264 176024 -1262
rect 327424 -1264 328024 -1262
rect 479424 -1264 480024 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 23606 -1286
rect 23842 -1522 175606 -1286
rect 175842 -1522 327606 -1286
rect 327842 -1522 479606 -1286
rect 479842 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 23606 -1606
rect 23842 -1842 175606 -1606
rect 175842 -1842 327606 -1606
rect 327842 -1842 479606 -1606
rect 479842 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 23424 -1866 24024 -1864
rect 175424 -1866 176024 -1864
rect 327424 -1866 328024 -1864
rect 479424 -1866 480024 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 99424 -2204 100024 -2202
rect 251424 -2204 252024 -2202
rect 403424 -2204 404024 -2202
rect 555424 -2204 556024 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 99606 -2226
rect 99842 -2462 251606 -2226
rect 251842 -2462 403606 -2226
rect 403842 -2462 555606 -2226
rect 555842 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 99606 -2546
rect 99842 -2782 251606 -2546
rect 251842 -2782 403606 -2546
rect 403842 -2782 555606 -2546
rect 555842 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 99424 -2806 100024 -2804
rect 251424 -2806 252024 -2804
rect 403424 -2806 404024 -2804
rect 555424 -2806 556024 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 23424 -3144 24024 -3142
rect 175424 -3144 176024 -3142
rect 327424 -3144 328024 -3142
rect 479424 -3144 480024 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 23606 -3166
rect 23842 -3402 175606 -3166
rect 175842 -3402 327606 -3166
rect 327842 -3402 479606 -3166
rect 479842 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 23606 -3486
rect 23842 -3722 175606 -3486
rect 175842 -3722 327606 -3486
rect 327842 -3722 479606 -3486
rect 479842 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 23424 -3746 24024 -3744
rect 175424 -3746 176024 -3744
rect 327424 -3746 328024 -3744
rect 479424 -3746 480024 -3744
rect 588140 -3746 588740 -3744
use fpga  fpga250
timestamp 1608086250
transform 1 0 7000 0 1 7000
box 0 0 570000 680000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 637 nsew default input
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 638 nsew default input
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 639 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1608015108
<< locali >>
rect 576041 634831 576075 647785
rect 6653 618307 6687 621061
rect 6561 608651 6595 618137
rect 576041 597567 576075 602361
rect 6745 572407 6779 572849
rect 575949 554795 575983 564349
rect 575949 518007 575983 522257
rect 575949 509507 575983 514709
rect 575949 485503 575983 492609
rect 576041 485639 576075 487781
rect 576133 417843 576167 428485
rect 576041 396083 576075 405569
rect 575949 379423 575983 390065
rect 576041 379627 576075 384353
rect 576041 366503 576075 371909
rect 576133 365891 576167 376669
rect 575949 359363 575983 361233
rect 576041 359023 576075 359465
rect 575949 347463 575983 352665
rect 575949 328015 575983 334577
rect 576041 331891 576075 338045
rect 575949 319107 575983 321929
rect 576041 316047 576075 319209
rect 575949 316013 576075 316047
rect 575949 315775 575983 316013
rect 576041 306391 576075 315945
rect 576133 315639 576167 319481
rect 575949 278783 575983 299149
rect 575949 262735 575983 272969
rect 576041 270351 576075 272289
rect 575949 249135 575983 257601
rect 576041 243151 576075 257465
rect 576225 225063 576259 236793
rect 576133 224927 576167 225029
rect 575949 212619 575983 220949
rect 576041 216019 576075 217481
rect 576133 215543 576167 217617
rect 575949 192559 575983 198849
rect 576041 197455 576075 203065
rect 576133 201535 576167 212449
rect 576317 198747 576351 199257
rect 576041 191131 576075 192729
rect 575949 173995 575983 182937
rect 576041 174811 576075 186881
rect 576225 186303 576259 191777
rect 575949 160803 575983 170697
rect 576041 157879 576075 170221
rect 576133 164951 576167 175661
rect 576225 172567 576259 177225
rect 575949 150467 575983 153425
rect 576133 153255 576167 157981
rect 575949 144415 575983 149345
rect 575949 132583 575983 140913
rect 576041 140335 576075 145265
rect 576133 137207 576167 149685
rect 576225 144891 576259 145945
rect 575949 118575 575983 132073
rect 576133 125579 576167 127653
rect 575949 104431 575983 118405
rect 576041 117759 576075 122553
rect 576225 120751 576259 130509
rect 576317 118439 576351 125545
rect 576041 104295 576075 113985
rect 576133 110959 576167 115821
rect 576133 102459 576167 108817
rect 576133 81379 576167 90593
rect 575949 72199 575983 81345
rect 576041 74783 576075 79441
rect 576225 70363 576259 93789
rect 575949 57851 575983 63325
rect 576041 57987 576075 67541
rect 576041 57953 576167 57987
rect 576133 57307 576167 57953
rect 575949 57273 576167 57307
rect 576317 57307 576351 58769
rect 575949 43503 575983 57273
rect 576041 39423 576075 51765
rect 575949 20315 575983 37213
rect 576041 33847 576075 35309
rect 576133 35207 576167 43605
rect 576041 28339 576075 33065
rect 576041 19363 576075 24157
rect 576133 16711 576167 21505
rect 69489 7531 69523 7769
rect 6929 2907 6963 4029
rect 8861 3791 8895 3825
rect 8861 3757 9045 3791
rect 9229 3723 9263 4029
rect 16497 2907 16531 3961
<< viali >>
rect 576041 647785 576075 647819
rect 576041 634797 576075 634831
rect 6653 621061 6687 621095
rect 6653 618273 6687 618307
rect 6561 618137 6595 618171
rect 6561 608617 6595 608651
rect 576041 602361 576075 602395
rect 576041 597533 576075 597567
rect 6745 572849 6779 572883
rect 6745 572373 6779 572407
rect 575949 564349 575983 564383
rect 575949 554761 575983 554795
rect 575949 522257 575983 522291
rect 575949 517973 575983 518007
rect 575949 514709 575983 514743
rect 575949 509473 575983 509507
rect 575949 492609 575983 492643
rect 576041 487781 576075 487815
rect 576041 485605 576075 485639
rect 575949 485469 575983 485503
rect 576133 428485 576167 428519
rect 576133 417809 576167 417843
rect 576041 405569 576075 405603
rect 576041 396049 576075 396083
rect 575949 390065 575983 390099
rect 576041 384353 576075 384387
rect 576041 379593 576075 379627
rect 575949 379389 575983 379423
rect 576133 376669 576167 376703
rect 576041 371909 576075 371943
rect 576041 366469 576075 366503
rect 576133 365857 576167 365891
rect 575949 361233 575983 361267
rect 575949 359329 575983 359363
rect 576041 359465 576075 359499
rect 576041 358989 576075 359023
rect 575949 352665 575983 352699
rect 575949 347429 575983 347463
rect 576041 338045 576075 338079
rect 575949 334577 575983 334611
rect 576041 331857 576075 331891
rect 575949 327981 575983 328015
rect 575949 321929 575983 321963
rect 576133 319481 576167 319515
rect 575949 319073 575983 319107
rect 576041 319209 576075 319243
rect 575949 315741 575983 315775
rect 576041 315945 576075 315979
rect 576133 315605 576167 315639
rect 576041 306357 576075 306391
rect 575949 299149 575983 299183
rect 575949 278749 575983 278783
rect 575949 272969 575983 273003
rect 576041 272289 576075 272323
rect 576041 270317 576075 270351
rect 575949 262701 575983 262735
rect 575949 257601 575983 257635
rect 575949 249101 575983 249135
rect 576041 257465 576075 257499
rect 576041 243117 576075 243151
rect 576225 236793 576259 236827
rect 576133 225029 576167 225063
rect 576225 225029 576259 225063
rect 576133 224893 576167 224927
rect 575949 220949 575983 220983
rect 576133 217617 576167 217651
rect 576041 217481 576075 217515
rect 576041 215985 576075 216019
rect 576133 215509 576167 215543
rect 575949 212585 575983 212619
rect 576133 212449 576167 212483
rect 576041 203065 576075 203099
rect 575949 198849 575983 198883
rect 576133 201501 576167 201535
rect 576317 199257 576351 199291
rect 576317 198713 576351 198747
rect 576041 197421 576075 197455
rect 575949 192525 575983 192559
rect 576041 192729 576075 192763
rect 576041 191097 576075 191131
rect 576225 191777 576259 191811
rect 576041 186881 576075 186915
rect 575949 182937 575983 182971
rect 576225 186269 576259 186303
rect 576225 177225 576259 177259
rect 576041 174777 576075 174811
rect 576133 175661 576167 175695
rect 575949 173961 575983 173995
rect 575949 170697 575983 170731
rect 575949 160769 575983 160803
rect 576041 170221 576075 170255
rect 576225 172533 576259 172567
rect 576133 164917 576167 164951
rect 576041 157845 576075 157879
rect 576133 157981 576167 158015
rect 575949 153425 575983 153459
rect 576133 153221 576167 153255
rect 575949 150433 575983 150467
rect 576133 149685 576167 149719
rect 575949 149345 575983 149379
rect 575949 144381 575983 144415
rect 576041 145265 576075 145299
rect 575949 140913 575983 140947
rect 576041 140301 576075 140335
rect 576225 145945 576259 145979
rect 576225 144857 576259 144891
rect 576133 137173 576167 137207
rect 575949 132549 575983 132583
rect 575949 132073 575983 132107
rect 576225 130509 576259 130543
rect 576133 127653 576167 127687
rect 576133 125545 576167 125579
rect 575949 118541 575983 118575
rect 576041 122553 576075 122587
rect 575949 118405 575983 118439
rect 576225 120717 576259 120751
rect 576317 125545 576351 125579
rect 576317 118405 576351 118439
rect 576041 117725 576075 117759
rect 576133 115821 576167 115855
rect 575949 104397 575983 104431
rect 576041 113985 576075 114019
rect 576133 110925 576167 110959
rect 576041 104261 576075 104295
rect 576133 108817 576167 108851
rect 576133 102425 576167 102459
rect 576225 93789 576259 93823
rect 576133 90593 576167 90627
rect 575949 81345 575983 81379
rect 576133 81345 576167 81379
rect 576041 79441 576075 79475
rect 576041 74749 576075 74783
rect 575949 72165 575983 72199
rect 576225 70329 576259 70363
rect 576041 67541 576075 67575
rect 575949 63325 575983 63359
rect 576317 58769 576351 58803
rect 575949 57817 575983 57851
rect 576317 57273 576351 57307
rect 575949 43469 575983 43503
rect 576041 51765 576075 51799
rect 576041 39389 576075 39423
rect 576133 43605 576167 43639
rect 575949 37213 575983 37247
rect 576041 35309 576075 35343
rect 576133 35173 576167 35207
rect 576041 33813 576075 33847
rect 576041 33065 576075 33099
rect 576041 28305 576075 28339
rect 575949 20281 575983 20315
rect 576041 24157 576075 24191
rect 576041 19329 576075 19363
rect 576133 21505 576167 21539
rect 576133 16677 576167 16711
rect 69489 7769 69523 7803
rect 69489 7497 69523 7531
rect 6929 4029 6963 4063
rect 9229 4029 9263 4063
rect 8861 3825 8895 3859
rect 9045 3757 9079 3791
rect 9229 3689 9263 3723
rect 16497 3961 16531 3995
rect 6929 2873 6963 2907
rect 16497 2873 16531 2907
<< metal1 >>
rect 150342 700680 150348 700732
rect 150400 700720 150406 700732
rect 170306 700720 170312 700732
rect 150400 700692 170312 700720
rect 150400 700680 150406 700692
rect 170306 700680 170312 700692
rect 170364 700680 170370 700732
rect 128262 700612 128268 700664
rect 128320 700652 128326 700664
rect 235166 700652 235172 700664
rect 128320 700624 235172 700652
rect 128320 700612 128326 700624
rect 235166 700612 235172 700624
rect 235224 700612 235230 700664
rect 106182 700544 106188 700596
rect 106240 700584 106246 700596
rect 300118 700584 300124 700596
rect 106240 700556 300124 700584
rect 106240 700544 106246 700556
rect 300118 700544 300124 700556
rect 300176 700544 300182 700596
rect 84102 700476 84108 700528
rect 84160 700516 84166 700528
rect 364978 700516 364984 700528
rect 84160 700488 364984 700516
rect 84160 700476 84166 700488
rect 364978 700476 364984 700488
rect 365036 700476 365042 700528
rect 40494 700408 40500 700460
rect 40552 700448 40558 700460
rect 41322 700448 41328 700460
rect 40552 700420 41328 700448
rect 40552 700408 40558 700420
rect 41322 700408 41328 700420
rect 41380 700408 41386 700460
rect 62022 700408 62028 700460
rect 62080 700448 62086 700460
rect 429838 700448 429844 700460
rect 62080 700420 429844 700448
rect 62080 700408 62086 700420
rect 429838 700408 429844 700420
rect 429896 700408 429902 700460
rect 39942 700340 39948 700392
rect 40000 700380 40006 700392
rect 494790 700380 494796 700392
rect 40000 700352 494796 700380
rect 40000 700340 40006 700352
rect 494790 700340 494796 700352
rect 494848 700340 494854 700392
rect 19242 700272 19248 700324
rect 19300 700312 19306 700324
rect 559650 700312 559656 700324
rect 19300 700284 559656 700312
rect 19300 700272 19306 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106090 699700 106096 699712
rect 105504 699672 106096 699700
rect 105504 699660 105510 699672
rect 106090 699660 106096 699672
rect 106148 699660 106154 699712
rect 17954 689936 17960 689988
rect 18012 689976 18018 689988
rect 19242 689976 19248 689988
rect 18012 689948 19248 689976
rect 18012 689936 18018 689948
rect 19242 689936 19248 689948
rect 19300 689936 19306 689988
rect 127526 689528 127532 689580
rect 127584 689568 127590 689580
rect 128262 689568 128268 689580
rect 127584 689540 128268 689568
rect 127584 689528 127590 689540
rect 128262 689528 128268 689540
rect 128320 689528 128326 689580
rect 149422 689528 149428 689580
rect 149480 689568 149486 689580
rect 150342 689568 150348 689580
rect 149480 689540 150348 689568
rect 149480 689528 149486 689540
rect 150342 689528 150348 689540
rect 150400 689528 150406 689580
rect 9490 689392 9496 689444
rect 9548 689432 9554 689444
rect 456426 689432 456432 689444
rect 9548 689404 456432 689432
rect 9548 689392 9554 689404
rect 456426 689392 456432 689404
rect 456484 689392 456490 689444
rect 106090 689324 106096 689376
rect 106148 689364 106154 689376
rect 171410 689364 171416 689376
rect 106148 689336 171416 689364
rect 106148 689324 106154 689336
rect 171410 689324 171416 689336
rect 171468 689324 171474 689376
rect 41322 689256 41328 689308
rect 41380 689296 41386 689308
rect 193306 689296 193312 689308
rect 41380 689268 193312 689296
rect 41380 689256 41386 689268
rect 193306 689256 193312 689268
rect 193364 689256 193370 689308
rect 9122 689188 9128 689240
rect 9180 689228 9186 689240
rect 237190 689228 237196 689240
rect 9180 689200 237196 689228
rect 9180 689188 9186 689200
rect 237190 689188 237196 689200
rect 237248 689188 237254 689240
rect 9030 689120 9036 689172
rect 9088 689160 9094 689172
rect 259086 689160 259092 689172
rect 9088 689132 259092 689160
rect 9088 689120 9094 689132
rect 259086 689120 259092 689132
rect 259144 689120 259150 689172
rect 9398 689052 9404 689104
rect 9456 689092 9462 689104
rect 280982 689092 280988 689104
rect 9456 689064 280988 689092
rect 9456 689052 9462 689064
rect 280982 689052 280988 689064
rect 281040 689052 281046 689104
rect 9766 688984 9772 689036
rect 9824 689024 9830 689036
rect 302970 689024 302976 689036
rect 9824 688996 302976 689024
rect 9824 688984 9830 688996
rect 302970 688984 302976 688996
rect 303028 688984 303034 689036
rect 215202 688916 215208 688968
rect 215260 688956 215266 688968
rect 576118 688956 576124 688968
rect 215260 688928 576124 688956
rect 215260 688916 215266 688928
rect 576118 688916 576124 688928
rect 576176 688916 576182 688968
rect 8938 688848 8944 688900
rect 8996 688888 9002 688900
rect 390646 688888 390652 688900
rect 8996 688860 390652 688888
rect 8996 688848 9002 688860
rect 390646 688848 390652 688860
rect 390704 688848 390710 688900
rect 9674 688780 9680 688832
rect 9732 688820 9738 688832
rect 412542 688820 412548 688832
rect 9732 688792 412548 688820
rect 9732 688780 9738 688792
rect 412542 688780 412548 688792
rect 412600 688780 412606 688832
rect 9582 688712 9588 688764
rect 9640 688752 9646 688764
rect 434438 688752 434444 688764
rect 9640 688724 434444 688752
rect 9640 688712 9646 688724
rect 434438 688712 434444 688724
rect 434496 688712 434502 688764
rect 9306 686468 9312 686520
rect 9364 686508 9370 686520
rect 368382 686508 368388 686520
rect 9364 686480 368388 686508
rect 9364 686468 9370 686480
rect 368382 686468 368388 686480
rect 368440 686468 368446 686520
rect 3326 681708 3332 681760
rect 3384 681748 3390 681760
rect 6178 681748 6184 681760
rect 3384 681720 6184 681748
rect 3384 681708 3390 681720
rect 6178 681708 6184 681720
rect 6236 681708 6242 681760
rect 575934 674908 575940 674960
rect 575992 674948 575998 674960
rect 576302 674948 576308 674960
rect 575992 674920 576308 674948
rect 575992 674908 575998 674920
rect 576302 674908 576308 674920
rect 576360 674908 576366 674960
rect 575934 652876 575940 652928
rect 575992 652916 575998 652928
rect 576302 652916 576308 652928
rect 575992 652888 576308 652916
rect 575992 652876 575998 652888
rect 576302 652876 576308 652888
rect 576360 652876 576366 652928
rect 575934 647776 575940 647828
rect 575992 647816 575998 647828
rect 576029 647819 576087 647825
rect 576029 647816 576041 647819
rect 575992 647788 576041 647816
rect 575992 647776 575998 647788
rect 576029 647785 576041 647788
rect 576075 647785 576087 647819
rect 576029 647779 576087 647785
rect 576026 634828 576032 634840
rect 575987 634800 576032 634828
rect 576026 634788 576032 634800
rect 576084 634788 576090 634840
rect 6730 627920 6736 627972
rect 6788 627960 6794 627972
rect 6914 627960 6920 627972
rect 6788 627932 6920 627960
rect 6788 627920 6794 627932
rect 6914 627920 6920 627932
rect 6972 627920 6978 627972
rect 3142 624180 3148 624232
rect 3200 624220 3206 624232
rect 6270 624220 6276 624232
rect 3200 624192 6276 624220
rect 3200 624180 3206 624192
rect 6270 624180 6276 624192
rect 6328 624180 6334 624232
rect 6641 621095 6699 621101
rect 6641 621061 6653 621095
rect 6687 621092 6699 621095
rect 6730 621092 6736 621104
rect 6687 621064 6736 621092
rect 6687 621061 6699 621064
rect 6641 621055 6699 621061
rect 6730 621052 6736 621064
rect 6788 621052 6794 621104
rect 6638 618304 6644 618316
rect 6599 618276 6644 618304
rect 6638 618264 6644 618276
rect 6696 618264 6702 618316
rect 6549 618171 6607 618177
rect 6549 618137 6561 618171
rect 6595 618168 6607 618171
rect 6638 618168 6644 618180
rect 6595 618140 6644 618168
rect 6595 618137 6607 618140
rect 6549 618131 6607 618137
rect 6638 618128 6644 618140
rect 6696 618128 6702 618180
rect 6546 608648 6552 608660
rect 6507 608620 6552 608648
rect 6546 608608 6552 608620
rect 6604 608608 6610 608660
rect 575934 602352 575940 602404
rect 575992 602392 575998 602404
rect 576029 602395 576087 602401
rect 576029 602392 576041 602395
rect 575992 602364 576041 602392
rect 575992 602352 575998 602364
rect 576029 602361 576041 602364
rect 576075 602361 576087 602395
rect 576029 602355 576087 602361
rect 6546 601740 6552 601792
rect 6604 601780 6610 601792
rect 6914 601780 6920 601792
rect 6604 601752 6920 601780
rect 6604 601740 6610 601752
rect 6914 601740 6920 601752
rect 6972 601740 6978 601792
rect 6546 601604 6552 601656
rect 6604 601644 6610 601656
rect 6914 601644 6920 601656
rect 6604 601616 6920 601644
rect 6604 601604 6610 601616
rect 6914 601604 6920 601616
rect 6972 601604 6978 601656
rect 6454 601536 6460 601588
rect 6512 601576 6518 601588
rect 6730 601576 6736 601588
rect 6512 601548 6736 601576
rect 6512 601536 6518 601548
rect 6730 601536 6736 601548
rect 6788 601536 6794 601588
rect 576026 597564 576032 597576
rect 575987 597536 576032 597564
rect 576026 597524 576032 597536
rect 576084 597524 576090 597576
rect 6546 592084 6552 592136
rect 6604 592084 6610 592136
rect 6564 592000 6592 592084
rect 6546 591948 6552 592000
rect 6604 591948 6610 592000
rect 6454 591880 6460 591932
rect 6512 591920 6518 591932
rect 6730 591920 6736 591932
rect 6512 591892 6736 591920
rect 6512 591880 6518 591892
rect 6730 591880 6736 591892
rect 6788 591880 6794 591932
rect 6546 582360 6552 582412
rect 6604 582400 6610 582412
rect 6914 582400 6920 582412
rect 6604 582372 6920 582400
rect 6604 582360 6610 582372
rect 6914 582360 6920 582372
rect 6972 582360 6978 582412
rect 6362 582224 6368 582276
rect 6420 582264 6426 582276
rect 6730 582264 6736 582276
rect 6420 582236 6736 582264
rect 6420 582224 6426 582236
rect 6730 582224 6736 582236
rect 6788 582224 6794 582276
rect 6730 572880 6736 572892
rect 6691 572852 6736 572880
rect 6730 572840 6736 572852
rect 6788 572840 6794 572892
rect 6362 572432 6368 572484
rect 6420 572472 6426 572484
rect 6822 572472 6828 572484
rect 6420 572444 6828 572472
rect 6420 572432 6426 572444
rect 6822 572432 6828 572444
rect 6880 572432 6886 572484
rect 6730 572404 6736 572416
rect 6691 572376 6736 572404
rect 6730 572364 6736 572376
rect 6788 572364 6794 572416
rect 4062 567264 4068 567316
rect 4120 567304 4126 567316
rect 7558 567304 7564 567316
rect 4120 567276 7564 567304
rect 4120 567264 4126 567276
rect 7558 567264 7564 567276
rect 7616 567264 7622 567316
rect 575934 567196 575940 567248
rect 575992 567196 575998 567248
rect 575952 567112 575980 567196
rect 575934 567060 575940 567112
rect 575992 567060 575998 567112
rect 575934 564380 575940 564392
rect 575895 564352 575940 564380
rect 575934 564340 575940 564352
rect 575992 564340 575998 564392
rect 6822 563224 6828 563236
rect 6472 563196 6828 563224
rect 6472 563100 6500 563196
rect 6822 563184 6828 563196
rect 6880 563184 6886 563236
rect 6454 563048 6460 563100
rect 6512 563048 6518 563100
rect 6362 562980 6368 563032
rect 6420 563020 6426 563032
rect 6914 563020 6920 563032
rect 6420 562992 6920 563020
rect 6420 562980 6426 562992
rect 6914 562980 6920 562992
rect 6972 562980 6978 563032
rect 575937 554795 575995 554801
rect 575937 554761 575949 554795
rect 575983 554792 575995 554795
rect 576026 554792 576032 554804
rect 575983 554764 576032 554792
rect 575983 554761 575995 554764
rect 575937 554755 575995 554761
rect 576026 554752 576032 554764
rect 576084 554752 576090 554804
rect 6362 553460 6368 553512
rect 6420 553500 6426 553512
rect 6420 553472 6868 553500
rect 6420 553460 6426 553472
rect 6840 553444 6868 553472
rect 6454 553392 6460 553444
rect 6512 553432 6518 553444
rect 6730 553432 6736 553444
rect 6512 553404 6736 553432
rect 6512 553392 6518 553404
rect 6730 553392 6736 553404
rect 6788 553392 6794 553444
rect 6822 553392 6828 553444
rect 6880 553392 6886 553444
rect 6454 553256 6460 553308
rect 6512 553296 6518 553308
rect 6822 553296 6828 553308
rect 6512 553268 6828 553296
rect 6512 553256 6518 553268
rect 6822 553256 6828 553268
rect 6880 553256 6886 553308
rect 6454 543804 6460 543856
rect 6512 543844 6518 543856
rect 6914 543844 6920 543856
rect 6512 543816 6920 543844
rect 6512 543804 6518 543816
rect 6914 543804 6920 543816
rect 6972 543804 6978 543856
rect 6362 543668 6368 543720
rect 6420 543708 6426 543720
rect 6914 543708 6920 543720
rect 6420 543680 6920 543708
rect 6420 543668 6426 543680
rect 6914 543668 6920 543680
rect 6972 543668 6978 543720
rect 575934 536800 575940 536852
rect 575992 536840 575998 536852
rect 576026 536840 576032 536852
rect 575992 536812 576032 536840
rect 575992 536800 575998 536812
rect 576026 536800 576032 536812
rect 576084 536800 576090 536852
rect 6362 534148 6368 534200
rect 6420 534188 6426 534200
rect 6420 534160 6868 534188
rect 6420 534148 6426 534160
rect 6840 534132 6868 534160
rect 6454 534080 6460 534132
rect 6512 534120 6518 534132
rect 6730 534120 6736 534132
rect 6512 534092 6736 534120
rect 6512 534080 6518 534092
rect 6730 534080 6736 534092
rect 6788 534080 6794 534132
rect 6822 534080 6828 534132
rect 6880 534080 6886 534132
rect 6454 533944 6460 533996
rect 6512 533984 6518 533996
rect 6822 533984 6828 533996
rect 6512 533956 6828 533984
rect 6512 533944 6518 533956
rect 6822 533944 6828 533956
rect 6880 533944 6886 533996
rect 6454 524424 6460 524476
rect 6512 524464 6518 524476
rect 6914 524464 6920 524476
rect 6512 524436 6920 524464
rect 6512 524424 6518 524436
rect 6914 524424 6920 524436
rect 6972 524424 6978 524476
rect 575934 522288 575940 522300
rect 575895 522260 575940 522288
rect 575934 522248 575940 522260
rect 575992 522248 575998 522300
rect 575934 519936 575940 519988
rect 575992 519976 575998 519988
rect 576302 519976 576308 519988
rect 575992 519948 576308 519976
rect 575992 519936 575998 519948
rect 576302 519936 576308 519948
rect 576360 519936 576366 519988
rect 575934 518004 575940 518016
rect 575895 517976 575940 518004
rect 575934 517964 575940 517976
rect 575992 517964 575998 518016
rect 6730 514904 6736 514956
rect 6788 514944 6794 514956
rect 6788 514916 6868 514944
rect 6788 514904 6794 514916
rect 6840 514820 6868 514916
rect 6454 514768 6460 514820
rect 6512 514808 6518 514820
rect 6730 514808 6736 514820
rect 6512 514780 6736 514808
rect 6512 514768 6518 514780
rect 6730 514768 6736 514780
rect 6788 514768 6794 514820
rect 6822 514768 6828 514820
rect 6880 514768 6886 514820
rect 575934 514740 575940 514752
rect 575895 514712 575940 514740
rect 575934 514700 575940 514712
rect 575992 514700 575998 514752
rect 576026 514700 576032 514752
rect 576084 514740 576090 514752
rect 576210 514740 576216 514752
rect 576084 514712 576216 514740
rect 576084 514700 576090 514712
rect 576210 514700 576216 514712
rect 576268 514700 576274 514752
rect 6454 514632 6460 514684
rect 6512 514672 6518 514684
rect 6822 514672 6828 514684
rect 6512 514644 6828 514672
rect 6512 514632 6518 514644
rect 6822 514632 6828 514644
rect 6880 514632 6886 514684
rect 575934 509504 575940 509516
rect 575895 509476 575940 509504
rect 575934 509464 575940 509476
rect 575992 509464 575998 509516
rect 575934 505316 575940 505368
rect 575992 505356 575998 505368
rect 576210 505356 576216 505368
rect 575992 505328 576216 505356
rect 575992 505316 575998 505328
rect 576210 505316 576216 505328
rect 576268 505316 576274 505368
rect 6454 505112 6460 505164
rect 6512 505152 6518 505164
rect 6914 505152 6920 505164
rect 6512 505124 6920 505152
rect 6512 505112 6518 505124
rect 6914 505112 6920 505124
rect 6972 505112 6978 505164
rect 6730 495592 6736 495644
rect 6788 495632 6794 495644
rect 6788 495604 6868 495632
rect 6788 495592 6794 495604
rect 6840 495508 6868 495604
rect 6454 495456 6460 495508
rect 6512 495496 6518 495508
rect 6730 495496 6736 495508
rect 6512 495468 6736 495496
rect 6512 495456 6518 495468
rect 6730 495456 6736 495468
rect 6788 495456 6794 495508
rect 6822 495456 6828 495508
rect 6880 495456 6886 495508
rect 6454 495320 6460 495372
rect 6512 495360 6518 495372
rect 6822 495360 6828 495372
rect 6512 495332 6828 495360
rect 6512 495320 6518 495332
rect 6822 495320 6828 495332
rect 6880 495320 6886 495372
rect 575937 492643 575995 492649
rect 575937 492609 575949 492643
rect 575983 492640 575995 492643
rect 576026 492640 576032 492652
rect 575983 492612 576032 492640
rect 575983 492609 575995 492612
rect 575937 492603 575995 492609
rect 576026 492600 576032 492612
rect 576084 492600 576090 492652
rect 575934 487772 575940 487824
rect 575992 487812 575998 487824
rect 576029 487815 576087 487821
rect 576029 487812 576041 487815
rect 575992 487784 576041 487812
rect 575992 487772 575998 487784
rect 576029 487781 576041 487784
rect 576075 487781 576087 487815
rect 576029 487775 576087 487781
rect 576118 487092 576124 487144
rect 576176 487132 576182 487144
rect 579614 487132 579620 487144
rect 576176 487104 579620 487132
rect 576176 487092 576182 487104
rect 579614 487092 579620 487104
rect 579672 487092 579678 487144
rect 6454 485800 6460 485852
rect 6512 485840 6518 485852
rect 6914 485840 6920 485852
rect 6512 485812 6920 485840
rect 6512 485800 6518 485812
rect 6914 485800 6920 485812
rect 6972 485800 6978 485852
rect 575934 485732 575940 485784
rect 575992 485772 575998 485784
rect 576026 485772 576032 485784
rect 575992 485744 576032 485772
rect 575992 485732 575998 485744
rect 576026 485732 576032 485744
rect 576084 485732 576090 485784
rect 575934 485596 575940 485648
rect 575992 485636 575998 485648
rect 576029 485639 576087 485645
rect 576029 485636 576041 485639
rect 575992 485608 576041 485636
rect 575992 485596 575998 485608
rect 576029 485605 576041 485608
rect 576075 485605 576087 485639
rect 576029 485599 576087 485605
rect 575934 485500 575940 485512
rect 575895 485472 575940 485500
rect 575934 485460 575940 485472
rect 575992 485460 575998 485512
rect 6730 476212 6736 476264
rect 6788 476252 6794 476264
rect 6788 476224 6868 476252
rect 6788 476212 6794 476224
rect 6840 476128 6868 476224
rect 6454 476076 6460 476128
rect 6512 476116 6518 476128
rect 6730 476116 6736 476128
rect 6512 476088 6736 476116
rect 6512 476076 6518 476088
rect 6730 476076 6736 476088
rect 6788 476076 6794 476128
rect 6822 476076 6828 476128
rect 6880 476076 6886 476128
rect 575934 466488 575940 466540
rect 575992 466528 575998 466540
rect 575992 466500 576164 466528
rect 575992 466488 575998 466500
rect 576026 466460 576032 466472
rect 575952 466432 576032 466460
rect 575952 466268 575980 466432
rect 576026 466420 576032 466432
rect 576084 466420 576090 466472
rect 576136 466268 576164 466500
rect 575934 466216 575940 466268
rect 575992 466216 575998 466268
rect 576118 466216 576124 466268
rect 576176 466216 576182 466268
rect 6730 456900 6736 456952
rect 6788 456940 6794 456952
rect 6788 456912 6868 456940
rect 6788 456900 6794 456912
rect 6840 456816 6868 456912
rect 6454 456764 6460 456816
rect 6512 456804 6518 456816
rect 6730 456804 6736 456816
rect 6512 456776 6736 456804
rect 6512 456764 6518 456776
rect 6730 456764 6736 456776
rect 6788 456764 6794 456816
rect 6822 456764 6828 456816
rect 6880 456764 6886 456816
rect 576026 447108 576032 447160
rect 576084 447108 576090 447160
rect 576044 447080 576072 447108
rect 576118 447080 576124 447092
rect 576044 447052 576124 447080
rect 576118 447040 576124 447052
rect 576176 447040 576182 447092
rect 6730 437588 6736 437640
rect 6788 437628 6794 437640
rect 6788 437600 6868 437628
rect 6788 437588 6794 437600
rect 6840 437504 6868 437600
rect 6454 437452 6460 437504
rect 6512 437492 6518 437504
rect 6730 437492 6736 437504
rect 6512 437464 6736 437492
rect 6512 437452 6518 437464
rect 6730 437452 6736 437464
rect 6788 437452 6794 437504
rect 6822 437452 6828 437504
rect 6880 437452 6886 437504
rect 576026 428476 576032 428528
rect 576084 428516 576090 428528
rect 576121 428519 576179 428525
rect 576121 428516 576133 428519
rect 576084 428488 576133 428516
rect 576084 428476 576090 428488
rect 576121 428485 576133 428488
rect 576167 428485 576179 428519
rect 576121 428479 576179 428485
rect 575934 427660 575940 427712
rect 575992 427660 575998 427712
rect 575952 427576 575980 427660
rect 575934 427524 575940 427576
rect 575992 427524 575998 427576
rect 576118 417840 576124 417852
rect 576079 417812 576124 417840
rect 576118 417800 576124 417812
rect 576176 417800 576182 417852
rect 575934 405560 575940 405612
rect 575992 405600 575998 405612
rect 576029 405603 576087 405609
rect 576029 405600 576041 405603
rect 575992 405572 576041 405600
rect 575992 405560 575998 405572
rect 576029 405569 576041 405572
rect 576075 405569 576087 405603
rect 576029 405563 576087 405569
rect 6454 398828 6460 398880
rect 6512 398868 6518 398880
rect 6730 398868 6736 398880
rect 6512 398840 6736 398868
rect 6512 398828 6518 398840
rect 6730 398828 6736 398840
rect 6788 398828 6794 398880
rect 575934 396992 575940 397044
rect 575992 397032 575998 397044
rect 576118 397032 576124 397044
rect 575992 397004 576124 397032
rect 575992 396992 575998 397004
rect 576118 396992 576124 397004
rect 576176 396992 576182 397044
rect 576026 396080 576032 396092
rect 575987 396052 576032 396080
rect 576026 396040 576032 396052
rect 576084 396040 576090 396092
rect 575934 390096 575940 390108
rect 575895 390068 575940 390096
rect 575934 390056 575940 390068
rect 575992 390056 575998 390108
rect 6454 389104 6460 389156
rect 6512 389144 6518 389156
rect 6730 389144 6736 389156
rect 6512 389116 6736 389144
rect 6512 389104 6518 389116
rect 6730 389104 6736 389116
rect 6788 389104 6794 389156
rect 6822 389104 6828 389156
rect 6880 389104 6886 389156
rect 6362 389036 6368 389088
rect 6420 389076 6426 389088
rect 6840 389076 6868 389104
rect 6420 389048 6868 389076
rect 6420 389036 6426 389048
rect 575934 384344 575940 384396
rect 575992 384384 575998 384396
rect 576029 384387 576087 384393
rect 576029 384384 576041 384387
rect 575992 384356 576041 384384
rect 575992 384344 575998 384356
rect 576029 384353 576041 384356
rect 576075 384353 576087 384387
rect 576029 384347 576087 384353
rect 6362 379584 6368 379636
rect 6420 379624 6426 379636
rect 576029 379627 576087 379633
rect 576029 379624 576041 379627
rect 6420 379596 6868 379624
rect 6420 379584 6426 379596
rect 6840 379568 6868 379596
rect 575952 379596 576041 379624
rect 6454 379516 6460 379568
rect 6512 379556 6518 379568
rect 6730 379556 6736 379568
rect 6512 379528 6736 379556
rect 6512 379516 6518 379528
rect 6730 379516 6736 379528
rect 6788 379516 6794 379568
rect 6822 379516 6828 379568
rect 6880 379516 6886 379568
rect 575952 379488 575980 379596
rect 576029 379593 576041 379596
rect 576075 379593 576087 379627
rect 576029 379587 576087 379593
rect 576026 379488 576032 379500
rect 575952 379460 576032 379488
rect 576026 379448 576032 379460
rect 576084 379448 576090 379500
rect 575937 379423 575995 379429
rect 575937 379389 575949 379423
rect 575983 379420 575995 379423
rect 576118 379420 576124 379432
rect 575983 379392 576124 379420
rect 575983 379389 575995 379392
rect 575937 379383 575995 379389
rect 576118 379380 576124 379392
rect 576176 379380 576182 379432
rect 576118 376700 576124 376712
rect 576079 376672 576124 376700
rect 576118 376660 576124 376672
rect 576176 376660 576182 376712
rect 576026 371940 576032 371952
rect 575987 371912 576032 371940
rect 576026 371900 576032 371912
rect 576084 371900 576090 371952
rect 6454 369792 6460 369844
rect 6512 369832 6518 369844
rect 6730 369832 6736 369844
rect 6512 369804 6736 369832
rect 6512 369792 6518 369804
rect 6730 369792 6736 369804
rect 6788 369792 6794 369844
rect 6822 369792 6828 369844
rect 6880 369792 6886 369844
rect 6362 369724 6368 369776
rect 6420 369764 6426 369776
rect 6840 369764 6868 369792
rect 6420 369736 6868 369764
rect 6420 369724 6426 369736
rect 575934 366460 575940 366512
rect 575992 366500 575998 366512
rect 576029 366503 576087 366509
rect 576029 366500 576041 366503
rect 575992 366472 576041 366500
rect 575992 366460 575998 366472
rect 576029 366469 576041 366472
rect 576075 366469 576087 366503
rect 576029 366463 576087 366469
rect 575934 365848 575940 365900
rect 575992 365888 575998 365900
rect 576121 365891 576179 365897
rect 576121 365888 576133 365891
rect 575992 365860 576133 365888
rect 575992 365848 575998 365860
rect 576121 365857 576133 365860
rect 576167 365857 576179 365891
rect 576121 365851 576179 365857
rect 575934 361264 575940 361276
rect 575895 361236 575940 361264
rect 575934 361224 575940 361236
rect 575992 361224 575998 361276
rect 6362 360272 6368 360324
rect 6420 360312 6426 360324
rect 6420 360284 6868 360312
rect 6420 360272 6426 360284
rect 6840 360256 6868 360284
rect 6454 360204 6460 360256
rect 6512 360244 6518 360256
rect 6730 360244 6736 360256
rect 6512 360216 6736 360244
rect 6512 360204 6518 360216
rect 6730 360204 6736 360216
rect 6788 360204 6794 360256
rect 6822 360204 6828 360256
rect 6880 360204 6886 360256
rect 575934 359456 575940 359508
rect 575992 359496 575998 359508
rect 576029 359499 576087 359505
rect 576029 359496 576041 359499
rect 575992 359468 576041 359496
rect 575992 359456 575998 359468
rect 576029 359465 576041 359468
rect 576075 359465 576087 359499
rect 576029 359459 576087 359465
rect 575934 359360 575940 359372
rect 575895 359332 575940 359360
rect 575934 359320 575940 359332
rect 575992 359320 575998 359372
rect 575934 358980 575940 359032
rect 575992 359020 575998 359032
rect 576029 359023 576087 359029
rect 576029 359020 576041 359023
rect 575992 358992 576041 359020
rect 575992 358980 575998 358992
rect 576029 358989 576041 358992
rect 576075 358989 576087 359023
rect 576029 358983 576087 358989
rect 575934 352696 575940 352708
rect 575895 352668 575940 352696
rect 575934 352656 575940 352668
rect 575992 352656 575998 352708
rect 6454 350480 6460 350532
rect 6512 350520 6518 350532
rect 6730 350520 6736 350532
rect 6512 350492 6736 350520
rect 6512 350480 6518 350492
rect 6730 350480 6736 350492
rect 6788 350480 6794 350532
rect 6822 350480 6828 350532
rect 6880 350480 6886 350532
rect 6362 350412 6368 350464
rect 6420 350452 6426 350464
rect 6840 350452 6868 350480
rect 6420 350424 6868 350452
rect 6420 350412 6426 350424
rect 575934 347460 575940 347472
rect 575895 347432 575940 347460
rect 575934 347420 575940 347432
rect 575992 347420 575998 347472
rect 6362 340960 6368 341012
rect 6420 341000 6426 341012
rect 6420 340972 6868 341000
rect 6420 340960 6426 340972
rect 6840 340944 6868 340972
rect 6454 340892 6460 340944
rect 6512 340932 6518 340944
rect 6730 340932 6736 340944
rect 6512 340904 6736 340932
rect 6512 340892 6518 340904
rect 6730 340892 6736 340904
rect 6788 340892 6794 340944
rect 6822 340892 6828 340944
rect 6880 340892 6886 340944
rect 575934 338036 575940 338088
rect 575992 338076 575998 338088
rect 576029 338079 576087 338085
rect 576029 338076 576041 338079
rect 575992 338048 576041 338076
rect 575992 338036 575998 338048
rect 576029 338045 576041 338048
rect 576075 338045 576087 338079
rect 576029 338039 576087 338045
rect 575934 334608 575940 334620
rect 575895 334580 575940 334608
rect 575934 334568 575940 334580
rect 575992 334568 575998 334620
rect 575934 331848 575940 331900
rect 575992 331888 575998 331900
rect 576029 331891 576087 331897
rect 576029 331888 576041 331891
rect 575992 331860 576041 331888
rect 575992 331848 575998 331860
rect 576029 331857 576041 331860
rect 576075 331857 576087 331891
rect 576029 331851 576087 331857
rect 6362 331168 6368 331220
rect 6420 331208 6426 331220
rect 6730 331208 6736 331220
rect 6420 331180 6736 331208
rect 6420 331168 6426 331180
rect 6730 331168 6736 331180
rect 6788 331168 6794 331220
rect 6822 331168 6828 331220
rect 6880 331168 6886 331220
rect 6086 331100 6092 331152
rect 6144 331140 6150 331152
rect 6840 331140 6868 331168
rect 6144 331112 6868 331140
rect 6144 331100 6150 331112
rect 575934 328012 575940 328024
rect 575895 327984 575940 328012
rect 575934 327972 575940 327984
rect 575992 327972 575998 328024
rect 576118 325660 576124 325712
rect 576176 325700 576182 325712
rect 576210 325700 576216 325712
rect 576176 325672 576216 325700
rect 576176 325660 576182 325672
rect 576210 325660 576216 325672
rect 576268 325660 576274 325712
rect 575934 321960 575940 321972
rect 575895 321932 575940 321960
rect 575934 321920 575940 321932
rect 575992 321920 575998 321972
rect 6086 321648 6092 321700
rect 6144 321688 6150 321700
rect 6144 321660 6868 321688
rect 6144 321648 6150 321660
rect 6840 321632 6868 321660
rect 6362 321580 6368 321632
rect 6420 321620 6426 321632
rect 6730 321620 6736 321632
rect 6420 321592 6736 321620
rect 6420 321580 6426 321592
rect 6730 321580 6736 321592
rect 6788 321580 6794 321632
rect 6822 321580 6828 321632
rect 6880 321580 6886 321632
rect 575934 319472 575940 319524
rect 575992 319512 575998 319524
rect 576121 319515 576179 319521
rect 576121 319512 576133 319515
rect 575992 319484 576133 319512
rect 575992 319472 575998 319484
rect 576121 319481 576133 319484
rect 576167 319481 576179 319515
rect 576121 319475 576179 319481
rect 575934 319200 575940 319252
rect 575992 319240 575998 319252
rect 576029 319243 576087 319249
rect 576029 319240 576041 319243
rect 575992 319212 576041 319240
rect 575992 319200 575998 319212
rect 576029 319209 576041 319212
rect 576075 319209 576087 319243
rect 576029 319203 576087 319209
rect 575934 319104 575940 319116
rect 575895 319076 575940 319104
rect 575934 319064 575940 319076
rect 575992 319064 575998 319116
rect 576029 315979 576087 315985
rect 576029 315945 576041 315979
rect 576075 315976 576087 315979
rect 576118 315976 576124 315988
rect 576075 315948 576124 315976
rect 576075 315945 576087 315948
rect 576029 315939 576087 315945
rect 576118 315936 576124 315948
rect 576176 315936 576182 315988
rect 575934 315772 575940 315784
rect 575895 315744 575940 315772
rect 575934 315732 575940 315744
rect 575992 315732 575998 315784
rect 575934 315596 575940 315648
rect 575992 315636 575998 315648
rect 576121 315639 576179 315645
rect 576121 315636 576133 315639
rect 575992 315608 576133 315636
rect 575992 315596 575998 315608
rect 576121 315605 576133 315608
rect 576167 315605 576179 315639
rect 576121 315599 576179 315605
rect 6086 311788 6092 311840
rect 6144 311828 6150 311840
rect 6730 311828 6736 311840
rect 6144 311800 6736 311828
rect 6144 311788 6150 311800
rect 6730 311788 6736 311800
rect 6788 311788 6794 311840
rect 6822 311788 6828 311840
rect 6880 311788 6886 311840
rect 6362 311720 6368 311772
rect 6420 311760 6426 311772
rect 6840 311760 6868 311788
rect 6420 311732 6868 311760
rect 6420 311720 6426 311732
rect 575934 307776 575940 307828
rect 575992 307816 575998 307828
rect 576302 307816 576308 307828
rect 575992 307788 576308 307816
rect 575992 307776 575998 307788
rect 576302 307776 576308 307788
rect 576360 307776 576366 307828
rect 576026 306388 576032 306400
rect 575987 306360 576032 306388
rect 576026 306348 576032 306360
rect 576084 306348 576090 306400
rect 6362 302744 6368 302796
rect 6420 302784 6426 302796
rect 6420 302756 6868 302784
rect 6420 302744 6426 302756
rect 6840 302252 6868 302756
rect 6086 302200 6092 302252
rect 6144 302240 6150 302252
rect 6730 302240 6736 302252
rect 6144 302212 6736 302240
rect 6144 302200 6150 302212
rect 6730 302200 6736 302212
rect 6788 302200 6794 302252
rect 6822 302200 6828 302252
rect 6880 302200 6886 302252
rect 575934 299180 575940 299192
rect 575895 299152 575940 299180
rect 575934 299140 575940 299152
rect 575992 299140 575998 299192
rect 6086 292476 6092 292528
rect 6144 292516 6150 292528
rect 6730 292516 6736 292528
rect 6144 292488 6736 292516
rect 6144 292476 6150 292488
rect 6730 292476 6736 292488
rect 6788 292476 6794 292528
rect 6822 292476 6828 292528
rect 6880 292476 6886 292528
rect 5994 292408 6000 292460
rect 6052 292448 6058 292460
rect 6840 292448 6868 292476
rect 6052 292420 6868 292448
rect 6052 292408 6058 292420
rect 575934 288464 575940 288516
rect 575992 288504 575998 288516
rect 576118 288504 576124 288516
rect 575992 288476 576124 288504
rect 575992 288464 575998 288476
rect 576118 288464 576124 288476
rect 576176 288464 576182 288516
rect 575934 286424 575940 286476
rect 575992 286424 575998 286476
rect 576026 286424 576032 286476
rect 576084 286424 576090 286476
rect 575952 286272 575980 286424
rect 576044 286272 576072 286424
rect 575934 286220 575940 286272
rect 575992 286220 575998 286272
rect 576026 286220 576032 286272
rect 576084 286220 576090 286272
rect 5994 282956 6000 283008
rect 6052 282996 6058 283008
rect 6052 282968 6868 282996
rect 6052 282956 6058 282968
rect 6840 282940 6868 282968
rect 6086 282888 6092 282940
rect 6144 282928 6150 282940
rect 6730 282928 6736 282940
rect 6144 282900 6736 282928
rect 6144 282888 6150 282900
rect 6730 282888 6736 282900
rect 6788 282888 6794 282940
rect 6822 282888 6828 282940
rect 6880 282888 6886 282940
rect 575934 278876 575940 278928
rect 575992 278916 575998 278928
rect 576118 278916 576124 278928
rect 575992 278888 576124 278916
rect 575992 278876 575998 278888
rect 576118 278876 576124 278888
rect 576176 278876 576182 278928
rect 575934 278780 575940 278792
rect 575895 278752 575940 278780
rect 575934 278740 575940 278752
rect 575992 278740 575998 278792
rect 6086 273164 6092 273216
rect 6144 273204 6150 273216
rect 6730 273204 6736 273216
rect 6144 273176 6736 273204
rect 6144 273164 6150 273176
rect 6730 273164 6736 273176
rect 6788 273164 6794 273216
rect 6822 273164 6828 273216
rect 6880 273164 6886 273216
rect 5994 273096 6000 273148
rect 6052 273136 6058 273148
rect 6840 273136 6868 273164
rect 6052 273108 6868 273136
rect 6052 273096 6058 273108
rect 575934 273000 575940 273012
rect 575895 272972 575940 273000
rect 575934 272960 575940 272972
rect 575992 272960 575998 273012
rect 576026 272280 576032 272332
rect 576084 272320 576090 272332
rect 576084 272292 576129 272320
rect 576084 272280 576090 272292
rect 576026 270308 576032 270360
rect 576084 270348 576090 270360
rect 576084 270320 576129 270348
rect 576084 270308 576090 270320
rect 5994 263644 6000 263696
rect 6052 263684 6058 263696
rect 6052 263656 6868 263684
rect 6052 263644 6058 263656
rect 6840 263628 6868 263656
rect 6086 263576 6092 263628
rect 6144 263616 6150 263628
rect 6730 263616 6736 263628
rect 6144 263588 6736 263616
rect 6144 263576 6150 263588
rect 6730 263576 6736 263588
rect 6788 263576 6794 263628
rect 6822 263576 6828 263628
rect 6880 263576 6886 263628
rect 575934 262896 575940 262948
rect 575992 262936 575998 262948
rect 576210 262936 576216 262948
rect 575992 262908 576216 262936
rect 575992 262896 575998 262908
rect 576210 262896 576216 262908
rect 576268 262896 576274 262948
rect 575934 262732 575940 262744
rect 575895 262704 575940 262732
rect 575934 262692 575940 262704
rect 575992 262692 575998 262744
rect 575934 257632 575940 257644
rect 575895 257604 575940 257632
rect 575934 257592 575940 257604
rect 575992 257592 575998 257644
rect 575934 257456 575940 257508
rect 575992 257496 575998 257508
rect 576029 257499 576087 257505
rect 576029 257496 576041 257499
rect 575992 257468 576041 257496
rect 575992 257456 575998 257468
rect 576029 257465 576041 257468
rect 576075 257465 576087 257499
rect 576029 257459 576087 257465
rect 6086 253852 6092 253904
rect 6144 253892 6150 253904
rect 6730 253892 6736 253904
rect 6144 253864 6736 253892
rect 6144 253852 6150 253864
rect 6730 253852 6736 253864
rect 6788 253852 6794 253904
rect 6822 253852 6828 253904
rect 6880 253852 6886 253904
rect 5994 253784 6000 253836
rect 6052 253824 6058 253836
rect 6840 253824 6868 253852
rect 6052 253796 6868 253824
rect 6052 253784 6058 253796
rect 575934 253240 575940 253292
rect 575992 253240 575998 253292
rect 575952 253088 575980 253240
rect 575934 253036 575940 253088
rect 575992 253036 575998 253088
rect 575934 249132 575940 249144
rect 575895 249104 575940 249132
rect 575934 249092 575940 249104
rect 575992 249092 575998 249144
rect 5994 244332 6000 244384
rect 6052 244372 6058 244384
rect 6052 244344 6868 244372
rect 6052 244332 6058 244344
rect 6840 244316 6868 244344
rect 6086 244264 6092 244316
rect 6144 244304 6150 244316
rect 6730 244304 6736 244316
rect 6144 244276 6736 244304
rect 6144 244264 6150 244276
rect 6730 244264 6736 244276
rect 6788 244264 6794 244316
rect 6822 244264 6828 244316
rect 6880 244264 6886 244316
rect 576026 243148 576032 243160
rect 575987 243120 576032 243148
rect 576026 243108 576032 243120
rect 576084 243108 576090 243160
rect 575934 241680 575940 241732
rect 575992 241720 575998 241732
rect 576302 241720 576308 241732
rect 575992 241692 576308 241720
rect 575992 241680 575998 241692
rect 576302 241680 576308 241692
rect 576360 241680 576366 241732
rect 576026 241408 576032 241460
rect 576084 241408 576090 241460
rect 576044 241244 576072 241408
rect 576118 241244 576124 241256
rect 576044 241216 576124 241244
rect 576118 241204 576124 241216
rect 576176 241204 576182 241256
rect 576210 236824 576216 236836
rect 576171 236796 576216 236824
rect 576210 236784 576216 236796
rect 576268 236784 576274 236836
rect 575934 236648 575940 236700
rect 575992 236688 575998 236700
rect 576210 236688 576216 236700
rect 575992 236660 576216 236688
rect 575992 236648 575998 236660
rect 576210 236648 576216 236660
rect 576268 236648 576274 236700
rect 575934 235016 575940 235068
rect 575992 235056 575998 235068
rect 576302 235056 576308 235068
rect 575992 235028 576308 235056
rect 575992 235016 575998 235028
rect 576302 235016 576308 235028
rect 576360 235016 576366 235068
rect 6086 234540 6092 234592
rect 6144 234580 6150 234592
rect 6730 234580 6736 234592
rect 6144 234552 6736 234580
rect 6144 234540 6150 234552
rect 6730 234540 6736 234552
rect 6788 234540 6794 234592
rect 6822 234540 6828 234592
rect 6880 234540 6886 234592
rect 5994 234472 6000 234524
rect 6052 234512 6058 234524
rect 6840 234512 6868 234540
rect 6052 234484 6868 234512
rect 6052 234472 6058 234484
rect 576026 234268 576032 234320
rect 576084 234308 576090 234320
rect 576394 234308 576400 234320
rect 576084 234280 576400 234308
rect 576084 234268 576090 234280
rect 576394 234268 576400 234280
rect 576452 234268 576458 234320
rect 5994 225020 6000 225072
rect 6052 225060 6058 225072
rect 576121 225063 576179 225069
rect 6052 225032 6868 225060
rect 6052 225020 6058 225032
rect 6840 225004 6868 225032
rect 576121 225029 576133 225063
rect 576167 225060 576179 225063
rect 576213 225063 576271 225069
rect 576213 225060 576225 225063
rect 576167 225032 576225 225060
rect 576167 225029 576179 225032
rect 576121 225023 576179 225029
rect 576213 225029 576225 225032
rect 576259 225029 576271 225063
rect 576213 225023 576271 225029
rect 6086 224952 6092 225004
rect 6144 224992 6150 225004
rect 6730 224992 6736 225004
rect 6144 224964 6736 224992
rect 6144 224952 6150 224964
rect 6730 224952 6736 224964
rect 6788 224952 6794 225004
rect 6822 224952 6828 225004
rect 6880 224952 6886 225004
rect 576118 224924 576124 224936
rect 576079 224896 576124 224924
rect 576118 224884 576124 224896
rect 576176 224884 576182 224936
rect 575934 220980 575940 220992
rect 575895 220952 575940 220980
rect 575934 220940 575940 220952
rect 575992 220940 575998 220992
rect 575934 217608 575940 217660
rect 575992 217648 575998 217660
rect 576121 217651 576179 217657
rect 576121 217648 576133 217651
rect 575992 217620 576133 217648
rect 575992 217608 575998 217620
rect 576121 217617 576133 217620
rect 576167 217617 576179 217651
rect 576121 217611 576179 217617
rect 576026 217512 576032 217524
rect 575987 217484 576032 217512
rect 576026 217472 576032 217484
rect 576084 217472 576090 217524
rect 576210 217472 576216 217524
rect 576268 217512 576274 217524
rect 576394 217512 576400 217524
rect 576268 217484 576400 217512
rect 576268 217472 576274 217484
rect 576394 217472 576400 217484
rect 576452 217472 576458 217524
rect 579062 216316 579068 216368
rect 579120 216356 579126 216368
rect 580626 216356 580632 216368
rect 579120 216328 580632 216356
rect 579120 216316 579126 216328
rect 580626 216316 580632 216328
rect 580684 216316 580690 216368
rect 575934 215976 575940 216028
rect 575992 216016 575998 216028
rect 576029 216019 576087 216025
rect 576029 216016 576041 216019
rect 575992 215988 576041 216016
rect 575992 215976 575998 215988
rect 576029 215985 576041 215988
rect 576075 215985 576087 216019
rect 576029 215979 576087 215985
rect 575934 215500 575940 215552
rect 575992 215540 575998 215552
rect 576121 215543 576179 215549
rect 576121 215540 576133 215543
rect 575992 215512 576133 215540
rect 575992 215500 575998 215512
rect 576121 215509 576133 215512
rect 576167 215509 576179 215543
rect 576121 215503 576179 215509
rect 6086 215228 6092 215280
rect 6144 215268 6150 215280
rect 6730 215268 6736 215280
rect 6144 215240 6736 215268
rect 6144 215228 6150 215240
rect 6730 215228 6736 215240
rect 6788 215228 6794 215280
rect 6822 215228 6828 215280
rect 6880 215228 6886 215280
rect 5994 215160 6000 215212
rect 6052 215200 6058 215212
rect 6840 215200 6868 215228
rect 6052 215172 6868 215200
rect 6052 215160 6058 215172
rect 575937 212619 575995 212625
rect 575937 212585 575949 212619
rect 575983 212616 575995 212619
rect 576118 212616 576124 212628
rect 575983 212588 576124 212616
rect 575983 212585 575995 212588
rect 575937 212579 575995 212585
rect 576118 212576 576124 212588
rect 576176 212576 576182 212628
rect 576118 212480 576124 212492
rect 576079 212452 576124 212480
rect 576118 212440 576124 212452
rect 576176 212440 576182 212492
rect 5994 205708 6000 205760
rect 6052 205748 6058 205760
rect 6052 205720 6868 205748
rect 6052 205708 6058 205720
rect 6840 205692 6868 205720
rect 6086 205640 6092 205692
rect 6144 205680 6150 205692
rect 6730 205680 6736 205692
rect 6144 205652 6736 205680
rect 6144 205640 6150 205652
rect 6730 205640 6736 205652
rect 6788 205640 6794 205692
rect 6822 205640 6828 205692
rect 6880 205640 6886 205692
rect 576026 203096 576032 203108
rect 575987 203068 576032 203096
rect 576026 203056 576032 203068
rect 576084 203056 576090 203108
rect 575934 202716 575940 202768
rect 575992 202756 575998 202768
rect 576210 202756 576216 202768
rect 575992 202728 576216 202756
rect 575992 202716 575998 202728
rect 576210 202716 576216 202728
rect 576268 202716 576274 202768
rect 576121 201535 576179 201541
rect 576121 201501 576133 201535
rect 576167 201532 576179 201535
rect 576210 201532 576216 201544
rect 576167 201504 576216 201532
rect 576167 201501 576179 201504
rect 576121 201495 576179 201501
rect 576210 201492 576216 201504
rect 576268 201492 576274 201544
rect 575934 199248 575940 199300
rect 575992 199288 575998 199300
rect 576305 199291 576363 199297
rect 576305 199288 576317 199291
rect 575992 199260 576317 199288
rect 575992 199248 575998 199260
rect 576305 199257 576317 199260
rect 576351 199257 576363 199291
rect 576305 199251 576363 199257
rect 575937 198883 575995 198889
rect 575937 198849 575949 198883
rect 575983 198880 575995 198883
rect 576302 198880 576308 198892
rect 575983 198852 576308 198880
rect 575983 198849 575995 198852
rect 575937 198843 575995 198849
rect 576302 198840 576308 198852
rect 576360 198840 576366 198892
rect 576302 198744 576308 198756
rect 576263 198716 576308 198744
rect 576302 198704 576308 198716
rect 576360 198704 576366 198756
rect 576029 197455 576087 197461
rect 576029 197421 576041 197455
rect 576075 197452 576087 197455
rect 576075 197424 576164 197452
rect 576075 197421 576087 197424
rect 576029 197415 576087 197421
rect 576136 197396 576164 197424
rect 576118 197344 576124 197396
rect 576176 197344 576182 197396
rect 6086 195916 6092 195968
rect 6144 195956 6150 195968
rect 6730 195956 6736 195968
rect 6144 195928 6736 195956
rect 6144 195916 6150 195928
rect 6730 195916 6736 195928
rect 6788 195916 6794 195968
rect 6822 195916 6828 195968
rect 6880 195916 6886 195968
rect 5994 195848 6000 195900
rect 6052 195888 6058 195900
rect 6840 195888 6868 195916
rect 6052 195860 6868 195888
rect 6052 195848 6058 195860
rect 579062 194012 579068 194064
rect 579120 194052 579126 194064
rect 580718 194052 580724 194064
rect 579120 194024 580724 194052
rect 579120 194012 579126 194024
rect 580718 194012 580724 194024
rect 580776 194012 580782 194064
rect 576026 192760 576032 192772
rect 575987 192732 576032 192760
rect 576026 192720 576032 192732
rect 576084 192720 576090 192772
rect 575937 192559 575995 192565
rect 575937 192525 575949 192559
rect 575983 192556 575995 192559
rect 576118 192556 576124 192568
rect 575983 192528 576124 192556
rect 575983 192525 575995 192528
rect 575937 192519 575995 192525
rect 576118 192516 576124 192528
rect 576176 192516 576182 192568
rect 576210 191808 576216 191820
rect 576171 191780 576216 191808
rect 576210 191768 576216 191780
rect 576268 191768 576274 191820
rect 576026 191128 576032 191140
rect 575987 191100 576032 191128
rect 576026 191088 576032 191100
rect 576084 191088 576090 191140
rect 575934 186872 575940 186924
rect 575992 186912 575998 186924
rect 576029 186915 576087 186921
rect 576029 186912 576041 186915
rect 575992 186884 576041 186912
rect 575992 186872 575998 186884
rect 576029 186881 576041 186884
rect 576075 186881 576087 186915
rect 576029 186875 576087 186881
rect 5994 186396 6000 186448
rect 6052 186436 6058 186448
rect 6052 186408 6868 186436
rect 6052 186396 6058 186408
rect 6840 186380 6868 186408
rect 6086 186328 6092 186380
rect 6144 186368 6150 186380
rect 6730 186368 6736 186380
rect 6144 186340 6736 186368
rect 6144 186328 6150 186340
rect 6730 186328 6736 186340
rect 6788 186328 6794 186380
rect 6822 186328 6828 186380
rect 6880 186328 6886 186380
rect 576210 186300 576216 186312
rect 576171 186272 576216 186300
rect 576210 186260 576216 186272
rect 576268 186260 576274 186312
rect 575934 184900 575940 184952
rect 575992 184940 575998 184952
rect 576302 184940 576308 184952
rect 575992 184912 576308 184940
rect 575992 184900 575998 184912
rect 576302 184900 576308 184912
rect 576360 184900 576366 184952
rect 575934 183336 575940 183388
rect 575992 183376 575998 183388
rect 576302 183376 576308 183388
rect 575992 183348 576308 183376
rect 575992 183336 575998 183348
rect 576302 183336 576308 183348
rect 576360 183336 576366 183388
rect 575937 182971 575995 182977
rect 575937 182937 575949 182971
rect 575983 182968 575995 182971
rect 576026 182968 576032 182980
rect 575983 182940 576032 182968
rect 575983 182937 575995 182940
rect 575937 182931 575995 182937
rect 576026 182928 576032 182940
rect 576084 182928 576090 182980
rect 575934 177216 575940 177268
rect 575992 177256 575998 177268
rect 576213 177259 576271 177265
rect 576213 177256 576225 177259
rect 575992 177228 576225 177256
rect 575992 177216 575998 177228
rect 576213 177225 576225 177228
rect 576259 177225 576271 177259
rect 576213 177219 576271 177225
rect 6086 176604 6092 176656
rect 6144 176644 6150 176656
rect 6730 176644 6736 176656
rect 6144 176616 6736 176644
rect 6144 176604 6150 176616
rect 6730 176604 6736 176616
rect 6788 176604 6794 176656
rect 6822 176604 6828 176656
rect 6880 176604 6886 176656
rect 5994 176536 6000 176588
rect 6052 176576 6058 176588
rect 6840 176576 6868 176604
rect 6052 176548 6868 176576
rect 6052 176536 6058 176548
rect 575934 175652 575940 175704
rect 575992 175692 575998 175704
rect 576121 175695 576179 175701
rect 576121 175692 576133 175695
rect 575992 175664 576133 175692
rect 575992 175652 575998 175664
rect 576121 175661 576133 175664
rect 576167 175661 576179 175695
rect 576121 175655 576179 175661
rect 575934 174768 575940 174820
rect 575992 174808 575998 174820
rect 576029 174811 576087 174817
rect 576029 174808 576041 174811
rect 575992 174780 576041 174808
rect 575992 174768 575998 174780
rect 576029 174777 576041 174780
rect 576075 174777 576087 174811
rect 576029 174771 576087 174777
rect 575934 173992 575940 174004
rect 575895 173964 575940 173992
rect 575934 173952 575940 173964
rect 575992 173952 575998 174004
rect 576118 172524 576124 172576
rect 576176 172564 576182 172576
rect 576213 172567 576271 172573
rect 576213 172564 576225 172567
rect 576176 172536 576225 172564
rect 576176 172524 576182 172536
rect 576213 172533 576225 172536
rect 576259 172533 576271 172567
rect 576213 172527 576271 172533
rect 579062 172116 579068 172168
rect 579120 172156 579126 172168
rect 580810 172156 580816 172168
rect 579120 172128 580816 172156
rect 579120 172116 579126 172128
rect 580810 172116 580816 172128
rect 580868 172116 580874 172168
rect 3234 171096 3240 171148
rect 3292 171136 3298 171148
rect 4706 171136 4712 171148
rect 3292 171108 4712 171136
rect 3292 171096 3298 171108
rect 4706 171096 4712 171108
rect 4764 171096 4770 171148
rect 575934 170728 575940 170740
rect 575895 170700 575940 170728
rect 575934 170688 575940 170700
rect 575992 170688 575998 170740
rect 575934 170212 575940 170264
rect 575992 170252 575998 170264
rect 576029 170255 576087 170261
rect 576029 170252 576041 170255
rect 575992 170224 576041 170252
rect 575992 170212 575998 170224
rect 576029 170221 576041 170224
rect 576075 170221 576087 170255
rect 576029 170215 576087 170221
rect 575934 170076 575940 170128
rect 575992 170116 575998 170128
rect 576118 170116 576124 170128
rect 575992 170088 576124 170116
rect 575992 170076 575998 170088
rect 576118 170076 576124 170088
rect 576176 170076 576182 170128
rect 5994 167084 6000 167136
rect 6052 167124 6058 167136
rect 6052 167096 6868 167124
rect 6052 167084 6058 167096
rect 6840 167068 6868 167096
rect 6086 167016 6092 167068
rect 6144 167056 6150 167068
rect 6730 167056 6736 167068
rect 6144 167028 6736 167056
rect 6144 167016 6150 167028
rect 6730 167016 6736 167028
rect 6788 167016 6794 167068
rect 6822 167016 6828 167068
rect 6880 167016 6886 167068
rect 575934 164908 575940 164960
rect 575992 164948 575998 164960
rect 576121 164951 576179 164957
rect 576121 164948 576133 164951
rect 575992 164920 576133 164948
rect 575992 164908 575998 164920
rect 576121 164917 576133 164920
rect 576167 164917 576179 164951
rect 576121 164911 576179 164917
rect 575934 160800 575940 160812
rect 575895 160772 575940 160800
rect 575934 160760 575940 160772
rect 575992 160760 575998 160812
rect 576118 158012 576124 158024
rect 576079 157984 576124 158012
rect 576118 157972 576124 157984
rect 576176 157972 576182 158024
rect 576029 157879 576087 157885
rect 576029 157845 576041 157879
rect 576075 157876 576087 157879
rect 576118 157876 576124 157888
rect 576075 157848 576124 157876
rect 576075 157845 576087 157848
rect 576029 157839 576087 157845
rect 576118 157836 576124 157848
rect 576176 157836 576182 157888
rect 6086 157292 6092 157344
rect 6144 157332 6150 157344
rect 6730 157332 6736 157344
rect 6144 157304 6736 157332
rect 6144 157292 6150 157304
rect 6730 157292 6736 157304
rect 6788 157292 6794 157344
rect 6822 157292 6828 157344
rect 6880 157292 6886 157344
rect 5994 157224 6000 157276
rect 6052 157264 6058 157276
rect 6840 157264 6868 157292
rect 6052 157236 6868 157264
rect 6052 157224 6058 157236
rect 575934 153456 575940 153468
rect 575895 153428 575940 153456
rect 575934 153416 575940 153428
rect 575992 153416 575998 153468
rect 575934 153212 575940 153264
rect 575992 153252 575998 153264
rect 576121 153255 576179 153261
rect 576121 153252 576133 153255
rect 575992 153224 576133 153252
rect 575992 153212 575998 153224
rect 576121 153221 576133 153224
rect 576167 153221 576179 153255
rect 576121 153215 576179 153221
rect 575934 150464 575940 150476
rect 575895 150436 575940 150464
rect 575934 150424 575940 150436
rect 575992 150424 575998 150476
rect 579062 150084 579068 150136
rect 579120 150124 579126 150136
rect 580902 150124 580908 150136
rect 579120 150096 580908 150124
rect 579120 150084 579126 150096
rect 580902 150084 580908 150096
rect 580960 150084 580966 150136
rect 576026 149676 576032 149728
rect 576084 149716 576090 149728
rect 576121 149719 576179 149725
rect 576121 149716 576133 149719
rect 576084 149688 576133 149716
rect 576084 149676 576090 149688
rect 576121 149685 576133 149688
rect 576167 149685 576179 149719
rect 576121 149679 576179 149685
rect 575934 149376 575940 149388
rect 575895 149348 575940 149376
rect 575934 149336 575940 149348
rect 575992 149336 575998 149388
rect 5994 147704 6000 147756
rect 6052 147744 6058 147756
rect 6052 147716 6868 147744
rect 6052 147704 6058 147716
rect 6840 147688 6868 147716
rect 6086 147636 6092 147688
rect 6144 147676 6150 147688
rect 6730 147676 6736 147688
rect 6144 147648 6736 147676
rect 6144 147636 6150 147648
rect 6730 147636 6736 147648
rect 6788 147636 6794 147688
rect 6822 147636 6828 147688
rect 6880 147636 6886 147688
rect 575934 145936 575940 145988
rect 575992 145976 575998 145988
rect 576213 145979 576271 145985
rect 576213 145976 576225 145979
rect 575992 145948 576225 145976
rect 575992 145936 575998 145948
rect 576213 145945 576225 145948
rect 576259 145945 576271 145979
rect 576213 145939 576271 145945
rect 575934 145256 575940 145308
rect 575992 145296 575998 145308
rect 576029 145299 576087 145305
rect 576029 145296 576041 145299
rect 575992 145268 576041 145296
rect 575992 145256 575998 145268
rect 576029 145265 576041 145268
rect 576075 145265 576087 145299
rect 576029 145259 576087 145265
rect 575934 144848 575940 144900
rect 575992 144888 575998 144900
rect 576213 144891 576271 144897
rect 576213 144888 576225 144891
rect 575992 144860 576225 144888
rect 575992 144848 575998 144860
rect 576213 144857 576225 144860
rect 576259 144857 576271 144891
rect 576213 144851 576271 144857
rect 576026 144508 576032 144560
rect 576084 144548 576090 144560
rect 576302 144548 576308 144560
rect 576084 144520 576308 144548
rect 576084 144508 576090 144520
rect 576302 144508 576308 144520
rect 576360 144508 576366 144560
rect 575934 144412 575940 144424
rect 575895 144384 575940 144412
rect 575934 144372 575940 144384
rect 575992 144372 575998 144424
rect 575934 140944 575940 140956
rect 575895 140916 575940 140944
rect 575934 140904 575940 140916
rect 575992 140904 575998 140956
rect 575934 140292 575940 140344
rect 575992 140332 575998 140344
rect 576029 140335 576087 140341
rect 576029 140332 576041 140335
rect 575992 140304 576041 140332
rect 575992 140292 575998 140304
rect 576029 140301 576041 140304
rect 576075 140301 576087 140335
rect 576029 140295 576087 140301
rect 575934 139884 575940 139936
rect 575992 139924 575998 139936
rect 576118 139924 576124 139936
rect 575992 139896 576124 139924
rect 575992 139884 575998 139896
rect 576118 139884 576124 139896
rect 576176 139884 576182 139936
rect 6086 137912 6092 137964
rect 6144 137952 6150 137964
rect 6730 137952 6736 137964
rect 6144 137924 6736 137952
rect 6144 137912 6150 137924
rect 6730 137912 6736 137924
rect 6788 137912 6794 137964
rect 6822 137912 6828 137964
rect 6880 137912 6886 137964
rect 5994 137844 6000 137896
rect 6052 137884 6058 137896
rect 6840 137884 6868 137912
rect 6052 137856 6868 137884
rect 6052 137844 6058 137856
rect 575934 137164 575940 137216
rect 575992 137204 575998 137216
rect 576121 137207 576179 137213
rect 576121 137204 576133 137207
rect 575992 137176 576133 137204
rect 575992 137164 575998 137176
rect 576121 137173 576133 137176
rect 576167 137173 576179 137207
rect 576121 137167 576179 137173
rect 576026 137068 576032 137080
rect 575952 137040 576032 137068
rect 575952 137012 575980 137040
rect 576026 137028 576032 137040
rect 576084 137028 576090 137080
rect 575934 136960 575940 137012
rect 575992 136960 575998 137012
rect 575934 132580 575940 132592
rect 575895 132552 575940 132580
rect 575934 132540 575940 132552
rect 575992 132540 575998 132592
rect 575934 132104 575940 132116
rect 575895 132076 575940 132104
rect 575934 132064 575940 132076
rect 575992 132064 575998 132116
rect 575934 130500 575940 130552
rect 575992 130540 575998 130552
rect 576213 130543 576271 130549
rect 576213 130540 576225 130543
rect 575992 130512 576225 130540
rect 575992 130500 575998 130512
rect 576213 130509 576225 130512
rect 576259 130509 576271 130543
rect 576213 130503 576271 130509
rect 5994 128392 6000 128444
rect 6052 128432 6058 128444
rect 6052 128404 6868 128432
rect 6052 128392 6058 128404
rect 6840 128376 6868 128404
rect 6086 128324 6092 128376
rect 6144 128364 6150 128376
rect 6730 128364 6736 128376
rect 6144 128336 6736 128364
rect 6144 128324 6150 128336
rect 6730 128324 6736 128336
rect 6788 128324 6794 128376
rect 6822 128324 6828 128376
rect 6880 128324 6886 128376
rect 3326 128256 3332 128308
rect 3384 128296 3390 128308
rect 4154 128296 4160 128308
rect 3384 128268 4160 128296
rect 3384 128256 3390 128268
rect 4154 128256 4160 128268
rect 4212 128256 4218 128308
rect 579062 127916 579068 127968
rect 579120 127956 579126 127968
rect 580166 127956 580172 127968
rect 579120 127928 580172 127956
rect 579120 127916 579126 127928
rect 580166 127916 580172 127928
rect 580224 127916 580230 127968
rect 575934 127644 575940 127696
rect 575992 127684 575998 127696
rect 576121 127687 576179 127693
rect 576121 127684 576133 127687
rect 575992 127656 576133 127684
rect 575992 127644 575998 127656
rect 576121 127653 576133 127656
rect 576167 127653 576179 127687
rect 576121 127647 576179 127653
rect 576121 125579 576179 125585
rect 576121 125545 576133 125579
rect 576167 125576 576179 125579
rect 576305 125579 576363 125585
rect 576305 125576 576317 125579
rect 576167 125548 576317 125576
rect 576167 125545 576179 125548
rect 576121 125539 576179 125545
rect 576305 125545 576317 125548
rect 576351 125545 576363 125579
rect 576305 125539 576363 125545
rect 575934 122544 575940 122596
rect 575992 122584 575998 122596
rect 576029 122587 576087 122593
rect 576029 122584 576041 122587
rect 575992 122556 576041 122584
rect 575992 122544 575998 122556
rect 576029 122553 576041 122556
rect 576075 122553 576087 122587
rect 576029 122547 576087 122553
rect 575934 121592 575940 121644
rect 575992 121632 575998 121644
rect 576118 121632 576124 121644
rect 575992 121604 576124 121632
rect 575992 121592 575998 121604
rect 576118 121592 576124 121604
rect 576176 121592 576182 121644
rect 576213 120751 576271 120757
rect 576213 120717 576225 120751
rect 576259 120748 576271 120751
rect 576302 120748 576308 120760
rect 576259 120720 576308 120748
rect 576259 120717 576271 120720
rect 576213 120711 576271 120717
rect 576302 120708 576308 120720
rect 576360 120708 576366 120760
rect 6086 118600 6092 118652
rect 6144 118640 6150 118652
rect 6730 118640 6736 118652
rect 6144 118612 6736 118640
rect 6144 118600 6150 118612
rect 6730 118600 6736 118612
rect 6788 118600 6794 118652
rect 6822 118600 6828 118652
rect 6880 118600 6886 118652
rect 5994 118532 6000 118584
rect 6052 118572 6058 118584
rect 6840 118572 6868 118600
rect 6052 118544 6868 118572
rect 575937 118575 575995 118581
rect 6052 118532 6058 118544
rect 575937 118541 575949 118575
rect 575983 118572 575995 118575
rect 576118 118572 576124 118584
rect 575983 118544 576124 118572
rect 575983 118541 575995 118544
rect 575937 118535 575995 118541
rect 576118 118532 576124 118544
rect 576176 118532 576182 118584
rect 575937 118439 575995 118445
rect 575937 118405 575949 118439
rect 575983 118436 575995 118439
rect 576305 118439 576363 118445
rect 576305 118436 576317 118439
rect 575983 118408 576317 118436
rect 575983 118405 575995 118408
rect 575937 118399 575995 118405
rect 576305 118405 576317 118408
rect 576351 118405 576363 118439
rect 576305 118399 576363 118405
rect 575934 117716 575940 117768
rect 575992 117756 575998 117768
rect 576029 117759 576087 117765
rect 576029 117756 576041 117759
rect 575992 117728 576041 117756
rect 575992 117716 575998 117728
rect 576029 117725 576041 117728
rect 576075 117725 576087 117759
rect 576029 117719 576087 117725
rect 576026 115880 576032 115932
rect 576084 115880 576090 115932
rect 576044 115852 576072 115880
rect 576121 115855 576179 115861
rect 576121 115852 576133 115855
rect 576044 115824 576133 115852
rect 576121 115821 576133 115824
rect 576167 115821 576179 115855
rect 576121 115815 576179 115821
rect 575934 113976 575940 114028
rect 575992 114016 575998 114028
rect 576029 114019 576087 114025
rect 576029 114016 576041 114019
rect 575992 113988 576041 114016
rect 575992 113976 575998 113988
rect 576029 113985 576041 113988
rect 576075 113985 576087 114019
rect 576029 113979 576087 113985
rect 575934 110916 575940 110968
rect 575992 110956 575998 110968
rect 576121 110959 576179 110965
rect 576121 110956 576133 110959
rect 575992 110928 576133 110956
rect 575992 110916 575998 110928
rect 576121 110925 576133 110928
rect 576167 110925 576179 110959
rect 576121 110919 576179 110925
rect 5994 109080 6000 109132
rect 6052 109120 6058 109132
rect 6052 109092 6868 109120
rect 6052 109080 6058 109092
rect 6840 109064 6868 109092
rect 6086 109012 6092 109064
rect 6144 109052 6150 109064
rect 6730 109052 6736 109064
rect 6144 109024 6736 109052
rect 6144 109012 6150 109024
rect 6730 109012 6736 109024
rect 6788 109012 6794 109064
rect 6822 109012 6828 109064
rect 6880 109012 6886 109064
rect 576118 108848 576124 108860
rect 576079 108820 576124 108848
rect 576118 108808 576124 108820
rect 576176 108808 576182 108860
rect 579062 106156 579068 106208
rect 579120 106196 579126 106208
rect 580626 106196 580632 106208
rect 579120 106168 580632 106196
rect 579120 106156 579126 106168
rect 580626 106156 580632 106168
rect 580684 106156 580690 106208
rect 575934 104428 575940 104440
rect 575895 104400 575940 104428
rect 575934 104388 575940 104400
rect 575992 104388 575998 104440
rect 575934 104252 575940 104304
rect 575992 104292 575998 104304
rect 576029 104295 576087 104301
rect 576029 104292 576041 104295
rect 575992 104264 576041 104292
rect 575992 104252 575998 104264
rect 576029 104261 576041 104264
rect 576075 104261 576087 104295
rect 576029 104255 576087 104261
rect 575934 104116 575940 104168
rect 575992 104156 575998 104168
rect 576394 104156 576400 104168
rect 575992 104128 576400 104156
rect 575992 104116 575998 104128
rect 576394 104116 576400 104128
rect 576452 104116 576458 104168
rect 575934 102416 575940 102468
rect 575992 102456 575998 102468
rect 576121 102459 576179 102465
rect 576121 102456 576133 102459
rect 575992 102428 576133 102456
rect 575992 102416 575998 102428
rect 576121 102425 576133 102428
rect 576167 102425 576179 102459
rect 576121 102419 576179 102425
rect 575934 100444 575940 100496
rect 575992 100444 575998 100496
rect 575952 100360 575980 100444
rect 575934 100308 575940 100360
rect 575992 100308 575998 100360
rect 6086 99288 6092 99340
rect 6144 99328 6150 99340
rect 6730 99328 6736 99340
rect 6144 99300 6736 99328
rect 6144 99288 6150 99300
rect 6730 99288 6736 99300
rect 6788 99288 6794 99340
rect 6822 99288 6828 99340
rect 6880 99288 6886 99340
rect 5994 99220 6000 99272
rect 6052 99260 6058 99272
rect 6840 99260 6868 99288
rect 6052 99232 6868 99260
rect 6052 99220 6058 99232
rect 575934 93780 575940 93832
rect 575992 93820 575998 93832
rect 576213 93823 576271 93829
rect 576213 93820 576225 93823
rect 575992 93792 576225 93820
rect 575992 93780 575998 93792
rect 576213 93789 576225 93792
rect 576259 93789 576271 93823
rect 576213 93783 576271 93789
rect 575934 90584 575940 90636
rect 575992 90624 575998 90636
rect 576121 90627 576179 90633
rect 576121 90624 576133 90627
rect 575992 90596 576133 90624
rect 575992 90584 575998 90596
rect 576121 90593 576133 90596
rect 576167 90593 576179 90627
rect 576121 90587 576179 90593
rect 5994 89768 6000 89820
rect 6052 89808 6058 89820
rect 6052 89780 6868 89808
rect 6052 89768 6058 89780
rect 6840 89752 6868 89780
rect 6086 89700 6092 89752
rect 6144 89740 6150 89752
rect 6730 89740 6736 89752
rect 6144 89712 6736 89740
rect 6144 89700 6150 89712
rect 6730 89700 6736 89712
rect 6788 89700 6794 89752
rect 6822 89700 6828 89752
rect 6880 89700 6886 89752
rect 576302 85620 576308 85672
rect 576360 85620 576366 85672
rect 576320 85536 576348 85620
rect 576302 85484 576308 85536
rect 576360 85484 576366 85536
rect 579062 84124 579068 84176
rect 579120 84164 579126 84176
rect 580718 84164 580724 84176
rect 579120 84136 580724 84164
rect 579120 84124 579126 84136
rect 580718 84124 580724 84136
rect 580776 84124 580782 84176
rect 575934 81376 575940 81388
rect 575895 81348 575940 81376
rect 575934 81336 575940 81348
rect 575992 81336 575998 81388
rect 576118 81376 576124 81388
rect 576079 81348 576124 81376
rect 576118 81336 576124 81348
rect 576176 81336 576182 81388
rect 6086 79976 6092 80028
rect 6144 80016 6150 80028
rect 6730 80016 6736 80028
rect 6144 79988 6736 80016
rect 6144 79976 6150 79988
rect 6730 79976 6736 79988
rect 6788 79976 6794 80028
rect 6822 79976 6828 80028
rect 6880 79976 6886 80028
rect 5994 79908 6000 79960
rect 6052 79948 6058 79960
rect 6840 79948 6868 79976
rect 6052 79920 6868 79948
rect 6052 79908 6058 79920
rect 575934 79432 575940 79484
rect 575992 79472 575998 79484
rect 576029 79475 576087 79481
rect 576029 79472 576041 79475
rect 575992 79444 576041 79472
rect 575992 79432 575998 79444
rect 576029 79441 576041 79444
rect 576075 79441 576087 79475
rect 576029 79435 576087 79441
rect 576026 74780 576032 74792
rect 575987 74752 576032 74780
rect 576026 74740 576032 74752
rect 576084 74740 576090 74792
rect 575934 72196 575940 72208
rect 575895 72168 575940 72196
rect 575934 72156 575940 72168
rect 575992 72156 575998 72208
rect 5994 70456 6000 70508
rect 6052 70496 6058 70508
rect 6052 70468 6868 70496
rect 6052 70456 6058 70468
rect 6840 70440 6868 70468
rect 6086 70388 6092 70440
rect 6144 70428 6150 70440
rect 6730 70428 6736 70440
rect 6144 70400 6736 70428
rect 6144 70388 6150 70400
rect 6730 70388 6736 70400
rect 6788 70388 6794 70440
rect 6822 70388 6828 70440
rect 6880 70388 6886 70440
rect 575934 70320 575940 70372
rect 575992 70360 575998 70372
rect 576213 70363 576271 70369
rect 576213 70360 576225 70363
rect 575992 70332 576225 70360
rect 575992 70320 575998 70332
rect 576213 70329 576225 70332
rect 576259 70329 576271 70363
rect 576213 70323 576271 70329
rect 576026 67572 576032 67584
rect 575987 67544 576032 67572
rect 576026 67532 576032 67544
rect 576084 67532 576090 67584
rect 575934 63356 575940 63368
rect 575895 63328 575940 63356
rect 575934 63316 575940 63328
rect 575992 63316 575998 63368
rect 579062 61956 579068 62008
rect 579120 61996 579126 62008
rect 580810 61996 580816 62008
rect 579120 61968 580816 61996
rect 579120 61956 579126 61968
rect 580810 61956 580816 61968
rect 580868 61956 580874 62008
rect 576118 61548 576124 61600
rect 576176 61588 576182 61600
rect 576394 61588 576400 61600
rect 576176 61560 576400 61588
rect 576176 61548 576182 61560
rect 576394 61548 576400 61560
rect 576452 61548 576458 61600
rect 6086 60664 6092 60716
rect 6144 60704 6150 60716
rect 6730 60704 6736 60716
rect 6144 60676 6736 60704
rect 6144 60664 6150 60676
rect 6730 60664 6736 60676
rect 6788 60664 6794 60716
rect 6822 60664 6828 60716
rect 6880 60664 6886 60716
rect 5994 60596 6000 60648
rect 6052 60636 6058 60648
rect 6840 60636 6868 60664
rect 6052 60608 6868 60636
rect 6052 60596 6058 60608
rect 575934 58760 575940 58812
rect 575992 58800 575998 58812
rect 576305 58803 576363 58809
rect 576305 58800 576317 58803
rect 575992 58772 576317 58800
rect 575992 58760 575998 58772
rect 576305 58769 576317 58772
rect 576351 58769 576363 58803
rect 576305 58763 576363 58769
rect 576210 57944 576216 57996
rect 576268 57984 576274 57996
rect 576302 57984 576308 57996
rect 576268 57956 576308 57984
rect 576268 57944 576274 57956
rect 576302 57944 576308 57956
rect 576360 57944 576366 57996
rect 575937 57851 575995 57857
rect 575937 57817 575949 57851
rect 575983 57848 575995 57851
rect 576118 57848 576124 57860
rect 575983 57820 576124 57848
rect 575983 57817 575995 57820
rect 575937 57811 575995 57817
rect 576118 57808 576124 57820
rect 576176 57808 576182 57860
rect 576302 57304 576308 57316
rect 576263 57276 576308 57304
rect 576302 57264 576308 57276
rect 576360 57264 576366 57316
rect 575934 52776 575940 52828
rect 575992 52776 575998 52828
rect 575952 52624 575980 52776
rect 575934 52572 575940 52624
rect 575992 52572 575998 52624
rect 576029 51799 576087 51805
rect 576029 51765 576041 51799
rect 576075 51796 576087 51799
rect 576118 51796 576124 51808
rect 576075 51768 576124 51796
rect 576075 51765 576087 51768
rect 576029 51759 576087 51765
rect 576118 51756 576124 51768
rect 576176 51756 576182 51808
rect 5994 51144 6000 51196
rect 6052 51184 6058 51196
rect 6052 51156 6868 51184
rect 6052 51144 6058 51156
rect 6840 51128 6868 51156
rect 6086 51076 6092 51128
rect 6144 51116 6150 51128
rect 6730 51116 6736 51128
rect 6144 51088 6736 51116
rect 6144 51076 6150 51088
rect 6730 51076 6736 51088
rect 6788 51076 6794 51128
rect 6822 51076 6828 51128
rect 6880 51076 6886 51128
rect 575934 46384 575940 46436
rect 575992 46384 575998 46436
rect 575952 46220 575980 46384
rect 576026 46220 576032 46232
rect 575952 46192 576032 46220
rect 576026 46180 576032 46192
rect 576084 46180 576090 46232
rect 575934 43596 575940 43648
rect 575992 43636 575998 43648
rect 576121 43639 576179 43645
rect 576121 43636 576133 43639
rect 575992 43608 576133 43636
rect 575992 43596 575998 43608
rect 576121 43605 576133 43608
rect 576167 43605 576179 43639
rect 576121 43599 576179 43605
rect 575934 43500 575940 43512
rect 575895 43472 575940 43500
rect 575934 43460 575940 43472
rect 575992 43460 575998 43512
rect 6086 41352 6092 41404
rect 6144 41392 6150 41404
rect 6730 41392 6736 41404
rect 6144 41364 6736 41392
rect 6144 41352 6150 41364
rect 6730 41352 6736 41364
rect 6788 41352 6794 41404
rect 6822 41352 6828 41404
rect 6880 41352 6886 41404
rect 5994 41284 6000 41336
rect 6052 41324 6058 41336
rect 6840 41324 6868 41352
rect 6052 41296 6868 41324
rect 6052 41284 6058 41296
rect 579062 39924 579068 39976
rect 579120 39964 579126 39976
rect 580626 39964 580632 39976
rect 579120 39936 580632 39964
rect 579120 39924 579126 39936
rect 580626 39924 580632 39936
rect 580684 39924 580690 39976
rect 575934 39380 575940 39432
rect 575992 39420 575998 39432
rect 576029 39423 576087 39429
rect 576029 39420 576041 39423
rect 575992 39392 576041 39420
rect 575992 39380 575998 39392
rect 576029 39389 576041 39392
rect 576075 39389 576087 39423
rect 576029 39383 576087 39389
rect 575934 37244 575940 37256
rect 575895 37216 575940 37244
rect 575934 37204 575940 37216
rect 575992 37204 575998 37256
rect 575934 35300 575940 35352
rect 575992 35340 575998 35352
rect 576029 35343 576087 35349
rect 576029 35340 576041 35343
rect 575992 35312 576041 35340
rect 575992 35300 575998 35312
rect 576029 35309 576041 35312
rect 576075 35309 576087 35343
rect 576029 35303 576087 35309
rect 575934 35164 575940 35216
rect 575992 35204 575998 35216
rect 576121 35207 576179 35213
rect 576121 35204 576133 35207
rect 575992 35176 576133 35204
rect 575992 35164 575998 35176
rect 576121 35173 576133 35176
rect 576167 35173 576179 35207
rect 576121 35167 576179 35173
rect 575934 33804 575940 33856
rect 575992 33844 575998 33856
rect 576029 33847 576087 33853
rect 576029 33844 576041 33847
rect 575992 33816 576041 33844
rect 575992 33804 575998 33816
rect 576029 33813 576041 33816
rect 576075 33813 576087 33847
rect 576029 33807 576087 33813
rect 576118 33804 576124 33856
rect 576176 33844 576182 33856
rect 576394 33844 576400 33856
rect 576176 33816 576400 33844
rect 576176 33804 576182 33816
rect 576394 33804 576400 33816
rect 576452 33804 576458 33856
rect 575934 33056 575940 33108
rect 575992 33096 575998 33108
rect 576029 33099 576087 33105
rect 576029 33096 576041 33099
rect 575992 33068 576041 33096
rect 575992 33056 575998 33068
rect 576029 33065 576041 33068
rect 576075 33065 576087 33099
rect 576029 33059 576087 33065
rect 5994 31832 6000 31884
rect 6052 31872 6058 31884
rect 6052 31844 6868 31872
rect 6052 31832 6058 31844
rect 6840 31816 6868 31844
rect 6086 31764 6092 31816
rect 6144 31804 6150 31816
rect 6730 31804 6736 31816
rect 6144 31776 6736 31804
rect 6144 31764 6150 31776
rect 6730 31764 6736 31776
rect 6788 31764 6794 31816
rect 6822 31764 6828 31816
rect 6880 31764 6886 31816
rect 576026 28636 576032 28688
rect 576084 28676 576090 28688
rect 576302 28676 576308 28688
rect 576084 28648 576308 28676
rect 576084 28636 576090 28648
rect 576302 28636 576308 28648
rect 576360 28636 576366 28688
rect 575934 28296 575940 28348
rect 575992 28336 575998 28348
rect 576029 28339 576087 28345
rect 576029 28336 576041 28339
rect 575992 28308 576041 28336
rect 575992 28296 575998 28308
rect 576029 28305 576041 28308
rect 576075 28305 576087 28339
rect 576029 28299 576087 28305
rect 576029 24191 576087 24197
rect 576029 24157 576041 24191
rect 576075 24188 576087 24191
rect 576210 24188 576216 24200
rect 576075 24160 576216 24188
rect 576075 24157 576087 24160
rect 576029 24151 576087 24157
rect 576210 24148 576216 24160
rect 576268 24148 576274 24200
rect 6086 22040 6092 22092
rect 6144 22080 6150 22092
rect 6730 22080 6736 22092
rect 6144 22052 6736 22080
rect 6144 22040 6150 22052
rect 6730 22040 6736 22052
rect 6788 22040 6794 22092
rect 6822 22040 6828 22092
rect 6880 22040 6886 22092
rect 5994 21972 6000 22024
rect 6052 22012 6058 22024
rect 6840 22012 6868 22040
rect 6052 21984 6868 22012
rect 6052 21972 6058 21984
rect 576118 21536 576124 21548
rect 576079 21508 576124 21536
rect 576118 21496 576124 21508
rect 576176 21496 576182 21548
rect 576026 21360 576032 21412
rect 576084 21400 576090 21412
rect 576302 21400 576308 21412
rect 576084 21372 576308 21400
rect 576084 21360 576090 21372
rect 576302 21360 576308 21372
rect 576360 21360 576366 21412
rect 575934 20544 575940 20596
rect 575992 20584 575998 20596
rect 576118 20584 576124 20596
rect 575992 20556 576124 20584
rect 575992 20544 575998 20556
rect 576118 20544 576124 20556
rect 576176 20544 576182 20596
rect 575934 20312 575940 20324
rect 575895 20284 575940 20312
rect 575934 20272 575940 20284
rect 575992 20272 575998 20324
rect 576026 19360 576032 19372
rect 575987 19332 576032 19360
rect 576026 19320 576032 19332
rect 576084 19320 576090 19372
rect 575934 17212 575940 17264
rect 575992 17252 575998 17264
rect 576302 17252 576308 17264
rect 575992 17224 576308 17252
rect 575992 17212 575998 17224
rect 576302 17212 576308 17224
rect 576360 17212 576366 17264
rect 575934 16668 575940 16720
rect 575992 16708 575998 16720
rect 576121 16711 576179 16717
rect 576121 16708 576133 16711
rect 575992 16680 576133 16708
rect 575992 16668 575998 16680
rect 576121 16677 576133 16680
rect 576167 16677 576179 16711
rect 576121 16671 576179 16677
rect 5994 12520 6000 12572
rect 6052 12560 6058 12572
rect 6052 12532 6868 12560
rect 6052 12520 6058 12532
rect 6840 12504 6868 12532
rect 6086 12452 6092 12504
rect 6144 12492 6150 12504
rect 6730 12492 6736 12504
rect 6144 12464 6736 12492
rect 6144 12452 6150 12464
rect 6730 12452 6736 12464
rect 6788 12452 6794 12504
rect 6822 12452 6828 12504
rect 6880 12452 6886 12504
rect 4798 11976 4804 12028
rect 4856 11976 4862 12028
rect 4816 11824 4844 11976
rect 4798 11772 4804 11824
rect 4856 11772 4862 11824
rect 69477 7803 69535 7809
rect 69477 7769 69489 7803
rect 69523 7800 69535 7803
rect 576118 7800 576124 7812
rect 69523 7772 576124 7800
rect 69523 7769 69535 7772
rect 69477 7763 69535 7769
rect 576118 7760 576124 7772
rect 576176 7760 576182 7812
rect 9398 7692 9404 7744
rect 9456 7732 9462 7744
rect 17218 7732 17224 7744
rect 9456 7704 17224 7732
rect 9456 7692 9462 7704
rect 17218 7692 17224 7704
rect 17276 7692 17282 7744
rect 58802 7692 58808 7744
rect 58860 7732 58866 7744
rect 576210 7732 576216 7744
rect 58860 7704 576216 7732
rect 58860 7692 58866 7704
rect 576210 7692 576216 7704
rect 576268 7692 576274 7744
rect 1670 7624 1676 7676
rect 1728 7664 1734 7676
rect 576302 7664 576308 7676
rect 1728 7636 576308 7664
rect 1728 7624 1734 7636
rect 576302 7624 576308 7636
rect 576360 7624 576366 7676
rect 566 7556 572 7608
rect 624 7596 630 7608
rect 575750 7596 575756 7608
rect 624 7568 575756 7596
rect 624 7556 630 7568
rect 575750 7556 575756 7568
rect 575808 7556 575814 7608
rect 69474 7528 69480 7540
rect 69435 7500 69480 7528
rect 69474 7488 69480 7500
rect 69532 7488 69538 7540
rect 575106 7488 575112 7540
rect 575164 7528 575170 7540
rect 575934 7528 575940 7540
rect 575164 7500 575940 7528
rect 575164 7488 575170 7500
rect 575934 7488 575940 7500
rect 575992 7488 575998 7540
rect 575014 7420 575020 7472
rect 575072 7460 575078 7472
rect 575474 7460 575480 7472
rect 575072 7432 575480 7460
rect 575072 7420 575078 7432
rect 575474 7420 575480 7432
rect 575532 7420 575538 7472
rect 52730 6808 52736 6860
rect 52788 6848 52794 6860
rect 580534 6848 580540 6860
rect 52788 6820 580540 6848
rect 52788 6808 52794 6820
rect 580534 6808 580540 6820
rect 580592 6808 580598 6860
rect 62942 6740 62948 6792
rect 63000 6780 63006 6792
rect 580442 6780 580448 6792
rect 63000 6752 580448 6780
rect 63000 6740 63006 6752
rect 580442 6740 580448 6752
rect 580500 6740 580506 6792
rect 73062 6672 73068 6724
rect 73120 6712 73126 6724
rect 580350 6712 580356 6724
rect 73120 6684 580356 6712
rect 73120 6672 73126 6684
rect 580350 6672 580356 6684
rect 580408 6672 580414 6724
rect 83274 6604 83280 6656
rect 83332 6644 83338 6656
rect 580258 6644 580264 6656
rect 83332 6616 580264 6644
rect 83332 6604 83338 6616
rect 580258 6604 580264 6616
rect 580316 6604 580322 6656
rect 90910 6536 90916 6588
rect 90968 6576 90974 6588
rect 577038 6576 577044 6588
rect 90968 6548 577044 6576
rect 90968 6536 90974 6548
rect 577038 6536 577044 6548
rect 577096 6536 577102 6588
rect 83826 6468 83832 6520
rect 83884 6508 83890 6520
rect 577130 6508 577136 6520
rect 83884 6480 577136 6508
rect 83884 6468 83890 6480
rect 577130 6468 577136 6480
rect 577188 6468 577194 6520
rect 77846 6400 77852 6452
rect 77904 6440 77910 6452
rect 578510 6440 578516 6452
rect 77904 6412 578516 6440
rect 77904 6400 77910 6412
rect 578510 6400 578516 6412
rect 578568 6400 578574 6452
rect 6454 6332 6460 6384
rect 6512 6372 6518 6384
rect 65978 6372 65984 6384
rect 6512 6344 65984 6372
rect 6512 6332 6518 6344
rect 65978 6332 65984 6344
rect 66036 6332 66042 6384
rect 73062 6332 73068 6384
rect 73120 6372 73126 6384
rect 577222 6372 577228 6384
rect 73120 6344 577228 6372
rect 73120 6332 73126 6344
rect 577222 6332 577228 6344
rect 577280 6332 577286 6384
rect 63586 6264 63592 6316
rect 63644 6304 63650 6316
rect 578602 6304 578608 6316
rect 63644 6276 578608 6304
rect 63644 6264 63650 6276
rect 578602 6264 578608 6276
rect 578660 6264 578666 6316
rect 30282 6196 30288 6248
rect 30340 6236 30346 6248
rect 578878 6236 578884 6248
rect 30340 6208 578884 6236
rect 30340 6196 30346 6208
rect 578878 6196 578884 6208
rect 578936 6196 578942 6248
rect 21910 6128 21916 6180
rect 21968 6168 21974 6180
rect 578970 6168 578976 6180
rect 21968 6140 578976 6168
rect 21968 6128 21974 6140
rect 578970 6128 578976 6140
rect 579028 6128 579034 6180
rect 94498 6060 94504 6112
rect 94556 6100 94562 6112
rect 576946 6100 576952 6112
rect 94556 6072 576952 6100
rect 94556 6060 94562 6072
rect 576946 6060 576952 6072
rect 577004 6060 577010 6112
rect 101582 5992 101588 6044
rect 101640 6032 101646 6044
rect 576854 6032 576860 6044
rect 101640 6004 576860 6032
rect 101640 5992 101646 6004
rect 576854 5992 576860 6004
rect 576912 5992 576918 6044
rect 106366 5924 106372 5976
rect 106424 5964 106430 5976
rect 578418 5964 578424 5976
rect 106424 5936 578424 5964
rect 106424 5924 106430 5936
rect 578418 5924 578424 5936
rect 578476 5924 578482 5976
rect 7098 5856 7104 5908
rect 7156 5896 7162 5908
rect 115934 5896 115940 5908
rect 7156 5868 115940 5896
rect 7156 5856 7162 5868
rect 115934 5856 115940 5868
rect 115992 5856 115998 5908
rect 119430 5856 119436 5908
rect 119488 5896 119494 5908
rect 578786 5896 578792 5908
rect 119488 5868 578792 5896
rect 119488 5856 119494 5868
rect 578786 5856 578792 5868
rect 578844 5856 578850 5908
rect 9306 5788 9312 5840
rect 9364 5828 9370 5840
rect 123018 5828 123024 5840
rect 9364 5800 123024 5828
rect 9364 5788 9370 5800
rect 123018 5788 123024 5800
rect 123076 5788 123082 5840
rect 7190 5720 7196 5772
rect 7248 5760 7254 5772
rect 108758 5760 108764 5772
rect 7248 5732 108764 5760
rect 7248 5720 7254 5732
rect 108758 5720 108764 5732
rect 108816 5720 108822 5772
rect 6178 5448 6184 5500
rect 6236 5488 6242 5500
rect 12066 5488 12072 5500
rect 6236 5460 12072 5488
rect 6236 5448 6242 5460
rect 12066 5448 12072 5460
rect 12124 5448 12130 5500
rect 96890 5448 96896 5500
rect 96948 5488 96954 5500
rect 327534 5488 327540 5500
rect 96948 5460 327540 5488
rect 96948 5448 96954 5460
rect 327534 5448 327540 5460
rect 327592 5448 327598 5500
rect 7558 5380 7564 5432
rect 7616 5420 7622 5432
rect 32398 5420 32404 5432
rect 7616 5392 32404 5420
rect 7616 5380 7622 5392
rect 32398 5380 32404 5392
rect 32456 5380 32462 5432
rect 103974 5380 103980 5432
rect 104032 5420 104038 5432
rect 347958 5420 347964 5432
rect 104032 5392 347964 5420
rect 104032 5380 104038 5392
rect 347958 5380 347964 5392
rect 348016 5380 348022 5432
rect 14182 5312 14188 5364
rect 14240 5352 14246 5364
rect 99374 5352 99380 5364
rect 14240 5324 99380 5352
rect 14240 5312 14246 5324
rect 99374 5312 99380 5324
rect 99432 5312 99438 5364
rect 111150 5312 111156 5364
rect 111208 5352 111214 5364
rect 368290 5352 368296 5364
rect 111208 5324 368296 5352
rect 111208 5312 111214 5324
rect 368290 5312 368296 5324
rect 368348 5312 368354 5364
rect 15194 5244 15200 5296
rect 15252 5284 15258 5296
rect 104250 5284 104256 5296
rect 15252 5256 104256 5284
rect 15252 5244 15258 5256
rect 104250 5244 104256 5256
rect 104308 5244 104314 5296
rect 118234 5244 118240 5296
rect 118292 5284 118298 5296
rect 388622 5284 388628 5296
rect 118292 5256 388628 5284
rect 118292 5244 118298 5256
rect 388622 5244 388628 5256
rect 388680 5244 388686 5296
rect 19518 5176 19524 5228
rect 19576 5216 19582 5228
rect 113818 5216 113824 5228
rect 19576 5188 113824 5216
rect 19576 5176 19582 5188
rect 113818 5176 113824 5188
rect 113876 5176 113882 5228
rect 125410 5176 125416 5228
rect 125468 5216 125474 5228
rect 409046 5216 409052 5228
rect 125468 5188 409052 5216
rect 125468 5176 125474 5188
rect 409046 5176 409052 5188
rect 409104 5176 409110 5228
rect 3418 5108 3424 5160
rect 3476 5148 3482 5160
rect 42518 5148 42524 5160
rect 3476 5120 42524 5148
rect 3476 5108 3482 5120
rect 42518 5108 42524 5120
rect 42576 5108 42582 5160
rect 51626 5108 51632 5160
rect 51684 5148 51690 5160
rect 439590 5148 439596 5160
rect 51684 5120 439596 5148
rect 51684 5108 51690 5120
rect 439590 5108 439596 5120
rect 439648 5108 439654 5160
rect 55214 5040 55220 5092
rect 55272 5080 55278 5092
rect 449710 5080 449716 5092
rect 55272 5052 449716 5080
rect 55272 5040 55278 5052
rect 449710 5040 449716 5052
rect 449768 5040 449774 5092
rect 7374 4972 7380 5024
rect 7432 5012 7438 5024
rect 26694 5012 26700 5024
rect 7432 4984 26700 5012
rect 7432 4972 7438 4984
rect 26694 4972 26700 4984
rect 26752 4972 26758 5024
rect 62390 4972 62396 5024
rect 62448 5012 62454 5024
rect 459922 5012 459928 5024
rect 62448 4984 459928 5012
rect 62448 4972 62454 4984
rect 459922 4972 459928 4984
rect 459980 4972 459986 5024
rect 7282 4904 7288 4956
rect 7340 4944 7346 4956
rect 33870 4944 33876 4956
rect 7340 4916 33876 4944
rect 7340 4904 7346 4916
rect 33870 4904 33876 4916
rect 33928 4904 33934 4956
rect 80238 4904 80244 4956
rect 80296 4944 80302 4956
rect 480254 4944 480260 4956
rect 80296 4916 480260 4944
rect 80296 4904 80302 4916
rect 480254 4904 480260 4916
rect 480312 4904 480318 4956
rect 6914 4836 6920 4888
rect 6972 4876 6978 4888
rect 67174 4876 67180 4888
rect 6972 4848 67180 4876
rect 6972 4836 6978 4848
rect 67174 4836 67180 4848
rect 67232 4836 67238 4888
rect 98086 4836 98092 4888
rect 98144 4876 98150 4888
rect 500586 4876 500592 4888
rect 98144 4848 500592 4876
rect 98144 4836 98150 4848
rect 500586 4836 500592 4848
rect 500644 4836 500650 4888
rect 6362 4768 6368 4820
rect 6420 4808 6426 4820
rect 40954 4808 40960 4820
rect 6420 4780 40960 4808
rect 6420 4768 6426 4780
rect 40954 4768 40960 4780
rect 41012 4768 41018 4820
rect 52822 4768 52828 4820
rect 52880 4808 52886 4820
rect 551554 4808 551560 4820
rect 52880 4780 551560 4808
rect 52880 4768 52886 4780
rect 551554 4768 551560 4780
rect 551612 4768 551618 4820
rect 6270 4700 6276 4752
rect 6328 4740 6334 4752
rect 22186 4740 22192 4752
rect 6328 4712 22192 4740
rect 6328 4700 6334 4712
rect 22186 4700 22192 4712
rect 22244 4700 22250 4752
rect 89714 4700 89720 4752
rect 89772 4740 89778 4752
rect 307202 4740 307208 4752
rect 89772 4712 307208 4740
rect 89772 4700 89778 4712
rect 307202 4700 307208 4712
rect 307260 4700 307266 4752
rect 82630 4632 82636 4684
rect 82688 4672 82694 4684
rect 286870 4672 286876 4684
rect 82688 4644 286876 4672
rect 82688 4632 82694 4644
rect 286870 4632 286876 4644
rect 286928 4632 286934 4684
rect 75454 4564 75460 4616
rect 75512 4604 75518 4616
rect 266538 4604 266544 4616
rect 75512 4576 266544 4604
rect 75512 4564 75518 4576
rect 266538 4564 266544 4576
rect 266596 4564 266602 4616
rect 68278 4496 68284 4548
rect 68336 4536 68342 4548
rect 246114 4536 246120 4548
rect 68336 4508 246120 4536
rect 68336 4496 68342 4508
rect 246114 4496 246120 4508
rect 246172 4496 246178 4548
rect 64782 4428 64788 4480
rect 64840 4468 64846 4480
rect 235994 4468 236000 4480
rect 64840 4440 236000 4468
rect 64840 4428 64846 4440
rect 235994 4428 236000 4440
rect 236052 4428 236058 4480
rect 57606 4360 57612 4412
rect 57664 4400 57670 4412
rect 215570 4400 215576 4412
rect 57664 4372 215576 4400
rect 57664 4360 57670 4372
rect 215570 4360 215576 4372
rect 215628 4360 215634 4412
rect 54018 4292 54024 4344
rect 54076 4332 54082 4344
rect 205450 4332 205456 4344
rect 54076 4304 205456 4332
rect 54076 4292 54082 4304
rect 205450 4292 205456 4304
rect 205508 4292 205514 4344
rect 43346 4224 43352 4276
rect 43404 4264 43410 4276
rect 174906 4264 174912 4276
rect 43404 4236 174912 4264
rect 43404 4224 43410 4236
rect 174906 4224 174912 4236
rect 174964 4224 174970 4276
rect 7466 4156 7472 4208
rect 7524 4196 7530 4208
rect 12434 4196 12440 4208
rect 7524 4168 12440 4196
rect 7524 4156 7530 4168
rect 12434 4156 12440 4168
rect 12492 4156 12498 4208
rect 36170 4156 36176 4208
rect 36228 4196 36234 4208
rect 154574 4196 154580 4208
rect 36228 4168 154580 4196
rect 36228 4156 36234 4168
rect 154574 4156 154580 4168
rect 154632 4156 154638 4208
rect 6546 4088 6552 4140
rect 6604 4128 6610 4140
rect 88518 4128 88524 4140
rect 6604 4100 88524 4128
rect 6604 4088 6610 4100
rect 88518 4088 88524 4100
rect 88576 4088 88582 4140
rect 93302 4088 93308 4140
rect 93360 4128 93366 4140
rect 317414 4128 317420 4140
rect 93360 4100 317420 4128
rect 93360 4088 93366 4100
rect 317414 4088 317420 4100
rect 317472 4088 317478 4140
rect 6638 4020 6644 4072
rect 6696 4060 6702 4072
rect 6917 4063 6975 4069
rect 6917 4060 6929 4063
rect 6696 4032 6929 4060
rect 6696 4020 6702 4032
rect 6917 4029 6929 4032
rect 6963 4029 6975 4063
rect 6917 4023 6975 4029
rect 7006 4020 7012 4072
rect 7064 4060 7070 4072
rect 9217 4063 9275 4069
rect 9217 4060 9229 4063
rect 7064 4032 9229 4060
rect 7064 4020 7070 4032
rect 9217 4029 9229 4032
rect 9263 4029 9275 4063
rect 9217 4023 9275 4029
rect 10042 4020 10048 4072
rect 10100 4060 10106 4072
rect 93486 4060 93492 4072
rect 10100 4032 93492 4060
rect 10100 4020 10106 4032
rect 93486 4020 93492 4032
rect 93544 4020 93550 4072
rect 100478 4020 100484 4072
rect 100536 4060 100542 4072
rect 337746 4060 337752 4072
rect 100536 4032 337752 4060
rect 100536 4020 100542 4032
rect 337746 4020 337752 4032
rect 337804 4020 337810 4072
rect 16485 3995 16543 4001
rect 16485 3961 16497 3995
rect 16531 3992 16543 3995
rect 92106 3992 92112 4004
rect 16531 3964 92112 3992
rect 16531 3961 16543 3964
rect 16485 3955 16543 3961
rect 92106 3952 92112 3964
rect 92164 3952 92170 4004
rect 107562 3952 107568 4004
rect 107620 3992 107626 4004
rect 358078 3992 358084 4004
rect 107620 3964 358084 3992
rect 107620 3952 107626 3964
rect 358078 3952 358084 3964
rect 358136 3952 358142 4004
rect 6730 3884 6736 3936
rect 6788 3924 6794 3936
rect 95694 3924 95700 3936
rect 6788 3896 95700 3924
rect 6788 3884 6794 3896
rect 95694 3884 95700 3896
rect 95752 3884 95758 3936
rect 99374 3884 99380 3936
rect 99432 3924 99438 3936
rect 112346 3924 112352 3936
rect 99432 3896 112352 3924
rect 99432 3884 99438 3896
rect 112346 3884 112352 3896
rect 112404 3884 112410 3936
rect 114738 3884 114744 3936
rect 114796 3924 114802 3936
rect 378502 3924 378508 3936
rect 114796 3896 378508 3924
rect 114796 3884 114802 3896
rect 378502 3884 378508 3896
rect 378560 3884 378566 3936
rect 5350 3816 5356 3868
rect 5408 3856 5414 3868
rect 8849 3859 8907 3865
rect 8849 3856 8861 3859
rect 5408 3828 8861 3856
rect 5408 3816 5414 3828
rect 8849 3825 8861 3828
rect 8895 3825 8907 3859
rect 9122 3856 9128 3868
rect 8849 3819 8907 3825
rect 8956 3828 9128 3856
rect 2866 3748 2872 3800
rect 2924 3788 2930 3800
rect 8956 3788 8984 3828
rect 9122 3816 9128 3828
rect 9180 3816 9186 3868
rect 14826 3816 14832 3868
rect 14884 3856 14890 3868
rect 103606 3856 103612 3868
rect 14884 3828 103612 3856
rect 14884 3816 14890 3828
rect 103606 3816 103612 3828
rect 103664 3816 103670 3868
rect 104250 3816 104256 3868
rect 104308 3856 104314 3868
rect 105170 3856 105176 3868
rect 104308 3828 105176 3856
rect 104308 3816 104314 3828
rect 105170 3816 105176 3828
rect 105228 3816 105234 3868
rect 121822 3816 121828 3868
rect 121880 3856 121886 3868
rect 398834 3856 398840 3868
rect 121880 3828 398840 3856
rect 121880 3816 121886 3828
rect 398834 3816 398840 3828
rect 398892 3816 398898 3868
rect 2924 3760 8984 3788
rect 9033 3791 9091 3797
rect 2924 3748 2930 3760
rect 9033 3757 9045 3791
rect 9079 3788 9091 3791
rect 16022 3788 16028 3800
rect 9079 3760 16028 3788
rect 9079 3757 9091 3760
rect 9033 3751 9091 3757
rect 16022 3748 16028 3760
rect 16080 3748 16086 3800
rect 37366 3748 37372 3800
rect 37424 3788 37430 3800
rect 419166 3788 419172 3800
rect 37424 3760 419172 3788
rect 37424 3748 37430 3760
rect 419166 3748 419172 3760
rect 419224 3748 419230 3800
rect 9217 3723 9275 3729
rect 9217 3689 9229 3723
rect 9263 3720 9275 3723
rect 27890 3720 27896 3732
rect 9263 3692 27896 3720
rect 9263 3689 9275 3692
rect 9217 3683 9275 3689
rect 27890 3680 27896 3692
rect 27948 3680 27954 3732
rect 44542 3680 44548 3732
rect 44600 3720 44606 3732
rect 429378 3720 429384 3732
rect 44600 3692 429384 3720
rect 44600 3680 44606 3692
rect 429378 3680 429384 3692
rect 429436 3680 429442 3732
rect 5074 3612 5080 3664
rect 5132 3652 5138 3664
rect 74258 3652 74264 3664
rect 5132 3624 74264 3652
rect 5132 3612 5138 3624
rect 74258 3612 74264 3624
rect 74316 3612 74322 3664
rect 76650 3612 76656 3664
rect 76708 3652 76714 3664
rect 470042 3652 470048 3664
rect 76708 3624 470048 3652
rect 76708 3612 76714 3624
rect 470042 3612 470048 3624
rect 470100 3612 470106 3664
rect 5166 3544 5172 3596
rect 5224 3584 5230 3596
rect 81434 3584 81440 3596
rect 5224 3556 81440 3584
rect 5224 3544 5230 3556
rect 81434 3544 81440 3556
rect 81492 3544 81498 3596
rect 87322 3544 87328 3596
rect 87380 3584 87386 3596
rect 490466 3584 490472 3596
rect 87380 3556 490472 3584
rect 87380 3544 87386 3556
rect 490466 3544 490472 3556
rect 490524 3544 490530 3596
rect 5442 3476 5448 3528
rect 5500 3516 5506 3528
rect 6454 3516 6460 3528
rect 5500 3488 6460 3516
rect 5500 3476 5506 3488
rect 6454 3476 6460 3488
rect 6512 3476 6518 3528
rect 18322 3516 18328 3528
rect 6564 3488 18328 3516
rect 4798 3408 4804 3460
rect 4856 3448 4862 3460
rect 6564 3448 6592 3488
rect 18322 3476 18328 3488
rect 18380 3476 18386 3528
rect 24302 3476 24308 3528
rect 24360 3516 24366 3528
rect 124030 3516 124036 3528
rect 24360 3488 124036 3516
rect 24360 3476 24366 3488
rect 124030 3476 124036 3488
rect 124088 3476 124094 3528
rect 124214 3476 124220 3528
rect 124272 3516 124278 3528
rect 578234 3516 578240 3528
rect 124272 3488 578240 3516
rect 124272 3476 124278 3488
rect 578234 3476 578240 3488
rect 578292 3476 578298 3528
rect 4856 3420 6592 3448
rect 4856 3408 4862 3420
rect 7650 3408 7656 3460
rect 7708 3448 7714 3460
rect 9030 3448 9036 3460
rect 7708 3420 9036 3448
rect 7708 3408 7714 3420
rect 9030 3408 9036 3420
rect 9088 3408 9094 3460
rect 13630 3408 13636 3460
rect 13688 3448 13694 3460
rect 521010 3448 521016 3460
rect 13688 3420 521016 3448
rect 13688 3408 13694 3420
rect 521010 3408 521016 3420
rect 521068 3408 521074 3460
rect 4982 3340 4988 3392
rect 5040 3380 5046 3392
rect 70670 3380 70676 3392
rect 5040 3352 70676 3380
rect 5040 3340 5046 3352
rect 70670 3340 70676 3352
rect 70728 3340 70734 3392
rect 86126 3340 86132 3392
rect 86184 3380 86190 3392
rect 297082 3380 297088 3392
rect 86184 3352 297088 3380
rect 86184 3340 86190 3352
rect 297082 3340 297088 3352
rect 297140 3340 297146 3392
rect 9490 3272 9496 3324
rect 9548 3312 9554 3324
rect 59998 3312 60004 3324
rect 9548 3284 60004 3312
rect 9548 3272 9554 3284
rect 59998 3272 60004 3284
rect 60056 3272 60062 3324
rect 79042 3272 79048 3324
rect 79100 3312 79106 3324
rect 276658 3312 276664 3324
rect 79100 3284 276664 3312
rect 79100 3272 79106 3284
rect 276658 3272 276664 3284
rect 276716 3272 276722 3324
rect 9582 3204 9588 3256
rect 9640 3244 9646 3256
rect 56410 3244 56416 3256
rect 9640 3216 56416 3244
rect 9640 3204 9646 3216
rect 56410 3204 56416 3216
rect 56468 3204 56474 3256
rect 71866 3204 71872 3256
rect 71924 3244 71930 3256
rect 256326 3244 256332 3256
rect 71924 3216 256332 3244
rect 71924 3204 71930 3216
rect 256326 3204 256332 3216
rect 256384 3204 256390 3256
rect 4890 3136 4896 3188
rect 4948 3176 4954 3188
rect 45738 3176 45744 3188
rect 4948 3148 45744 3176
rect 4948 3136 4954 3148
rect 45738 3136 45744 3148
rect 45796 3136 45802 3188
rect 46934 3136 46940 3188
rect 46992 3176 46998 3188
rect 46992 3148 49464 3176
rect 46992 3136 46998 3148
rect 4062 3068 4068 3120
rect 4120 3108 4126 3120
rect 8938 3108 8944 3120
rect 4120 3080 8944 3108
rect 4120 3068 4126 3080
rect 8938 3068 8944 3080
rect 8996 3068 9002 3120
rect 9674 3068 9680 3120
rect 9732 3108 9738 3120
rect 49326 3108 49332 3120
rect 9732 3080 49332 3108
rect 9732 3068 9738 3080
rect 49326 3068 49332 3080
rect 49384 3068 49390 3120
rect 9766 3000 9772 3052
rect 9824 3040 9830 3052
rect 48130 3040 48136 3052
rect 9824 3012 48136 3040
rect 9824 3000 9830 3012
rect 48130 3000 48136 3012
rect 48188 3000 48194 3052
rect 49436 3040 49464 3148
rect 61194 3136 61200 3188
rect 61252 3176 61258 3188
rect 225782 3176 225788 3188
rect 61252 3148 225788 3176
rect 61252 3136 61258 3148
rect 225782 3136 225788 3148
rect 225840 3136 225846 3188
rect 50522 3068 50528 3120
rect 50580 3108 50586 3120
rect 195238 3108 195244 3120
rect 50580 3080 195244 3108
rect 50580 3068 50586 3080
rect 195238 3068 195244 3080
rect 195296 3068 195302 3120
rect 185026 3040 185032 3052
rect 49436 3012 185032 3040
rect 185026 3000 185032 3012
rect 185084 3000 185090 3052
rect 4706 2932 4712 2984
rect 4764 2972 4770 2984
rect 38562 2972 38568 2984
rect 4764 2944 38568 2972
rect 4764 2932 4770 2944
rect 38562 2932 38568 2944
rect 38620 2932 38626 2984
rect 39758 2932 39764 2984
rect 39816 2972 39822 2984
rect 164694 2972 164700 2984
rect 39816 2944 164700 2972
rect 39816 2932 39822 2944
rect 164694 2932 164700 2944
rect 164752 2932 164758 2984
rect 6917 2907 6975 2913
rect 6917 2873 6929 2907
rect 6963 2904 6975 2907
rect 16485 2907 16543 2913
rect 16485 2904 16497 2907
rect 6963 2876 16497 2904
rect 6963 2873 6975 2876
rect 6917 2867 6975 2873
rect 16485 2873 16497 2876
rect 16531 2873 16543 2907
rect 16485 2867 16543 2873
rect 32674 2864 32680 2916
rect 32732 2904 32738 2916
rect 144362 2904 144368 2916
rect 32732 2876 144368 2904
rect 32732 2864 32738 2876
rect 144362 2864 144368 2876
rect 144420 2864 144426 2916
rect 29086 2796 29092 2848
rect 29144 2836 29150 2848
rect 134150 2836 134156 2848
rect 29144 2808 134156 2836
rect 29144 2796 29150 2808
rect 134150 2796 134156 2808
rect 134208 2796 134214 2848
<< via1 >>
rect 150348 700680 150400 700732
rect 170312 700680 170364 700732
rect 128268 700612 128320 700664
rect 235172 700612 235224 700664
rect 106188 700544 106240 700596
rect 300124 700544 300176 700596
rect 84108 700476 84160 700528
rect 364984 700476 365036 700528
rect 40500 700408 40552 700460
rect 41328 700408 41380 700460
rect 62028 700408 62080 700460
rect 429844 700408 429896 700460
rect 39948 700340 40000 700392
rect 494796 700340 494848 700392
rect 19248 700272 19300 700324
rect 559656 700272 559708 700324
rect 105452 699660 105504 699712
rect 106096 699660 106148 699712
rect 17960 689936 18012 689988
rect 19248 689936 19300 689988
rect 127532 689528 127584 689580
rect 128268 689528 128320 689580
rect 149428 689528 149480 689580
rect 150348 689528 150400 689580
rect 9496 689392 9548 689444
rect 456432 689392 456484 689444
rect 106096 689324 106148 689376
rect 171416 689324 171468 689376
rect 41328 689256 41380 689308
rect 193312 689256 193364 689308
rect 9128 689188 9180 689240
rect 237196 689188 237248 689240
rect 9036 689120 9088 689172
rect 259092 689120 259144 689172
rect 9404 689052 9456 689104
rect 280988 689052 281040 689104
rect 9772 688984 9824 689036
rect 302976 688984 303028 689036
rect 215208 688916 215260 688968
rect 576124 688916 576176 688968
rect 8944 688848 8996 688900
rect 390652 688848 390704 688900
rect 9680 688780 9732 688832
rect 412548 688780 412600 688832
rect 9588 688712 9640 688764
rect 434444 688712 434496 688764
rect 9312 686468 9364 686520
rect 368388 686468 368440 686520
rect 3332 681708 3384 681760
rect 6184 681708 6236 681760
rect 575940 674908 575992 674960
rect 576308 674908 576360 674960
rect 575940 652876 575992 652928
rect 576308 652876 576360 652928
rect 575940 647776 575992 647828
rect 576032 634831 576084 634840
rect 576032 634797 576041 634831
rect 576041 634797 576075 634831
rect 576075 634797 576084 634831
rect 576032 634788 576084 634797
rect 6736 627920 6788 627972
rect 6920 627920 6972 627972
rect 3148 624180 3200 624232
rect 6276 624180 6328 624232
rect 6736 621052 6788 621104
rect 6644 618307 6696 618316
rect 6644 618273 6653 618307
rect 6653 618273 6687 618307
rect 6687 618273 6696 618307
rect 6644 618264 6696 618273
rect 6644 618128 6696 618180
rect 6552 608651 6604 608660
rect 6552 608617 6561 608651
rect 6561 608617 6595 608651
rect 6595 608617 6604 608651
rect 6552 608608 6604 608617
rect 575940 602352 575992 602404
rect 6552 601740 6604 601792
rect 6920 601740 6972 601792
rect 6552 601604 6604 601656
rect 6920 601604 6972 601656
rect 6460 601536 6512 601588
rect 6736 601536 6788 601588
rect 576032 597567 576084 597576
rect 576032 597533 576041 597567
rect 576041 597533 576075 597567
rect 576075 597533 576084 597567
rect 576032 597524 576084 597533
rect 6552 592084 6604 592136
rect 6552 591948 6604 592000
rect 6460 591880 6512 591932
rect 6736 591880 6788 591932
rect 6552 582360 6604 582412
rect 6920 582360 6972 582412
rect 6368 582224 6420 582276
rect 6736 582224 6788 582276
rect 6736 572883 6788 572892
rect 6736 572849 6745 572883
rect 6745 572849 6779 572883
rect 6779 572849 6788 572883
rect 6736 572840 6788 572849
rect 6368 572432 6420 572484
rect 6828 572432 6880 572484
rect 6736 572407 6788 572416
rect 6736 572373 6745 572407
rect 6745 572373 6779 572407
rect 6779 572373 6788 572407
rect 6736 572364 6788 572373
rect 4068 567264 4120 567316
rect 7564 567264 7616 567316
rect 575940 567196 575992 567248
rect 575940 567060 575992 567112
rect 575940 564383 575992 564392
rect 575940 564349 575949 564383
rect 575949 564349 575983 564383
rect 575983 564349 575992 564383
rect 575940 564340 575992 564349
rect 6828 563184 6880 563236
rect 6460 563048 6512 563100
rect 6368 562980 6420 563032
rect 6920 562980 6972 563032
rect 576032 554752 576084 554804
rect 6368 553460 6420 553512
rect 6460 553392 6512 553444
rect 6736 553392 6788 553444
rect 6828 553392 6880 553444
rect 6460 553256 6512 553308
rect 6828 553256 6880 553308
rect 6460 543804 6512 543856
rect 6920 543804 6972 543856
rect 6368 543668 6420 543720
rect 6920 543668 6972 543720
rect 575940 536800 575992 536852
rect 576032 536800 576084 536852
rect 6368 534148 6420 534200
rect 6460 534080 6512 534132
rect 6736 534080 6788 534132
rect 6828 534080 6880 534132
rect 6460 533944 6512 533996
rect 6828 533944 6880 533996
rect 6460 524424 6512 524476
rect 6920 524424 6972 524476
rect 575940 522291 575992 522300
rect 575940 522257 575949 522291
rect 575949 522257 575983 522291
rect 575983 522257 575992 522291
rect 575940 522248 575992 522257
rect 575940 519936 575992 519988
rect 576308 519936 576360 519988
rect 575940 518007 575992 518016
rect 575940 517973 575949 518007
rect 575949 517973 575983 518007
rect 575983 517973 575992 518007
rect 575940 517964 575992 517973
rect 6736 514904 6788 514956
rect 6460 514768 6512 514820
rect 6736 514768 6788 514820
rect 6828 514768 6880 514820
rect 575940 514743 575992 514752
rect 575940 514709 575949 514743
rect 575949 514709 575983 514743
rect 575983 514709 575992 514743
rect 575940 514700 575992 514709
rect 576032 514700 576084 514752
rect 576216 514700 576268 514752
rect 6460 514632 6512 514684
rect 6828 514632 6880 514684
rect 575940 509507 575992 509516
rect 575940 509473 575949 509507
rect 575949 509473 575983 509507
rect 575983 509473 575992 509507
rect 575940 509464 575992 509473
rect 575940 505316 575992 505368
rect 576216 505316 576268 505368
rect 6460 505112 6512 505164
rect 6920 505112 6972 505164
rect 6736 495592 6788 495644
rect 6460 495456 6512 495508
rect 6736 495456 6788 495508
rect 6828 495456 6880 495508
rect 6460 495320 6512 495372
rect 6828 495320 6880 495372
rect 576032 492600 576084 492652
rect 575940 487772 575992 487824
rect 576124 487092 576176 487144
rect 579620 487092 579672 487144
rect 6460 485800 6512 485852
rect 6920 485800 6972 485852
rect 575940 485732 575992 485784
rect 576032 485732 576084 485784
rect 575940 485596 575992 485648
rect 575940 485503 575992 485512
rect 575940 485469 575949 485503
rect 575949 485469 575983 485503
rect 575983 485469 575992 485503
rect 575940 485460 575992 485469
rect 6736 476212 6788 476264
rect 6460 476076 6512 476128
rect 6736 476076 6788 476128
rect 6828 476076 6880 476128
rect 575940 466488 575992 466540
rect 576032 466420 576084 466472
rect 575940 466216 575992 466268
rect 576124 466216 576176 466268
rect 6736 456900 6788 456952
rect 6460 456764 6512 456816
rect 6736 456764 6788 456816
rect 6828 456764 6880 456816
rect 576032 447108 576084 447160
rect 576124 447040 576176 447092
rect 6736 437588 6788 437640
rect 6460 437452 6512 437504
rect 6736 437452 6788 437504
rect 6828 437452 6880 437504
rect 576032 428476 576084 428528
rect 575940 427660 575992 427712
rect 575940 427524 575992 427576
rect 576124 417843 576176 417852
rect 576124 417809 576133 417843
rect 576133 417809 576167 417843
rect 576167 417809 576176 417843
rect 576124 417800 576176 417809
rect 575940 405560 575992 405612
rect 6460 398828 6512 398880
rect 6736 398828 6788 398880
rect 575940 396992 575992 397044
rect 576124 396992 576176 397044
rect 576032 396083 576084 396092
rect 576032 396049 576041 396083
rect 576041 396049 576075 396083
rect 576075 396049 576084 396083
rect 576032 396040 576084 396049
rect 575940 390099 575992 390108
rect 575940 390065 575949 390099
rect 575949 390065 575983 390099
rect 575983 390065 575992 390099
rect 575940 390056 575992 390065
rect 6460 389104 6512 389156
rect 6736 389104 6788 389156
rect 6828 389104 6880 389156
rect 6368 389036 6420 389088
rect 575940 384344 575992 384396
rect 6368 379584 6420 379636
rect 6460 379516 6512 379568
rect 6736 379516 6788 379568
rect 6828 379516 6880 379568
rect 576032 379448 576084 379500
rect 576124 379380 576176 379432
rect 576124 376703 576176 376712
rect 576124 376669 576133 376703
rect 576133 376669 576167 376703
rect 576167 376669 576176 376703
rect 576124 376660 576176 376669
rect 576032 371943 576084 371952
rect 576032 371909 576041 371943
rect 576041 371909 576075 371943
rect 576075 371909 576084 371943
rect 576032 371900 576084 371909
rect 6460 369792 6512 369844
rect 6736 369792 6788 369844
rect 6828 369792 6880 369844
rect 6368 369724 6420 369776
rect 575940 366460 575992 366512
rect 575940 365848 575992 365900
rect 575940 361267 575992 361276
rect 575940 361233 575949 361267
rect 575949 361233 575983 361267
rect 575983 361233 575992 361267
rect 575940 361224 575992 361233
rect 6368 360272 6420 360324
rect 6460 360204 6512 360256
rect 6736 360204 6788 360256
rect 6828 360204 6880 360256
rect 575940 359456 575992 359508
rect 575940 359363 575992 359372
rect 575940 359329 575949 359363
rect 575949 359329 575983 359363
rect 575983 359329 575992 359363
rect 575940 359320 575992 359329
rect 575940 358980 575992 359032
rect 575940 352699 575992 352708
rect 575940 352665 575949 352699
rect 575949 352665 575983 352699
rect 575983 352665 575992 352699
rect 575940 352656 575992 352665
rect 6460 350480 6512 350532
rect 6736 350480 6788 350532
rect 6828 350480 6880 350532
rect 6368 350412 6420 350464
rect 575940 347463 575992 347472
rect 575940 347429 575949 347463
rect 575949 347429 575983 347463
rect 575983 347429 575992 347463
rect 575940 347420 575992 347429
rect 6368 340960 6420 341012
rect 6460 340892 6512 340944
rect 6736 340892 6788 340944
rect 6828 340892 6880 340944
rect 575940 338036 575992 338088
rect 575940 334611 575992 334620
rect 575940 334577 575949 334611
rect 575949 334577 575983 334611
rect 575983 334577 575992 334611
rect 575940 334568 575992 334577
rect 575940 331848 575992 331900
rect 6368 331168 6420 331220
rect 6736 331168 6788 331220
rect 6828 331168 6880 331220
rect 6092 331100 6144 331152
rect 575940 328015 575992 328024
rect 575940 327981 575949 328015
rect 575949 327981 575983 328015
rect 575983 327981 575992 328015
rect 575940 327972 575992 327981
rect 576124 325660 576176 325712
rect 576216 325660 576268 325712
rect 575940 321963 575992 321972
rect 575940 321929 575949 321963
rect 575949 321929 575983 321963
rect 575983 321929 575992 321963
rect 575940 321920 575992 321929
rect 6092 321648 6144 321700
rect 6368 321580 6420 321632
rect 6736 321580 6788 321632
rect 6828 321580 6880 321632
rect 575940 319472 575992 319524
rect 575940 319200 575992 319252
rect 575940 319107 575992 319116
rect 575940 319073 575949 319107
rect 575949 319073 575983 319107
rect 575983 319073 575992 319107
rect 575940 319064 575992 319073
rect 576124 315936 576176 315988
rect 575940 315775 575992 315784
rect 575940 315741 575949 315775
rect 575949 315741 575983 315775
rect 575983 315741 575992 315775
rect 575940 315732 575992 315741
rect 575940 315596 575992 315648
rect 6092 311788 6144 311840
rect 6736 311788 6788 311840
rect 6828 311788 6880 311840
rect 6368 311720 6420 311772
rect 575940 307776 575992 307828
rect 576308 307776 576360 307828
rect 576032 306391 576084 306400
rect 576032 306357 576041 306391
rect 576041 306357 576075 306391
rect 576075 306357 576084 306391
rect 576032 306348 576084 306357
rect 6368 302744 6420 302796
rect 6092 302200 6144 302252
rect 6736 302200 6788 302252
rect 6828 302200 6880 302252
rect 575940 299183 575992 299192
rect 575940 299149 575949 299183
rect 575949 299149 575983 299183
rect 575983 299149 575992 299183
rect 575940 299140 575992 299149
rect 6092 292476 6144 292528
rect 6736 292476 6788 292528
rect 6828 292476 6880 292528
rect 6000 292408 6052 292460
rect 575940 288464 575992 288516
rect 576124 288464 576176 288516
rect 575940 286424 575992 286476
rect 576032 286424 576084 286476
rect 575940 286220 575992 286272
rect 576032 286220 576084 286272
rect 6000 282956 6052 283008
rect 6092 282888 6144 282940
rect 6736 282888 6788 282940
rect 6828 282888 6880 282940
rect 575940 278876 575992 278928
rect 576124 278876 576176 278928
rect 575940 278783 575992 278792
rect 575940 278749 575949 278783
rect 575949 278749 575983 278783
rect 575983 278749 575992 278783
rect 575940 278740 575992 278749
rect 6092 273164 6144 273216
rect 6736 273164 6788 273216
rect 6828 273164 6880 273216
rect 6000 273096 6052 273148
rect 575940 273003 575992 273012
rect 575940 272969 575949 273003
rect 575949 272969 575983 273003
rect 575983 272969 575992 273003
rect 575940 272960 575992 272969
rect 576032 272323 576084 272332
rect 576032 272289 576041 272323
rect 576041 272289 576075 272323
rect 576075 272289 576084 272323
rect 576032 272280 576084 272289
rect 576032 270351 576084 270360
rect 576032 270317 576041 270351
rect 576041 270317 576075 270351
rect 576075 270317 576084 270351
rect 576032 270308 576084 270317
rect 6000 263644 6052 263696
rect 6092 263576 6144 263628
rect 6736 263576 6788 263628
rect 6828 263576 6880 263628
rect 575940 262896 575992 262948
rect 576216 262896 576268 262948
rect 575940 262735 575992 262744
rect 575940 262701 575949 262735
rect 575949 262701 575983 262735
rect 575983 262701 575992 262735
rect 575940 262692 575992 262701
rect 575940 257635 575992 257644
rect 575940 257601 575949 257635
rect 575949 257601 575983 257635
rect 575983 257601 575992 257635
rect 575940 257592 575992 257601
rect 575940 257456 575992 257508
rect 6092 253852 6144 253904
rect 6736 253852 6788 253904
rect 6828 253852 6880 253904
rect 6000 253784 6052 253836
rect 575940 253240 575992 253292
rect 575940 253036 575992 253088
rect 575940 249135 575992 249144
rect 575940 249101 575949 249135
rect 575949 249101 575983 249135
rect 575983 249101 575992 249135
rect 575940 249092 575992 249101
rect 6000 244332 6052 244384
rect 6092 244264 6144 244316
rect 6736 244264 6788 244316
rect 6828 244264 6880 244316
rect 576032 243151 576084 243160
rect 576032 243117 576041 243151
rect 576041 243117 576075 243151
rect 576075 243117 576084 243151
rect 576032 243108 576084 243117
rect 575940 241680 575992 241732
rect 576308 241680 576360 241732
rect 576032 241408 576084 241460
rect 576124 241204 576176 241256
rect 576216 236827 576268 236836
rect 576216 236793 576225 236827
rect 576225 236793 576259 236827
rect 576259 236793 576268 236827
rect 576216 236784 576268 236793
rect 575940 236648 575992 236700
rect 576216 236648 576268 236700
rect 575940 235016 575992 235068
rect 576308 235016 576360 235068
rect 6092 234540 6144 234592
rect 6736 234540 6788 234592
rect 6828 234540 6880 234592
rect 6000 234472 6052 234524
rect 576032 234268 576084 234320
rect 576400 234268 576452 234320
rect 6000 225020 6052 225072
rect 6092 224952 6144 225004
rect 6736 224952 6788 225004
rect 6828 224952 6880 225004
rect 576124 224927 576176 224936
rect 576124 224893 576133 224927
rect 576133 224893 576167 224927
rect 576167 224893 576176 224927
rect 576124 224884 576176 224893
rect 575940 220983 575992 220992
rect 575940 220949 575949 220983
rect 575949 220949 575983 220983
rect 575983 220949 575992 220983
rect 575940 220940 575992 220949
rect 575940 217608 575992 217660
rect 576032 217515 576084 217524
rect 576032 217481 576041 217515
rect 576041 217481 576075 217515
rect 576075 217481 576084 217515
rect 576032 217472 576084 217481
rect 576216 217472 576268 217524
rect 576400 217472 576452 217524
rect 579068 216316 579120 216368
rect 580632 216316 580684 216368
rect 575940 215976 575992 216028
rect 575940 215500 575992 215552
rect 6092 215228 6144 215280
rect 6736 215228 6788 215280
rect 6828 215228 6880 215280
rect 6000 215160 6052 215212
rect 576124 212576 576176 212628
rect 576124 212483 576176 212492
rect 576124 212449 576133 212483
rect 576133 212449 576167 212483
rect 576167 212449 576176 212483
rect 576124 212440 576176 212449
rect 6000 205708 6052 205760
rect 6092 205640 6144 205692
rect 6736 205640 6788 205692
rect 6828 205640 6880 205692
rect 576032 203099 576084 203108
rect 576032 203065 576041 203099
rect 576041 203065 576075 203099
rect 576075 203065 576084 203099
rect 576032 203056 576084 203065
rect 575940 202716 575992 202768
rect 576216 202716 576268 202768
rect 576216 201492 576268 201544
rect 575940 199248 575992 199300
rect 576308 198840 576360 198892
rect 576308 198747 576360 198756
rect 576308 198713 576317 198747
rect 576317 198713 576351 198747
rect 576351 198713 576360 198747
rect 576308 198704 576360 198713
rect 576124 197344 576176 197396
rect 6092 195916 6144 195968
rect 6736 195916 6788 195968
rect 6828 195916 6880 195968
rect 6000 195848 6052 195900
rect 579068 194012 579120 194064
rect 580724 194012 580776 194064
rect 576032 192763 576084 192772
rect 576032 192729 576041 192763
rect 576041 192729 576075 192763
rect 576075 192729 576084 192763
rect 576032 192720 576084 192729
rect 576124 192516 576176 192568
rect 576216 191811 576268 191820
rect 576216 191777 576225 191811
rect 576225 191777 576259 191811
rect 576259 191777 576268 191811
rect 576216 191768 576268 191777
rect 576032 191131 576084 191140
rect 576032 191097 576041 191131
rect 576041 191097 576075 191131
rect 576075 191097 576084 191131
rect 576032 191088 576084 191097
rect 575940 186872 575992 186924
rect 6000 186396 6052 186448
rect 6092 186328 6144 186380
rect 6736 186328 6788 186380
rect 6828 186328 6880 186380
rect 576216 186303 576268 186312
rect 576216 186269 576225 186303
rect 576225 186269 576259 186303
rect 576259 186269 576268 186303
rect 576216 186260 576268 186269
rect 575940 184900 575992 184952
rect 576308 184900 576360 184952
rect 575940 183336 575992 183388
rect 576308 183336 576360 183388
rect 576032 182928 576084 182980
rect 575940 177216 575992 177268
rect 6092 176604 6144 176656
rect 6736 176604 6788 176656
rect 6828 176604 6880 176656
rect 6000 176536 6052 176588
rect 575940 175652 575992 175704
rect 575940 174768 575992 174820
rect 575940 173995 575992 174004
rect 575940 173961 575949 173995
rect 575949 173961 575983 173995
rect 575983 173961 575992 173995
rect 575940 173952 575992 173961
rect 576124 172524 576176 172576
rect 579068 172116 579120 172168
rect 580816 172116 580868 172168
rect 3240 171096 3292 171148
rect 4712 171096 4764 171148
rect 575940 170731 575992 170740
rect 575940 170697 575949 170731
rect 575949 170697 575983 170731
rect 575983 170697 575992 170731
rect 575940 170688 575992 170697
rect 575940 170212 575992 170264
rect 575940 170076 575992 170128
rect 576124 170076 576176 170128
rect 6000 167084 6052 167136
rect 6092 167016 6144 167068
rect 6736 167016 6788 167068
rect 6828 167016 6880 167068
rect 575940 164908 575992 164960
rect 575940 160803 575992 160812
rect 575940 160769 575949 160803
rect 575949 160769 575983 160803
rect 575983 160769 575992 160803
rect 575940 160760 575992 160769
rect 576124 158015 576176 158024
rect 576124 157981 576133 158015
rect 576133 157981 576167 158015
rect 576167 157981 576176 158015
rect 576124 157972 576176 157981
rect 576124 157836 576176 157888
rect 6092 157292 6144 157344
rect 6736 157292 6788 157344
rect 6828 157292 6880 157344
rect 6000 157224 6052 157276
rect 575940 153459 575992 153468
rect 575940 153425 575949 153459
rect 575949 153425 575983 153459
rect 575983 153425 575992 153459
rect 575940 153416 575992 153425
rect 575940 153212 575992 153264
rect 575940 150467 575992 150476
rect 575940 150433 575949 150467
rect 575949 150433 575983 150467
rect 575983 150433 575992 150467
rect 575940 150424 575992 150433
rect 579068 150084 579120 150136
rect 580908 150084 580960 150136
rect 576032 149676 576084 149728
rect 575940 149379 575992 149388
rect 575940 149345 575949 149379
rect 575949 149345 575983 149379
rect 575983 149345 575992 149379
rect 575940 149336 575992 149345
rect 6000 147704 6052 147756
rect 6092 147636 6144 147688
rect 6736 147636 6788 147688
rect 6828 147636 6880 147688
rect 575940 145936 575992 145988
rect 575940 145256 575992 145308
rect 575940 144848 575992 144900
rect 576032 144508 576084 144560
rect 576308 144508 576360 144560
rect 575940 144415 575992 144424
rect 575940 144381 575949 144415
rect 575949 144381 575983 144415
rect 575983 144381 575992 144415
rect 575940 144372 575992 144381
rect 575940 140947 575992 140956
rect 575940 140913 575949 140947
rect 575949 140913 575983 140947
rect 575983 140913 575992 140947
rect 575940 140904 575992 140913
rect 575940 140292 575992 140344
rect 575940 139884 575992 139936
rect 576124 139884 576176 139936
rect 6092 137912 6144 137964
rect 6736 137912 6788 137964
rect 6828 137912 6880 137964
rect 6000 137844 6052 137896
rect 575940 137164 575992 137216
rect 576032 137028 576084 137080
rect 575940 136960 575992 137012
rect 575940 132583 575992 132592
rect 575940 132549 575949 132583
rect 575949 132549 575983 132583
rect 575983 132549 575992 132583
rect 575940 132540 575992 132549
rect 575940 132107 575992 132116
rect 575940 132073 575949 132107
rect 575949 132073 575983 132107
rect 575983 132073 575992 132107
rect 575940 132064 575992 132073
rect 575940 130500 575992 130552
rect 6000 128392 6052 128444
rect 6092 128324 6144 128376
rect 6736 128324 6788 128376
rect 6828 128324 6880 128376
rect 3332 128256 3384 128308
rect 4160 128256 4212 128308
rect 579068 127916 579120 127968
rect 580172 127916 580224 127968
rect 575940 127644 575992 127696
rect 575940 122544 575992 122596
rect 575940 121592 575992 121644
rect 576124 121592 576176 121644
rect 576308 120708 576360 120760
rect 6092 118600 6144 118652
rect 6736 118600 6788 118652
rect 6828 118600 6880 118652
rect 6000 118532 6052 118584
rect 576124 118532 576176 118584
rect 575940 117716 575992 117768
rect 576032 115880 576084 115932
rect 575940 113976 575992 114028
rect 575940 110916 575992 110968
rect 6000 109080 6052 109132
rect 6092 109012 6144 109064
rect 6736 109012 6788 109064
rect 6828 109012 6880 109064
rect 576124 108851 576176 108860
rect 576124 108817 576133 108851
rect 576133 108817 576167 108851
rect 576167 108817 576176 108851
rect 576124 108808 576176 108817
rect 579068 106156 579120 106208
rect 580632 106156 580684 106208
rect 575940 104431 575992 104440
rect 575940 104397 575949 104431
rect 575949 104397 575983 104431
rect 575983 104397 575992 104431
rect 575940 104388 575992 104397
rect 575940 104252 575992 104304
rect 575940 104116 575992 104168
rect 576400 104116 576452 104168
rect 575940 102416 575992 102468
rect 575940 100444 575992 100496
rect 575940 100308 575992 100360
rect 6092 99288 6144 99340
rect 6736 99288 6788 99340
rect 6828 99288 6880 99340
rect 6000 99220 6052 99272
rect 575940 93780 575992 93832
rect 575940 90584 575992 90636
rect 6000 89768 6052 89820
rect 6092 89700 6144 89752
rect 6736 89700 6788 89752
rect 6828 89700 6880 89752
rect 576308 85620 576360 85672
rect 576308 85484 576360 85536
rect 579068 84124 579120 84176
rect 580724 84124 580776 84176
rect 575940 81379 575992 81388
rect 575940 81345 575949 81379
rect 575949 81345 575983 81379
rect 575983 81345 575992 81379
rect 575940 81336 575992 81345
rect 576124 81379 576176 81388
rect 576124 81345 576133 81379
rect 576133 81345 576167 81379
rect 576167 81345 576176 81379
rect 576124 81336 576176 81345
rect 6092 79976 6144 80028
rect 6736 79976 6788 80028
rect 6828 79976 6880 80028
rect 6000 79908 6052 79960
rect 575940 79432 575992 79484
rect 576032 74783 576084 74792
rect 576032 74749 576041 74783
rect 576041 74749 576075 74783
rect 576075 74749 576084 74783
rect 576032 74740 576084 74749
rect 575940 72199 575992 72208
rect 575940 72165 575949 72199
rect 575949 72165 575983 72199
rect 575983 72165 575992 72199
rect 575940 72156 575992 72165
rect 6000 70456 6052 70508
rect 6092 70388 6144 70440
rect 6736 70388 6788 70440
rect 6828 70388 6880 70440
rect 575940 70320 575992 70372
rect 576032 67575 576084 67584
rect 576032 67541 576041 67575
rect 576041 67541 576075 67575
rect 576075 67541 576084 67575
rect 576032 67532 576084 67541
rect 575940 63359 575992 63368
rect 575940 63325 575949 63359
rect 575949 63325 575983 63359
rect 575983 63325 575992 63359
rect 575940 63316 575992 63325
rect 579068 61956 579120 62008
rect 580816 61956 580868 62008
rect 576124 61548 576176 61600
rect 576400 61548 576452 61600
rect 6092 60664 6144 60716
rect 6736 60664 6788 60716
rect 6828 60664 6880 60716
rect 6000 60596 6052 60648
rect 575940 58760 575992 58812
rect 576216 57944 576268 57996
rect 576308 57944 576360 57996
rect 576124 57808 576176 57860
rect 576308 57307 576360 57316
rect 576308 57273 576317 57307
rect 576317 57273 576351 57307
rect 576351 57273 576360 57307
rect 576308 57264 576360 57273
rect 575940 52776 575992 52828
rect 575940 52572 575992 52624
rect 576124 51756 576176 51808
rect 6000 51144 6052 51196
rect 6092 51076 6144 51128
rect 6736 51076 6788 51128
rect 6828 51076 6880 51128
rect 575940 46384 575992 46436
rect 576032 46180 576084 46232
rect 575940 43596 575992 43648
rect 575940 43503 575992 43512
rect 575940 43469 575949 43503
rect 575949 43469 575983 43503
rect 575983 43469 575992 43503
rect 575940 43460 575992 43469
rect 6092 41352 6144 41404
rect 6736 41352 6788 41404
rect 6828 41352 6880 41404
rect 6000 41284 6052 41336
rect 579068 39924 579120 39976
rect 580632 39924 580684 39976
rect 575940 39380 575992 39432
rect 575940 37247 575992 37256
rect 575940 37213 575949 37247
rect 575949 37213 575983 37247
rect 575983 37213 575992 37247
rect 575940 37204 575992 37213
rect 575940 35300 575992 35352
rect 575940 35164 575992 35216
rect 575940 33804 575992 33856
rect 576124 33804 576176 33856
rect 576400 33804 576452 33856
rect 575940 33056 575992 33108
rect 6000 31832 6052 31884
rect 6092 31764 6144 31816
rect 6736 31764 6788 31816
rect 6828 31764 6880 31816
rect 576032 28636 576084 28688
rect 576308 28636 576360 28688
rect 575940 28296 575992 28348
rect 576216 24148 576268 24200
rect 6092 22040 6144 22092
rect 6736 22040 6788 22092
rect 6828 22040 6880 22092
rect 6000 21972 6052 22024
rect 576124 21539 576176 21548
rect 576124 21505 576133 21539
rect 576133 21505 576167 21539
rect 576167 21505 576176 21539
rect 576124 21496 576176 21505
rect 576032 21360 576084 21412
rect 576308 21360 576360 21412
rect 575940 20544 575992 20596
rect 576124 20544 576176 20596
rect 575940 20315 575992 20324
rect 575940 20281 575949 20315
rect 575949 20281 575983 20315
rect 575983 20281 575992 20315
rect 575940 20272 575992 20281
rect 576032 19363 576084 19372
rect 576032 19329 576041 19363
rect 576041 19329 576075 19363
rect 576075 19329 576084 19363
rect 576032 19320 576084 19329
rect 575940 17212 575992 17264
rect 576308 17212 576360 17264
rect 575940 16668 575992 16720
rect 6000 12520 6052 12572
rect 6092 12452 6144 12504
rect 6736 12452 6788 12504
rect 6828 12452 6880 12504
rect 4804 11976 4856 12028
rect 4804 11772 4856 11824
rect 576124 7760 576176 7812
rect 9404 7692 9456 7744
rect 17224 7692 17276 7744
rect 58808 7692 58860 7744
rect 576216 7692 576268 7744
rect 1676 7624 1728 7676
rect 576308 7624 576360 7676
rect 572 7556 624 7608
rect 575756 7556 575808 7608
rect 69480 7531 69532 7540
rect 69480 7497 69489 7531
rect 69489 7497 69523 7531
rect 69523 7497 69532 7531
rect 69480 7488 69532 7497
rect 575112 7488 575164 7540
rect 575940 7488 575992 7540
rect 575020 7420 575072 7472
rect 575480 7420 575532 7472
rect 52736 6808 52788 6860
rect 580540 6808 580592 6860
rect 62948 6740 63000 6792
rect 580448 6740 580500 6792
rect 73068 6672 73120 6724
rect 580356 6672 580408 6724
rect 83280 6604 83332 6656
rect 580264 6604 580316 6656
rect 90916 6536 90968 6588
rect 577044 6536 577096 6588
rect 83832 6468 83884 6520
rect 577136 6468 577188 6520
rect 77852 6400 77904 6452
rect 578516 6400 578568 6452
rect 6460 6332 6512 6384
rect 65984 6332 66036 6384
rect 73068 6332 73120 6384
rect 577228 6332 577280 6384
rect 63592 6264 63644 6316
rect 578608 6264 578660 6316
rect 30288 6196 30340 6248
rect 578884 6196 578936 6248
rect 21916 6128 21968 6180
rect 578976 6128 579028 6180
rect 94504 6060 94556 6112
rect 576952 6060 577004 6112
rect 101588 5992 101640 6044
rect 576860 5992 576912 6044
rect 106372 5924 106424 5976
rect 578424 5924 578476 5976
rect 7104 5856 7156 5908
rect 115940 5856 115992 5908
rect 119436 5856 119488 5908
rect 578792 5856 578844 5908
rect 9312 5788 9364 5840
rect 123024 5788 123076 5840
rect 7196 5720 7248 5772
rect 108764 5720 108816 5772
rect 6184 5448 6236 5500
rect 12072 5448 12124 5500
rect 96896 5448 96948 5500
rect 327540 5448 327592 5500
rect 7564 5380 7616 5432
rect 32404 5380 32456 5432
rect 103980 5380 104032 5432
rect 347964 5380 348016 5432
rect 14188 5312 14240 5364
rect 99380 5312 99432 5364
rect 111156 5312 111208 5364
rect 368296 5312 368348 5364
rect 15200 5244 15252 5296
rect 104256 5244 104308 5296
rect 118240 5244 118292 5296
rect 388628 5244 388680 5296
rect 19524 5176 19576 5228
rect 113824 5176 113876 5228
rect 125416 5176 125468 5228
rect 409052 5176 409104 5228
rect 3424 5108 3476 5160
rect 42524 5108 42576 5160
rect 51632 5108 51684 5160
rect 439596 5108 439648 5160
rect 55220 5040 55272 5092
rect 449716 5040 449768 5092
rect 7380 4972 7432 5024
rect 26700 4972 26752 5024
rect 62396 4972 62448 5024
rect 459928 4972 459980 5024
rect 7288 4904 7340 4956
rect 33876 4904 33928 4956
rect 80244 4904 80296 4956
rect 480260 4904 480312 4956
rect 6920 4836 6972 4888
rect 67180 4836 67232 4888
rect 98092 4836 98144 4888
rect 500592 4836 500644 4888
rect 6368 4768 6420 4820
rect 40960 4768 41012 4820
rect 52828 4768 52880 4820
rect 551560 4768 551612 4820
rect 6276 4700 6328 4752
rect 22192 4700 22244 4752
rect 89720 4700 89772 4752
rect 307208 4700 307260 4752
rect 82636 4632 82688 4684
rect 286876 4632 286928 4684
rect 75460 4564 75512 4616
rect 266544 4564 266596 4616
rect 68284 4496 68336 4548
rect 246120 4496 246172 4548
rect 64788 4428 64840 4480
rect 236000 4428 236052 4480
rect 57612 4360 57664 4412
rect 215576 4360 215628 4412
rect 54024 4292 54076 4344
rect 205456 4292 205508 4344
rect 43352 4224 43404 4276
rect 174912 4224 174964 4276
rect 7472 4156 7524 4208
rect 12440 4156 12492 4208
rect 36176 4156 36228 4208
rect 154580 4156 154632 4208
rect 6552 4088 6604 4140
rect 88524 4088 88576 4140
rect 93308 4088 93360 4140
rect 317420 4088 317472 4140
rect 6644 4020 6696 4072
rect 7012 4020 7064 4072
rect 10048 4020 10100 4072
rect 93492 4020 93544 4072
rect 100484 4020 100536 4072
rect 337752 4020 337804 4072
rect 92112 3952 92164 4004
rect 107568 3952 107620 4004
rect 358084 3952 358136 4004
rect 6736 3884 6788 3936
rect 95700 3884 95752 3936
rect 99380 3884 99432 3936
rect 112352 3884 112404 3936
rect 114744 3884 114796 3936
rect 378508 3884 378560 3936
rect 5356 3816 5408 3868
rect 2872 3748 2924 3800
rect 9128 3816 9180 3868
rect 14832 3816 14884 3868
rect 103612 3816 103664 3868
rect 104256 3816 104308 3868
rect 105176 3816 105228 3868
rect 121828 3816 121880 3868
rect 398840 3816 398892 3868
rect 16028 3748 16080 3800
rect 37372 3748 37424 3800
rect 419172 3748 419224 3800
rect 27896 3680 27948 3732
rect 44548 3680 44600 3732
rect 429384 3680 429436 3732
rect 5080 3612 5132 3664
rect 74264 3612 74316 3664
rect 76656 3612 76708 3664
rect 470048 3612 470100 3664
rect 5172 3544 5224 3596
rect 81440 3544 81492 3596
rect 87328 3544 87380 3596
rect 490472 3544 490524 3596
rect 5448 3476 5500 3528
rect 6460 3476 6512 3528
rect 4804 3408 4856 3460
rect 18328 3476 18380 3528
rect 24308 3476 24360 3528
rect 124036 3476 124088 3528
rect 124220 3476 124272 3528
rect 578240 3476 578292 3528
rect 7656 3408 7708 3460
rect 9036 3408 9088 3460
rect 13636 3408 13688 3460
rect 521016 3408 521068 3460
rect 4988 3340 5040 3392
rect 70676 3340 70728 3392
rect 86132 3340 86184 3392
rect 297088 3340 297140 3392
rect 9496 3272 9548 3324
rect 60004 3272 60056 3324
rect 79048 3272 79100 3324
rect 276664 3272 276716 3324
rect 9588 3204 9640 3256
rect 56416 3204 56468 3256
rect 71872 3204 71924 3256
rect 256332 3204 256384 3256
rect 4896 3136 4948 3188
rect 45744 3136 45796 3188
rect 46940 3136 46992 3188
rect 4068 3068 4120 3120
rect 8944 3068 8996 3120
rect 9680 3068 9732 3120
rect 49332 3068 49384 3120
rect 9772 3000 9824 3052
rect 48136 3000 48188 3052
rect 61200 3136 61252 3188
rect 225788 3136 225840 3188
rect 50528 3068 50580 3120
rect 195244 3068 195296 3120
rect 185032 3000 185084 3052
rect 4712 2932 4764 2984
rect 38568 2932 38620 2984
rect 39764 2932 39816 2984
rect 164700 2932 164752 2984
rect 32680 2864 32732 2916
rect 144368 2864 144420 2916
rect 29092 2796 29144 2848
rect 134156 2796 134208 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 40512 700466 40540 703520
rect 84108 700528 84160 700534
rect 84108 700470 84160 700476
rect 40500 700460 40552 700466
rect 40500 700402 40552 700408
rect 41328 700460 41380 700466
rect 41328 700402 41380 700408
rect 62028 700460 62080 700466
rect 62028 700402 62080 700408
rect 39948 700392 40000 700398
rect 39948 700334 40000 700340
rect 19248 700324 19300 700330
rect 19248 700266 19300 700272
rect 19260 689994 19288 700266
rect 17960 689988 18012 689994
rect 17960 689930 18012 689936
rect 19248 689988 19300 689994
rect 19248 689930 19300 689936
rect 9496 689444 9548 689450
rect 9496 689386 9548 689392
rect 9128 689240 9180 689246
rect 9128 689182 9180 689188
rect 9036 689172 9088 689178
rect 9036 689114 9088 689120
rect 8944 688900 8996 688906
rect 8944 688842 8996 688848
rect 3330 682272 3386 682281
rect 3330 682207 3386 682216
rect 3344 681766 3372 682207
rect 3332 681760 3384 681766
rect 3332 681702 3384 681708
rect 6184 681760 6236 681766
rect 6184 681702 6236 681708
rect 5446 675336 5502 675345
rect 5446 675271 5502 675280
rect 5354 653440 5410 653449
rect 5354 653375 5410 653384
rect 3146 624880 3202 624889
rect 3146 624815 3202 624824
rect 3160 624238 3188 624815
rect 3148 624232 3200 624238
rect 3148 624174 3200 624180
rect 4066 567352 4122 567361
rect 4066 567287 4068 567296
rect 4120 567287 4122 567296
rect 4068 567258 4120 567264
rect 5262 543960 5318 543969
rect 5262 543895 5318 543904
rect 5170 521792 5226 521801
rect 5170 521727 5226 521736
rect 3422 509960 3478 509969
rect 3422 509895 3478 509904
rect 3330 208176 3386 208185
rect 3330 208111 3386 208120
rect 3240 171148 3292 171154
rect 3240 171090 3292 171096
rect 3252 122097 3280 171090
rect 3344 128314 3372 208111
rect 3332 128308 3384 128314
rect 3332 128250 3384 128256
rect 3238 122088 3294 122097
rect 3238 122023 3294 122032
rect 1676 7676 1728 7682
rect 1676 7618 1728 7624
rect 572 7608 624 7614
rect 572 7550 624 7556
rect 584 480 612 7550
rect 1688 480 1716 7618
rect 3436 5166 3464 509895
rect 5078 499896 5134 499905
rect 5078 499831 5134 499840
rect 4986 455968 5042 455977
rect 4986 455903 5042 455912
rect 3514 452432 3570 452441
rect 3514 452367 3570 452376
rect 3528 18601 3556 452367
rect 4894 434072 4950 434081
rect 4894 434007 4950 434016
rect 3606 395040 3662 395049
rect 3606 394975 3662 394984
rect 3620 39953 3648 394975
rect 4802 390688 4858 390697
rect 4802 390623 4858 390632
rect 3698 337512 3754 337521
rect 3698 337447 3754 337456
rect 3712 62121 3740 337447
rect 3790 294400 3846 294409
rect 3790 294335 3846 294344
rect 3804 84153 3832 294335
rect 3974 251288 4030 251297
rect 3974 251223 4030 251232
rect 3882 215384 3938 215393
rect 3882 215319 3938 215328
rect 3790 84144 3846 84153
rect 3790 84079 3846 84088
rect 3698 62112 3754 62121
rect 3698 62047 3754 62056
rect 3606 39944 3662 39953
rect 3606 39879 3662 39888
rect 3896 35873 3924 215319
rect 3988 106049 4016 251223
rect 4066 193352 4122 193361
rect 4066 193287 4122 193296
rect 3974 106040 4030 106049
rect 3974 105975 4030 105984
rect 4080 78985 4108 193287
rect 4710 171184 4766 171193
rect 4710 171119 4712 171128
rect 4764 171119 4766 171128
rect 4712 171090 4764 171096
rect 4710 165064 4766 165073
rect 4710 164999 4766 165008
rect 4724 150113 4752 164999
rect 4710 150104 4766 150113
rect 4710 150039 4766 150048
rect 4160 128308 4212 128314
rect 4160 128250 4212 128256
rect 4172 128217 4200 128250
rect 4158 128208 4214 128217
rect 4158 128143 4214 128152
rect 4066 78976 4122 78985
rect 4066 78911 4122 78920
rect 3882 35864 3938 35873
rect 3882 35799 3938 35808
rect 3514 18592 3570 18601
rect 3514 18527 3570 18536
rect 4816 12034 4844 390623
rect 4804 12028 4856 12034
rect 4804 11970 4856 11976
rect 4908 11914 4936 434007
rect 4724 11886 4936 11914
rect 3424 5160 3476 5166
rect 3424 5102 3476 5108
rect 2872 3800 2924 3806
rect 2872 3742 2924 3748
rect 2884 480 2912 3742
rect 4068 3120 4120 3126
rect 4068 3062 4120 3068
rect 4080 480 4108 3062
rect 4724 2990 4752 11886
rect 4804 11824 4856 11830
rect 5000 11778 5028 455903
rect 4804 11766 4856 11772
rect 4816 3466 4844 11766
rect 4908 11750 5028 11778
rect 4804 3460 4856 3466
rect 4804 3402 4856 3408
rect 4908 3194 4936 11750
rect 5092 5522 5120 499831
rect 5000 5494 5120 5522
rect 5000 3398 5028 5494
rect 5184 5386 5212 521727
rect 5092 5358 5212 5386
rect 5092 3670 5120 5358
rect 5276 5250 5304 543895
rect 5184 5222 5304 5250
rect 5080 3664 5132 3670
rect 5080 3606 5132 3612
rect 5184 3602 5212 5222
rect 5262 4856 5318 4865
rect 5262 4791 5318 4800
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 4896 3188 4948 3194
rect 4896 3130 4948 3136
rect 4712 2984 4764 2990
rect 4712 2926 4764 2932
rect 5276 480 5304 4791
rect 5368 3874 5396 653375
rect 5356 3868 5408 3874
rect 5356 3810 5408 3816
rect 5460 3534 5488 675271
rect 6092 331152 6144 331158
rect 6092 331094 6144 331100
rect 6104 321706 6132 331094
rect 6092 321700 6144 321706
rect 6092 321642 6144 321648
rect 6092 311840 6144 311846
rect 6092 311782 6144 311788
rect 6104 302258 6132 311782
rect 6092 302252 6144 302258
rect 6092 302194 6144 302200
rect 6092 292528 6144 292534
rect 6092 292470 6144 292476
rect 6000 292460 6052 292466
rect 6000 292402 6052 292408
rect 6012 283014 6040 292402
rect 6000 283008 6052 283014
rect 6000 282950 6052 282956
rect 6104 282946 6132 292470
rect 6092 282940 6144 282946
rect 6092 282882 6144 282888
rect 6092 273216 6144 273222
rect 6092 273158 6144 273164
rect 6000 273148 6052 273154
rect 6000 273090 6052 273096
rect 6012 263702 6040 273090
rect 6000 263696 6052 263702
rect 6000 263638 6052 263644
rect 6104 263634 6132 273158
rect 6092 263628 6144 263634
rect 6092 263570 6144 263576
rect 6092 253904 6144 253910
rect 6092 253846 6144 253852
rect 6000 253836 6052 253842
rect 6000 253778 6052 253784
rect 6012 244390 6040 253778
rect 6000 244384 6052 244390
rect 6000 244326 6052 244332
rect 6104 244322 6132 253846
rect 6092 244316 6144 244322
rect 6092 244258 6144 244264
rect 6092 234592 6144 234598
rect 6092 234534 6144 234540
rect 6000 234524 6052 234530
rect 6000 234466 6052 234472
rect 6012 225078 6040 234466
rect 6000 225072 6052 225078
rect 6000 225014 6052 225020
rect 6104 225010 6132 234534
rect 6092 225004 6144 225010
rect 6092 224946 6144 224952
rect 6092 215280 6144 215286
rect 6092 215222 6144 215228
rect 6000 215212 6052 215218
rect 6000 215154 6052 215160
rect 6012 205766 6040 215154
rect 6000 205760 6052 205766
rect 6000 205702 6052 205708
rect 6104 205698 6132 215222
rect 6092 205692 6144 205698
rect 6092 205634 6144 205640
rect 6092 195968 6144 195974
rect 6092 195910 6144 195916
rect 6000 195900 6052 195906
rect 6000 195842 6052 195848
rect 6012 186454 6040 195842
rect 6000 186448 6052 186454
rect 6000 186390 6052 186396
rect 6104 186386 6132 195910
rect 6092 186380 6144 186386
rect 6092 186322 6144 186328
rect 6092 176656 6144 176662
rect 6092 176598 6144 176604
rect 6000 176588 6052 176594
rect 6000 176530 6052 176536
rect 6012 167142 6040 176530
rect 6000 167136 6052 167142
rect 6000 167078 6052 167084
rect 6104 167074 6132 176598
rect 6092 167068 6144 167074
rect 6092 167010 6144 167016
rect 6092 157344 6144 157350
rect 6092 157286 6144 157292
rect 6000 157276 6052 157282
rect 6000 157218 6052 157224
rect 6012 147762 6040 157218
rect 6000 147756 6052 147762
rect 6000 147698 6052 147704
rect 6104 147694 6132 157286
rect 6092 147688 6144 147694
rect 6092 147630 6144 147636
rect 6092 137964 6144 137970
rect 6092 137906 6144 137912
rect 6000 137896 6052 137902
rect 6000 137838 6052 137844
rect 6012 128450 6040 137838
rect 6000 128444 6052 128450
rect 6000 128386 6052 128392
rect 6104 128382 6132 137906
rect 6092 128376 6144 128382
rect 6092 128318 6144 128324
rect 6092 118652 6144 118658
rect 6092 118594 6144 118600
rect 6000 118584 6052 118590
rect 6000 118526 6052 118532
rect 6012 109138 6040 118526
rect 6000 109132 6052 109138
rect 6000 109074 6052 109080
rect 6104 109070 6132 118594
rect 6092 109064 6144 109070
rect 6092 109006 6144 109012
rect 6092 99340 6144 99346
rect 6092 99282 6144 99288
rect 6000 99272 6052 99278
rect 6000 99214 6052 99220
rect 6012 89826 6040 99214
rect 6000 89820 6052 89826
rect 6000 89762 6052 89768
rect 6104 89758 6132 99282
rect 6092 89752 6144 89758
rect 6092 89694 6144 89700
rect 6092 80028 6144 80034
rect 6092 79970 6144 79976
rect 6000 79960 6052 79966
rect 6000 79902 6052 79908
rect 6012 70514 6040 79902
rect 6000 70508 6052 70514
rect 6000 70450 6052 70456
rect 6104 70446 6132 79970
rect 6092 70440 6144 70446
rect 6092 70382 6144 70388
rect 6092 60716 6144 60722
rect 6092 60658 6144 60664
rect 6000 60648 6052 60654
rect 6000 60590 6052 60596
rect 6012 51202 6040 60590
rect 6000 51196 6052 51202
rect 6000 51138 6052 51144
rect 6104 51134 6132 60658
rect 6092 51128 6144 51134
rect 6092 51070 6144 51076
rect 6092 41404 6144 41410
rect 6092 41346 6144 41352
rect 6000 41336 6052 41342
rect 6000 41278 6052 41284
rect 6012 31890 6040 41278
rect 6000 31884 6052 31890
rect 6000 31826 6052 31832
rect 6104 31822 6132 41346
rect 6092 31816 6144 31822
rect 6092 31758 6144 31764
rect 6092 22092 6144 22098
rect 6092 22034 6144 22040
rect 6000 22024 6052 22030
rect 6000 21966 6052 21972
rect 6012 12578 6040 21966
rect 6000 12572 6052 12578
rect 6000 12514 6052 12520
rect 6104 12510 6132 22034
rect 6092 12504 6144 12510
rect 6092 12446 6144 12452
rect 6196 5506 6224 681702
rect 6918 631544 6974 631553
rect 6918 631479 6974 631488
rect 6932 627978 6960 631479
rect 6736 627972 6788 627978
rect 6736 627914 6788 627920
rect 6920 627972 6972 627978
rect 6920 627914 6972 627920
rect 6276 624232 6328 624238
rect 6276 624174 6328 624180
rect 6184 5500 6236 5506
rect 6184 5442 6236 5448
rect 6288 4758 6316 624174
rect 6748 621110 6776 627914
rect 6736 621104 6788 621110
rect 6736 621046 6788 621052
rect 6644 618316 6696 618322
rect 6644 618258 6696 618264
rect 6656 618186 6684 618258
rect 6644 618180 6696 618186
rect 6644 618122 6696 618128
rect 6734 610124 6790 610133
rect 6734 610059 6790 610068
rect 6552 608660 6604 608666
rect 6552 608602 6604 608608
rect 6564 601798 6592 608602
rect 6552 601792 6604 601798
rect 6552 601734 6604 601740
rect 6552 601656 6604 601662
rect 6552 601598 6604 601604
rect 6460 601588 6512 601594
rect 6460 601530 6512 601536
rect 6472 591938 6500 601530
rect 6564 592142 6592 601598
rect 6748 601594 6776 610059
rect 6920 601792 6972 601798
rect 6920 601734 6972 601740
rect 6932 601662 6960 601734
rect 6920 601656 6972 601662
rect 6920 601598 6972 601604
rect 6736 601588 6788 601594
rect 6736 601530 6788 601536
rect 6552 592136 6604 592142
rect 6552 592078 6604 592084
rect 6552 592000 6604 592006
rect 6552 591942 6604 591948
rect 6460 591932 6512 591938
rect 6460 591874 6512 591880
rect 6564 582418 6592 591942
rect 6736 591932 6788 591938
rect 6736 591874 6788 591880
rect 6642 588228 6698 588237
rect 6642 588163 6698 588172
rect 6552 582412 6604 582418
rect 6552 582354 6604 582360
rect 6368 582276 6420 582282
rect 6368 582218 6420 582224
rect 6380 572490 6408 582218
rect 6368 572484 6420 572490
rect 6368 572426 6420 572432
rect 6550 566332 6606 566341
rect 6550 566267 6606 566276
rect 6460 563100 6512 563106
rect 6460 563042 6512 563048
rect 6368 563032 6420 563038
rect 6368 562974 6420 562980
rect 6380 553518 6408 562974
rect 6368 553512 6420 553518
rect 6368 553454 6420 553460
rect 6472 553450 6500 563042
rect 6460 553444 6512 553450
rect 6460 553386 6512 553392
rect 6460 553308 6512 553314
rect 6460 553250 6512 553256
rect 6472 543862 6500 553250
rect 6460 543856 6512 543862
rect 6460 543798 6512 543804
rect 6368 543720 6420 543726
rect 6368 543662 6420 543668
rect 6458 543688 6514 543697
rect 6380 534206 6408 543662
rect 6458 543623 6514 543632
rect 6368 534200 6420 534206
rect 6368 534142 6420 534148
rect 6472 534138 6500 543623
rect 6460 534132 6512 534138
rect 6460 534074 6512 534080
rect 6460 533996 6512 534002
rect 6460 533938 6512 533944
rect 6472 524482 6500 533938
rect 6460 524476 6512 524482
rect 6460 524418 6512 524424
rect 6458 524376 6514 524385
rect 6458 524311 6514 524320
rect 6472 514826 6500 524311
rect 6460 514820 6512 514826
rect 6460 514762 6512 514768
rect 6460 514684 6512 514690
rect 6460 514626 6512 514632
rect 6472 505170 6500 514626
rect 6460 505164 6512 505170
rect 6460 505106 6512 505112
rect 6458 505064 6514 505073
rect 6458 504999 6514 505008
rect 6472 495514 6500 504999
rect 6460 495508 6512 495514
rect 6460 495450 6512 495456
rect 6460 495372 6512 495378
rect 6460 495314 6512 495320
rect 6472 485858 6500 495314
rect 6460 485852 6512 485858
rect 6460 485794 6512 485800
rect 6458 485752 6514 485761
rect 6458 485687 6514 485696
rect 6472 476134 6500 485687
rect 6460 476128 6512 476134
rect 6460 476070 6512 476076
rect 6458 466440 6514 466449
rect 6458 466375 6514 466384
rect 6472 456822 6500 466375
rect 6460 456816 6512 456822
rect 6460 456758 6512 456764
rect 6458 447128 6514 447137
rect 6458 447063 6514 447072
rect 6472 437510 6500 447063
rect 6460 437504 6512 437510
rect 6460 437446 6512 437452
rect 6458 408504 6514 408513
rect 6458 408439 6514 408448
rect 6472 398886 6500 408439
rect 6460 398880 6512 398886
rect 6460 398822 6512 398828
rect 6460 389156 6512 389162
rect 6460 389098 6512 389104
rect 6368 389088 6420 389094
rect 6368 389030 6420 389036
rect 6380 379642 6408 389030
rect 6368 379636 6420 379642
rect 6368 379578 6420 379584
rect 6472 379574 6500 389098
rect 6460 379568 6512 379574
rect 6460 379510 6512 379516
rect 6460 369844 6512 369850
rect 6460 369786 6512 369792
rect 6368 369776 6420 369782
rect 6368 369718 6420 369724
rect 6380 360330 6408 369718
rect 6368 360324 6420 360330
rect 6368 360266 6420 360272
rect 6472 360262 6500 369786
rect 6460 360256 6512 360262
rect 6460 360198 6512 360204
rect 6460 350532 6512 350538
rect 6460 350474 6512 350480
rect 6368 350464 6420 350470
rect 6368 350406 6420 350412
rect 6380 341018 6408 350406
rect 6368 341012 6420 341018
rect 6368 340954 6420 340960
rect 6472 340950 6500 350474
rect 6460 340944 6512 340950
rect 6460 340886 6512 340892
rect 6368 331220 6420 331226
rect 6368 331162 6420 331168
rect 6380 321638 6408 331162
rect 6458 324456 6514 324465
rect 6458 324391 6514 324400
rect 6368 321632 6420 321638
rect 6368 321574 6420 321580
rect 6368 311772 6420 311778
rect 6368 311714 6420 311720
rect 6380 302802 6408 311714
rect 6368 302796 6420 302802
rect 6368 302738 6420 302744
rect 6366 302696 6422 302705
rect 6366 302631 6422 302640
rect 6380 4826 6408 302631
rect 6472 6390 6500 324391
rect 6460 6384 6512 6390
rect 6460 6326 6512 6332
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 6276 4752 6328 4758
rect 6276 4694 6328 4700
rect 6564 4146 6592 566267
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 6656 4078 6684 588163
rect 6748 582282 6776 591874
rect 6920 582412 6972 582418
rect 6920 582354 6972 582360
rect 6736 582276 6788 582282
rect 6736 582218 6788 582224
rect 6932 582162 6960 582354
rect 6748 582134 6960 582162
rect 6748 572898 6776 582134
rect 6736 572892 6788 572898
rect 6736 572834 6788 572840
rect 6828 572484 6880 572490
rect 6828 572426 6880 572432
rect 6736 572416 6788 572422
rect 6736 572358 6788 572364
rect 6748 563122 6776 572358
rect 6840 563242 6868 572426
rect 7564 567316 7616 567322
rect 7564 567258 7616 567264
rect 6828 563236 6880 563242
rect 6828 563178 6880 563184
rect 6748 563094 6960 563122
rect 6932 563038 6960 563094
rect 6920 563032 6972 563038
rect 6920 562974 6972 562980
rect 6736 553444 6788 553450
rect 6736 553386 6788 553392
rect 6828 553444 6880 553450
rect 6828 553386 6880 553392
rect 6748 543697 6776 553386
rect 6840 553314 6868 553386
rect 6828 553308 6880 553314
rect 6828 553250 6880 553256
rect 6920 543856 6972 543862
rect 6920 543798 6972 543804
rect 6932 543726 6960 543798
rect 6920 543720 6972 543726
rect 6734 543688 6790 543697
rect 6920 543662 6972 543668
rect 6734 543623 6790 543632
rect 6736 534132 6788 534138
rect 6736 534074 6788 534080
rect 6828 534132 6880 534138
rect 6828 534074 6880 534080
rect 6748 524385 6776 534074
rect 6840 534002 6868 534074
rect 6828 533996 6880 534002
rect 6828 533938 6880 533944
rect 6920 524476 6972 524482
rect 6920 524418 6972 524424
rect 6734 524376 6790 524385
rect 6734 524311 6790 524320
rect 6932 524226 6960 524418
rect 6748 524198 6960 524226
rect 6748 514962 6776 524198
rect 6736 514956 6788 514962
rect 6736 514898 6788 514904
rect 6736 514820 6788 514826
rect 6736 514762 6788 514768
rect 6828 514820 6880 514826
rect 6828 514762 6880 514768
rect 6748 505073 6776 514762
rect 6840 514690 6868 514762
rect 6828 514684 6880 514690
rect 6828 514626 6880 514632
rect 6920 505164 6972 505170
rect 6920 505106 6972 505112
rect 6734 505064 6790 505073
rect 6734 504999 6790 505008
rect 6932 504914 6960 505106
rect 6748 504886 6960 504914
rect 6748 495650 6776 504886
rect 6736 495644 6788 495650
rect 6736 495586 6788 495592
rect 6736 495508 6788 495514
rect 6736 495450 6788 495456
rect 6828 495508 6880 495514
rect 6828 495450 6880 495456
rect 6748 485761 6776 495450
rect 6840 495378 6868 495450
rect 6828 495372 6880 495378
rect 6828 495314 6880 495320
rect 6920 485852 6972 485858
rect 6920 485794 6972 485800
rect 6734 485752 6790 485761
rect 6734 485687 6790 485696
rect 6932 485602 6960 485794
rect 6748 485574 6960 485602
rect 6748 476270 6776 485574
rect 6918 478000 6974 478009
rect 6918 477935 6974 477944
rect 6736 476264 6788 476270
rect 6736 476206 6788 476212
rect 6736 476128 6788 476134
rect 6736 476070 6788 476076
rect 6828 476128 6880 476134
rect 6828 476070 6880 476076
rect 6748 466449 6776 476070
rect 6734 466440 6790 466449
rect 6734 466375 6790 466384
rect 6840 466290 6868 476070
rect 6748 466262 6868 466290
rect 6748 456958 6776 466262
rect 6736 456952 6788 456958
rect 6736 456894 6788 456900
rect 6736 456816 6788 456822
rect 6736 456758 6788 456764
rect 6828 456816 6880 456822
rect 6828 456758 6880 456764
rect 6748 447137 6776 456758
rect 6734 447128 6790 447137
rect 6734 447063 6790 447072
rect 6840 446978 6868 456758
rect 6748 446950 6868 446978
rect 6748 437646 6776 446950
rect 6736 437640 6788 437646
rect 6736 437582 6788 437588
rect 6736 437504 6788 437510
rect 6736 437446 6788 437452
rect 6828 437504 6880 437510
rect 6828 437446 6880 437452
rect 6748 408513 6776 437446
rect 6734 408504 6790 408513
rect 6734 408439 6790 408448
rect 6736 398880 6788 398886
rect 6736 398822 6788 398828
rect 6748 389162 6776 398822
rect 6840 389162 6868 437446
rect 6736 389156 6788 389162
rect 6736 389098 6788 389104
rect 6828 389156 6880 389162
rect 6828 389098 6880 389104
rect 6736 379568 6788 379574
rect 6736 379510 6788 379516
rect 6828 379568 6880 379574
rect 6828 379510 6880 379516
rect 6748 369850 6776 379510
rect 6840 369850 6868 379510
rect 6736 369844 6788 369850
rect 6736 369786 6788 369792
rect 6828 369844 6880 369850
rect 6828 369786 6880 369792
rect 6736 360256 6788 360262
rect 6736 360198 6788 360204
rect 6828 360256 6880 360262
rect 6828 360198 6880 360204
rect 6748 350538 6776 360198
rect 6840 350538 6868 360198
rect 6736 350532 6788 350538
rect 6736 350474 6788 350480
rect 6828 350532 6880 350538
rect 6828 350474 6880 350480
rect 6736 340944 6788 340950
rect 6736 340886 6788 340892
rect 6828 340944 6880 340950
rect 6828 340886 6880 340892
rect 6748 331226 6776 340886
rect 6840 331226 6868 340886
rect 6736 331220 6788 331226
rect 6736 331162 6788 331168
rect 6828 331220 6880 331226
rect 6828 331162 6880 331168
rect 6736 321632 6788 321638
rect 6736 321574 6788 321580
rect 6828 321632 6880 321638
rect 6828 321574 6880 321580
rect 6748 311846 6776 321574
rect 6840 311846 6868 321574
rect 6736 311840 6788 311846
rect 6736 311782 6788 311788
rect 6828 311840 6880 311846
rect 6828 311782 6880 311788
rect 6736 302252 6788 302258
rect 6736 302194 6788 302200
rect 6828 302252 6880 302258
rect 6828 302194 6880 302200
rect 6748 292534 6776 302194
rect 6840 292534 6868 302194
rect 6736 292528 6788 292534
rect 6736 292470 6788 292476
rect 6828 292528 6880 292534
rect 6828 292470 6880 292476
rect 6736 282940 6788 282946
rect 6736 282882 6788 282888
rect 6828 282940 6880 282946
rect 6828 282882 6880 282888
rect 6748 273222 6776 282882
rect 6840 273222 6868 282882
rect 6736 273216 6788 273222
rect 6736 273158 6788 273164
rect 6828 273216 6880 273222
rect 6828 273158 6880 273164
rect 6736 263628 6788 263634
rect 6736 263570 6788 263576
rect 6828 263628 6880 263634
rect 6828 263570 6880 263576
rect 6748 253910 6776 263570
rect 6840 253910 6868 263570
rect 6736 253904 6788 253910
rect 6736 253846 6788 253852
rect 6828 253904 6880 253910
rect 6828 253846 6880 253852
rect 6736 244316 6788 244322
rect 6736 244258 6788 244264
rect 6828 244316 6880 244322
rect 6828 244258 6880 244264
rect 6748 234598 6776 244258
rect 6840 234598 6868 244258
rect 6736 234592 6788 234598
rect 6736 234534 6788 234540
rect 6828 234592 6880 234598
rect 6828 234534 6880 234540
rect 6736 225004 6788 225010
rect 6736 224946 6788 224952
rect 6828 225004 6880 225010
rect 6828 224946 6880 224952
rect 6748 215286 6776 224946
rect 6840 215286 6868 224946
rect 6736 215280 6788 215286
rect 6736 215222 6788 215228
rect 6828 215280 6880 215286
rect 6828 215222 6880 215228
rect 6736 205692 6788 205698
rect 6736 205634 6788 205640
rect 6828 205692 6880 205698
rect 6828 205634 6880 205640
rect 6748 195974 6776 205634
rect 6840 195974 6868 205634
rect 6736 195968 6788 195974
rect 6736 195910 6788 195916
rect 6828 195968 6880 195974
rect 6828 195910 6880 195916
rect 6736 186380 6788 186386
rect 6736 186322 6788 186328
rect 6828 186380 6880 186386
rect 6828 186322 6880 186328
rect 6748 176662 6776 186322
rect 6840 176662 6868 186322
rect 6736 176656 6788 176662
rect 6736 176598 6788 176604
rect 6828 176656 6880 176662
rect 6828 176598 6880 176604
rect 6736 167068 6788 167074
rect 6736 167010 6788 167016
rect 6828 167068 6880 167074
rect 6828 167010 6880 167016
rect 6748 157350 6776 167010
rect 6840 157350 6868 167010
rect 6736 157344 6788 157350
rect 6736 157286 6788 157292
rect 6828 157344 6880 157350
rect 6828 157286 6880 157292
rect 6736 147688 6788 147694
rect 6736 147630 6788 147636
rect 6828 147688 6880 147694
rect 6828 147630 6880 147636
rect 6748 137970 6776 147630
rect 6840 137970 6868 147630
rect 6736 137964 6788 137970
rect 6736 137906 6788 137912
rect 6828 137964 6880 137970
rect 6828 137906 6880 137912
rect 6736 128376 6788 128382
rect 6736 128318 6788 128324
rect 6828 128376 6880 128382
rect 6828 128318 6880 128324
rect 6748 118658 6776 128318
rect 6840 118658 6868 128318
rect 6736 118652 6788 118658
rect 6736 118594 6788 118600
rect 6828 118652 6880 118658
rect 6828 118594 6880 118600
rect 6736 109064 6788 109070
rect 6736 109006 6788 109012
rect 6828 109064 6880 109070
rect 6828 109006 6880 109012
rect 6748 99346 6776 109006
rect 6840 99346 6868 109006
rect 6736 99340 6788 99346
rect 6736 99282 6788 99288
rect 6828 99340 6880 99346
rect 6828 99282 6880 99288
rect 6736 89752 6788 89758
rect 6736 89694 6788 89700
rect 6828 89752 6880 89758
rect 6828 89694 6880 89700
rect 6748 80034 6776 89694
rect 6840 80034 6868 89694
rect 6736 80028 6788 80034
rect 6736 79970 6788 79976
rect 6828 80028 6880 80034
rect 6828 79970 6880 79976
rect 6736 70440 6788 70446
rect 6736 70382 6788 70388
rect 6828 70440 6880 70446
rect 6828 70382 6880 70388
rect 6748 60722 6776 70382
rect 6840 60722 6868 70382
rect 6736 60716 6788 60722
rect 6736 60658 6788 60664
rect 6828 60716 6880 60722
rect 6828 60658 6880 60664
rect 6736 51128 6788 51134
rect 6736 51070 6788 51076
rect 6828 51128 6880 51134
rect 6828 51070 6880 51076
rect 6748 41410 6776 51070
rect 6840 41410 6868 51070
rect 6736 41404 6788 41410
rect 6736 41346 6788 41352
rect 6828 41404 6880 41410
rect 6828 41346 6880 41352
rect 6736 31816 6788 31822
rect 6736 31758 6788 31764
rect 6828 31816 6880 31822
rect 6828 31758 6880 31764
rect 6748 22098 6776 31758
rect 6840 22098 6868 31758
rect 6736 22092 6788 22098
rect 6736 22034 6788 22040
rect 6828 22092 6880 22098
rect 6828 22034 6880 22040
rect 6736 12504 6788 12510
rect 6736 12446 6788 12452
rect 6828 12504 6880 12510
rect 6828 12446 6880 12452
rect 6644 4072 6696 4078
rect 6644 4014 6696 4020
rect 6748 3942 6776 12446
rect 6736 3936 6788 3942
rect 6840 3913 6868 12446
rect 6932 4894 6960 477935
rect 7010 412584 7066 412593
rect 7010 412519 7066 412528
rect 6920 4888 6972 4894
rect 6920 4830 6972 4836
rect 7024 4078 7052 412519
rect 7102 368520 7158 368529
rect 7102 368455 7158 368464
rect 7116 5914 7144 368455
rect 7194 346488 7250 346497
rect 7194 346423 7250 346432
rect 7104 5908 7156 5914
rect 7104 5850 7156 5856
rect 7208 5778 7236 346423
rect 7286 280528 7342 280537
rect 7286 280463 7342 280472
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 7300 4962 7328 280463
rect 7378 258632 7434 258641
rect 7378 258567 7434 258576
rect 7392 5030 7420 258567
rect 7470 236600 7526 236609
rect 7470 236535 7526 236544
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 7288 4956 7340 4962
rect 7288 4898 7340 4904
rect 7484 4214 7512 236535
rect 7576 5438 7604 567258
rect 7564 5432 7616 5438
rect 7564 5374 7616 5380
rect 8850 5128 8906 5137
rect 8850 5063 8906 5072
rect 7472 4208 7524 4214
rect 7472 4150 7524 4156
rect 7012 4072 7064 4078
rect 7012 4014 7064 4020
rect 6736 3878 6788 3884
rect 6826 3904 6882 3913
rect 6826 3839 6882 3848
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 6472 480 6500 3470
rect 7656 3460 7708 3466
rect 7656 3402 7708 3408
rect 7668 480 7696 3402
rect 8864 480 8892 5063
rect 8956 3126 8984 688842
rect 9048 3466 9076 689114
rect 9140 3874 9168 689182
rect 9404 689104 9456 689110
rect 9404 689046 9456 689052
rect 9312 686520 9364 686526
rect 9312 686462 9364 686468
rect 9324 5846 9352 686462
rect 9416 7750 9444 689046
rect 9404 7744 9456 7750
rect 9404 7686 9456 7692
rect 9312 5840 9364 5846
rect 9312 5782 9364 5788
rect 9128 3868 9180 3874
rect 9128 3810 9180 3816
rect 9036 3460 9088 3466
rect 9036 3402 9088 3408
rect 9508 3330 9536 689386
rect 9772 689036 9824 689042
rect 9772 688978 9824 688984
rect 9680 688832 9732 688838
rect 9680 688774 9732 688780
rect 9588 688764 9640 688770
rect 9588 688706 9640 688712
rect 9496 3324 9548 3330
rect 9496 3266 9548 3272
rect 9600 3262 9628 688706
rect 9588 3256 9640 3262
rect 9588 3198 9640 3204
rect 9692 3126 9720 688774
rect 8944 3120 8996 3126
rect 8944 3062 8996 3068
rect 9680 3120 9732 3126
rect 9680 3062 9732 3068
rect 9784 3058 9812 688978
rect 17972 686868 18000 689930
rect 39960 686882 39988 700334
rect 41340 689314 41368 700402
rect 41328 689308 41380 689314
rect 41328 689250 41380 689256
rect 62040 686882 62068 700402
rect 84120 686882 84148 700470
rect 105464 699718 105492 703520
rect 170324 700738 170352 703520
rect 150348 700732 150400 700738
rect 150348 700674 150400 700680
rect 170312 700732 170364 700738
rect 170312 700674 170364 700680
rect 128268 700664 128320 700670
rect 128268 700606 128320 700612
rect 106188 700596 106240 700602
rect 106188 700538 106240 700544
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106096 699712 106148 699718
rect 106096 699654 106148 699660
rect 106108 689382 106136 699654
rect 106096 689376 106148 689382
rect 106096 689318 106148 689324
rect 106200 687018 106228 700538
rect 128280 689586 128308 700606
rect 150360 689586 150388 700674
rect 235184 700670 235212 703520
rect 235172 700664 235224 700670
rect 235172 700606 235224 700612
rect 300136 700602 300164 703520
rect 300124 700596 300176 700602
rect 300124 700538 300176 700544
rect 364996 700534 365024 703520
rect 364984 700528 365036 700534
rect 364984 700470 365036 700476
rect 429856 700466 429884 703520
rect 429844 700460 429896 700466
rect 429844 700402 429896 700408
rect 494808 700398 494836 703520
rect 494796 700392 494848 700398
rect 494796 700334 494848 700340
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 127532 689580 127584 689586
rect 127532 689522 127584 689528
rect 128268 689580 128320 689586
rect 128268 689522 128320 689528
rect 149428 689580 149480 689586
rect 149428 689522 149480 689528
rect 150348 689580 150400 689586
rect 150348 689522 150400 689528
rect 105924 686990 106228 687018
rect 105924 686882 105952 686990
rect 39882 686854 39988 686882
rect 61778 686854 62068 686882
rect 83674 686854 84148 686882
rect 105662 686854 105952 686882
rect 127544 686868 127572 689522
rect 149440 686868 149468 689522
rect 456432 689444 456484 689450
rect 456432 689386 456484 689392
rect 171416 689376 171468 689382
rect 171416 689318 171468 689324
rect 171428 686868 171456 689318
rect 193312 689308 193364 689314
rect 193312 689250 193364 689256
rect 193324 686868 193352 689250
rect 237196 689240 237248 689246
rect 237196 689182 237248 689188
rect 215208 688968 215260 688974
rect 215208 688910 215260 688916
rect 215220 686868 215248 688910
rect 237208 686868 237236 689182
rect 259092 689172 259144 689178
rect 259092 689114 259144 689120
rect 259104 686868 259132 689114
rect 280988 689104 281040 689110
rect 280988 689046 281040 689052
rect 281000 686868 281028 689046
rect 302976 689036 303028 689042
rect 302976 688978 303028 688984
rect 302988 686868 303016 688978
rect 390652 688900 390704 688906
rect 390652 688842 390704 688848
rect 346766 688800 346822 688809
rect 346766 688735 346822 688744
rect 346780 686868 346808 688735
rect 390664 686868 390692 688842
rect 412548 688832 412600 688838
rect 412548 688774 412600 688780
rect 412560 686868 412588 688774
rect 434444 688764 434496 688770
rect 434444 688706 434496 688712
rect 434456 686868 434484 688706
rect 456444 686868 456472 689386
rect 576124 688968 576176 688974
rect 544106 688936 544162 688945
rect 576124 688910 576176 688916
rect 544106 688871 544162 688880
rect 522210 688800 522266 688809
rect 522210 688735 522266 688744
rect 478326 688664 478382 688673
rect 478326 688599 478382 688608
rect 500222 688664 500278 688673
rect 500222 688599 500278 688608
rect 478340 686868 478368 688599
rect 500236 686868 500264 688599
rect 522224 686868 522252 688735
rect 544120 686868 544148 688871
rect 368388 686520 368440 686526
rect 324594 686488 324650 686497
rect 324650 686446 324898 686474
rect 368440 686468 368690 686474
rect 368388 686462 368690 686468
rect 368400 686446 368690 686462
rect 324594 686423 324650 686432
rect 565910 686352 565966 686361
rect 565966 686310 566030 686338
rect 565910 686287 565966 686296
rect 575940 674960 575992 674966
rect 575860 674908 575940 674914
rect 575860 674902 575992 674908
rect 575860 674886 575980 674902
rect 575860 669338 575888 674886
rect 575768 669310 575888 669338
rect 575768 652610 575796 669310
rect 575940 652928 575992 652934
rect 575584 652582 575796 652610
rect 575860 652888 575940 652916
rect 575584 652338 575612 652582
rect 575308 652310 575612 652338
rect 575308 647306 575336 652310
rect 575860 647850 575888 652888
rect 575940 652870 575992 652876
rect 575860 647834 575980 647850
rect 575860 647828 575992 647834
rect 575860 647822 575940 647828
rect 575940 647770 575992 647776
rect 575308 647278 575612 647306
rect 575584 644314 575612 647278
rect 575584 644286 575796 644314
rect 575768 625274 575796 644286
rect 576032 634840 576084 634846
rect 576032 634782 576084 634788
rect 576044 630578 576072 634782
rect 575584 625246 575796 625274
rect 575952 630550 576072 630578
rect 575584 623098 575612 625246
rect 575308 623070 575612 623098
rect 575308 608546 575336 623070
rect 575952 621738 575980 630550
rect 575860 621710 575980 621738
rect 575860 608546 575888 621710
rect 575308 608518 575704 608546
rect 575676 602290 575704 608518
rect 575768 608518 575888 608546
rect 575768 607186 575796 608518
rect 575768 607158 575888 607186
rect 575860 606914 575888 607158
rect 575860 606886 575980 606914
rect 575952 602410 575980 606886
rect 575940 602404 575992 602410
rect 575940 602346 575992 602352
rect 575676 602262 575796 602290
rect 575768 591682 575796 602262
rect 576032 597576 576084 597582
rect 576032 597518 576084 597524
rect 575584 591654 575796 591682
rect 575584 581618 575612 591654
rect 575492 581590 575612 581618
rect 575492 562986 575520 581590
rect 576044 576994 576072 597518
rect 575952 576966 576072 576994
rect 575952 567254 575980 576966
rect 575940 567248 575992 567254
rect 575940 567190 575992 567196
rect 575940 567112 575992 567118
rect 575940 567054 575992 567060
rect 575952 564398 575980 567054
rect 575940 564392 575992 564398
rect 575940 564334 575992 564340
rect 575492 562958 575796 562986
rect 575768 556050 575796 562958
rect 575492 556022 575796 556050
rect 575492 543674 575520 556022
rect 576032 554804 576084 554810
rect 576032 554746 576084 554752
rect 576044 551154 576072 554746
rect 575952 551126 576072 551154
rect 575952 546394 575980 551126
rect 575952 546366 576072 546394
rect 575492 543646 575612 543674
rect 575584 540954 575612 543646
rect 575584 540926 575704 540954
rect 575676 522322 575704 540926
rect 576044 536858 576072 546366
rect 575940 536852 575992 536858
rect 575940 536794 575992 536800
rect 576032 536852 576084 536858
rect 576032 536794 576084 536800
rect 575952 528578 575980 536794
rect 575952 528550 576072 528578
rect 575676 522306 575980 522322
rect 575676 522300 575992 522306
rect 575676 522294 575940 522300
rect 575940 522242 575992 522248
rect 575940 519988 575992 519994
rect 575940 519930 575992 519936
rect 575952 518242 575980 519930
rect 575584 518214 575980 518242
rect 575584 514842 575612 518214
rect 575940 518016 575992 518022
rect 575860 517964 575940 517970
rect 575860 517958 575992 517964
rect 575860 517942 575980 517958
rect 575584 514814 575704 514842
rect 575676 510218 575704 514814
rect 575860 514740 575888 517942
rect 576044 514758 576072 528550
rect 575940 514752 575992 514758
rect 575860 514712 575940 514740
rect 575940 514694 575992 514700
rect 576032 514752 576084 514758
rect 576032 514694 576084 514700
rect 575676 510190 576072 510218
rect 575940 509516 575992 509522
rect 575940 509458 575992 509464
rect 575952 509402 575980 509458
rect 575492 509374 575980 509402
rect 575492 505050 575520 509374
rect 575940 505368 575992 505374
rect 575400 505022 575520 505050
rect 575860 505328 575940 505356
rect 575400 504778 575428 505022
rect 575400 504750 575520 504778
rect 575492 495122 575520 504750
rect 575860 503418 575888 505328
rect 575940 505310 575992 505316
rect 575584 503390 575888 503418
rect 575584 495258 575612 503390
rect 576044 503146 576072 510190
rect 575676 503118 576072 503146
rect 575676 495394 575704 503118
rect 575676 495366 576072 495394
rect 575584 495230 575980 495258
rect 575492 495094 575612 495122
rect 575584 486962 575612 495094
rect 575952 487830 575980 495230
rect 576044 492658 576072 495366
rect 576032 492652 576084 492658
rect 576032 492594 576084 492600
rect 575940 487824 575992 487830
rect 575940 487766 575992 487772
rect 576136 487150 576164 688910
rect 576306 675336 576362 675345
rect 576306 675271 576362 675280
rect 576320 674966 576348 675271
rect 576308 674960 576360 674966
rect 576308 674902 576360 674908
rect 580262 674656 580318 674665
rect 580262 674591 580318 674600
rect 576306 653440 576362 653449
rect 576306 653375 576362 653384
rect 576320 652934 576348 653375
rect 576308 652928 576360 652934
rect 576308 652870 576360 652876
rect 578238 632088 578294 632097
rect 578238 632023 578294 632032
rect 576306 521792 576362 521801
rect 576306 521727 576362 521736
rect 576320 519994 576348 521727
rect 576308 519988 576360 519994
rect 576308 519930 576360 519936
rect 576216 514752 576268 514758
rect 576216 514694 576268 514700
rect 576228 505374 576256 514694
rect 576216 505368 576268 505374
rect 576216 505310 576268 505316
rect 576124 487144 576176 487150
rect 576124 487086 576176 487092
rect 575584 486934 575980 486962
rect 575952 485790 575980 486934
rect 575940 485784 575992 485790
rect 575940 485726 575992 485732
rect 576032 485784 576084 485790
rect 576032 485726 576084 485732
rect 575940 485648 575992 485654
rect 575768 485596 575940 485602
rect 575768 485590 575992 485596
rect 575768 485574 575980 485590
rect 575768 483018 575796 485574
rect 575940 485512 575992 485518
rect 575940 485454 575992 485460
rect 575584 482990 575796 483018
rect 575584 475946 575612 482990
rect 575952 476218 575980 485454
rect 575676 476190 575980 476218
rect 575676 476082 575704 476190
rect 575676 476054 575888 476082
rect 575584 475918 575704 475946
rect 575676 456770 575704 475918
rect 575860 468466 575888 476054
rect 575860 468438 575980 468466
rect 575952 466546 575980 468438
rect 575940 466540 575992 466546
rect 575940 466482 575992 466488
rect 576044 466478 576072 485726
rect 576032 466472 576084 466478
rect 576032 466414 576084 466420
rect 575860 466274 575980 466290
rect 575860 466268 575992 466274
rect 575860 466262 575940 466268
rect 575860 463706 575888 466262
rect 575940 466210 575992 466216
rect 576124 466268 576176 466274
rect 576124 466210 576176 466216
rect 576136 463706 576164 466210
rect 575216 456742 575704 456770
rect 575768 463678 575888 463706
rect 576044 463678 576164 463706
rect 575216 444530 575244 456742
rect 575768 449290 575796 463678
rect 575768 449262 575980 449290
rect 575952 446978 575980 449262
rect 576044 447166 576072 463678
rect 576858 455968 576914 455977
rect 576858 455903 576914 455912
rect 576032 447160 576084 447166
rect 576032 447102 576084 447108
rect 576124 447092 576176 447098
rect 576124 447034 576176 447040
rect 575768 446950 575980 446978
rect 575216 444502 575428 444530
rect 575400 444394 575428 444502
rect 575400 444366 575612 444394
rect 575584 439498 575612 444366
rect 575768 442218 575796 446950
rect 575768 442190 575888 442218
rect 575584 439470 575796 439498
rect 575768 437322 575796 439470
rect 575676 437294 575796 437322
rect 575676 428346 575704 437294
rect 575860 433242 575888 442190
rect 576136 437458 576164 447034
rect 576044 437430 576164 437458
rect 575860 433214 575980 433242
rect 575492 428318 575704 428346
rect 575492 427394 575520 428318
rect 575952 427718 575980 433214
rect 576044 428534 576072 437430
rect 576032 428528 576084 428534
rect 576032 428470 576084 428476
rect 575940 427712 575992 427718
rect 575940 427654 575992 427660
rect 575940 427576 575992 427582
rect 575940 427518 575992 427524
rect 575492 427366 575612 427394
rect 575584 415426 575612 427366
rect 575952 423722 575980 427518
rect 575768 423694 575980 423722
rect 575768 422906 575796 423694
rect 575768 422878 575888 422906
rect 575584 415398 575704 415426
rect 575676 409170 575704 415398
rect 575400 409142 575704 409170
rect 575400 396114 575428 409142
rect 575860 405600 575888 422878
rect 576124 417852 576176 417858
rect 576124 417794 576176 417800
rect 575940 405612 575992 405618
rect 575860 405572 575940 405600
rect 575940 405554 575992 405560
rect 576136 397050 576164 417794
rect 575940 397044 575992 397050
rect 575940 396986 575992 396992
rect 576124 397044 576176 397050
rect 576124 396986 576176 396992
rect 575400 396086 575520 396114
rect 575492 390130 575520 396086
rect 575492 390102 575704 390130
rect 575952 390114 575980 396986
rect 576032 396092 576084 396098
rect 576032 396034 576084 396040
rect 575676 389314 575704 390102
rect 575940 390108 575992 390114
rect 575940 390050 575992 390056
rect 575584 389286 575704 389314
rect 575584 388634 575612 389286
rect 575584 388606 575704 388634
rect 575676 388498 575704 388606
rect 575676 388470 575980 388498
rect 575952 384402 575980 388470
rect 575940 384396 575992 384402
rect 575940 384338 575992 384344
rect 576044 384282 576072 396034
rect 575400 384254 576072 384282
rect 575400 379114 575428 384254
rect 576032 379500 576084 379506
rect 576032 379442 576084 379448
rect 575400 379086 575796 379114
rect 575768 372178 575796 379086
rect 575768 372150 575980 372178
rect 575952 369594 575980 372150
rect 576044 371958 576072 379442
rect 576124 379432 576176 379438
rect 576124 379374 576176 379380
rect 576136 376718 576164 379374
rect 576124 376712 576176 376718
rect 576124 376654 576176 376660
rect 576032 371952 576084 371958
rect 576032 371894 576084 371900
rect 575492 369566 575980 369594
rect 575492 360074 575520 369566
rect 575940 366512 575992 366518
rect 575860 366460 575940 366466
rect 575860 366454 575992 366460
rect 575860 366438 575980 366454
rect 575860 361026 575888 366438
rect 575940 365900 575992 365906
rect 575940 365842 575992 365848
rect 575952 361282 575980 365842
rect 575940 361276 575992 361282
rect 575940 361218 575992 361224
rect 575860 360998 575980 361026
rect 575308 360046 575520 360074
rect 575308 356402 575336 360046
rect 575952 359514 575980 360998
rect 575940 359508 575992 359514
rect 575940 359450 575992 359456
rect 575940 359372 575992 359378
rect 575940 359314 575992 359320
rect 575952 359122 575980 359314
rect 575676 359094 575980 359122
rect 575308 356374 575428 356402
rect 575400 350282 575428 356374
rect 575676 352594 575704 359094
rect 575940 359032 575992 359038
rect 575940 358974 575992 358980
rect 575952 358850 575980 358974
rect 575860 358822 575980 358850
rect 575860 352730 575888 358822
rect 575860 352714 575980 352730
rect 575860 352708 575992 352714
rect 575860 352702 575940 352708
rect 575940 352650 575992 352656
rect 575676 352566 576164 352594
rect 575400 350254 575704 350282
rect 575676 350010 575704 350254
rect 575676 349982 576072 350010
rect 575940 347472 575992 347478
rect 575584 347420 575940 347426
rect 575584 347414 575992 347420
rect 575584 347398 575980 347414
rect 575584 332738 575612 347398
rect 576044 347290 576072 349982
rect 575860 347262 576072 347290
rect 575860 347154 575888 347262
rect 575676 347126 575888 347154
rect 575676 336818 575704 347126
rect 576136 347018 576164 352566
rect 575952 346990 576164 347018
rect 575952 338094 575980 346990
rect 576306 346352 576362 346361
rect 576228 346310 576306 346338
rect 575940 338088 575992 338094
rect 575940 338030 575992 338036
rect 575676 336790 575796 336818
rect 575768 336682 575796 336790
rect 575768 336654 575980 336682
rect 575952 334626 575980 336654
rect 575940 334620 575992 334626
rect 575940 334562 575992 334568
rect 575308 332710 575612 332738
rect 575308 327570 575336 332710
rect 575940 331900 575992 331906
rect 575940 331842 575992 331848
rect 575952 328250 575980 331842
rect 575584 328222 575980 328250
rect 575584 327842 575612 328222
rect 575940 328024 575992 328030
rect 575940 327966 575992 327972
rect 575584 327814 575704 327842
rect 575308 327542 575612 327570
rect 575584 319410 575612 327542
rect 575676 319546 575704 327814
rect 575952 321978 575980 327966
rect 576228 325718 576256 346310
rect 576306 346287 576362 346296
rect 576124 325712 576176 325718
rect 576124 325654 576176 325660
rect 576216 325712 576268 325718
rect 576216 325654 576268 325660
rect 575940 321972 575992 321978
rect 575940 321914 575992 321920
rect 575676 319530 575980 319546
rect 575676 319524 575992 319530
rect 575676 319518 575940 319524
rect 575940 319466 575992 319472
rect 575584 319382 575980 319410
rect 575952 319258 575980 319382
rect 575940 319252 575992 319258
rect 575940 319194 575992 319200
rect 575940 319116 575992 319122
rect 575940 319058 575992 319064
rect 575952 319002 575980 319058
rect 575492 318974 575980 319002
rect 575492 296698 575520 318974
rect 576136 315994 576164 325654
rect 576306 324456 576362 324465
rect 576306 324391 576362 324400
rect 576124 315988 576176 315994
rect 576124 315930 576176 315936
rect 575940 315784 575992 315790
rect 575216 296670 575520 296698
rect 575584 315732 575940 315738
rect 575584 315726 575992 315732
rect 575584 315710 575980 315726
rect 575216 287994 575244 296670
rect 575584 292482 575612 315710
rect 575940 315648 575992 315654
rect 575860 315596 575940 315602
rect 575860 315590 575992 315596
rect 575860 315574 575980 315590
rect 575860 312610 575888 315574
rect 575492 292454 575612 292482
rect 575676 312582 575888 312610
rect 575492 288402 575520 292454
rect 575676 292346 575704 312582
rect 576320 307834 576348 324391
rect 575940 307828 575992 307834
rect 575940 307770 575992 307776
rect 576308 307828 576360 307834
rect 576308 307770 576360 307776
rect 575952 299198 575980 307770
rect 576032 306400 576084 306406
rect 576032 306342 576084 306348
rect 575940 299192 575992 299198
rect 575940 299134 575992 299140
rect 575676 292318 575796 292346
rect 575768 288674 575796 292318
rect 575768 288646 575980 288674
rect 575952 288522 575980 288646
rect 575940 288516 575992 288522
rect 575940 288458 575992 288464
rect 575492 288374 575980 288402
rect 575216 287966 575612 287994
rect 575584 287722 575612 287966
rect 575492 287694 575612 287722
rect 575492 279970 575520 287694
rect 575952 286482 575980 288374
rect 576044 286482 576072 306342
rect 576124 288516 576176 288522
rect 576124 288458 576176 288464
rect 575940 286476 575992 286482
rect 575940 286418 575992 286424
rect 576032 286476 576084 286482
rect 576032 286418 576084 286424
rect 576136 286362 576164 288458
rect 575216 279942 575520 279970
rect 575584 286334 576164 286362
rect 575216 261474 575244 279942
rect 575584 279834 575612 286334
rect 575940 286272 575992 286278
rect 575940 286214 575992 286220
rect 576032 286272 576084 286278
rect 576032 286214 576084 286220
rect 575492 279806 575612 279834
rect 575492 279562 575520 279806
rect 575400 279534 575520 279562
rect 575400 273442 575428 279534
rect 575952 278934 575980 286214
rect 575940 278928 575992 278934
rect 575940 278870 575992 278876
rect 575940 278792 575992 278798
rect 575860 278752 575940 278780
rect 575400 273414 575520 273442
rect 575492 273170 575520 273414
rect 575400 273142 575520 273170
rect 575400 269770 575428 273142
rect 575860 273034 575888 278752
rect 575940 278734 575992 278740
rect 575860 273018 575980 273034
rect 575860 273012 575992 273018
rect 575860 273006 575940 273012
rect 575940 272954 575992 272960
rect 576044 272338 576072 286214
rect 576124 278928 576176 278934
rect 576124 278870 576176 278876
rect 576032 272332 576084 272338
rect 576032 272274 576084 272280
rect 576032 270360 576084 270366
rect 576032 270302 576084 270308
rect 575400 269742 575520 269770
rect 575492 262970 575520 269742
rect 575492 262954 575980 262970
rect 575492 262948 575992 262954
rect 575492 262942 575940 262948
rect 575940 262890 575992 262896
rect 576044 262834 576072 270302
rect 575768 262806 576072 262834
rect 575216 261446 575520 261474
rect 575492 253314 575520 261446
rect 575768 257530 575796 262806
rect 575940 262744 575992 262750
rect 575940 262686 575992 262692
rect 575952 262290 575980 262686
rect 575860 262262 575980 262290
rect 575860 257666 575888 262262
rect 575860 257650 575980 257666
rect 575860 257644 575992 257650
rect 575860 257638 575940 257644
rect 575940 257586 575992 257592
rect 575768 257514 575980 257530
rect 575768 257508 575992 257514
rect 575768 257502 575940 257508
rect 575940 257450 575992 257456
rect 575492 253298 575980 253314
rect 575492 253292 575992 253298
rect 575492 253286 575940 253292
rect 575940 253234 575992 253240
rect 575676 253150 576072 253178
rect 575676 249132 575704 253150
rect 575940 253088 575992 253094
rect 575400 249104 575704 249132
rect 575860 253036 575940 253042
rect 575860 253030 575992 253036
rect 576044 253042 576072 253150
rect 576136 253042 576164 278870
rect 576216 262948 576268 262954
rect 576216 262890 576268 262896
rect 575860 253014 575980 253030
rect 576044 253014 576164 253042
rect 575400 246650 575428 249104
rect 575860 246650 575888 253014
rect 575940 249144 575992 249150
rect 575940 249086 575992 249092
rect 575308 246622 575428 246650
rect 575768 246622 575888 246650
rect 575308 229786 575336 246622
rect 575768 234546 575796 246622
rect 575952 246378 575980 249086
rect 575860 246350 575980 246378
rect 575860 235090 575888 246350
rect 576032 243160 576084 243166
rect 576032 243102 576084 243108
rect 575940 241732 575992 241738
rect 575940 241674 575992 241680
rect 575952 236706 575980 241674
rect 576044 241466 576072 243102
rect 576032 241460 576084 241466
rect 576032 241402 576084 241408
rect 576124 241256 576176 241262
rect 576124 241198 576176 241204
rect 575940 236700 575992 236706
rect 575940 236642 575992 236648
rect 575860 235074 575980 235090
rect 575860 235068 575992 235074
rect 575860 235062 575940 235068
rect 575940 235010 575992 235016
rect 575676 234518 575796 234546
rect 575308 229758 575612 229786
rect 575584 217682 575612 229758
rect 575032 217654 575612 217682
rect 575032 202314 575060 217654
rect 575676 217648 575704 234518
rect 576032 234320 576084 234326
rect 576032 234262 576084 234268
rect 576044 225162 576072 234262
rect 575952 225134 576072 225162
rect 575952 220998 575980 225134
rect 576136 225026 576164 241198
rect 576228 236842 576256 262890
rect 576306 258632 576362 258641
rect 576306 258567 576362 258576
rect 576320 241738 576348 258567
rect 576308 241732 576360 241738
rect 576308 241674 576360 241680
rect 576216 236836 576268 236842
rect 576216 236778 576268 236784
rect 576216 236700 576268 236706
rect 576216 236642 576268 236648
rect 576044 224998 576164 225026
rect 575940 220992 575992 220998
rect 575940 220934 575992 220940
rect 575940 217660 575992 217666
rect 575676 217620 575940 217648
rect 575940 217602 575992 217608
rect 576044 217530 576072 224998
rect 576124 224936 576176 224942
rect 576124 224878 576176 224884
rect 576032 217524 576084 217530
rect 576032 217466 576084 217472
rect 576136 217410 576164 224878
rect 576228 217530 576256 236642
rect 576398 236600 576454 236609
rect 576398 236535 576454 236544
rect 576308 235068 576360 235074
rect 576308 235010 576360 235016
rect 576216 217524 576268 217530
rect 576216 217466 576268 217472
rect 576320 217410 576348 235010
rect 576412 234326 576440 236535
rect 576400 234320 576452 234326
rect 576400 234262 576452 234268
rect 576400 217524 576452 217530
rect 576400 217466 576452 217472
rect 576044 217382 576164 217410
rect 576228 217382 576348 217410
rect 575940 216028 575992 216034
rect 575940 215970 575992 215976
rect 575952 215642 575980 215970
rect 575492 215614 575980 215642
rect 575492 215506 575520 215614
rect 575308 215478 575520 215506
rect 575940 215552 575992 215558
rect 575940 215494 575992 215500
rect 575308 203946 575336 215478
rect 575952 212242 575980 215494
rect 575768 212214 575980 212242
rect 575308 203918 575612 203946
rect 575032 202286 575336 202314
rect 575308 195378 575336 202286
rect 574848 195350 575336 195378
rect 574848 176474 574876 195350
rect 575584 186402 575612 203918
rect 575768 202960 575796 212214
rect 576044 203114 576072 217382
rect 576124 212628 576176 212634
rect 576124 212570 576176 212576
rect 576136 212498 576164 212570
rect 576124 212492 576176 212498
rect 576124 212434 576176 212440
rect 576032 203108 576084 203114
rect 576032 203050 576084 203056
rect 575768 202932 576072 202960
rect 575940 202768 575992 202774
rect 575940 202710 575992 202716
rect 575952 199306 575980 202710
rect 575940 199300 575992 199306
rect 575940 199242 575992 199248
rect 576044 192778 576072 202932
rect 576228 202774 576256 217382
rect 576412 217274 576440 217466
rect 576320 217246 576440 217274
rect 576216 202768 576268 202774
rect 576216 202710 576268 202716
rect 576216 201544 576268 201550
rect 576216 201486 576268 201492
rect 576124 197396 576176 197402
rect 576124 197338 576176 197344
rect 576032 192772 576084 192778
rect 576032 192714 576084 192720
rect 576136 192658 576164 197338
rect 576044 192630 576164 192658
rect 576044 192250 576072 192630
rect 576124 192568 576176 192574
rect 576124 192510 576176 192516
rect 575860 192222 576072 192250
rect 575860 186946 575888 192222
rect 576032 191140 576084 191146
rect 576032 191082 576084 191088
rect 575860 186930 575980 186946
rect 575860 186924 575992 186930
rect 575860 186918 575940 186924
rect 575940 186866 575992 186872
rect 575308 186374 575612 186402
rect 575308 177426 575336 186374
rect 576044 186266 576072 191082
rect 575676 186238 576072 186266
rect 575308 177398 575520 177426
rect 575492 177018 575520 177398
rect 575676 177290 575704 186238
rect 576136 186130 576164 192510
rect 576228 191826 576256 201486
rect 576320 198898 576348 217246
rect 576308 198892 576360 198898
rect 576308 198834 576360 198840
rect 576308 198756 576360 198762
rect 576308 198698 576360 198704
rect 576216 191820 576268 191826
rect 576216 191762 576268 191768
rect 576216 186312 576268 186318
rect 576216 186254 576268 186260
rect 576044 186102 576164 186130
rect 575940 184952 575992 184958
rect 575860 184900 575940 184906
rect 575860 184894 575992 184900
rect 575860 184878 575980 184894
rect 575860 183410 575888 184878
rect 575860 183394 575980 183410
rect 575860 183388 575992 183394
rect 575860 183382 575940 183388
rect 575940 183330 575992 183336
rect 576044 182986 576072 186102
rect 576032 182980 576084 182986
rect 576032 182922 576084 182928
rect 575676 177274 575980 177290
rect 575676 177268 575992 177274
rect 575676 177262 575940 177268
rect 575940 177210 575992 177216
rect 575492 176990 576072 177018
rect 574848 176446 575796 176474
rect 575768 175692 575796 176446
rect 575940 175704 575992 175710
rect 575768 175664 575940 175692
rect 575940 175646 575992 175652
rect 576044 175386 576072 176990
rect 575492 175358 576072 175386
rect 575492 165322 575520 175358
rect 575940 174820 575992 174826
rect 575940 174762 575992 174768
rect 575952 174706 575980 174762
rect 575860 174678 575980 174706
rect 575860 170354 575888 174678
rect 575940 174004 575992 174010
rect 575940 173946 575992 173952
rect 575952 170746 575980 173946
rect 576124 172576 576176 172582
rect 576124 172518 576176 172524
rect 575940 170740 575992 170746
rect 575940 170682 575992 170688
rect 575860 170326 575980 170354
rect 575952 170270 575980 170326
rect 575940 170264 575992 170270
rect 575940 170206 575992 170212
rect 576136 170134 576164 172518
rect 575940 170128 575992 170134
rect 575940 170070 575992 170076
rect 576124 170128 576176 170134
rect 576124 170070 576176 170076
rect 575952 169810 575980 170070
rect 575676 169782 575980 169810
rect 575676 166002 575704 169782
rect 575676 165974 576164 166002
rect 575492 165294 576072 165322
rect 575940 164960 575992 164966
rect 575768 164920 575940 164948
rect 575768 163554 575796 164920
rect 575940 164902 575992 164908
rect 575400 163526 575796 163554
rect 575400 145296 575428 163526
rect 575940 160812 575992 160818
rect 575940 160754 575992 160760
rect 575952 153474 575980 160754
rect 575940 153468 575992 153474
rect 575940 153410 575992 153416
rect 575940 153264 575992 153270
rect 575860 153212 575940 153218
rect 575860 153206 575992 153212
rect 575860 153190 575980 153206
rect 575860 146146 575888 153190
rect 575940 150476 575992 150482
rect 575940 150418 575992 150424
rect 575952 149394 575980 150418
rect 576044 149734 576072 165294
rect 576136 158030 576164 165974
rect 576124 158024 576176 158030
rect 576124 157966 576176 157972
rect 576124 157888 576176 157894
rect 576124 157830 576176 157836
rect 576032 149728 576084 149734
rect 576032 149670 576084 149676
rect 575940 149388 575992 149394
rect 575940 149330 575992 149336
rect 575860 146118 575980 146146
rect 575952 145994 575980 146118
rect 575940 145988 575992 145994
rect 575940 145930 575992 145936
rect 575940 145308 575992 145314
rect 575400 145268 575940 145296
rect 575940 145250 575992 145256
rect 574756 144906 575980 144922
rect 574756 144900 575992 144906
rect 574756 144894 575940 144900
rect 574756 135946 574784 144894
rect 575940 144842 575992 144848
rect 576032 144560 576084 144566
rect 575860 144508 576032 144514
rect 575860 144502 576084 144508
rect 575860 144486 576072 144502
rect 575860 140434 575888 144486
rect 575940 144424 575992 144430
rect 575940 144366 575992 144372
rect 575952 140962 575980 144366
rect 575940 140956 575992 140962
rect 575940 140898 575992 140904
rect 575860 140406 576072 140434
rect 575940 140344 575992 140350
rect 575584 140304 575940 140332
rect 575400 136190 575520 136218
rect 575400 135946 575428 136190
rect 574756 135918 575428 135946
rect 575492 129010 575520 136190
rect 575216 128982 575520 129010
rect 575216 127956 575244 128982
rect 575584 128874 575612 140304
rect 575940 140286 575992 140292
rect 575940 139936 575992 139942
rect 575940 139878 575992 139884
rect 575952 137306 575980 139878
rect 575400 128846 575612 128874
rect 575676 137278 575980 137306
rect 575400 128092 575428 128846
rect 575400 128064 575612 128092
rect 575216 127928 575520 127956
rect 575492 125474 575520 127928
rect 575400 125446 575520 125474
rect 575400 124148 575428 125446
rect 575584 124930 575612 128064
rect 575676 127786 575704 137278
rect 575940 137216 575992 137222
rect 575768 137164 575940 137170
rect 575768 137158 575992 137164
rect 575768 137142 575980 137158
rect 575768 128194 575796 137142
rect 576044 137086 576072 140406
rect 576136 139942 576164 157830
rect 576124 139936 576176 139942
rect 576124 139878 576176 139884
rect 576032 137080 576084 137086
rect 576032 137022 576084 137028
rect 575940 137012 575992 137018
rect 575940 136954 575992 136960
rect 575952 136898 575980 136954
rect 575860 136870 575980 136898
rect 575860 131968 575888 136870
rect 576228 136762 576256 186254
rect 576320 184958 576348 198698
rect 576308 184952 576360 184958
rect 576308 184894 576360 184900
rect 576308 183388 576360 183394
rect 576308 183330 576360 183336
rect 576320 144566 576348 183330
rect 576308 144560 576360 144566
rect 576308 144502 576360 144508
rect 576136 136734 576256 136762
rect 575940 132592 575992 132598
rect 575940 132534 575992 132540
rect 575952 132122 575980 132534
rect 575940 132116 575992 132122
rect 575940 132058 575992 132064
rect 575860 131940 575980 131968
rect 575952 130558 575980 131940
rect 575940 130552 575992 130558
rect 575940 130494 575992 130500
rect 576136 128330 576164 136734
rect 576136 128302 576256 128330
rect 575768 128166 576164 128194
rect 575676 127758 575980 127786
rect 575952 127702 575980 127758
rect 575940 127696 575992 127702
rect 575940 127638 575992 127644
rect 575584 124902 576072 124930
rect 575400 124120 575980 124148
rect 575952 122602 575980 124120
rect 575940 122596 575992 122602
rect 575940 122538 575992 122544
rect 575940 121644 575992 121650
rect 574940 121604 575940 121632
rect 574940 114050 574968 121604
rect 575940 121586 575992 121592
rect 575940 117768 575992 117774
rect 575860 117716 575940 117722
rect 575860 117710 575992 117716
rect 575860 117694 575980 117710
rect 575860 115954 575888 117694
rect 575768 115926 575888 115954
rect 576044 115938 576072 124902
rect 576136 121650 576164 128166
rect 576124 121644 576176 121650
rect 576124 121586 576176 121592
rect 576124 118584 576176 118590
rect 576124 118526 576176 118532
rect 576032 115932 576084 115938
rect 575768 114186 575796 115926
rect 576032 115874 576084 115880
rect 575768 114158 576072 114186
rect 574940 114034 575980 114050
rect 574940 114028 575992 114034
rect 574940 114022 575940 114028
rect 575940 113970 575992 113976
rect 576044 111058 576072 114158
rect 575124 111030 576072 111058
rect 575124 101402 575152 111030
rect 575940 110968 575992 110974
rect 575940 110910 575992 110916
rect 575952 106298 575980 110910
rect 576136 108866 576164 118526
rect 576228 109052 576256 128302
rect 576308 120760 576360 120766
rect 576308 120702 576360 120708
rect 576320 109120 576348 120702
rect 576320 109092 576440 109120
rect 576228 109024 576348 109052
rect 576124 108860 576176 108866
rect 576124 108802 576176 108808
rect 575032 101374 575152 101402
rect 575400 106270 575980 106298
rect 575032 92018 575060 101374
rect 575400 96642 575428 106270
rect 575940 104440 575992 104446
rect 575676 104388 575940 104394
rect 575676 104382 575992 104388
rect 575676 104366 575980 104382
rect 575400 96614 575612 96642
rect 575032 91990 575336 92018
rect 575308 84266 575336 91990
rect 575584 89026 575612 96614
rect 575676 92290 575704 104366
rect 575940 104304 575992 104310
rect 575768 104252 575940 104258
rect 575768 104246 575992 104252
rect 575768 104230 575980 104246
rect 575768 93378 575796 104230
rect 575940 104168 575992 104174
rect 575860 104116 575940 104122
rect 575860 104110 575992 104116
rect 575860 104094 575980 104110
rect 575860 93514 575888 104094
rect 575940 102468 575992 102474
rect 575940 102410 575992 102416
rect 575952 100502 575980 102410
rect 575940 100496 575992 100502
rect 575940 100438 575992 100444
rect 575940 100360 575992 100366
rect 575940 100302 575992 100308
rect 575952 93838 575980 100302
rect 575940 93832 575992 93838
rect 575940 93774 575992 93780
rect 575860 93486 576164 93514
rect 575768 93350 576072 93378
rect 575676 92262 575980 92290
rect 575952 90642 575980 92262
rect 575940 90636 575992 90642
rect 575940 90578 575992 90584
rect 576044 90522 576072 93350
rect 575768 90494 576072 90522
rect 575584 88998 575704 89026
rect 575216 84238 575336 84266
rect 575216 62098 575244 84238
rect 575676 81410 575704 88998
rect 575584 81382 575704 81410
rect 575584 79370 575612 81382
rect 575768 79506 575796 90494
rect 576136 88618 576164 93486
rect 575860 88590 576164 88618
rect 575860 81376 575888 88590
rect 576320 85678 576348 109024
rect 576412 104174 576440 109092
rect 576400 104168 576452 104174
rect 576400 104110 576452 104116
rect 576308 85672 576360 85678
rect 576308 85614 576360 85620
rect 576308 85536 576360 85542
rect 576228 85484 576308 85490
rect 576228 85478 576360 85484
rect 576228 85462 576348 85478
rect 575940 81388 575992 81394
rect 575860 81348 575940 81376
rect 575940 81330 575992 81336
rect 576124 81388 576176 81394
rect 576124 81330 576176 81336
rect 575768 79490 575980 79506
rect 575768 79484 575992 79490
rect 575768 79478 575940 79484
rect 575940 79426 575992 79432
rect 575584 79342 575796 79370
rect 575216 62070 575336 62098
rect 575308 52442 575336 62070
rect 575768 58562 575796 79342
rect 576032 74792 576084 74798
rect 576032 74734 576084 74740
rect 575940 72208 575992 72214
rect 575860 72156 575940 72162
rect 575860 72150 575992 72156
rect 575860 72134 575980 72150
rect 575860 58800 575888 72134
rect 575940 70372 575992 70378
rect 575940 70314 575992 70320
rect 575952 63374 575980 70314
rect 576044 67590 576072 74734
rect 576032 67584 576084 67590
rect 576032 67526 576084 67532
rect 575940 63368 575992 63374
rect 575940 63310 575992 63316
rect 576136 61606 576164 81330
rect 576228 79506 576256 85462
rect 576228 79478 576348 79506
rect 576124 61600 576176 61606
rect 576124 61542 576176 61548
rect 575940 58812 575992 58818
rect 575860 58772 575940 58800
rect 575940 58754 575992 58760
rect 575768 58534 575888 58562
rect 575860 53258 575888 58534
rect 576320 58002 576348 79478
rect 576400 61600 576452 61606
rect 576400 61542 576452 61548
rect 576216 57996 576268 58002
rect 576216 57938 576268 57944
rect 576308 57996 576360 58002
rect 576308 57938 576360 57944
rect 576124 57860 576176 57866
rect 576124 57802 576176 57808
rect 575860 53230 576072 53258
rect 575584 52958 575980 52986
rect 575584 52442 575612 52958
rect 575952 52834 575980 52958
rect 575940 52828 575992 52834
rect 575940 52770 575992 52776
rect 576044 52714 576072 53230
rect 575308 52414 575612 52442
rect 575768 52686 576072 52714
rect 575768 52306 575796 52686
rect 575940 52624 575992 52630
rect 575940 52566 575992 52572
rect 575584 52278 575796 52306
rect 575584 52034 575612 52278
rect 575492 52006 575612 52034
rect 575492 46594 575520 52006
rect 575952 51490 575980 52566
rect 576136 51814 576164 57802
rect 576124 51808 576176 51814
rect 576124 51750 576176 51756
rect 575952 51462 576072 51490
rect 575492 46566 575980 46594
rect 575492 46430 575888 46458
rect 575952 46442 575980 46566
rect 575492 43738 575520 46430
rect 575860 46322 575888 46430
rect 575940 46436 575992 46442
rect 575940 46378 575992 46384
rect 576044 46322 576072 51462
rect 575860 46294 576072 46322
rect 576032 46232 576084 46238
rect 576032 46174 576084 46180
rect 575492 43710 575980 43738
rect 575952 43654 575980 43710
rect 575940 43648 575992 43654
rect 575940 43590 575992 43596
rect 575940 43512 575992 43518
rect 575768 43472 575940 43500
rect 575768 41562 575796 43472
rect 575940 43454 575992 43460
rect 575492 41534 575796 41562
rect 575492 37210 575520 41534
rect 576044 41426 576072 46174
rect 575676 41398 576072 41426
rect 575676 39522 575704 41398
rect 575676 39494 576072 39522
rect 575940 39432 575992 39438
rect 575940 39374 575992 39380
rect 575952 37262 575980 39374
rect 575940 37256 575992 37262
rect 575492 37182 575796 37210
rect 575940 37198 575992 37204
rect 575768 36938 575796 37182
rect 575768 36910 575980 36938
rect 575952 35358 575980 36910
rect 575940 35352 575992 35358
rect 575940 35294 575992 35300
rect 575940 35216 575992 35222
rect 575940 35158 575992 35164
rect 575952 35034 575980 35158
rect 575768 35006 575980 35034
rect 575768 21570 575796 35006
rect 575940 33856 575992 33862
rect 575400 21542 575796 21570
rect 575860 33816 575940 33844
rect 575400 21434 575428 21542
rect 575308 21406 575428 21434
rect 575308 16538 575336 21406
rect 575860 21026 575888 33816
rect 575940 33798 575992 33804
rect 576044 33402 576072 39494
rect 576124 33856 576176 33862
rect 576124 33798 576176 33804
rect 575952 33374 576072 33402
rect 575952 33114 575980 33374
rect 575940 33108 575992 33114
rect 575940 33050 575992 33056
rect 576032 28688 576084 28694
rect 576032 28630 576084 28636
rect 575940 28348 575992 28354
rect 575940 28290 575992 28296
rect 575952 21298 575980 28290
rect 576044 21418 576072 28630
rect 576136 21554 576164 33798
rect 576228 24206 576256 57938
rect 576308 57316 576360 57322
rect 576308 57258 576360 57264
rect 576320 28694 576348 57258
rect 576412 33862 576440 61542
rect 576400 33856 576452 33862
rect 576400 33798 576452 33804
rect 576308 28688 576360 28694
rect 576308 28630 576360 28636
rect 576216 24200 576268 24206
rect 576216 24142 576268 24148
rect 576124 21548 576176 21554
rect 576124 21490 576176 21496
rect 576032 21412 576084 21418
rect 576032 21354 576084 21360
rect 576308 21412 576360 21418
rect 576308 21354 576360 21360
rect 575952 21270 576072 21298
rect 575860 20998 575980 21026
rect 575952 20602 575980 20998
rect 575940 20596 575992 20602
rect 575940 20538 575992 20544
rect 576044 20482 576072 21270
rect 576124 20596 576176 20602
rect 576124 20538 576176 20544
rect 575032 16510 575336 16538
rect 575400 20454 576072 20482
rect 17224 7744 17276 7750
rect 14186 7712 14242 7721
rect 17224 7686 17276 7692
rect 58808 7744 58860 7750
rect 58808 7686 58860 7692
rect 113546 7712 113602 7721
rect 14186 7647 14242 7656
rect 12084 5506 12112 7004
rect 12072 5500 12124 5506
rect 12072 5442 12124 5448
rect 14200 5370 14228 7647
rect 15198 7440 15254 7449
rect 15198 7375 15254 7384
rect 14188 5364 14240 5370
rect 14188 5306 14240 5312
rect 15212 5302 15240 7375
rect 15200 5296 15252 5302
rect 15200 5238 15252 5244
rect 12440 4208 12492 4214
rect 12440 4150 12492 4156
rect 10048 4072 10100 4078
rect 10048 4014 10100 4020
rect 9772 3052 9824 3058
rect 9772 2994 9824 3000
rect 10060 480 10088 4014
rect 11242 3360 11298 3369
rect 11242 3295 11298 3304
rect 11256 480 11284 3295
rect 12452 480 12480 4150
rect 14832 3868 14884 3874
rect 14832 3810 14884 3816
rect 13636 3460 13688 3466
rect 13636 3402 13688 3408
rect 13648 480 13676 3402
rect 14844 480 14872 3810
rect 16028 3800 16080 3806
rect 16028 3742 16080 3748
rect 16040 480 16068 3742
rect 17236 480 17264 7686
rect 21916 6180 21968 6186
rect 21916 6122 21968 6128
rect 19524 5228 19576 5234
rect 19524 5170 19576 5176
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 18340 480 18368 3470
rect 19536 480 19564 5170
rect 20718 3632 20774 3641
rect 20718 3567 20774 3576
rect 20732 480 20760 3567
rect 21928 480 21956 6122
rect 22204 4758 22232 7004
rect 30288 6248 30340 6254
rect 30288 6190 30340 6196
rect 26700 5024 26752 5030
rect 25502 4992 25558 5001
rect 26700 4966 26752 4972
rect 25502 4927 25558 4936
rect 22192 4752 22244 4758
rect 22192 4694 22244 4700
rect 24308 3528 24360 3534
rect 23110 3496 23166 3505
rect 24308 3470 24360 3476
rect 23110 3431 23166 3440
rect 23124 480 23152 3431
rect 24320 480 24348 3470
rect 25516 480 25544 4927
rect 26712 480 26740 4966
rect 27896 3732 27948 3738
rect 27896 3674 27948 3680
rect 27908 480 27936 3674
rect 29092 2848 29144 2854
rect 29092 2790 29144 2796
rect 29104 480 29132 2790
rect 30300 480 30328 6190
rect 32416 5438 32444 7004
rect 32404 5432 32456 5438
rect 31482 5400 31538 5409
rect 32404 5374 32456 5380
rect 31482 5335 31538 5344
rect 31496 480 31524 5335
rect 42154 5264 42210 5273
rect 42154 5199 42210 5208
rect 33876 4956 33928 4962
rect 33876 4898 33928 4904
rect 32680 2916 32732 2922
rect 32680 2858 32732 2864
rect 32692 480 32720 2858
rect 33888 480 33916 4898
rect 40960 4820 41012 4826
rect 40960 4762 41012 4768
rect 36176 4208 36228 4214
rect 36176 4150 36228 4156
rect 34978 3768 35034 3777
rect 34978 3703 35034 3712
rect 34992 480 35020 3703
rect 36188 480 36216 4150
rect 37372 3800 37424 3806
rect 37372 3742 37424 3748
rect 37384 480 37412 3742
rect 38568 2984 38620 2990
rect 38568 2926 38620 2932
rect 39764 2984 39816 2990
rect 39764 2926 39816 2932
rect 38580 480 38608 2926
rect 39776 480 39804 2926
rect 40972 480 41000 4762
rect 42168 480 42196 5199
rect 42536 5166 42564 7004
rect 52748 6866 52776 7004
rect 52736 6860 52788 6866
rect 52736 6802 52788 6808
rect 42524 5160 42576 5166
rect 42524 5102 42576 5108
rect 51632 5160 51684 5166
rect 51632 5102 51684 5108
rect 43352 4276 43404 4282
rect 43352 4218 43404 4224
rect 43364 480 43392 4218
rect 44548 3732 44600 3738
rect 44548 3674 44600 3680
rect 44560 480 44588 3674
rect 45744 3188 45796 3194
rect 45744 3130 45796 3136
rect 46940 3188 46992 3194
rect 46940 3130 46992 3136
rect 45756 480 45784 3130
rect 46952 480 46980 3130
rect 49332 3120 49384 3126
rect 49332 3062 49384 3068
rect 50528 3120 50580 3126
rect 50528 3062 50580 3068
rect 48136 3052 48188 3058
rect 48136 2994 48188 3000
rect 48148 480 48176 2994
rect 49344 480 49372 3062
rect 50540 480 50568 3062
rect 51644 480 51672 5102
rect 55220 5092 55272 5098
rect 55220 5034 55272 5040
rect 52828 4820 52880 4826
rect 52828 4762 52880 4768
rect 52840 480 52868 4762
rect 54024 4344 54076 4350
rect 54024 4286 54076 4292
rect 54036 480 54064 4286
rect 55232 480 55260 5034
rect 57612 4412 57664 4418
rect 57612 4354 57664 4360
rect 56416 3256 56468 3262
rect 56416 3198 56468 3204
rect 56428 480 56456 3198
rect 57624 480 57652 4354
rect 58820 480 58848 7686
rect 113546 7647 113602 7656
rect 84934 7576 84990 7585
rect 69480 7540 69532 7546
rect 84934 7511 84990 7520
rect 109958 7576 110014 7585
rect 109958 7511 110014 7520
rect 69480 7482 69532 7488
rect 62960 6798 62988 7004
rect 62948 6792 63000 6798
rect 62948 6734 63000 6740
rect 65984 6384 66036 6390
rect 65984 6326 66036 6332
rect 63592 6316 63644 6322
rect 63592 6258 63644 6264
rect 62396 5024 62448 5030
rect 62396 4966 62448 4972
rect 60004 3324 60056 3330
rect 60004 3266 60056 3272
rect 60016 480 60044 3266
rect 61200 3188 61252 3194
rect 61200 3130 61252 3136
rect 61212 480 61240 3130
rect 62408 480 62436 4966
rect 63604 480 63632 6258
rect 64788 4480 64840 4486
rect 64788 4422 64840 4428
rect 64800 480 64828 4422
rect 65996 480 66024 6326
rect 67180 4888 67232 4894
rect 67180 4830 67232 4836
rect 67192 480 67220 4830
rect 68284 4548 68336 4554
rect 68284 4490 68336 4496
rect 68296 480 68324 4490
rect 69492 480 69520 7482
rect 73080 6730 73108 7004
rect 73068 6724 73120 6730
rect 73068 6666 73120 6672
rect 83292 6662 83320 7004
rect 83280 6656 83332 6662
rect 83280 6598 83332 6604
rect 83832 6520 83884 6526
rect 83832 6462 83884 6468
rect 77852 6452 77904 6458
rect 77852 6394 77904 6400
rect 73068 6384 73120 6390
rect 73068 6326 73120 6332
rect 70676 3392 70728 3398
rect 70676 3334 70728 3340
rect 70688 480 70716 3334
rect 71872 3256 71924 3262
rect 71872 3198 71924 3204
rect 71884 480 71912 3198
rect 73080 480 73108 6326
rect 75460 4616 75512 4622
rect 75460 4558 75512 4564
rect 74264 3664 74316 3670
rect 74264 3606 74316 3612
rect 74276 480 74304 3606
rect 75472 480 75500 4558
rect 76656 3664 76708 3670
rect 76656 3606 76708 3612
rect 76668 480 76696 3606
rect 77864 480 77892 6394
rect 80244 4956 80296 4962
rect 80244 4898 80296 4904
rect 79048 3324 79100 3330
rect 79048 3266 79100 3272
rect 79060 480 79088 3266
rect 80256 480 80284 4898
rect 82636 4684 82688 4690
rect 82636 4626 82688 4632
rect 81440 3596 81492 3602
rect 81440 3538 81492 3544
rect 81452 480 81480 3538
rect 82648 480 82676 4626
rect 83844 480 83872 6462
rect 84948 480 84976 7511
rect 90916 6588 90968 6594
rect 90916 6530 90968 6536
rect 89720 4752 89772 4758
rect 89720 4694 89772 4700
rect 88524 4140 88576 4146
rect 88524 4082 88576 4088
rect 87328 3596 87380 3602
rect 87328 3538 87380 3544
rect 86132 3392 86184 3398
rect 86132 3334 86184 3340
rect 86144 480 86172 3334
rect 87340 480 87368 3538
rect 88536 480 88564 4082
rect 89732 480 89760 4694
rect 90928 480 90956 6530
rect 93308 4140 93360 4146
rect 93308 4082 93360 4088
rect 92112 4004 92164 4010
rect 92112 3946 92164 3952
rect 92124 480 92152 3946
rect 93320 480 93348 4082
rect 93504 4078 93532 7004
rect 94504 6112 94556 6118
rect 94504 6054 94556 6060
rect 93492 4072 93544 4078
rect 93492 4014 93544 4020
rect 94516 480 94544 6054
rect 101588 6044 101640 6050
rect 101588 5986 101640 5992
rect 96896 5500 96948 5506
rect 96896 5442 96948 5448
rect 95700 3936 95752 3942
rect 95700 3878 95752 3884
rect 95712 480 95740 3878
rect 96908 480 96936 5442
rect 99380 5364 99432 5370
rect 99380 5306 99432 5312
rect 98092 4888 98144 4894
rect 98092 4830 98144 4836
rect 98104 480 98132 4830
rect 99392 3942 99420 5306
rect 100484 4072 100536 4078
rect 100484 4014 100536 4020
rect 99380 3936 99432 3942
rect 99286 3904 99342 3913
rect 99380 3878 99432 3884
rect 99286 3839 99342 3848
rect 99300 480 99328 3839
rect 100496 480 100524 4014
rect 101600 480 101628 5986
rect 102782 3904 102838 3913
rect 103624 3874 103652 7004
rect 106372 5976 106424 5982
rect 106372 5918 106424 5924
rect 103980 5432 104032 5438
rect 103980 5374 104032 5380
rect 102782 3839 102838 3848
rect 103612 3868 103664 3874
rect 102796 480 102824 3839
rect 103612 3810 103664 3816
rect 103992 480 104020 5374
rect 104256 5296 104308 5302
rect 104256 5238 104308 5244
rect 104268 3874 104296 5238
rect 104256 3868 104308 3874
rect 104256 3810 104308 3816
rect 105176 3868 105228 3874
rect 105176 3810 105228 3816
rect 105188 480 105216 3810
rect 106384 480 106412 5918
rect 108764 5772 108816 5778
rect 108764 5714 108816 5720
rect 107568 4004 107620 4010
rect 107568 3946 107620 3952
rect 107580 480 107608 3946
rect 108776 480 108804 5714
rect 109972 480 110000 7511
rect 111156 5364 111208 5370
rect 111156 5306 111208 5312
rect 111168 480 111196 5306
rect 112352 3936 112404 3942
rect 112352 3878 112404 3884
rect 112364 480 112392 3878
rect 113560 480 113588 7647
rect 575032 7478 575060 16510
rect 575400 15314 575428 20454
rect 575940 20324 575992 20330
rect 575940 20266 575992 20272
rect 575952 17270 575980 20266
rect 576032 19372 576084 19378
rect 576032 19314 576084 19320
rect 575940 17264 575992 17270
rect 575940 17206 575992 17212
rect 575940 16720 575992 16726
rect 575124 15286 575428 15314
rect 575492 16668 575940 16674
rect 575492 16662 575992 16668
rect 575492 16646 575980 16662
rect 575124 7546 575152 15286
rect 575492 15178 575520 16646
rect 575400 15150 575520 15178
rect 575400 14906 575428 15150
rect 575400 14878 575520 14906
rect 575492 11778 575520 14878
rect 575492 11750 575612 11778
rect 575112 7540 575164 7546
rect 575112 7482 575164 7488
rect 575020 7472 575072 7478
rect 575020 7414 575072 7420
rect 575480 7472 575532 7478
rect 575480 7414 575532 7420
rect 113836 5234 113864 7004
rect 115940 5908 115992 5914
rect 115940 5850 115992 5856
rect 119436 5908 119488 5914
rect 119436 5850 119488 5856
rect 113824 5228 113876 5234
rect 113824 5170 113876 5176
rect 114744 3936 114796 3942
rect 114744 3878 114796 3884
rect 114756 480 114784 3878
rect 115952 480 115980 5850
rect 118240 5296 118292 5302
rect 118240 5238 118292 5244
rect 117134 3224 117190 3233
rect 117134 3159 117190 3168
rect 117148 480 117176 3159
rect 118252 480 118280 5238
rect 119448 480 119476 5850
rect 123024 5840 123076 5846
rect 123024 5782 123076 5788
rect 120630 4040 120686 4049
rect 120630 3975 120686 3984
rect 120644 480 120672 3975
rect 121828 3868 121880 3874
rect 121828 3810 121880 3816
rect 121840 480 121868 3810
rect 123036 480 123064 5782
rect 124048 3534 124076 7004
rect 125416 5228 125468 5234
rect 125416 5170 125468 5176
rect 124036 3528 124088 3534
rect 124036 3470 124088 3476
rect 124220 3528 124272 3534
rect 124220 3470 124272 3476
rect 124232 480 124260 3470
rect 125428 480 125456 5170
rect 134168 2854 134196 7004
rect 144380 2922 144408 7004
rect 154592 4214 154620 7004
rect 154580 4208 154632 4214
rect 154580 4150 154632 4156
rect 164712 2990 164740 7004
rect 174924 4282 174952 7004
rect 174912 4276 174964 4282
rect 174912 4218 174964 4224
rect 185044 3058 185072 7004
rect 195256 3126 195284 7004
rect 205468 4350 205496 7004
rect 215588 4418 215616 7004
rect 215576 4412 215628 4418
rect 215576 4354 215628 4360
rect 205456 4344 205508 4350
rect 205456 4286 205508 4292
rect 225800 3194 225828 7004
rect 236012 4486 236040 7004
rect 246132 4554 246160 7004
rect 246120 4548 246172 4554
rect 246120 4490 246172 4496
rect 236000 4480 236052 4486
rect 236000 4422 236052 4428
rect 256344 3262 256372 7004
rect 266556 4622 266584 7004
rect 266544 4616 266596 4622
rect 266544 4558 266596 4564
rect 276676 3330 276704 7004
rect 286888 4690 286916 7004
rect 286876 4684 286928 4690
rect 286876 4626 286928 4632
rect 297100 3398 297128 7004
rect 307220 4758 307248 7004
rect 307208 4752 307260 4758
rect 307208 4694 307260 4700
rect 317432 4146 317460 7004
rect 327552 5506 327580 7004
rect 327540 5500 327592 5506
rect 327540 5442 327592 5448
rect 317420 4140 317472 4146
rect 317420 4082 317472 4088
rect 337764 4078 337792 7004
rect 347976 5438 348004 7004
rect 347964 5432 348016 5438
rect 347964 5374 348016 5380
rect 337752 4072 337804 4078
rect 337752 4014 337804 4020
rect 358096 4010 358124 7004
rect 368308 5370 368336 7004
rect 368296 5364 368348 5370
rect 368296 5306 368348 5312
rect 358084 4004 358136 4010
rect 358084 3946 358136 3952
rect 378520 3942 378548 7004
rect 388640 5302 388668 7004
rect 388628 5296 388680 5302
rect 388628 5238 388680 5244
rect 378508 3936 378560 3942
rect 378508 3878 378560 3884
rect 398852 3874 398880 7004
rect 409064 5234 409092 7004
rect 409052 5228 409104 5234
rect 409052 5170 409104 5176
rect 398840 3868 398892 3874
rect 398840 3810 398892 3816
rect 419184 3806 419212 7004
rect 419172 3800 419224 3806
rect 419172 3742 419224 3748
rect 429396 3738 429424 7004
rect 439608 5166 439636 7004
rect 439596 5160 439648 5166
rect 439596 5102 439648 5108
rect 449728 5098 449756 7004
rect 449716 5092 449768 5098
rect 449716 5034 449768 5040
rect 459940 5030 459968 7004
rect 459928 5024 459980 5030
rect 459928 4966 459980 4972
rect 429384 3732 429436 3738
rect 429384 3674 429436 3680
rect 470060 3670 470088 7004
rect 480272 4962 480300 7004
rect 480260 4956 480312 4962
rect 480260 4898 480312 4904
rect 470048 3664 470100 3670
rect 470048 3606 470100 3612
rect 490484 3602 490512 7004
rect 500604 4894 500632 7004
rect 510816 5137 510844 7004
rect 510802 5128 510858 5137
rect 510802 5063 510858 5072
rect 500592 4888 500644 4894
rect 500592 4830 500644 4836
rect 490472 3596 490524 3602
rect 490472 3538 490524 3544
rect 521028 3466 521056 7004
rect 531148 5409 531176 7004
rect 531134 5400 531190 5409
rect 531134 5335 531190 5344
rect 541360 5273 541388 7004
rect 541346 5264 541402 5273
rect 541346 5199 541402 5208
rect 551572 4826 551600 7004
rect 561692 5001 561720 7004
rect 561678 4992 561734 5001
rect 561678 4927 561734 4936
rect 571904 4865 571932 7004
rect 571890 4856 571946 4865
rect 551560 4820 551612 4826
rect 571890 4791 571946 4800
rect 551560 4762 551612 4768
rect 575492 3641 575520 7414
rect 575584 3777 575612 11750
rect 576044 11642 576072 19314
rect 575768 11614 576072 11642
rect 575768 7614 575796 11614
rect 576136 7818 576164 20538
rect 576320 20346 576348 21354
rect 576228 20318 576348 20346
rect 576124 7812 576176 7818
rect 576124 7754 576176 7760
rect 576228 7750 576256 20318
rect 576308 17264 576360 17270
rect 576308 17206 576360 17212
rect 576216 7744 576268 7750
rect 576216 7686 576268 7692
rect 576320 7682 576348 17206
rect 576308 7676 576360 7682
rect 576308 7618 576360 7624
rect 575756 7608 575808 7614
rect 575756 7550 575808 7556
rect 575940 7540 575992 7546
rect 575940 7482 575992 7488
rect 575570 3768 575626 3777
rect 575570 3703 575626 3712
rect 575478 3632 575534 3641
rect 575478 3567 575534 3576
rect 521016 3460 521068 3466
rect 521016 3402 521068 3408
rect 297088 3392 297140 3398
rect 575952 3369 575980 7482
rect 576872 6050 576900 455903
rect 576950 434072 577006 434081
rect 576950 434007 577006 434016
rect 576964 6118 576992 434007
rect 577042 412584 577098 412593
rect 577042 412519 577098 412528
rect 577056 6594 577084 412519
rect 577134 390756 577190 390765
rect 577134 390691 577190 390700
rect 577044 6588 577096 6594
rect 577044 6530 577096 6536
rect 577148 6526 577176 390691
rect 577226 368860 577282 368869
rect 577226 368795 577282 368804
rect 577136 6520 577188 6526
rect 577136 6462 577188 6468
rect 577240 6390 577268 368795
rect 577228 6384 577280 6390
rect 577228 6326 577280 6332
rect 576952 6112 577004 6118
rect 576952 6054 577004 6060
rect 576860 6044 576912 6050
rect 576860 5986 576912 5992
rect 578252 3534 578280 632023
rect 578330 610056 578386 610065
rect 578330 609991 578386 610000
rect 578344 4049 578372 609991
rect 578422 588024 578478 588033
rect 578422 587959 578478 587968
rect 578436 5982 578464 587959
rect 578514 565856 578570 565865
rect 578514 565791 578570 565800
rect 578528 6458 578556 565791
rect 578606 543960 578662 543969
rect 578606 543895 578662 543904
rect 578516 6452 578568 6458
rect 578516 6394 578568 6400
rect 578620 6322 578648 543895
rect 578698 500032 578754 500041
rect 578698 499967 578754 499976
rect 578608 6316 578660 6322
rect 578608 6258 578660 6264
rect 578424 5976 578476 5982
rect 578424 5918 578476 5924
rect 578330 4040 578386 4049
rect 578330 3975 578386 3984
rect 578240 3528 578292 3534
rect 578712 3505 578740 499967
rect 579620 487144 579672 487150
rect 579620 487086 579672 487092
rect 579632 486849 579660 487086
rect 579618 486840 579674 486849
rect 579618 486775 579674 486784
rect 578790 478000 578846 478009
rect 578790 477935 578846 477944
rect 578804 5914 578832 477935
rect 578882 302696 578938 302705
rect 578882 302631 578938 302640
rect 578896 6254 578924 302631
rect 578974 280528 579030 280537
rect 578974 280463 579030 280472
rect 578884 6248 578936 6254
rect 578884 6190 578936 6196
rect 578988 6186 579016 280463
rect 580170 252240 580226 252249
rect 580170 252175 580226 252184
rect 579068 216368 579120 216374
rect 579068 216310 579120 216316
rect 579080 215937 579108 216310
rect 579066 215928 579122 215937
rect 579066 215863 579122 215872
rect 579068 194064 579120 194070
rect 579066 194032 579068 194041
rect 579120 194032 579122 194041
rect 579066 193967 579122 193976
rect 579068 172168 579120 172174
rect 579066 172136 579068 172145
rect 579120 172136 579122 172145
rect 579066 172071 579122 172080
rect 579068 150136 579120 150142
rect 579066 150104 579068 150113
rect 579120 150104 579122 150113
rect 579066 150039 579122 150048
rect 580184 127974 580212 252175
rect 579068 127968 579120 127974
rect 579066 127936 579068 127945
rect 580172 127968 580224 127974
rect 579120 127936 579122 127945
rect 580172 127910 580224 127916
rect 579066 127871 579122 127880
rect 579068 106208 579120 106214
rect 579066 106176 579068 106185
rect 579120 106176 579122 106185
rect 579066 106111 579122 106120
rect 579068 84176 579120 84182
rect 579066 84144 579068 84153
rect 579120 84144 579122 84153
rect 579066 84079 579122 84088
rect 579068 62008 579120 62014
rect 579066 61976 579068 61985
rect 579120 61976 579122 61985
rect 579066 61911 579122 61920
rect 579068 39976 579120 39982
rect 579066 39944 579068 39953
rect 579120 39944 579122 39953
rect 579066 39879 579122 39888
rect 580276 6662 580304 674591
rect 580354 627736 580410 627745
rect 580354 627671 580410 627680
rect 580368 6730 580396 627671
rect 580446 580816 580502 580825
rect 580446 580751 580502 580760
rect 580460 6798 580488 580751
rect 580538 533896 580594 533905
rect 580538 533831 580594 533840
rect 580552 6866 580580 533831
rect 580630 439920 580686 439929
rect 580630 439855 580686 439864
rect 580644 216374 580672 439855
rect 580722 393000 580778 393009
rect 580722 392935 580778 392944
rect 580632 216368 580684 216374
rect 580632 216310 580684 216316
rect 580630 205320 580686 205329
rect 580630 205255 580686 205264
rect 580644 106214 580672 205255
rect 580736 194070 580764 392935
rect 580814 346080 580870 346089
rect 580814 346015 580870 346024
rect 580724 194064 580776 194070
rect 580724 194006 580776 194012
rect 580828 172174 580856 346015
rect 580906 299160 580962 299169
rect 580906 299095 580962 299104
rect 580816 172168 580868 172174
rect 580816 172110 580868 172116
rect 580722 158400 580778 158409
rect 580722 158335 580778 158344
rect 580632 106208 580684 106214
rect 580632 106150 580684 106156
rect 580736 84182 580764 158335
rect 580920 150142 580948 299095
rect 580908 150136 580960 150142
rect 580908 150078 580960 150084
rect 580814 111480 580870 111489
rect 580814 111415 580870 111424
rect 580724 84176 580776 84182
rect 580724 84118 580776 84124
rect 580630 64560 580686 64569
rect 580630 64495 580686 64504
rect 580644 39982 580672 64495
rect 580828 62014 580856 111415
rect 580816 62008 580868 62014
rect 580816 61950 580868 61956
rect 580632 39976 580684 39982
rect 580632 39918 580684 39924
rect 580540 6860 580592 6866
rect 580540 6802 580592 6808
rect 580448 6792 580500 6798
rect 580448 6734 580500 6740
rect 580356 6724 580408 6730
rect 580356 6666 580408 6672
rect 580264 6656 580316 6662
rect 580264 6598 580316 6604
rect 578976 6180 579028 6186
rect 578976 6122 579028 6128
rect 578792 5908 578844 5914
rect 578792 5850 578844 5856
rect 578240 3470 578292 3476
rect 578698 3496 578754 3505
rect 578698 3431 578754 3440
rect 297088 3334 297140 3340
rect 575938 3360 575994 3369
rect 276664 3324 276716 3330
rect 575938 3295 575994 3304
rect 276664 3266 276716 3272
rect 256332 3256 256384 3262
rect 256332 3198 256384 3204
rect 225788 3188 225840 3194
rect 225788 3130 225840 3136
rect 195244 3120 195296 3126
rect 195244 3062 195296 3068
rect 185032 3052 185084 3058
rect 185032 2994 185084 3000
rect 164700 2984 164752 2990
rect 164700 2926 164752 2932
rect 144368 2916 144420 2922
rect 144368 2858 144420 2864
rect 134156 2848 134208 2854
rect 134156 2790 134208 2796
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3330 682216 3386 682272
rect 5446 675280 5502 675336
rect 5354 653384 5410 653440
rect 3146 624824 3202 624880
rect 4066 567316 4122 567352
rect 4066 567296 4068 567316
rect 4068 567296 4120 567316
rect 4120 567296 4122 567316
rect 5262 543904 5318 543960
rect 5170 521736 5226 521792
rect 3422 509904 3478 509960
rect 3330 208120 3386 208176
rect 3238 122032 3294 122088
rect 5078 499840 5134 499896
rect 4986 455912 5042 455968
rect 3514 452376 3570 452432
rect 4894 434016 4950 434072
rect 3606 394984 3662 395040
rect 4802 390632 4858 390688
rect 3698 337456 3754 337512
rect 3790 294344 3846 294400
rect 3974 251232 4030 251288
rect 3882 215328 3938 215384
rect 3790 84088 3846 84144
rect 3698 62056 3754 62112
rect 3606 39888 3662 39944
rect 4066 193296 4122 193352
rect 3974 105984 4030 106040
rect 4710 171148 4766 171184
rect 4710 171128 4712 171148
rect 4712 171128 4764 171148
rect 4764 171128 4766 171148
rect 4710 165008 4766 165064
rect 4710 150048 4766 150104
rect 4158 128152 4214 128208
rect 4066 78920 4122 78976
rect 3882 35808 3938 35864
rect 3514 18536 3570 18592
rect 5262 4800 5318 4856
rect 6918 631488 6974 631544
rect 6734 610068 6790 610124
rect 6642 588172 6698 588228
rect 6550 566276 6606 566332
rect 6458 543632 6514 543688
rect 6458 524320 6514 524376
rect 6458 505008 6514 505064
rect 6458 485696 6514 485752
rect 6458 466384 6514 466440
rect 6458 447072 6514 447128
rect 6458 408448 6514 408504
rect 6458 324400 6514 324456
rect 6366 302640 6422 302696
rect 6734 543632 6790 543688
rect 6734 524320 6790 524376
rect 6734 505008 6790 505064
rect 6734 485696 6790 485752
rect 6918 477944 6974 478000
rect 6734 466384 6790 466440
rect 6734 447072 6790 447128
rect 6734 408448 6790 408504
rect 7010 412528 7066 412584
rect 7102 368464 7158 368520
rect 7194 346432 7250 346488
rect 7286 280472 7342 280528
rect 7378 258576 7434 258632
rect 7470 236544 7526 236600
rect 8850 5072 8906 5128
rect 6826 3848 6882 3904
rect 346766 688744 346822 688800
rect 544106 688880 544162 688936
rect 522210 688744 522266 688800
rect 478326 688608 478382 688664
rect 500222 688608 500278 688664
rect 324594 686432 324650 686488
rect 565910 686296 565966 686352
rect 576306 675280 576362 675336
rect 580262 674600 580318 674656
rect 576306 653384 576362 653440
rect 578238 632032 578294 632088
rect 576306 521736 576362 521792
rect 576858 455912 576914 455968
rect 576306 346296 576362 346352
rect 576306 324400 576362 324456
rect 576306 258576 576362 258632
rect 576398 236544 576454 236600
rect 14186 7656 14242 7712
rect 15198 7384 15254 7440
rect 11242 3304 11298 3360
rect 20718 3576 20774 3632
rect 25502 4936 25558 4992
rect 23110 3440 23166 3496
rect 31482 5344 31538 5400
rect 42154 5208 42210 5264
rect 34978 3712 35034 3768
rect 113546 7656 113602 7712
rect 84934 7520 84990 7576
rect 109958 7520 110014 7576
rect 99286 3848 99342 3904
rect 102782 3848 102838 3904
rect 117134 3168 117190 3224
rect 120630 3984 120686 4040
rect 510802 5072 510858 5128
rect 531134 5344 531190 5400
rect 541346 5208 541402 5264
rect 561678 4936 561734 4992
rect 571890 4800 571946 4856
rect 575570 3712 575626 3768
rect 575478 3576 575534 3632
rect 576950 434016 577006 434072
rect 577042 412528 577098 412584
rect 577134 390700 577190 390756
rect 577226 368804 577282 368860
rect 578330 610000 578386 610056
rect 578422 587968 578478 588024
rect 578514 565800 578570 565856
rect 578606 543904 578662 543960
rect 578698 499976 578754 500032
rect 578330 3984 578386 4040
rect 579618 486784 579674 486840
rect 578790 477944 578846 478000
rect 578882 302640 578938 302696
rect 578974 280472 579030 280528
rect 580170 252184 580226 252240
rect 579066 215872 579122 215928
rect 579066 194012 579068 194032
rect 579068 194012 579120 194032
rect 579120 194012 579122 194032
rect 579066 193976 579122 194012
rect 579066 172116 579068 172136
rect 579068 172116 579120 172136
rect 579120 172116 579122 172136
rect 579066 172080 579122 172116
rect 579066 150084 579068 150104
rect 579068 150084 579120 150104
rect 579120 150084 579122 150104
rect 579066 150048 579122 150084
rect 579066 127916 579068 127936
rect 579068 127916 579120 127936
rect 579120 127916 579122 127936
rect 579066 127880 579122 127916
rect 579066 106156 579068 106176
rect 579068 106156 579120 106176
rect 579120 106156 579122 106176
rect 579066 106120 579122 106156
rect 579066 84124 579068 84144
rect 579068 84124 579120 84144
rect 579120 84124 579122 84144
rect 579066 84088 579122 84124
rect 579066 61956 579068 61976
rect 579068 61956 579120 61976
rect 579120 61956 579122 61976
rect 579066 61920 579122 61956
rect 579066 39924 579068 39944
rect 579068 39924 579120 39944
rect 579120 39924 579122 39944
rect 579066 39888 579122 39924
rect 580354 627680 580410 627736
rect 580446 580760 580502 580816
rect 580538 533840 580594 533896
rect 580630 439864 580686 439920
rect 580722 392944 580778 393000
rect 580630 205264 580686 205320
rect 580814 346024 580870 346080
rect 580906 299104 580962 299160
rect 580722 158344 580778 158400
rect 580814 111424 580870 111480
rect 580630 64504 580686 64560
rect 578698 3440 578754 3496
rect 575938 3304 575994 3360
<< metal3 >>
rect 583520 697900 584960 698140
rect -960 696540 480 696780
rect 544101 688938 544167 688941
rect 564750 688938 564756 688940
rect 544101 688936 564756 688938
rect 544101 688880 544106 688936
rect 544162 688880 564756 688936
rect 544101 688878 564756 688880
rect 544101 688875 544167 688878
rect 564750 688876 564756 688878
rect 564820 688876 564826 688940
rect 340822 688740 340828 688804
rect 340892 688802 340898 688804
rect 346761 688802 346827 688805
rect 340892 688800 346827 688802
rect 340892 688744 346766 688800
rect 346822 688744 346827 688800
rect 340892 688742 346827 688744
rect 340892 688740 340898 688742
rect 346761 688739 346827 688742
rect 522205 688802 522271 688805
rect 566038 688802 566044 688804
rect 522205 688800 566044 688802
rect 522205 688744 522210 688800
rect 522266 688744 566044 688800
rect 522205 688742 566044 688744
rect 522205 688739 522271 688742
rect 566038 688740 566044 688742
rect 566108 688740 566114 688804
rect 10910 688604 10916 688668
rect 10980 688666 10986 688668
rect 478321 688666 478387 688669
rect 10980 688664 478387 688666
rect 10980 688608 478326 688664
rect 478382 688608 478387 688664
rect 10980 688606 478387 688608
rect 10980 688604 10986 688606
rect 478321 688603 478387 688606
rect 500217 688666 500283 688669
rect 564566 688666 564572 688668
rect 500217 688664 564572 688666
rect 500217 688608 500222 688664
rect 500278 688608 564572 688664
rect 500217 688606 564572 688608
rect 500217 688603 500283 688606
rect 564566 688604 564572 688606
rect 564636 688604 564642 688668
rect 166390 687108 166396 687172
rect 166460 687170 166466 687172
rect 177614 687170 177620 687172
rect 166460 687110 177620 687170
rect 166460 687108 166466 687110
rect 177614 687108 177620 687110
rect 177684 687108 177690 687172
rect 202822 687108 202828 687172
rect 202892 687170 202898 687172
rect 212390 687170 212396 687172
rect 202892 687110 212396 687170
rect 202892 687108 202898 687110
rect 212390 687108 212396 687110
rect 212460 687108 212466 687172
rect 230422 687108 230428 687172
rect 230492 687170 230498 687172
rect 235206 687170 235212 687172
rect 230492 687110 235212 687170
rect 230492 687108 230498 687110
rect 235206 687108 235212 687110
rect 235276 687108 235282 687172
rect 10174 686428 10180 686492
rect 10244 686490 10250 686492
rect 12566 686490 12572 686492
rect 10244 686430 12572 686490
rect 10244 686428 10250 686430
rect 12566 686428 12572 686430
rect 12636 686428 12642 686492
rect 95182 686428 95188 686492
rect 95252 686490 95258 686492
rect 99966 686490 99972 686492
rect 95252 686430 99972 686490
rect 95252 686428 95258 686430
rect 99966 686428 99972 686430
rect 100036 686428 100042 686492
rect 240174 686428 240180 686492
rect 240244 686490 240250 686492
rect 249558 686490 249564 686492
rect 240244 686430 249564 686490
rect 240244 686428 240250 686430
rect 249558 686428 249564 686430
rect 249628 686428 249634 686492
rect 324446 686428 324452 686492
rect 324516 686490 324522 686492
rect 324589 686490 324655 686493
rect 324516 686488 324655 686490
rect 324516 686432 324594 686488
rect 324650 686432 324655 686488
rect 324516 686430 324655 686432
rect 324516 686428 324522 686430
rect 324589 686427 324655 686430
rect 565905 686356 565971 686357
rect 93894 686292 93900 686356
rect 93964 686354 93970 686356
rect 103278 686354 103284 686356
rect 93964 686294 103284 686354
rect 93964 686292 93970 686294
rect 103278 686292 103284 686294
rect 103348 686292 103354 686356
rect 108246 686292 108252 686356
rect 108316 686354 108322 686356
rect 113030 686354 113036 686356
rect 108316 686294 113036 686354
rect 108316 686292 108322 686294
rect 113030 686292 113036 686294
rect 113100 686292 113106 686356
rect 182214 686292 182220 686356
rect 182284 686354 182290 686356
rect 186262 686354 186268 686356
rect 182284 686294 186268 686354
rect 182284 686292 182290 686294
rect 186262 686292 186268 686294
rect 186332 686292 186338 686356
rect 340638 686292 340644 686356
rect 340708 686354 340714 686356
rect 340822 686354 340828 686356
rect 340708 686294 340828 686354
rect 340708 686292 340714 686294
rect 340822 686292 340828 686294
rect 340892 686292 340898 686356
rect 565854 686354 565860 686356
rect 565814 686294 565860 686354
rect 565924 686352 565971 686356
rect 565966 686296 565971 686352
rect 565854 686292 565860 686294
rect 565924 686292 565971 686296
rect 565905 686291 565971 686292
rect 583520 686204 584960 686444
rect -960 682274 480 682364
rect 3325 682274 3391 682277
rect -960 682272 3391 682274
rect -960 682216 3330 682272
rect 3386 682216 3391 682272
rect -960 682214 3391 682216
rect -960 682124 480 682214
rect 3325 682211 3391 682214
rect 5441 675338 5507 675341
rect 7054 675338 7114 675920
rect 576350 675341 576410 675920
rect 5441 675336 7114 675338
rect 5441 675280 5446 675336
rect 5502 675280 7114 675336
rect 5441 675278 7114 675280
rect 576301 675336 576410 675341
rect 576301 675280 576306 675336
rect 576362 675280 576410 675336
rect 576301 675278 576410 675280
rect 5441 675275 5507 675278
rect 576301 675275 576367 675278
rect 580257 674658 580323 674661
rect 583520 674658 584960 674748
rect 580257 674656 584960 674658
rect 580257 674600 580262 674656
rect 580318 674600 584960 674656
rect 580257 674598 584960 674600
rect 580257 674595 580323 674598
rect 583520 674508 584960 674598
rect -960 667844 480 668084
rect 583520 662676 584960 662916
rect -960 653428 480 653668
rect 5349 653442 5415 653445
rect 7054 653442 7114 654024
rect 576350 653445 576410 654024
rect 5349 653440 7114 653442
rect 5349 653384 5354 653440
rect 5410 653384 7114 653440
rect 5349 653382 7114 653384
rect 576301 653440 576410 653445
rect 576301 653384 576306 653440
rect 576362 653384 576410 653440
rect 576301 653382 576410 653384
rect 5349 653379 5415 653382
rect 576301 653379 576367 653382
rect 583520 650980 584960 651220
rect 583520 639284 584960 639524
rect -960 639012 480 639252
rect 6913 631546 6979 631549
rect 7054 631546 7114 632128
rect 576902 632090 576962 632128
rect 578233 632090 578299 632093
rect 576902 632088 578299 632090
rect 576902 632032 578238 632088
rect 578294 632032 578299 632088
rect 576902 632030 578299 632032
rect 578233 632027 578299 632030
rect 6913 631544 7114 631546
rect 6913 631488 6918 631544
rect 6974 631488 7114 631544
rect 6913 631486 7114 631488
rect 6913 631483 6979 631486
rect 580349 627738 580415 627741
rect 583520 627738 584960 627828
rect 580349 627736 584960 627738
rect 580349 627680 580354 627736
rect 580410 627680 584960 627736
rect 580349 627678 584960 627680
rect 580349 627675 580415 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 3141 624882 3207 624885
rect -960 624880 3207 624882
rect -960 624824 3146 624880
rect 3202 624824 3207 624880
rect -960 624822 3207 624824
rect -960 624732 480 624822
rect 3141 624819 3207 624822
rect 583520 615756 584960 615996
rect -960 610316 480 610556
rect 6729 610126 6795 610129
rect 6729 610124 7084 610126
rect 6729 610068 6734 610124
rect 6790 610068 7084 610124
rect 6729 610066 7084 610068
rect 6729 610063 6795 610066
rect 576902 610058 576962 610096
rect 578325 610058 578391 610061
rect 576902 610056 578391 610058
rect 576902 610000 578330 610056
rect 578386 610000 578391 610056
rect 576902 609998 578391 610000
rect 578325 609995 578391 609998
rect 583520 604060 584960 604300
rect -960 595900 480 596140
rect 583520 592364 584960 592604
rect 6637 588230 6703 588233
rect 6637 588228 7084 588230
rect 6637 588172 6642 588228
rect 6698 588172 7084 588228
rect 6637 588170 7084 588172
rect 6637 588167 6703 588170
rect 576902 588026 576962 588200
rect 578417 588026 578483 588029
rect 576902 588024 578483 588026
rect 576902 587968 578422 588024
rect 578478 587968 578483 588024
rect 576902 587966 578483 587968
rect 578417 587963 578483 587966
rect -960 581620 480 581860
rect 580441 580818 580507 580821
rect 583520 580818 584960 580908
rect 580441 580816 584960 580818
rect 580441 580760 580446 580816
rect 580502 580760 584960 580816
rect 580441 580758 584960 580760
rect 580441 580755 580507 580758
rect 583520 580668 584960 580758
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 4061 567354 4127 567357
rect -960 567352 4127 567354
rect -960 567296 4066 567352
rect 4122 567296 4127 567352
rect -960 567294 4127 567296
rect -960 567204 480 567294
rect 4061 567291 4127 567294
rect 6545 566334 6611 566337
rect 6545 566332 7084 566334
rect 6545 566276 6550 566332
rect 6606 566276 7084 566332
rect 6545 566274 7084 566276
rect 6545 566271 6611 566274
rect 576902 565858 576962 566304
rect 578509 565858 578575 565861
rect 576902 565856 578575 565858
rect 576902 565800 578514 565856
rect 578570 565800 578575 565856
rect 576902 565798 578575 565800
rect 578509 565795 578575 565798
rect 583520 557140 584960 557380
rect -960 552924 480 553164
rect 583520 545444 584960 545684
rect 5257 543962 5323 543965
rect 7054 543962 7114 544272
rect 5257 543960 7114 543962
rect 5257 543904 5262 543960
rect 5318 543904 7114 543960
rect 5257 543902 7114 543904
rect 576902 543962 576962 544272
rect 578601 543962 578667 543965
rect 576902 543960 578667 543962
rect 576902 543904 578606 543960
rect 578662 543904 578667 543960
rect 576902 543902 578667 543904
rect 5257 543899 5323 543902
rect 578601 543899 578667 543902
rect 6453 543690 6519 543693
rect 6729 543690 6795 543693
rect 6453 543688 6795 543690
rect 6453 543632 6458 543688
rect 6514 543632 6734 543688
rect 6790 543632 6795 543688
rect 6453 543630 6795 543632
rect 6453 543627 6519 543630
rect 6729 543627 6795 543630
rect -960 538508 480 538748
rect 580533 533898 580599 533901
rect 583520 533898 584960 533988
rect 580533 533896 584960 533898
rect 580533 533840 580538 533896
rect 580594 533840 584960 533896
rect 580533 533838 584960 533840
rect 580533 533835 580599 533838
rect 583520 533748 584960 533838
rect 6453 524378 6519 524381
rect 6729 524378 6795 524381
rect 6453 524376 6795 524378
rect -960 524092 480 524332
rect 6453 524320 6458 524376
rect 6514 524320 6734 524376
rect 6790 524320 6795 524376
rect 6453 524318 6795 524320
rect 6453 524315 6519 524318
rect 6729 524315 6795 524318
rect 5165 521794 5231 521797
rect 7054 521794 7114 522376
rect 576350 521797 576410 522376
rect 583520 521916 584960 522156
rect 5165 521792 7114 521794
rect 5165 521736 5170 521792
rect 5226 521736 7114 521792
rect 5165 521734 7114 521736
rect 576301 521792 576410 521797
rect 576301 521736 576306 521792
rect 576362 521736 576410 521792
rect 576301 521734 576410 521736
rect 5165 521731 5231 521734
rect 576301 521731 576367 521734
rect 583520 510220 584960 510460
rect -960 509962 480 510052
rect 3417 509962 3483 509965
rect -960 509960 3483 509962
rect -960 509904 3422 509960
rect 3478 509904 3483 509960
rect -960 509902 3483 509904
rect -960 509812 480 509902
rect 3417 509899 3483 509902
rect 6453 505066 6519 505069
rect 6729 505066 6795 505069
rect 6453 505064 6795 505066
rect 6453 505008 6458 505064
rect 6514 505008 6734 505064
rect 6790 505008 6795 505064
rect 6453 505006 6795 505008
rect 6453 505003 6519 505006
rect 6729 505003 6795 505006
rect 5073 499898 5139 499901
rect 7054 499898 7114 500480
rect 576902 500034 576962 500480
rect 578693 500034 578759 500037
rect 576902 500032 578759 500034
rect 576902 499976 578698 500032
rect 578754 499976 578759 500032
rect 576902 499974 578759 499976
rect 578693 499971 578759 499974
rect 5073 499896 7114 499898
rect 5073 499840 5078 499896
rect 5134 499840 7114 499896
rect 5073 499838 7114 499840
rect 5073 499835 5139 499838
rect 583520 498524 584960 498764
rect -960 495396 480 495636
rect 579613 486842 579679 486845
rect 583520 486842 584960 486932
rect 579613 486840 584960 486842
rect 579613 486784 579618 486840
rect 579674 486784 584960 486840
rect 579613 486782 584960 486784
rect 579613 486779 579679 486782
rect 583520 486692 584960 486782
rect 6453 485754 6519 485757
rect 6729 485754 6795 485757
rect 6453 485752 6795 485754
rect 6453 485696 6458 485752
rect 6514 485696 6734 485752
rect 6790 485696 6795 485752
rect 6453 485694 6795 485696
rect 6453 485691 6519 485694
rect 6729 485691 6795 485694
rect -960 480980 480 481220
rect 6913 478002 6979 478005
rect 7054 478002 7114 478584
rect 6913 478000 7114 478002
rect 6913 477944 6918 478000
rect 6974 477944 7114 478000
rect 6913 477942 7114 477944
rect 576902 478002 576962 478584
rect 578785 478002 578851 478005
rect 576902 478000 578851 478002
rect 576902 477944 578790 478000
rect 578846 477944 578851 478000
rect 576902 477942 578851 477944
rect 6913 477939 6979 477942
rect 578785 477939 578851 477942
rect 583520 474996 584960 475236
rect -960 466700 480 466940
rect 6453 466442 6519 466445
rect 6729 466442 6795 466445
rect 6453 466440 6795 466442
rect 6453 466384 6458 466440
rect 6514 466384 6734 466440
rect 6790 466384 6795 466440
rect 6453 466382 6795 466384
rect 6453 466379 6519 466382
rect 6729 466379 6795 466382
rect 583520 463300 584960 463540
rect 4981 455970 5047 455973
rect 7054 455970 7114 456552
rect 576902 455973 576962 456552
rect 4981 455968 7114 455970
rect 4981 455912 4986 455968
rect 5042 455912 7114 455968
rect 4981 455910 7114 455912
rect 576853 455968 576962 455973
rect 576853 455912 576858 455968
rect 576914 455912 576962 455968
rect 576853 455910 576962 455912
rect 4981 455907 5047 455910
rect 576853 455907 576919 455910
rect -960 452434 480 452524
rect 3509 452434 3575 452437
rect -960 452432 3575 452434
rect -960 452376 3514 452432
rect 3570 452376 3575 452432
rect -960 452374 3575 452376
rect -960 452284 480 452374
rect 3509 452371 3575 452374
rect 583520 451604 584960 451844
rect 6453 447130 6519 447133
rect 6729 447130 6795 447133
rect 6453 447128 6795 447130
rect 6453 447072 6458 447128
rect 6514 447072 6734 447128
rect 6790 447072 6795 447128
rect 6453 447070 6795 447072
rect 6453 447067 6519 447070
rect 6729 447067 6795 447070
rect 580625 439922 580691 439925
rect 583520 439922 584960 440012
rect 580625 439920 584960 439922
rect 580625 439864 580630 439920
rect 580686 439864 584960 439920
rect 580625 439862 584960 439864
rect 580625 439859 580691 439862
rect 583520 439772 584960 439862
rect -960 437868 480 438108
rect 4889 434074 4955 434077
rect 7054 434074 7114 434656
rect 4889 434072 7114 434074
rect 4889 434016 4894 434072
rect 4950 434016 7114 434072
rect 4889 434014 7114 434016
rect 576902 434077 576962 434656
rect 576902 434072 577011 434077
rect 576902 434016 576950 434072
rect 577006 434016 577011 434072
rect 576902 434014 577011 434016
rect 4889 434011 4955 434014
rect 576945 434011 577011 434014
rect 583520 428076 584960 428316
rect -960 423588 480 423828
rect 583520 416380 584960 416620
rect 7054 412589 7114 412760
rect 7005 412584 7114 412589
rect 7005 412528 7010 412584
rect 7066 412528 7114 412584
rect 7005 412526 7114 412528
rect 576902 412586 576962 412760
rect 577037 412586 577103 412589
rect 576902 412584 577103 412586
rect 576902 412528 577042 412584
rect 577098 412528 577103 412584
rect 576902 412526 577103 412528
rect 7005 412523 7071 412526
rect 577037 412523 577103 412526
rect -960 409172 480 409412
rect 6453 408506 6519 408509
rect 6729 408506 6795 408509
rect 6453 408504 6795 408506
rect 6453 408448 6458 408504
rect 6514 408448 6734 408504
rect 6790 408448 6795 408504
rect 6453 408446 6795 408448
rect 6453 408443 6519 408446
rect 6729 408443 6795 408446
rect 583520 404684 584960 404924
rect -960 395042 480 395132
rect 3601 395042 3667 395045
rect -960 395040 3667 395042
rect -960 394984 3606 395040
rect 3662 394984 3667 395040
rect -960 394982 3667 394984
rect -960 394892 480 394982
rect 3601 394979 3667 394982
rect 580717 393002 580783 393005
rect 583520 393002 584960 393092
rect 580717 393000 584960 393002
rect 580717 392944 580722 393000
rect 580778 392944 584960 393000
rect 580717 392942 584960 392944
rect 580717 392939 580783 392942
rect 583520 392852 584960 392942
rect 577129 390758 577195 390761
rect 576932 390756 577195 390758
rect 4797 390690 4863 390693
rect 7054 390690 7114 390728
rect 576932 390700 577134 390756
rect 577190 390700 577195 390756
rect 576932 390698 577195 390700
rect 577129 390695 577195 390698
rect 4797 390688 7114 390690
rect 4797 390632 4802 390688
rect 4858 390632 7114 390688
rect 4797 390630 7114 390632
rect 4797 390627 4863 390630
rect 583520 381156 584960 381396
rect -960 380476 480 380716
rect 583520 369460 584960 369700
rect 577221 368862 577287 368865
rect 576932 368860 577287 368862
rect 7054 368525 7114 368832
rect 576932 368804 577226 368860
rect 577282 368804 577287 368860
rect 576932 368802 577287 368804
rect 577221 368799 577287 368802
rect 7054 368520 7163 368525
rect 7054 368464 7102 368520
rect 7158 368464 7163 368520
rect 7054 368462 7163 368464
rect 7097 368459 7163 368462
rect -960 366060 480 366300
rect 583520 357764 584960 358004
rect -960 351780 480 352020
rect 7238 346493 7298 346936
rect 7189 346488 7298 346493
rect 7189 346432 7194 346488
rect 7250 346432 7298 346488
rect 7189 346430 7298 346432
rect 7189 346427 7255 346430
rect 576350 346357 576410 346936
rect 576301 346352 576410 346357
rect 576301 346296 576306 346352
rect 576362 346296 576410 346352
rect 576301 346294 576410 346296
rect 576301 346291 576367 346294
rect 580809 346082 580875 346085
rect 583520 346082 584960 346172
rect 580809 346080 584960 346082
rect 580809 346024 580814 346080
rect 580870 346024 584960 346080
rect 580809 346022 584960 346024
rect 580809 346019 580875 346022
rect 583520 345932 584960 346022
rect -960 337514 480 337604
rect 3693 337514 3759 337517
rect -960 337512 3759 337514
rect -960 337456 3698 337512
rect 3754 337456 3759 337512
rect -960 337454 3759 337456
rect -960 337364 480 337454
rect 3693 337451 3759 337454
rect 583520 334236 584960 334476
rect 6453 324458 6519 324461
rect 7054 324458 7114 325040
rect 576350 324461 576410 325040
rect 6453 324456 7114 324458
rect 6453 324400 6458 324456
rect 6514 324400 7114 324456
rect 6453 324398 7114 324400
rect 576301 324456 576410 324461
rect 576301 324400 576306 324456
rect 576362 324400 576410 324456
rect 576301 324398 576410 324400
rect 6453 324395 6519 324398
rect 576301 324395 576367 324398
rect -960 322948 480 323188
rect 583520 322540 584960 322780
rect 583520 310708 584960 310948
rect -960 308668 480 308908
rect 6361 302698 6427 302701
rect 7054 302698 7114 303008
rect 6361 302696 7114 302698
rect 6361 302640 6366 302696
rect 6422 302640 7114 302696
rect 6361 302638 7114 302640
rect 576902 302698 576962 303008
rect 578877 302698 578943 302701
rect 576902 302696 578943 302698
rect 576902 302640 578882 302696
rect 578938 302640 578943 302696
rect 576902 302638 578943 302640
rect 6361 302635 6427 302638
rect 578877 302635 578943 302638
rect 580901 299162 580967 299165
rect 583520 299162 584960 299252
rect 580901 299160 584960 299162
rect 580901 299104 580906 299160
rect 580962 299104 584960 299160
rect 580901 299102 584960 299104
rect 580901 299099 580967 299102
rect 583520 299012 584960 299102
rect -960 294402 480 294492
rect 3785 294402 3851 294405
rect -960 294400 3851 294402
rect -960 294344 3790 294400
rect 3846 294344 3851 294400
rect -960 294342 3851 294344
rect -960 294252 480 294342
rect 3785 294339 3851 294342
rect 583520 287316 584960 287556
rect 7238 280533 7298 281112
rect 7238 280528 7347 280533
rect 7238 280472 7286 280528
rect 7342 280472 7347 280528
rect 7238 280470 7347 280472
rect 576902 280530 576962 281112
rect 578969 280530 579035 280533
rect 576902 280528 579035 280530
rect 576902 280472 578974 280528
rect 579030 280472 579035 280528
rect 576902 280470 579035 280472
rect 7281 280467 7347 280470
rect 578969 280467 579035 280470
rect -960 279972 480 280212
rect 583520 275620 584960 275860
rect -960 265556 480 265796
rect 583520 263788 584960 264028
rect 7422 258637 7482 259216
rect 576350 258637 576410 259216
rect 7373 258632 7482 258637
rect 7373 258576 7378 258632
rect 7434 258576 7482 258632
rect 7373 258574 7482 258576
rect 576301 258632 576410 258637
rect 576301 258576 576306 258632
rect 576362 258576 576410 258632
rect 576301 258574 576410 258576
rect 7373 258571 7439 258574
rect 576301 258571 576367 258574
rect 580165 252242 580231 252245
rect 583520 252242 584960 252332
rect 580165 252240 584960 252242
rect 580165 252184 580170 252240
rect 580226 252184 584960 252240
rect 580165 252182 584960 252184
rect 580165 252179 580231 252182
rect 583520 252092 584960 252182
rect -960 251290 480 251380
rect 3969 251290 4035 251293
rect -960 251288 4035 251290
rect -960 251232 3974 251288
rect 4030 251232 4035 251288
rect -960 251230 4035 251232
rect -960 251140 480 251230
rect 3969 251227 4035 251230
rect 583520 240396 584960 240636
rect -960 236860 480 237100
rect 7422 236605 7482 237184
rect 576350 236605 576410 237184
rect 7422 236600 7531 236605
rect 7422 236544 7470 236600
rect 7526 236544 7531 236600
rect 7422 236542 7531 236544
rect 576350 236600 576459 236605
rect 576350 236544 576398 236600
rect 576454 236544 576459 236600
rect 576350 236542 576459 236544
rect 7465 236539 7531 236542
rect 576393 236539 576459 236542
rect 583520 228700 584960 228940
rect -960 222444 480 222684
rect 583520 216868 584960 217108
rect 579061 215930 579127 215933
rect 576902 215928 579127 215930
rect 576902 215872 579066 215928
rect 579122 215872 579127 215928
rect 576902 215870 579127 215872
rect 3877 215386 3943 215389
rect 3877 215384 7114 215386
rect 3877 215328 3882 215384
rect 3938 215328 7114 215384
rect 3877 215326 7114 215328
rect 3877 215323 3943 215326
rect 7054 215288 7114 215326
rect 576902 215288 576962 215870
rect 579061 215867 579127 215870
rect -960 208178 480 208268
rect 3325 208178 3391 208181
rect -960 208176 3391 208178
rect -960 208120 3330 208176
rect 3386 208120 3391 208176
rect -960 208118 3391 208120
rect -960 208028 480 208118
rect 3325 208115 3391 208118
rect 580625 205322 580691 205325
rect 583520 205322 584960 205412
rect 580625 205320 584960 205322
rect 580625 205264 580630 205320
rect 580686 205264 584960 205320
rect 580625 205262 584960 205264
rect 580625 205259 580691 205262
rect 583520 205172 584960 205262
rect 579061 194034 579127 194037
rect 576902 194032 579127 194034
rect -960 193748 480 193988
rect 576902 193976 579066 194032
rect 579122 193976 579127 194032
rect 576902 193974 579127 193976
rect 576902 193392 576962 193974
rect 579061 193971 579127 193974
rect 583520 193476 584960 193716
rect 4061 193354 4127 193357
rect 7054 193354 7114 193392
rect 4061 193352 7114 193354
rect 4061 193296 4066 193352
rect 4122 193296 7114 193352
rect 4061 193294 7114 193296
rect 4061 193291 4127 193294
rect 583520 181780 584960 182020
rect -960 179332 480 179572
rect 579061 172138 579127 172141
rect 576902 172136 579127 172138
rect 576902 172080 579066 172136
rect 579122 172080 579127 172136
rect 576902 172078 579127 172080
rect 576902 171496 576962 172078
rect 579061 172075 579127 172078
rect 4705 171186 4771 171189
rect 7054 171186 7114 171496
rect 4705 171184 7114 171186
rect 4705 171128 4710 171184
rect 4766 171128 7114 171184
rect 4705 171126 7114 171128
rect 4705 171123 4771 171126
rect 583520 169948 584960 170188
rect -960 165066 480 165156
rect 4705 165066 4771 165069
rect -960 165064 4771 165066
rect -960 165008 4710 165064
rect 4766 165008 4771 165064
rect -960 165006 4771 165008
rect -960 164916 480 165006
rect 4705 165003 4771 165006
rect 580717 158402 580783 158405
rect 583520 158402 584960 158492
rect 580717 158400 584960 158402
rect 580717 158344 580722 158400
rect 580778 158344 584960 158400
rect 580717 158342 584960 158344
rect 580717 158339 580783 158342
rect 583520 158252 584960 158342
rect -960 150636 480 150876
rect 4705 150106 4771 150109
rect 579061 150106 579127 150109
rect 4705 150104 7114 150106
rect 4705 150048 4710 150104
rect 4766 150048 7114 150104
rect 4705 150046 7114 150048
rect 4705 150043 4771 150046
rect 7054 149464 7114 150046
rect 576902 150104 579127 150106
rect 576902 150048 579066 150104
rect 579122 150048 579127 150104
rect 576902 150046 579127 150048
rect 576902 149464 576962 150046
rect 579061 150043 579127 150046
rect 583520 146556 584960 146796
rect -960 136220 480 136460
rect 583520 134724 584960 134964
rect 4153 128210 4219 128213
rect 4153 128208 7114 128210
rect 4153 128152 4158 128208
rect 4214 128152 7114 128208
rect 4153 128150 7114 128152
rect 4153 128147 4219 128150
rect 7054 127568 7114 128150
rect 579061 127938 579127 127941
rect 576902 127936 579127 127938
rect 576902 127880 579066 127936
rect 579122 127880 579127 127936
rect 576902 127878 579127 127880
rect 576902 127568 576962 127878
rect 579061 127875 579127 127878
rect 583520 123028 584960 123268
rect -960 122090 480 122180
rect 3233 122090 3299 122093
rect -960 122088 3299 122090
rect -960 122032 3238 122088
rect 3294 122032 3299 122088
rect -960 122030 3299 122032
rect -960 121940 480 122030
rect 3233 122027 3299 122030
rect 580809 111482 580875 111485
rect 583520 111482 584960 111572
rect 580809 111480 584960 111482
rect 580809 111424 580814 111480
rect 580870 111424 584960 111480
rect 580809 111422 584960 111424
rect 580809 111419 580875 111422
rect 583520 111332 584960 111422
rect -960 107524 480 107764
rect 579061 106178 579127 106181
rect 576902 106176 579127 106178
rect 576902 106120 579066 106176
rect 579122 106120 579127 106176
rect 576902 106118 579127 106120
rect 3969 106042 4035 106045
rect 3969 106040 7114 106042
rect 3969 105984 3974 106040
rect 4030 105984 7114 106040
rect 3969 105982 7114 105984
rect 3969 105979 4035 105982
rect 7054 105672 7114 105982
rect 576902 105672 576962 106118
rect 579061 106115 579127 106118
rect 583520 99636 584960 99876
rect -960 93108 480 93348
rect 583520 87804 584960 88044
rect 3785 84146 3851 84149
rect 579061 84146 579127 84149
rect 3785 84144 7114 84146
rect 3785 84088 3790 84144
rect 3846 84088 7114 84144
rect 3785 84086 7114 84088
rect 3785 84083 3851 84086
rect 7054 83640 7114 84086
rect 576902 84144 579127 84146
rect 576902 84088 579066 84144
rect 579122 84088 579127 84144
rect 576902 84086 579127 84088
rect 576902 83640 576962 84086
rect 579061 84083 579127 84086
rect -960 78978 480 79068
rect 4061 78978 4127 78981
rect -960 78976 4127 78978
rect -960 78920 4066 78976
rect 4122 78920 4127 78976
rect -960 78918 4127 78920
rect -960 78828 480 78918
rect 4061 78915 4127 78918
rect 583520 76108 584960 76348
rect -960 64412 480 64652
rect 580625 64562 580691 64565
rect 583520 64562 584960 64652
rect 580625 64560 584960 64562
rect 580625 64504 580630 64560
rect 580686 64504 584960 64560
rect 580625 64502 584960 64504
rect 580625 64499 580691 64502
rect 583520 64412 584960 64502
rect 3693 62114 3759 62117
rect 3693 62112 7114 62114
rect 3693 62056 3698 62112
rect 3754 62056 7114 62112
rect 3693 62054 7114 62056
rect 3693 62051 3759 62054
rect 7054 61744 7114 62054
rect 579061 61978 579127 61981
rect 576902 61976 579127 61978
rect 576902 61920 579066 61976
rect 579122 61920 579127 61976
rect 576902 61918 579127 61920
rect 576902 61744 576962 61918
rect 579061 61915 579127 61918
rect 583520 52716 584960 52956
rect -960 49996 480 50236
rect 583520 40884 584960 41124
rect 3601 39946 3667 39949
rect 579061 39946 579127 39949
rect 3601 39944 7114 39946
rect 3601 39888 3606 39944
rect 3662 39888 7114 39944
rect 3601 39886 7114 39888
rect 3601 39883 3667 39886
rect 7054 39848 7114 39886
rect 576902 39944 579127 39946
rect 576902 39888 579066 39944
rect 579122 39888 579127 39944
rect 576902 39886 579127 39888
rect 576902 39848 576962 39886
rect 579061 39883 579127 39886
rect -960 35866 480 35956
rect 3877 35866 3943 35869
rect -960 35864 3943 35866
rect -960 35808 3882 35864
rect 3938 35808 3943 35864
rect -960 35806 3943 35808
rect -960 35716 480 35806
rect 3877 35803 3943 35806
rect 583520 29188 584960 29428
rect -960 21300 480 21540
rect 3509 18594 3575 18597
rect 3509 18592 7114 18594
rect 3509 18536 3514 18592
rect 3570 18536 7114 18592
rect 3509 18534 7114 18536
rect 3509 18531 3575 18534
rect 7054 17952 7114 18534
rect 576902 17990 579538 18050
rect 576902 17952 576962 17990
rect 579478 17778 579538 17990
rect 579478 17718 579722 17778
rect 579662 17642 579722 17718
rect 583520 17642 584960 17732
rect 579662 17582 584960 17642
rect 583520 17492 584960 17582
rect 10542 7652 10548 7716
rect 10612 7714 10618 7716
rect 14181 7714 14247 7717
rect 10612 7712 14247 7714
rect 10612 7656 14186 7712
rect 14242 7656 14247 7712
rect 10612 7654 14247 7656
rect 10612 7652 10618 7654
rect 14181 7651 14247 7654
rect 113541 7714 113607 7717
rect 564750 7714 564756 7716
rect 113541 7712 564756 7714
rect 113541 7656 113546 7712
rect 113602 7656 564756 7712
rect 113541 7654 564756 7656
rect 113541 7651 113607 7654
rect 564750 7652 564756 7654
rect 564820 7652 564826 7716
rect 10910 7516 10916 7580
rect 10980 7578 10986 7580
rect 84929 7578 84995 7581
rect 10980 7576 84995 7578
rect 10980 7520 84934 7576
rect 84990 7520 84995 7576
rect 10980 7518 84995 7520
rect 10980 7516 10986 7518
rect 84929 7515 84995 7518
rect 109953 7578 110019 7581
rect 566038 7578 566044 7580
rect 109953 7576 566044 7578
rect 109953 7520 109958 7576
rect 110014 7520 566044 7576
rect 109953 7518 566044 7520
rect 109953 7515 110019 7518
rect 566038 7516 566044 7518
rect 566108 7516 566114 7580
rect 10174 7380 10180 7444
rect 10244 7442 10250 7444
rect 15193 7442 15259 7445
rect 10244 7440 15259 7442
rect 10244 7384 15198 7440
rect 15254 7384 15259 7440
rect 10244 7382 15259 7384
rect 10244 7380 10250 7382
rect 15193 7379 15259 7382
rect -960 7020 480 7260
rect 583520 5796 584960 6036
rect 31477 5402 31543 5405
rect 531129 5402 531195 5405
rect 31477 5400 531195 5402
rect 31477 5344 31482 5400
rect 31538 5344 531134 5400
rect 531190 5344 531195 5400
rect 31477 5342 531195 5344
rect 31477 5339 31543 5342
rect 531129 5339 531195 5342
rect 42149 5266 42215 5269
rect 541341 5266 541407 5269
rect 42149 5264 541407 5266
rect 42149 5208 42154 5264
rect 42210 5208 541346 5264
rect 541402 5208 541407 5264
rect 42149 5206 541407 5208
rect 42149 5203 42215 5206
rect 541341 5203 541407 5206
rect 8845 5130 8911 5133
rect 510797 5130 510863 5133
rect 8845 5128 510863 5130
rect 8845 5072 8850 5128
rect 8906 5072 510802 5128
rect 510858 5072 510863 5128
rect 8845 5070 510863 5072
rect 8845 5067 8911 5070
rect 510797 5067 510863 5070
rect 25497 4994 25563 4997
rect 561673 4994 561739 4997
rect 25497 4992 561739 4994
rect 25497 4936 25502 4992
rect 25558 4936 561678 4992
rect 561734 4936 561739 4992
rect 25497 4934 561739 4936
rect 25497 4931 25563 4934
rect 561673 4931 561739 4934
rect 5257 4858 5323 4861
rect 571885 4858 571951 4861
rect 5257 4856 571951 4858
rect 5257 4800 5262 4856
rect 5318 4800 571890 4856
rect 571946 4800 571951 4856
rect 5257 4798 571951 4800
rect 5257 4795 5323 4798
rect 571885 4795 571951 4798
rect 120625 4042 120691 4045
rect 578325 4042 578391 4045
rect 120625 4040 578391 4042
rect 120625 3984 120630 4040
rect 120686 3984 578330 4040
rect 578386 3984 578391 4040
rect 120625 3982 578391 3984
rect 120625 3979 120691 3982
rect 578325 3979 578391 3982
rect 6821 3906 6887 3909
rect 99281 3906 99347 3909
rect 6821 3904 99347 3906
rect 6821 3848 6826 3904
rect 6882 3848 99286 3904
rect 99342 3848 99347 3904
rect 6821 3846 99347 3848
rect 6821 3843 6887 3846
rect 99281 3843 99347 3846
rect 102777 3906 102843 3909
rect 564566 3906 564572 3908
rect 102777 3904 564572 3906
rect 102777 3848 102782 3904
rect 102838 3848 564572 3904
rect 102777 3846 564572 3848
rect 102777 3843 102843 3846
rect 564566 3844 564572 3846
rect 564636 3844 564642 3908
rect 34973 3770 35039 3773
rect 575565 3770 575631 3773
rect 34973 3768 575631 3770
rect 34973 3712 34978 3768
rect 35034 3712 575570 3768
rect 575626 3712 575631 3768
rect 34973 3710 575631 3712
rect 34973 3707 35039 3710
rect 575565 3707 575631 3710
rect 20713 3634 20779 3637
rect 575473 3634 575539 3637
rect 20713 3632 575539 3634
rect 20713 3576 20718 3632
rect 20774 3576 575478 3632
rect 575534 3576 575539 3632
rect 20713 3574 575539 3576
rect 20713 3571 20779 3574
rect 575473 3571 575539 3574
rect 23105 3498 23171 3501
rect 578693 3498 578759 3501
rect 23105 3496 578759 3498
rect 23105 3440 23110 3496
rect 23166 3440 578698 3496
rect 578754 3440 578759 3496
rect 23105 3438 578759 3440
rect 23105 3435 23171 3438
rect 578693 3435 578759 3438
rect 11237 3362 11303 3365
rect 575933 3362 575999 3365
rect 11237 3360 575999 3362
rect 11237 3304 11242 3360
rect 11298 3304 575938 3360
rect 575994 3304 575999 3360
rect 11237 3302 575999 3304
rect 11237 3299 11303 3302
rect 575933 3299 575999 3302
rect 117129 3226 117195 3229
rect 565854 3226 565860 3228
rect 117129 3224 565860 3226
rect 117129 3168 117134 3224
rect 117190 3168 565860 3224
rect 117129 3166 565860 3168
rect 117129 3163 117195 3166
rect 565854 3164 565860 3166
rect 565924 3164 565930 3228
<< via3 >>
rect 564756 688876 564820 688940
rect 340828 688740 340892 688804
rect 566044 688740 566108 688804
rect 10916 688604 10980 688668
rect 564572 688604 564636 688668
rect 166396 687108 166460 687172
rect 177620 687108 177684 687172
rect 202828 687108 202892 687172
rect 212396 687108 212460 687172
rect 230428 687108 230492 687172
rect 235212 687108 235276 687172
rect 10180 686428 10244 686492
rect 12572 686428 12636 686492
rect 95188 686428 95252 686492
rect 99972 686428 100036 686492
rect 240180 686428 240244 686492
rect 249564 686428 249628 686492
rect 324452 686428 324516 686492
rect 93900 686292 93964 686356
rect 103284 686292 103348 686356
rect 108252 686292 108316 686356
rect 113036 686292 113100 686356
rect 182220 686292 182284 686356
rect 186268 686292 186332 686356
rect 340644 686292 340708 686356
rect 340828 686292 340892 686356
rect 565860 686352 565924 686356
rect 565860 686296 565910 686352
rect 565910 686296 565924 686352
rect 565860 686292 565924 686296
rect 10548 7652 10612 7716
rect 564756 7652 564820 7716
rect 10916 7516 10980 7580
rect 566044 7516 566108 7580
rect 10180 7380 10244 7444
rect 564572 3844 564636 3908
rect 565860 3164 565924 3228
<< metal4 >>
rect -8436 711278 -7836 711300
rect -8436 711042 -8254 711278
rect -8018 711042 -7836 711278
rect -8436 710958 -7836 711042
rect -8436 710722 -8254 710958
rect -8018 710722 -7836 710958
rect -8436 -6786 -7836 710722
rect 591760 711278 592360 711300
rect 591760 711042 591942 711278
rect 592178 711042 592360 711278
rect 591760 710958 592360 711042
rect 591760 710722 591942 710958
rect 592178 710722 592360 710958
rect -7516 710358 -6916 710380
rect -7516 710122 -7334 710358
rect -7098 710122 -6916 710358
rect -7516 710038 -6916 710122
rect -7516 709802 -7334 710038
rect -7098 709802 -6916 710038
rect -7516 -5866 -6916 709802
rect 590840 710358 591440 710380
rect 590840 710122 591022 710358
rect 591258 710122 591440 710358
rect 590840 710038 591440 710122
rect 590840 709802 591022 710038
rect 591258 709802 591440 710038
rect -6596 709438 -5996 709460
rect -6596 709202 -6414 709438
rect -6178 709202 -5996 709438
rect -6596 709118 -5996 709202
rect -6596 708882 -6414 709118
rect -6178 708882 -5996 709118
rect -6596 -4946 -5996 708882
rect 589920 709438 590520 709460
rect 589920 709202 590102 709438
rect 590338 709202 590520 709438
rect 589920 709118 590520 709202
rect 589920 708882 590102 709118
rect 590338 708882 590520 709118
rect -5676 708518 -5076 708540
rect -5676 708282 -5494 708518
rect -5258 708282 -5076 708518
rect -5676 708198 -5076 708282
rect -5676 707962 -5494 708198
rect -5258 707962 -5076 708198
rect -5676 -4026 -5076 707962
rect 589000 708518 589600 708540
rect 589000 708282 589182 708518
rect 589418 708282 589600 708518
rect 589000 708198 589600 708282
rect 589000 707962 589182 708198
rect 589418 707962 589600 708198
rect -4756 707598 -4156 707620
rect -4756 707362 -4574 707598
rect -4338 707362 -4156 707598
rect -4756 707278 -4156 707362
rect -4756 707042 -4574 707278
rect -4338 707042 -4156 707278
rect -4756 -3106 -4156 707042
rect 588080 707598 588680 707620
rect 588080 707362 588262 707598
rect 588498 707362 588680 707598
rect 588080 707278 588680 707362
rect 588080 707042 588262 707278
rect 588498 707042 588680 707278
rect -3836 706678 -3236 706700
rect -3836 706442 -3654 706678
rect -3418 706442 -3236 706678
rect -3836 706358 -3236 706442
rect -3836 706122 -3654 706358
rect -3418 706122 -3236 706358
rect -3836 -2186 -3236 706122
rect 587160 706678 587760 706700
rect 587160 706442 587342 706678
rect 587578 706442 587760 706678
rect 587160 706358 587760 706442
rect 587160 706122 587342 706358
rect 587578 706122 587760 706358
rect -2916 705758 -2316 705780
rect -2916 705522 -2734 705758
rect -2498 705522 -2316 705758
rect -2916 705438 -2316 705522
rect -2916 705202 -2734 705438
rect -2498 705202 -2316 705438
rect -2916 -1266 -2316 705202
rect 586240 705758 586840 705780
rect 586240 705522 586422 705758
rect 586658 705522 586840 705758
rect 586240 705438 586840 705522
rect 586240 705202 586422 705438
rect 586658 705202 586840 705438
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 -346 -1396 704282
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 564755 688940 564821 688941
rect 564755 688876 564756 688940
rect 564820 688876 564821 688940
rect 564755 688875 564821 688876
rect 340827 688804 340893 688805
rect 340827 688740 340828 688804
rect 340892 688740 340893 688804
rect 340827 688739 340893 688740
rect 10915 688668 10981 688669
rect 10915 688604 10916 688668
rect 10980 688604 10981 688668
rect 10915 688603 10981 688604
rect 10179 686492 10245 686493
rect 10179 686428 10180 686492
rect 10244 686428 10245 686492
rect 10179 686427 10245 686428
rect 10182 7445 10242 686427
rect 10550 7717 10610 684302
rect 10547 7716 10613 7717
rect 10547 7652 10548 7716
rect 10612 7652 10613 7716
rect 10547 7651 10613 7652
rect 10918 7581 10978 688603
rect 166395 687172 166461 687173
rect 166395 687108 166396 687172
rect 166460 687108 166461 687172
rect 166395 687107 166461 687108
rect 177619 687172 177685 687173
rect 177619 687108 177620 687172
rect 177684 687108 177685 687172
rect 177619 687107 177685 687108
rect 13090 685750 19110 685810
rect 10915 7580 10981 7581
rect 10915 7516 10916 7580
rect 10980 7516 10981 7580
rect 10915 7515 10981 7516
rect 10179 7444 10245 7445
rect 10179 7380 10180 7444
rect 10244 7380 10245 7444
rect 10179 7379 10245 7380
rect 24700 7000 25300 687000
rect 62700 7000 63300 687000
rect 95187 686492 95253 686493
rect 95187 686428 95188 686492
rect 95252 686428 95253 686492
rect 95187 686427 95253 686428
rect 93899 686356 93965 686357
rect 93899 686292 93900 686356
rect 93964 686292 93965 686356
rect 93899 686291 93965 686292
rect 93902 685218 93962 686291
rect 95190 685898 95250 686427
rect 100700 7000 101300 687000
rect 103283 686356 103349 686357
rect 103283 686292 103284 686356
rect 103348 686292 103349 686356
rect 103283 686291 103349 686292
rect 108251 686356 108317 686357
rect 108251 686292 108252 686356
rect 108316 686292 108317 686356
rect 108251 686291 108317 686292
rect 113035 686356 113101 686357
rect 113035 686292 113036 686356
rect 113100 686292 113101 686356
rect 113035 686291 113101 686292
rect 103286 685218 103346 686291
rect 108254 685898 108314 686291
rect 113038 685218 113098 686291
rect 138700 7000 139300 687000
rect 166398 686578 166458 687107
rect 164190 685750 167046 685810
rect 164190 685218 164250 685750
rect 176700 7000 177300 687000
rect 177622 685898 177682 687107
rect 212395 687172 212461 687173
rect 212395 687108 212396 687172
rect 212460 687108 212461 687172
rect 212395 687107 212461 687108
rect 212398 686578 212458 687107
rect 235211 687172 235277 687173
rect 235211 687108 235212 687172
rect 235276 687108 235277 687172
rect 235211 687107 235277 687108
rect 182219 686356 182285 686357
rect 182219 686292 182220 686356
rect 182284 686292 182285 686356
rect 182219 686291 182285 686292
rect 186267 686356 186333 686357
rect 186267 686292 186268 686356
rect 186332 686292 186333 686356
rect 186267 686291 186333 686292
rect 182222 685898 182282 686291
rect 186270 685898 186330 686291
rect 195434 685750 195934 685810
rect 214700 7000 215300 687000
rect 235214 685898 235274 687107
rect 240179 686492 240245 686493
rect 240179 686428 240180 686492
rect 240244 686428 240245 686492
rect 240179 686427 240245 686428
rect 240182 685898 240242 686427
rect 252700 7000 253300 687000
rect 290700 7000 291300 687000
rect 328700 7000 329300 687000
rect 340830 686357 340890 688739
rect 564571 688668 564637 688669
rect 564571 688604 564572 688668
rect 564636 688604 564637 688668
rect 564571 688603 564637 688604
rect 340643 686356 340709 686357
rect 340643 686292 340644 686356
rect 340708 686292 340709 686356
rect 340643 686291 340709 686292
rect 340827 686356 340893 686357
rect 340827 686292 340828 686356
rect 340892 686292 340893 686356
rect 340827 686291 340893 686292
rect 340646 685898 340706 686291
rect 366700 7000 367300 687000
rect 404700 7000 405300 687000
rect 442700 7000 443300 687000
rect 480700 7000 481300 687000
rect 518700 7000 519300 687000
rect 556700 7000 557300 687000
rect 564574 3909 564634 688603
rect 564758 7717 564818 688875
rect 566043 688804 566109 688805
rect 566043 688740 566044 688804
rect 566108 688740 566109 688804
rect 566043 688739 566109 688740
rect 565859 686356 565925 686357
rect 565859 686292 565860 686356
rect 565924 686292 565925 686356
rect 565859 686291 565925 686292
rect 564755 7716 564821 7717
rect 564755 7652 564756 7716
rect 564820 7652 564821 7716
rect 564755 7651 564821 7652
rect 564571 3908 564637 3909
rect 564571 3844 564572 3908
rect 564636 3844 564637 3908
rect 564571 3843 564637 3844
rect 565862 3229 565922 686291
rect 566046 7581 566106 688739
rect 566043 7580 566109 7581
rect 566043 7516 566044 7580
rect 566108 7516 566109 7580
rect 566043 7515 566109 7516
rect 565859 3228 565925 3229
rect 565859 3164 565860 3228
rect 565924 3164 565925 3228
rect 565859 3163 565925 3164
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 585320 -346 585920 704282
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect -2916 -1502 -2734 -1266
rect -2498 -1502 -2316 -1266
rect -2916 -1586 -2316 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 -2316 -1586
rect -2916 -1844 -2316 -1822
rect 586240 -1266 586840 705202
rect 586240 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect 586240 -1586 586840 -1502
rect 586240 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect 586240 -1844 586840 -1822
rect -3836 -2422 -3654 -2186
rect -3418 -2422 -3236 -2186
rect -3836 -2506 -3236 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 -3236 -2506
rect -3836 -2764 -3236 -2742
rect 587160 -2186 587760 706122
rect 587160 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect 587160 -2506 587760 -2422
rect 587160 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect 587160 -2764 587760 -2742
rect -4756 -3342 -4574 -3106
rect -4338 -3342 -4156 -3106
rect -4756 -3426 -4156 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 -4156 -3426
rect -4756 -3684 -4156 -3662
rect 588080 -3106 588680 707042
rect 588080 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect 588080 -3426 588680 -3342
rect 588080 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect 588080 -3684 588680 -3662
rect -5676 -4262 -5494 -4026
rect -5258 -4262 -5076 -4026
rect -5676 -4346 -5076 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 -5076 -4346
rect -5676 -4604 -5076 -4582
rect 589000 -4026 589600 707962
rect 589000 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect 589000 -4346 589600 -4262
rect 589000 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect 589000 -4604 589600 -4582
rect -6596 -5182 -6414 -4946
rect -6178 -5182 -5996 -4946
rect -6596 -5266 -5996 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 -5996 -5266
rect -6596 -5524 -5996 -5502
rect 589920 -4946 590520 708882
rect 589920 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect 589920 -5266 590520 -5182
rect 589920 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect 589920 -5524 590520 -5502
rect -7516 -6102 -7334 -5866
rect -7098 -6102 -6916 -5866
rect -7516 -6186 -6916 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 -6916 -6186
rect -7516 -6444 -6916 -6422
rect 590840 -5866 591440 709802
rect 590840 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect 590840 -6186 591440 -6102
rect 590840 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect 590840 -6444 591440 -6422
rect -8436 -7022 -8254 -6786
rect -8018 -7022 -7836 -6786
rect -8436 -7106 -7836 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 -7836 -7106
rect -8436 -7364 -7836 -7342
rect 591760 -6786 592360 710722
rect 591760 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect 591760 -7106 592360 -7022
rect 591760 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect 591760 -7364 592360 -7342
<< via4 >>
rect -8254 711042 -8018 711278
rect -8254 710722 -8018 710958
rect 591942 711042 592178 711278
rect 591942 710722 592178 710958
rect -7334 710122 -7098 710358
rect -7334 709802 -7098 710038
rect 591022 710122 591258 710358
rect 591022 709802 591258 710038
rect -6414 709202 -6178 709438
rect -6414 708882 -6178 709118
rect 590102 709202 590338 709438
rect 590102 708882 590338 709118
rect -5494 708282 -5258 708518
rect -5494 707962 -5258 708198
rect 589182 708282 589418 708518
rect 589182 707962 589418 708198
rect -4574 707362 -4338 707598
rect -4574 707042 -4338 707278
rect 588262 707362 588498 707598
rect 588262 707042 588498 707278
rect -3654 706442 -3418 706678
rect -3654 706122 -3418 706358
rect 587342 706442 587578 706678
rect 587342 706122 587578 706358
rect -2734 705522 -2498 705758
rect -2734 705202 -2498 705438
rect 586422 705522 586658 705758
rect 586422 705202 586658 705438
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 10462 684302 10698 684538
rect 202742 687172 202978 687258
rect 202742 687108 202828 687172
rect 202828 687108 202892 687172
rect 202892 687108 202978 687172
rect 12486 686492 12722 686578
rect 12486 686428 12572 686492
rect 12572 686428 12636 686492
rect 12636 686428 12722 686492
rect 12486 686342 12722 686428
rect 12854 685662 13090 685898
rect 19110 685662 19346 685898
rect 99886 686492 100122 686578
rect 99886 686428 99972 686492
rect 99972 686428 100036 686492
rect 100036 686428 100122 686492
rect 99886 686342 100122 686428
rect 95102 685662 95338 685898
rect 93814 684982 94050 685218
rect 108166 685662 108402 685898
rect 103198 684982 103434 685218
rect 112950 684982 113186 685218
rect 166310 686342 166546 686578
rect 167046 685662 167282 685898
rect 164102 684982 164338 685218
rect 202742 687022 202978 687108
rect 230342 687172 230578 687258
rect 230342 687108 230428 687172
rect 230428 687108 230492 687172
rect 230492 687108 230578 687172
rect 230342 687022 230578 687108
rect 212310 686342 212546 686578
rect 177534 685662 177770 685898
rect 182134 685662 182370 685898
rect 186182 685662 186418 685898
rect 195198 685662 195434 685898
rect 195934 685662 196170 685898
rect 249478 686492 249714 686578
rect 249478 686428 249564 686492
rect 249564 686428 249628 686492
rect 249628 686428 249714 686492
rect 249478 686342 249714 686428
rect 235126 685662 235362 685898
rect 240094 685662 240330 685898
rect 324366 686492 324602 686578
rect 324366 686428 324452 686492
rect 324452 686428 324516 686492
rect 324516 686428 324602 686492
rect 324366 686342 324602 686428
rect 340558 685662 340794 685898
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect -2734 -1502 -2498 -1266
rect -2734 -1822 -2498 -1586
rect 586422 -1502 586658 -1266
rect 586422 -1822 586658 -1586
rect -3654 -2422 -3418 -2186
rect -3654 -2742 -3418 -2506
rect 587342 -2422 587578 -2186
rect 587342 -2742 587578 -2506
rect -4574 -3342 -4338 -3106
rect -4574 -3662 -4338 -3426
rect 588262 -3342 588498 -3106
rect 588262 -3662 588498 -3426
rect -5494 -4262 -5258 -4026
rect -5494 -4582 -5258 -4346
rect 589182 -4262 589418 -4026
rect 589182 -4582 589418 -4346
rect -6414 -5182 -6178 -4946
rect -6414 -5502 -6178 -5266
rect 590102 -5182 590338 -4946
rect 590102 -5502 590338 -5266
rect -7334 -6102 -7098 -5866
rect -7334 -6422 -7098 -6186
rect 591022 -6102 591258 -5866
rect 591022 -6422 591258 -6186
rect -8254 -7022 -8018 -6786
rect -8254 -7342 -8018 -7106
rect 591942 -7022 592178 -6786
rect 591942 -7342 592178 -7106
<< metal5 >>
rect -8436 711300 -7836 711302
rect 591760 711300 592360 711302
rect -8436 711278 592360 711300
rect -8436 711042 -8254 711278
rect -8018 711042 591942 711278
rect 592178 711042 592360 711278
rect -8436 710958 592360 711042
rect -8436 710722 -8254 710958
rect -8018 710722 591942 710958
rect 592178 710722 592360 710958
rect -8436 710700 592360 710722
rect -8436 710698 -7836 710700
rect 591760 710698 592360 710700
rect -7516 710380 -6916 710382
rect 590840 710380 591440 710382
rect -7516 710358 591440 710380
rect -7516 710122 -7334 710358
rect -7098 710122 591022 710358
rect 591258 710122 591440 710358
rect -7516 710038 591440 710122
rect -7516 709802 -7334 710038
rect -7098 709802 591022 710038
rect 591258 709802 591440 710038
rect -7516 709780 591440 709802
rect -7516 709778 -6916 709780
rect 590840 709778 591440 709780
rect -6596 709460 -5996 709462
rect 589920 709460 590520 709462
rect -6596 709438 590520 709460
rect -6596 709202 -6414 709438
rect -6178 709202 590102 709438
rect 590338 709202 590520 709438
rect -6596 709118 590520 709202
rect -6596 708882 -6414 709118
rect -6178 708882 590102 709118
rect 590338 708882 590520 709118
rect -6596 708860 590520 708882
rect -6596 708858 -5996 708860
rect 589920 708858 590520 708860
rect -5676 708540 -5076 708542
rect 589000 708540 589600 708542
rect -5676 708518 589600 708540
rect -5676 708282 -5494 708518
rect -5258 708282 589182 708518
rect 589418 708282 589600 708518
rect -5676 708198 589600 708282
rect -5676 707962 -5494 708198
rect -5258 707962 589182 708198
rect 589418 707962 589600 708198
rect -5676 707940 589600 707962
rect -5676 707938 -5076 707940
rect 589000 707938 589600 707940
rect -4756 707620 -4156 707622
rect 588080 707620 588680 707622
rect -4756 707598 588680 707620
rect -4756 707362 -4574 707598
rect -4338 707362 588262 707598
rect 588498 707362 588680 707598
rect -4756 707278 588680 707362
rect -4756 707042 -4574 707278
rect -4338 707042 588262 707278
rect 588498 707042 588680 707278
rect -4756 707020 588680 707042
rect -4756 707018 -4156 707020
rect 588080 707018 588680 707020
rect -3836 706700 -3236 706702
rect 587160 706700 587760 706702
rect -3836 706678 587760 706700
rect -3836 706442 -3654 706678
rect -3418 706442 587342 706678
rect 587578 706442 587760 706678
rect -3836 706358 587760 706442
rect -3836 706122 -3654 706358
rect -3418 706122 587342 706358
rect 587578 706122 587760 706358
rect -3836 706100 587760 706122
rect -3836 706098 -3236 706100
rect 587160 706098 587760 706100
rect -2916 705780 -2316 705782
rect 586240 705780 586840 705782
rect -2916 705758 586840 705780
rect -2916 705522 -2734 705758
rect -2498 705522 586422 705758
rect 586658 705522 586840 705758
rect -2916 705438 586840 705522
rect -2916 705202 -2734 705438
rect -2498 705202 586422 705438
rect 586658 705202 586840 705438
rect -2916 705180 586840 705202
rect -2916 705178 -2316 705180
rect 586240 705178 586840 705180
rect -1996 704860 -1396 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 585320 704258 585920 704260
rect 195892 687258 203020 687300
rect 195892 687022 202742 687258
rect 202978 687022 203020 687258
rect 195892 686980 203020 687022
rect 224596 687258 230620 687300
rect 224596 687022 230342 687258
rect 230578 687022 230620 687258
rect 224596 686980 230620 687022
rect 12260 686578 12764 686620
rect 12260 686342 12486 686578
rect 12722 686342 12764 686578
rect 12260 686300 12764 686342
rect 12260 685940 12580 686300
rect 31396 685940 31900 686620
rect 50716 685940 51220 686620
rect 70036 685940 70540 686620
rect 89356 685940 89860 686620
rect 99844 686578 109180 686620
rect 99844 686342 99886 686578
rect 100122 686342 109180 686578
rect 99844 686300 109180 686342
rect 108860 685940 109180 686300
rect 127996 685940 128500 686620
rect 147316 685940 147820 686620
rect 166268 686578 166588 686620
rect 166268 686342 166310 686578
rect 166546 686342 166588 686578
rect 166268 685940 166588 686342
rect 12260 685898 13132 685940
rect 12260 685662 12854 685898
rect 13090 685662 13132 685898
rect 12260 685620 13132 685662
rect 19068 685898 95380 685940
rect 19068 685662 19110 685898
rect 19346 685662 95102 685898
rect 95338 685662 95380 685898
rect 19068 685620 95380 685662
rect 103340 685898 108444 685940
rect 103340 685662 108166 685898
rect 108402 685662 108444 685898
rect 103340 685620 108444 685662
rect 108860 685620 166588 685940
rect 167004 685898 173764 685940
rect 167004 685662 167046 685898
rect 167282 685662 173764 685898
rect 167004 685620 173764 685662
rect 177492 685898 182412 685940
rect 177492 685662 177534 685898
rect 177770 685662 182134 685898
rect 182370 685662 182412 685898
rect 177492 685620 182412 685662
rect 186140 685898 195476 685940
rect 186140 685662 186182 685898
rect 186418 685662 195198 685898
rect 195434 685662 195476 685898
rect 186140 685620 195476 685662
rect 195892 685898 196212 686980
rect 224596 686620 224916 686980
rect 212268 686578 215532 686620
rect 212268 686342 212310 686578
rect 212546 686342 215532 686578
rect 212268 686300 215532 686342
rect 215212 685940 215532 686300
rect 224228 686300 224916 686620
rect 249436 686578 254172 686620
rect 249436 686342 249478 686578
rect 249714 686342 254172 686578
rect 249436 686300 254172 686342
rect 224228 685940 224548 686300
rect 253852 685940 254172 686300
rect 263236 686300 273492 686620
rect 263236 685940 263556 686300
rect 195892 685662 195934 685898
rect 196170 685662 196212 685898
rect 195892 685620 196212 685662
rect 196812 685620 205412 685940
rect 215212 685620 224548 685940
rect 235084 685898 240372 685940
rect 235084 685662 235126 685898
rect 235362 685662 240094 685898
rect 240330 685662 240372 685898
rect 235084 685620 240372 685662
rect 253852 685620 263556 685940
rect 273172 685940 273492 686300
rect 282556 686300 292812 686620
rect 282556 685940 282876 686300
rect 273172 685620 282876 685940
rect 292492 685940 292812 686300
rect 301876 686300 312132 686620
rect 301876 685940 302196 686300
rect 292492 685620 302196 685940
rect 311812 685940 312132 686300
rect 320828 686578 324644 686620
rect 320828 686342 324366 686578
rect 324602 686342 324644 686578
rect 320828 686300 324644 686342
rect 320828 685940 321148 686300
rect 311812 685620 321148 685940
rect 322116 685898 340836 685940
rect 322116 685662 340558 685898
rect 340794 685662 340836 685898
rect 322116 685620 340836 685662
rect 103340 685260 103660 685620
rect 12260 685218 94092 685260
rect 12260 684982 93814 685218
rect 94050 684982 94092 685218
rect 12260 684940 94092 684982
rect 103156 685218 103660 685260
rect 103156 684982 103198 685218
rect 103434 684982 103660 685218
rect 12260 684580 12580 684940
rect 10420 684538 12580 684580
rect 10420 684302 10462 684538
rect 10698 684302 12580 684538
rect 10420 684260 12580 684302
rect 31396 684260 31900 684940
rect 50716 684260 51220 684940
rect 70036 684260 70540 684940
rect 89356 684260 89860 684940
rect 103156 684260 103660 684982
rect 112908 685218 113228 685260
rect 112908 684982 112950 685218
rect 113186 684982 113228 685218
rect 112908 684580 113228 684982
rect 122476 685218 164380 685260
rect 122476 684982 164102 685218
rect 164338 684982 164380 685218
rect 122476 684940 164380 684982
rect 122476 684580 122796 684940
rect 112908 684260 122796 684580
rect 147316 684260 147820 684940
rect 173444 683900 173764 685620
rect 177124 684940 185908 685260
rect 177124 684580 177444 684940
rect 176572 684260 177444 684580
rect 185588 684580 185908 684940
rect 186692 684940 193452 685260
rect 186692 684580 187012 684940
rect 185588 684260 187012 684580
rect 176572 683900 176892 684260
rect 173444 683580 176892 683900
rect 185956 683580 186460 684260
rect 193132 683900 193452 684940
rect 196812 683900 197132 685620
rect 205092 685260 205412 685620
rect 205092 684940 205780 685260
rect 205460 684580 205780 684940
rect 215212 684940 224916 685260
rect 215212 684580 215532 684940
rect 205460 684260 215532 684580
rect 224596 684580 224916 684940
rect 234532 684940 244236 685260
rect 234532 684580 234852 684940
rect 224596 684260 234852 684580
rect 243916 684580 244236 684940
rect 260476 684940 263556 685260
rect 243916 684260 251412 684580
rect 193132 683580 197132 683900
rect 251092 683220 251412 684260
rect 260476 683220 260796 684940
rect 263236 684580 263556 684940
rect 279796 684940 282876 685260
rect 263236 684260 270732 684580
rect 251092 682900 260796 683220
rect 270412 683220 270732 684260
rect 279796 683220 280116 684940
rect 282556 684580 282876 684940
rect 299116 684940 302196 685260
rect 282556 684260 290052 684580
rect 270412 682900 280116 683220
rect 289732 683220 290052 684260
rect 299116 683220 299436 684940
rect 301876 684580 302196 684940
rect 318436 684940 321148 685260
rect 301876 684260 309372 684580
rect 289732 682900 299436 683220
rect 309052 683220 309372 684260
rect 318436 683220 318756 684940
rect 320828 684580 321148 684940
rect 322116 684580 322436 685620
rect 320828 684260 322436 684580
rect 309052 682900 318756 683220
rect -1996 -324 -1396 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 585320 -926 585920 -924
rect -2916 -1244 -2316 -1242
rect 586240 -1244 586840 -1242
rect -2916 -1266 586840 -1244
rect -2916 -1502 -2734 -1266
rect -2498 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect -2916 -1586 586840 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect -2916 -1844 586840 -1822
rect -2916 -1846 -2316 -1844
rect 586240 -1846 586840 -1844
rect -3836 -2164 -3236 -2162
rect 587160 -2164 587760 -2162
rect -3836 -2186 587760 -2164
rect -3836 -2422 -3654 -2186
rect -3418 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect -3836 -2506 587760 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect -3836 -2764 587760 -2742
rect -3836 -2766 -3236 -2764
rect 587160 -2766 587760 -2764
rect -4756 -3084 -4156 -3082
rect 588080 -3084 588680 -3082
rect -4756 -3106 588680 -3084
rect -4756 -3342 -4574 -3106
rect -4338 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect -4756 -3426 588680 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect -4756 -3684 588680 -3662
rect -4756 -3686 -4156 -3684
rect 588080 -3686 588680 -3684
rect -5676 -4004 -5076 -4002
rect 589000 -4004 589600 -4002
rect -5676 -4026 589600 -4004
rect -5676 -4262 -5494 -4026
rect -5258 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect -5676 -4346 589600 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect -5676 -4604 589600 -4582
rect -5676 -4606 -5076 -4604
rect 589000 -4606 589600 -4604
rect -6596 -4924 -5996 -4922
rect 589920 -4924 590520 -4922
rect -6596 -4946 590520 -4924
rect -6596 -5182 -6414 -4946
rect -6178 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect -6596 -5266 590520 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect -6596 -5524 590520 -5502
rect -6596 -5526 -5996 -5524
rect 589920 -5526 590520 -5524
rect -7516 -5844 -6916 -5842
rect 590840 -5844 591440 -5842
rect -7516 -5866 591440 -5844
rect -7516 -6102 -7334 -5866
rect -7098 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect -7516 -6186 591440 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect -7516 -6444 591440 -6422
rect -7516 -6446 -6916 -6444
rect 590840 -6446 591440 -6444
rect -8436 -6764 -7836 -6762
rect 591760 -6764 592360 -6762
rect -8436 -6786 592360 -6764
rect -8436 -7022 -8254 -6786
rect -8018 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect -8436 -7106 592360 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect -8436 -7364 592360 -7342
rect -8436 -7366 -7836 -7364
rect 591760 -7366 592360 -7364
use fpga  fpga250
timestamp 1608015108
transform 1 0 7000 0 1 7000
box 0 0 570000 680000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2916 -1844 586840 -1244 8 vssd1
port 637 nsew default input
rlabel metal5 s -3836 -2764 587760 -2164 8 vccd2
port 638 nsew default input
rlabel metal5 s -4756 -3684 588680 -3084 8 vssd2
port 639 nsew default input
rlabel metal5 s -5676 -4604 589600 -4004 8 vdda1
port 640 nsew default input
rlabel metal5 s -6596 -5524 590520 -4924 8 vssa1
port 641 nsew default input
rlabel metal5 s -7516 -6444 591440 -5844 8 vdda2
port 642 nsew default input
rlabel metal5 s -8436 -7364 592360 -6764 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>

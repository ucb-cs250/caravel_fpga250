VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga
  CLASS BLOCK ;
  FOREIGN fpga ;
  ORIGIN 0.000 0.000 ;
  SIZE 2745.000 BY 3320.000 ;
  PIN gpio_east[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 66.000 2745.000 66.600 ;
    END
  END gpio_east[0]
  PIN gpio_east[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 198.600 2745.000 199.200 ;
    END
  END gpio_east[1]
  PIN gpio_east[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 331.200 2745.000 331.800 ;
    END
  END gpio_east[2]
  PIN gpio_east[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 463.800 2745.000 464.400 ;
    END
  END gpio_east[3]
  PIN gpio_east[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 597.080 2745.000 597.680 ;
    END
  END gpio_east[4]
  PIN gpio_east[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 729.680 2745.000 730.280 ;
    END
  END gpio_east[5]
  PIN gpio_east[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 862.280 2745.000 862.880 ;
    END
  END gpio_east[6]
  PIN gpio_east[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 994.880 2745.000 995.480 ;
    END
  END gpio_east[7]
  PIN gpio_east[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 1128.160 2745.000 1128.760 ;
    END
  END gpio_east[8]
  PIN gpio_east[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 1260.760 2745.000 1261.360 ;
    END
  END gpio_east[9]
  PIN gpio_north[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 54.830 3316.000 55.110 3320.000 ;
    END
  END gpio_north[0]
  PIN gpio_north[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 164.310 3316.000 164.590 3320.000 ;
    END
  END gpio_north[1]
  PIN gpio_north[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 274.250 3316.000 274.530 3320.000 ;
    END
  END gpio_north[2]
  PIN gpio_north[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 384.190 3316.000 384.470 3320.000 ;
    END
  END gpio_north[3]
  PIN gpio_north[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 493.670 3316.000 493.950 3320.000 ;
    END
  END gpio_north[4]
  PIN gpio_north[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 603.610 3316.000 603.890 3320.000 ;
    END
  END gpio_north[5]
  PIN gpio_north[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 713.550 3316.000 713.830 3320.000 ;
    END
  END gpio_north[6]
  PIN gpio_north[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 823.030 3316.000 823.310 3320.000 ;
    END
  END gpio_north[7]
  PIN gpio_north[8]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.970 3316.000 933.250 3320.000 ;
    END
  END gpio_north[8]
  PIN gpio_north[9]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1042.910 3316.000 1043.190 3320.000 ;
    END
  END gpio_north[9]
  PIN gpio_south[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END gpio_south[0]
  PIN gpio_south[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END gpio_south[1]
  PIN gpio_south[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END gpio_south[2]
  PIN gpio_south[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 162.470 0.000 162.750 4.000 ;
    END
  END gpio_south[3]
  PIN gpio_south[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 208.930 0.000 209.210 4.000 ;
    END
  END gpio_south[4]
  PIN gpio_south[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 255.390 0.000 255.670 4.000 ;
    END
  END gpio_south[5]
  PIN gpio_south[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END gpio_south[6]
  PIN gpio_south[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 348.310 0.000 348.590 4.000 ;
    END
  END gpio_south[7]
  PIN gpio_west[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 4.000 47.560 ;
    END
  END gpio_west[0]
  PIN gpio_west[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END gpio_west[1]
  PIN gpio_west[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.000 4.000 236.600 ;
    END
  END gpio_west[2]
  PIN gpio_west[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.200 4.000 331.800 ;
    END
  END gpio_west[3]
  PIN gpio_west[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 4.000 426.320 ;
    END
  END gpio_west[4]
  PIN gpio_west[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.920 4.000 521.520 ;
    END
  END gpio_west[5]
  PIN gpio_west[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 615.440 4.000 616.040 ;
    END
  END gpio_west[6]
  PIN gpio_west[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 710.640 4.000 711.240 ;
    END
  END gpio_west[7]
  PIN gpio_west[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 805.160 4.000 805.760 ;
    END
  END gpio_west[8]
  PIN gpio_west[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 900.360 4.000 900.960 ;
    END
  END gpio_west[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 994.880 4.000 995.480 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1152.390 3316.000 1152.670 3320.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2741.000 1393.360 2745.000 1393.960 ;
    END
  END wbs_ack_o
  PIN wbs_addr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1090.080 4.000 1090.680 ;
    END
  END wbs_addr_i[0]
  PIN wbs_addr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1883.790 0.000 1884.070 4.000 ;
    END
  END wbs_addr_i[10]
  PIN wbs_addr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1469.520 4.000 1470.120 ;
    END
  END wbs_addr_i[11]
  PIN wbs_addr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1930.250 0.000 1930.530 4.000 ;
    END
  END wbs_addr_i[12]
  PIN wbs_addr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1481.750 3316.000 1482.030 3320.000 ;
    END
  END wbs_addr_i[13]
  PIN wbs_addr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1591.690 3316.000 1591.970 3320.000 ;
    END
  END wbs_addr_i[14]
  PIN wbs_addr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1564.040 4.000 1564.640 ;
    END
  END wbs_addr_i[15]
  PIN wbs_addr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 2057.720 2745.000 2058.320 ;
    END
  END wbs_addr_i[16]
  PIN wbs_addr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1659.240 4.000 1659.840 ;
    END
  END wbs_addr_i[17]
  PIN wbs_addr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1701.630 3316.000 1701.910 3320.000 ;
    END
  END wbs_addr_i[18]
  PIN wbs_addr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1976.710 0.000 1976.990 4.000 ;
    END
  END wbs_addr_i[19]
  PIN wbs_addr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 1526.640 2745.000 1527.240 ;
    END
  END wbs_addr_i[1]
  PIN wbs_addr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1753.760 4.000 1754.360 ;
    END
  END wbs_addr_i[20]
  PIN wbs_addr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2023.170 0.000 2023.450 4.000 ;
    END
  END wbs_addr_i[21]
  PIN wbs_addr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2069.630 0.000 2069.910 4.000 ;
    END
  END wbs_addr_i[22]
  PIN wbs_addr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 2190.320 2745.000 2190.920 ;
    END
  END wbs_addr_i[23]
  PIN wbs_addr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2116.550 0.000 2116.830 4.000 ;
    END
  END wbs_addr_i[24]
  PIN wbs_addr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1848.960 4.000 1849.560 ;
    END
  END wbs_addr_i[25]
  PIN wbs_addr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2163.010 0.000 2163.290 4.000 ;
    END
  END wbs_addr_i[26]
  PIN wbs_addr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2209.470 0.000 2209.750 4.000 ;
    END
  END wbs_addr_i[27]
  PIN wbs_addr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2255.930 0.000 2256.210 4.000 ;
    END
  END wbs_addr_i[28]
  PIN wbs_addr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1943.480 4.000 1944.080 ;
    END
  END wbs_addr_i[29]
  PIN wbs_addr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1262.330 3316.000 1262.610 3320.000 ;
    END
  END wbs_addr_i[2]
  PIN wbs_addr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2038.680 4.000 2039.280 ;
    END
  END wbs_addr_i[30]
  PIN wbs_addr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2302.390 0.000 2302.670 4.000 ;
    END
  END wbs_addr_i[31]
  PIN wbs_addr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 1659.240 2745.000 1659.840 ;
    END
  END wbs_addr_i[3]
  PIN wbs_addr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1184.600 4.000 1185.200 ;
    END
  END wbs_addr_i[4]
  PIN wbs_addr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1279.800 4.000 1280.400 ;
    END
  END wbs_addr_i[5]
  PIN wbs_addr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1372.270 3316.000 1372.550 3320.000 ;
    END
  END wbs_addr_i[6]
  PIN wbs_addr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1374.320 4.000 1374.920 ;
    END
  END wbs_addr_i[7]
  PIN wbs_addr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 1791.840 2745.000 1792.440 ;
    END
  END wbs_addr_i[8]
  PIN wbs_addr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 1924.440 2745.000 1925.040 ;
    END
  END wbs_addr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1811.110 3316.000 1811.390 3320.000 ;
    END
  END wbs_cyc_i
  PIN wbs_data_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1921.050 3316.000 1921.330 3320.000 ;
    END
  END wbs_data_i[0]
  PIN wbs_data_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2133.200 4.000 2133.800 ;
    END
  END wbs_data_i[10]
  PIN wbs_data_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2250.410 3316.000 2250.690 3320.000 ;
    END
  END wbs_data_i[11]
  PIN wbs_data_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2228.400 4.000 2229.000 ;
    END
  END wbs_data_i[12]
  PIN wbs_data_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2360.350 3316.000 2360.630 3320.000 ;
    END
  END wbs_data_i[13]
  PIN wbs_data_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2322.920 4.000 2323.520 ;
    END
  END wbs_data_i[14]
  PIN wbs_data_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2469.830 3316.000 2470.110 3320.000 ;
    END
  END wbs_data_i[15]
  PIN wbs_data_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2418.120 4.000 2418.720 ;
    END
  END wbs_data_i[16]
  PIN wbs_data_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2579.770 3316.000 2580.050 3320.000 ;
    END
  END wbs_data_i[17]
  PIN wbs_data_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 2854.000 2745.000 2854.600 ;
    END
  END wbs_data_i[18]
  PIN wbs_data_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 2987.280 2745.000 2987.880 ;
    END
  END wbs_data_i[19]
  PIN wbs_data_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 2322.920 2745.000 2323.520 ;
    END
  END wbs_data_i[1]
  PIN wbs_data_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2512.640 4.000 2513.240 ;
    END
  END wbs_data_i[20]
  PIN wbs_data_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2488.690 0.000 2488.970 4.000 ;
    END
  END wbs_data_i[21]
  PIN wbs_data_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 3119.880 2745.000 3120.480 ;
    END
  END wbs_data_i[22]
  PIN wbs_data_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2689.710 3316.000 2689.990 3320.000 ;
    END
  END wbs_data_i[23]
  PIN wbs_data_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2535.150 0.000 2535.430 4.000 ;
    END
  END wbs_data_i[24]
  PIN wbs_data_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2581.610 0.000 2581.890 4.000 ;
    END
  END wbs_data_i[25]
  PIN wbs_data_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2607.840 4.000 2608.440 ;
    END
  END wbs_data_i[26]
  PIN wbs_data_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2702.360 4.000 2702.960 ;
    END
  END wbs_data_i[27]
  PIN wbs_data_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2628.070 0.000 2628.350 4.000 ;
    END
  END wbs_data_i[28]
  PIN wbs_data_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2797.560 4.000 2798.160 ;
    END
  END wbs_data_i[29]
  PIN wbs_data_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2030.990 3316.000 2031.270 3320.000 ;
    END
  END wbs_data_i[2]
  PIN wbs_data_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2674.530 0.000 2674.810 4.000 ;
    END
  END wbs_data_i[30]
  PIN wbs_data_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 3252.480 2745.000 3253.080 ;
    END
  END wbs_data_i[31]
  PIN wbs_data_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2348.850 0.000 2349.130 4.000 ;
    END
  END wbs_data_i[3]
  PIN wbs_data_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2395.310 0.000 2395.590 4.000 ;
    END
  END wbs_data_i[4]
  PIN wbs_data_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 2456.200 2745.000 2456.800 ;
    END
  END wbs_data_i[5]
  PIN wbs_data_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2442.230 0.000 2442.510 4.000 ;
    END
  END wbs_data_i[6]
  PIN wbs_data_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 2588.800 2745.000 2589.400 ;
    END
  END wbs_data_i[7]
  PIN wbs_data_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2140.470 3316.000 2140.750 3320.000 ;
    END
  END wbs_data_i[8]
  PIN wbs_data_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 2721.400 2745.000 2722.000 ;
    END
  END wbs_data_i[9]
  PIN wbs_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 395.230 0.000 395.510 4.000 ;
    END
  END wbs_data_o[0]
  PIN wbs_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 860.290 0.000 860.570 4.000 ;
    END
  END wbs_data_o[10]
  PIN wbs_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 906.750 0.000 907.030 4.000 ;
    END
  END wbs_data_o[11]
  PIN wbs_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 953.210 0.000 953.490 4.000 ;
    END
  END wbs_data_o[12]
  PIN wbs_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 999.670 0.000 999.950 4.000 ;
    END
  END wbs_data_o[13]
  PIN wbs_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1046.130 0.000 1046.410 4.000 ;
    END
  END wbs_data_o[14]
  PIN wbs_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1093.050 0.000 1093.330 4.000 ;
    END
  END wbs_data_o[15]
  PIN wbs_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1139.510 0.000 1139.790 4.000 ;
    END
  END wbs_data_o[16]
  PIN wbs_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1185.970 0.000 1186.250 4.000 ;
    END
  END wbs_data_o[17]
  PIN wbs_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1232.430 0.000 1232.710 4.000 ;
    END
  END wbs_data_o[18]
  PIN wbs_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1278.890 0.000 1279.170 4.000 ;
    END
  END wbs_data_o[19]
  PIN wbs_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 441.690 0.000 441.970 4.000 ;
    END
  END wbs_data_o[1]
  PIN wbs_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1325.350 0.000 1325.630 4.000 ;
    END
  END wbs_data_o[20]
  PIN wbs_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1371.810 0.000 1372.090 4.000 ;
    END
  END wbs_data_o[21]
  PIN wbs_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1418.730 0.000 1419.010 4.000 ;
    END
  END wbs_data_o[22]
  PIN wbs_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1465.190 0.000 1465.470 4.000 ;
    END
  END wbs_data_o[23]
  PIN wbs_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1511.650 0.000 1511.930 4.000 ;
    END
  END wbs_data_o[24]
  PIN wbs_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1558.110 0.000 1558.390 4.000 ;
    END
  END wbs_data_o[25]
  PIN wbs_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1604.570 0.000 1604.850 4.000 ;
    END
  END wbs_data_o[26]
  PIN wbs_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1651.030 0.000 1651.310 4.000 ;
    END
  END wbs_data_o[27]
  PIN wbs_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1697.490 0.000 1697.770 4.000 ;
    END
  END wbs_data_o[28]
  PIN wbs_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1744.410 0.000 1744.690 4.000 ;
    END
  END wbs_data_o[29]
  PIN wbs_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 488.150 0.000 488.430 4.000 ;
    END
  END wbs_data_o[2]
  PIN wbs_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1790.870 0.000 1791.150 4.000 ;
    END
  END wbs_data_o[30]
  PIN wbs_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1837.330 0.000 1837.610 4.000 ;
    END
  END wbs_data_o[31]
  PIN wbs_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 534.610 0.000 534.890 4.000 ;
    END
  END wbs_data_o[3]
  PIN wbs_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 581.070 0.000 581.350 4.000 ;
    END
  END wbs_data_o[4]
  PIN wbs_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 627.530 0.000 627.810 4.000 ;
    END
  END wbs_data_o[5]
  PIN wbs_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 673.990 0.000 674.270 4.000 ;
    END
  END wbs_data_o[6]
  PIN wbs_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 720.910 0.000 721.190 4.000 ;
    END
  END wbs_data_o[7]
  PIN wbs_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 767.370 0.000 767.650 4.000 ;
    END
  END wbs_data_o[8]
  PIN wbs_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 813.830 0.000 814.110 4.000 ;
    END
  END wbs_data_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2720.990 0.000 2721.270 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2892.080 4.000 2892.680 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2987.280 4.000 2987.880 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3081.800 4.000 3082.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3177.000 4.000 3177.600 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3271.520 4.000 3272.120 ;
    END
  END wbs_we_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 2739.300 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 64.785 2739.300 66.385 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2739.300 3307.605 ;
      LAYER met1 ;
        RECT 5.520 4.460 2739.300 3315.640 ;
      LAYER met2 ;
        RECT 13.890 3315.720 54.550 3316.000 ;
        RECT 55.390 3315.720 164.030 3316.000 ;
        RECT 164.870 3315.720 273.970 3316.000 ;
        RECT 274.810 3315.720 383.910 3316.000 ;
        RECT 384.750 3315.720 493.390 3316.000 ;
        RECT 494.230 3315.720 603.330 3316.000 ;
        RECT 604.170 3315.720 713.270 3316.000 ;
        RECT 714.110 3315.720 822.750 3316.000 ;
        RECT 823.590 3315.720 932.690 3316.000 ;
        RECT 933.530 3315.720 1042.630 3316.000 ;
        RECT 1043.470 3315.720 1152.110 3316.000 ;
        RECT 1152.950 3315.720 1262.050 3316.000 ;
        RECT 1262.890 3315.720 1371.990 3316.000 ;
        RECT 1372.830 3315.720 1481.470 3316.000 ;
        RECT 1482.310 3315.720 1591.410 3316.000 ;
        RECT 1592.250 3315.720 1701.350 3316.000 ;
        RECT 1702.190 3315.720 1810.830 3316.000 ;
        RECT 1811.670 3315.720 1920.770 3316.000 ;
        RECT 1921.610 3315.720 2030.710 3316.000 ;
        RECT 2031.550 3315.720 2140.190 3316.000 ;
        RECT 2141.030 3315.720 2250.130 3316.000 ;
        RECT 2250.970 3315.720 2360.070 3316.000 ;
        RECT 2360.910 3315.720 2469.550 3316.000 ;
        RECT 2470.390 3315.720 2579.490 3316.000 ;
        RECT 2580.330 3315.720 2689.430 3316.000 ;
        RECT 2690.270 3315.720 2725.410 3316.000 ;
        RECT 13.890 4.280 2725.410 3315.720 ;
        RECT 13.890 4.000 22.810 4.280 ;
        RECT 23.650 4.000 69.270 4.280 ;
        RECT 70.110 4.000 115.730 4.280 ;
        RECT 116.570 4.000 162.190 4.280 ;
        RECT 163.030 4.000 208.650 4.280 ;
        RECT 209.490 4.000 255.110 4.280 ;
        RECT 255.950 4.000 301.570 4.280 ;
        RECT 302.410 4.000 348.030 4.280 ;
        RECT 348.870 4.000 394.950 4.280 ;
        RECT 395.790 4.000 441.410 4.280 ;
        RECT 442.250 4.000 487.870 4.280 ;
        RECT 488.710 4.000 534.330 4.280 ;
        RECT 535.170 4.000 580.790 4.280 ;
        RECT 581.630 4.000 627.250 4.280 ;
        RECT 628.090 4.000 673.710 4.280 ;
        RECT 674.550 4.000 720.630 4.280 ;
        RECT 721.470 4.000 767.090 4.280 ;
        RECT 767.930 4.000 813.550 4.280 ;
        RECT 814.390 4.000 860.010 4.280 ;
        RECT 860.850 4.000 906.470 4.280 ;
        RECT 907.310 4.000 952.930 4.280 ;
        RECT 953.770 4.000 999.390 4.280 ;
        RECT 1000.230 4.000 1045.850 4.280 ;
        RECT 1046.690 4.000 1092.770 4.280 ;
        RECT 1093.610 4.000 1139.230 4.280 ;
        RECT 1140.070 4.000 1185.690 4.280 ;
        RECT 1186.530 4.000 1232.150 4.280 ;
        RECT 1232.990 4.000 1278.610 4.280 ;
        RECT 1279.450 4.000 1325.070 4.280 ;
        RECT 1325.910 4.000 1371.530 4.280 ;
        RECT 1372.370 4.000 1418.450 4.280 ;
        RECT 1419.290 4.000 1464.910 4.280 ;
        RECT 1465.750 4.000 1511.370 4.280 ;
        RECT 1512.210 4.000 1557.830 4.280 ;
        RECT 1558.670 4.000 1604.290 4.280 ;
        RECT 1605.130 4.000 1650.750 4.280 ;
        RECT 1651.590 4.000 1697.210 4.280 ;
        RECT 1698.050 4.000 1744.130 4.280 ;
        RECT 1744.970 4.000 1790.590 4.280 ;
        RECT 1791.430 4.000 1837.050 4.280 ;
        RECT 1837.890 4.000 1883.510 4.280 ;
        RECT 1884.350 4.000 1929.970 4.280 ;
        RECT 1930.810 4.000 1976.430 4.280 ;
        RECT 1977.270 4.000 2022.890 4.280 ;
        RECT 2023.730 4.000 2069.350 4.280 ;
        RECT 2070.190 4.000 2116.270 4.280 ;
        RECT 2117.110 4.000 2162.730 4.280 ;
        RECT 2163.570 4.000 2209.190 4.280 ;
        RECT 2210.030 4.000 2255.650 4.280 ;
        RECT 2256.490 4.000 2302.110 4.280 ;
        RECT 2302.950 4.000 2348.570 4.280 ;
        RECT 2349.410 4.000 2395.030 4.280 ;
        RECT 2395.870 4.000 2441.950 4.280 ;
        RECT 2442.790 4.000 2488.410 4.280 ;
        RECT 2489.250 4.000 2534.870 4.280 ;
        RECT 2535.710 4.000 2581.330 4.280 ;
        RECT 2582.170 4.000 2627.790 4.280 ;
        RECT 2628.630 4.000 2674.250 4.280 ;
        RECT 2675.090 4.000 2720.710 4.280 ;
        RECT 2721.550 4.000 2725.410 4.280 ;
      LAYER met3 ;
        RECT 4.000 3272.520 2741.000 3307.685 ;
        RECT 4.400 3271.120 2741.000 3272.520 ;
        RECT 4.000 3253.480 2741.000 3271.120 ;
        RECT 4.000 3252.080 2740.600 3253.480 ;
        RECT 4.000 3178.000 2741.000 3252.080 ;
        RECT 4.400 3176.600 2741.000 3178.000 ;
        RECT 4.000 3120.880 2741.000 3176.600 ;
        RECT 4.000 3119.480 2740.600 3120.880 ;
        RECT 4.000 3082.800 2741.000 3119.480 ;
        RECT 4.400 3081.400 2741.000 3082.800 ;
        RECT 4.000 2988.280 2741.000 3081.400 ;
        RECT 4.400 2986.880 2740.600 2988.280 ;
        RECT 4.000 2893.080 2741.000 2986.880 ;
        RECT 4.400 2891.680 2741.000 2893.080 ;
        RECT 4.000 2855.000 2741.000 2891.680 ;
        RECT 4.000 2853.600 2740.600 2855.000 ;
        RECT 4.000 2798.560 2741.000 2853.600 ;
        RECT 4.400 2797.160 2741.000 2798.560 ;
        RECT 4.000 2722.400 2741.000 2797.160 ;
        RECT 4.000 2721.000 2740.600 2722.400 ;
        RECT 4.000 2703.360 2741.000 2721.000 ;
        RECT 4.400 2701.960 2741.000 2703.360 ;
        RECT 4.000 2608.840 2741.000 2701.960 ;
        RECT 4.400 2607.440 2741.000 2608.840 ;
        RECT 4.000 2589.800 2741.000 2607.440 ;
        RECT 4.000 2588.400 2740.600 2589.800 ;
        RECT 4.000 2513.640 2741.000 2588.400 ;
        RECT 4.400 2512.240 2741.000 2513.640 ;
        RECT 4.000 2457.200 2741.000 2512.240 ;
        RECT 4.000 2455.800 2740.600 2457.200 ;
        RECT 4.000 2419.120 2741.000 2455.800 ;
        RECT 4.400 2417.720 2741.000 2419.120 ;
        RECT 4.000 2323.920 2741.000 2417.720 ;
        RECT 4.400 2322.520 2740.600 2323.920 ;
        RECT 4.000 2229.400 2741.000 2322.520 ;
        RECT 4.400 2228.000 2741.000 2229.400 ;
        RECT 4.000 2191.320 2741.000 2228.000 ;
        RECT 4.000 2189.920 2740.600 2191.320 ;
        RECT 4.000 2134.200 2741.000 2189.920 ;
        RECT 4.400 2132.800 2741.000 2134.200 ;
        RECT 4.000 2058.720 2741.000 2132.800 ;
        RECT 4.000 2057.320 2740.600 2058.720 ;
        RECT 4.000 2039.680 2741.000 2057.320 ;
        RECT 4.400 2038.280 2741.000 2039.680 ;
        RECT 4.000 1944.480 2741.000 2038.280 ;
        RECT 4.400 1943.080 2741.000 1944.480 ;
        RECT 4.000 1925.440 2741.000 1943.080 ;
        RECT 4.000 1924.040 2740.600 1925.440 ;
        RECT 4.000 1849.960 2741.000 1924.040 ;
        RECT 4.400 1848.560 2741.000 1849.960 ;
        RECT 4.000 1792.840 2741.000 1848.560 ;
        RECT 4.000 1791.440 2740.600 1792.840 ;
        RECT 4.000 1754.760 2741.000 1791.440 ;
        RECT 4.400 1753.360 2741.000 1754.760 ;
        RECT 4.000 1660.240 2741.000 1753.360 ;
        RECT 4.400 1658.840 2740.600 1660.240 ;
        RECT 4.000 1565.040 2741.000 1658.840 ;
        RECT 4.400 1563.640 2741.000 1565.040 ;
        RECT 4.000 1527.640 2741.000 1563.640 ;
        RECT 4.000 1526.240 2740.600 1527.640 ;
        RECT 4.000 1470.520 2741.000 1526.240 ;
        RECT 4.400 1469.120 2741.000 1470.520 ;
        RECT 4.000 1394.360 2741.000 1469.120 ;
        RECT 4.000 1392.960 2740.600 1394.360 ;
        RECT 4.000 1375.320 2741.000 1392.960 ;
        RECT 4.400 1373.920 2741.000 1375.320 ;
        RECT 4.000 1280.800 2741.000 1373.920 ;
        RECT 4.400 1279.400 2741.000 1280.800 ;
        RECT 4.000 1261.760 2741.000 1279.400 ;
        RECT 4.000 1260.360 2740.600 1261.760 ;
        RECT 4.000 1185.600 2741.000 1260.360 ;
        RECT 4.400 1184.200 2741.000 1185.600 ;
        RECT 4.000 1129.160 2741.000 1184.200 ;
        RECT 4.000 1127.760 2740.600 1129.160 ;
        RECT 4.000 1091.080 2741.000 1127.760 ;
        RECT 4.400 1089.680 2741.000 1091.080 ;
        RECT 4.000 995.880 2741.000 1089.680 ;
        RECT 4.400 994.480 2740.600 995.880 ;
        RECT 4.000 901.360 2741.000 994.480 ;
        RECT 4.400 899.960 2741.000 901.360 ;
        RECT 4.000 863.280 2741.000 899.960 ;
        RECT 4.000 861.880 2740.600 863.280 ;
        RECT 4.000 806.160 2741.000 861.880 ;
        RECT 4.400 804.760 2741.000 806.160 ;
        RECT 4.000 730.680 2741.000 804.760 ;
        RECT 4.000 729.280 2740.600 730.680 ;
        RECT 4.000 711.640 2741.000 729.280 ;
        RECT 4.400 710.240 2741.000 711.640 ;
        RECT 4.000 616.440 2741.000 710.240 ;
        RECT 4.400 615.040 2741.000 616.440 ;
        RECT 4.000 598.080 2741.000 615.040 ;
        RECT 4.000 596.680 2740.600 598.080 ;
        RECT 4.000 521.920 2741.000 596.680 ;
        RECT 4.400 520.520 2741.000 521.920 ;
        RECT 4.000 464.800 2741.000 520.520 ;
        RECT 4.000 463.400 2740.600 464.800 ;
        RECT 4.000 426.720 2741.000 463.400 ;
        RECT 4.400 425.320 2741.000 426.720 ;
        RECT 4.000 332.200 2741.000 425.320 ;
        RECT 4.400 330.800 2740.600 332.200 ;
        RECT 4.000 237.000 2741.000 330.800 ;
        RECT 4.400 235.600 2741.000 237.000 ;
        RECT 4.000 199.600 2741.000 235.600 ;
        RECT 4.000 198.200 2740.600 199.600 ;
        RECT 4.000 142.480 2741.000 198.200 ;
        RECT 4.400 141.080 2741.000 142.480 ;
        RECT 4.000 67.000 2741.000 141.080 ;
        RECT 4.000 65.600 2740.600 67.000 ;
        RECT 4.000 47.960 2741.000 65.600 ;
        RECT 4.400 46.560 2741.000 47.960 ;
        RECT 4.000 10.715 2741.000 46.560 ;
      LAYER met4 ;
        RECT 18.905 10.640 2706.705 3307.760 ;
      LAYER met5 ;
        RECT 5.520 92.700 2739.300 3283.165 ;
  END
END fpga
END LIBRARY


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2858.050 75.720 2858.370 75.780 ;
        RECT 2900.830 75.720 2901.150 75.780 ;
        RECT 2858.050 75.580 2901.150 75.720 ;
        RECT 2858.050 75.520 2858.370 75.580 ;
        RECT 2900.830 75.520 2901.150 75.580 ;
      LAYER via ;
        RECT 2858.080 75.520 2858.340 75.780 ;
        RECT 2900.860 75.520 2901.120 75.780 ;
      LAYER met2 ;
        RECT 2900.850 87.875 2901.130 88.245 ;
        RECT 2900.920 75.810 2901.060 87.875 ;
        RECT 2858.080 75.490 2858.340 75.810 ;
        RECT 2900.860 75.490 2901.120 75.810 ;
        RECT 2858.140 73.285 2858.280 75.490 ;
        RECT 2858.070 72.915 2858.350 73.285 ;
      LAYER via2 ;
        RECT 2900.850 87.920 2901.130 88.200 ;
        RECT 2858.070 72.960 2858.350 73.240 ;
      LAYER met3 ;
        RECT 2900.825 88.210 2901.155 88.225 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2900.825 87.910 2924.800 88.210 ;
        RECT 2900.825 87.895 2901.155 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
        RECT 2851.000 73.250 2855.000 73.640 ;
        RECT 2858.045 73.250 2858.375 73.265 ;
        RECT 2851.000 73.040 2858.375 73.250 ;
        RECT 2854.300 72.950 2858.375 73.040 ;
        RECT 2858.045 72.935 2858.375 72.950 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2849.845 3270.205 2850.015 3296.215 ;
        RECT 2849.845 2644.265 2850.015 2654.975 ;
        RECT 2850.305 2605.165 2850.475 2612.475 ;
        RECT 2850.305 2515.745 2850.475 2521.015 ;
      LAYER mcon ;
        RECT 2849.845 3296.045 2850.015 3296.215 ;
        RECT 2849.845 2654.805 2850.015 2654.975 ;
        RECT 2850.305 2612.305 2850.475 2612.475 ;
        RECT 2850.305 2520.845 2850.475 2521.015 ;
      LAYER met1 ;
        RECT 938.010 3415.880 938.330 3415.940 ;
        RECT 2849.310 3415.880 2849.630 3415.940 ;
        RECT 938.010 3415.740 2849.630 3415.880 ;
        RECT 938.010 3415.680 938.330 3415.740 ;
        RECT 2849.310 3415.680 2849.630 3415.740 ;
        RECT 2849.770 3296.200 2850.090 3296.260 ;
        RECT 2849.575 3296.060 2850.090 3296.200 ;
        RECT 2849.770 3296.000 2850.090 3296.060 ;
        RECT 2849.770 3270.360 2850.090 3270.420 ;
        RECT 2849.575 3270.220 2850.090 3270.360 ;
        RECT 2849.770 3270.160 2850.090 3270.220 ;
        RECT 2849.770 3046.300 2850.090 3046.360 ;
        RECT 2850.230 3046.300 2850.550 3046.360 ;
        RECT 2849.770 3046.160 2850.550 3046.300 ;
        RECT 2849.770 3046.100 2850.090 3046.160 ;
        RECT 2850.230 3046.100 2850.550 3046.160 ;
        RECT 2849.770 2654.960 2850.090 2655.020 ;
        RECT 2849.575 2654.820 2850.090 2654.960 ;
        RECT 2849.770 2654.760 2850.090 2654.820 ;
        RECT 2849.770 2644.420 2850.090 2644.480 ;
        RECT 2849.575 2644.280 2850.090 2644.420 ;
        RECT 2849.770 2644.220 2850.090 2644.280 ;
        RECT 2849.770 2612.460 2850.090 2612.520 ;
        RECT 2850.245 2612.460 2850.535 2612.505 ;
        RECT 2849.770 2612.320 2850.535 2612.460 ;
        RECT 2849.770 2612.260 2850.090 2612.320 ;
        RECT 2850.245 2612.275 2850.535 2612.320 ;
        RECT 2849.770 2605.320 2850.090 2605.380 ;
        RECT 2850.245 2605.320 2850.535 2605.365 ;
        RECT 2849.770 2605.180 2850.535 2605.320 ;
        RECT 2849.770 2605.120 2850.090 2605.180 ;
        RECT 2850.245 2605.135 2850.535 2605.180 ;
        RECT 2849.770 2521.000 2850.090 2521.060 ;
        RECT 2850.245 2521.000 2850.535 2521.045 ;
        RECT 2849.770 2520.860 2850.535 2521.000 ;
        RECT 2849.770 2520.800 2850.090 2520.860 ;
        RECT 2850.245 2520.815 2850.535 2520.860 ;
        RECT 2849.770 2515.900 2850.090 2515.960 ;
        RECT 2850.245 2515.900 2850.535 2515.945 ;
        RECT 2849.770 2515.760 2850.535 2515.900 ;
        RECT 2849.770 2515.700 2850.090 2515.760 ;
        RECT 2850.245 2515.715 2850.535 2515.760 ;
        RECT 2849.770 2435.660 2850.090 2435.720 ;
        RECT 2898.990 2435.660 2899.310 2435.720 ;
        RECT 2849.770 2435.520 2899.310 2435.660 ;
        RECT 2849.770 2435.460 2850.090 2435.520 ;
        RECT 2898.990 2435.460 2899.310 2435.520 ;
      LAYER via ;
        RECT 938.040 3415.680 938.300 3415.940 ;
        RECT 2849.340 3415.680 2849.600 3415.940 ;
        RECT 2849.800 3296.000 2850.060 3296.260 ;
        RECT 2849.800 3270.160 2850.060 3270.420 ;
        RECT 2849.800 3046.100 2850.060 3046.360 ;
        RECT 2850.260 3046.100 2850.520 3046.360 ;
        RECT 2849.800 2654.760 2850.060 2655.020 ;
        RECT 2849.800 2644.220 2850.060 2644.480 ;
        RECT 2849.800 2612.260 2850.060 2612.520 ;
        RECT 2849.800 2605.120 2850.060 2605.380 ;
        RECT 2849.800 2520.800 2850.060 2521.060 ;
        RECT 2849.800 2515.700 2850.060 2515.960 ;
        RECT 2849.800 2435.460 2850.060 2435.720 ;
        RECT 2899.020 2435.460 2899.280 2435.720 ;
      LAYER met2 ;
        RECT 938.040 3415.650 938.300 3415.970 ;
        RECT 2849.340 3415.650 2849.600 3415.970 ;
        RECT 938.100 3405.000 938.240 3415.650 ;
        RECT 937.970 3401.000 938.250 3405.000 ;
        RECT 2849.400 3374.060 2849.540 3415.650 ;
        RECT 2848.940 3373.920 2849.540 3374.060 ;
        RECT 2848.940 3318.810 2849.080 3373.920 ;
        RECT 2848.940 3318.670 2849.540 3318.810 ;
        RECT 2849.400 3296.370 2849.540 3318.670 ;
        RECT 2849.400 3296.290 2850.000 3296.370 ;
        RECT 2849.400 3296.230 2850.060 3296.290 ;
        RECT 2849.800 3295.970 2850.060 3296.230 ;
        RECT 2849.800 3270.130 2850.060 3270.450 ;
        RECT 2849.860 3269.850 2850.000 3270.130 ;
        RECT 2848.480 3269.710 2850.000 3269.850 ;
        RECT 2848.480 3235.850 2848.620 3269.710 ;
        RECT 2848.020 3235.710 2848.620 3235.850 ;
        RECT 2848.020 3152.210 2848.160 3235.710 ;
        RECT 2848.020 3152.070 2850.460 3152.210 ;
        RECT 2850.320 3126.370 2850.460 3152.070 ;
        RECT 2848.940 3126.230 2850.460 3126.370 ;
        RECT 2848.940 3065.170 2849.080 3126.230 ;
        RECT 2848.940 3065.030 2850.460 3065.170 ;
        RECT 2850.320 3046.390 2850.460 3065.030 ;
        RECT 2849.800 3046.130 2850.060 3046.390 ;
        RECT 2848.940 3046.070 2850.060 3046.130 ;
        RECT 2850.260 3046.070 2850.520 3046.390 ;
        RECT 2848.940 3045.990 2850.000 3046.070 ;
        RECT 2848.940 3022.330 2849.080 3045.990 ;
        RECT 2848.940 3022.190 2849.540 3022.330 ;
        RECT 2849.400 2940.050 2849.540 3022.190 ;
        RECT 2848.480 2939.910 2849.540 2940.050 ;
        RECT 2848.480 2874.770 2848.620 2939.910 ;
        RECT 2848.480 2874.630 2850.460 2874.770 ;
        RECT 2850.320 2847.570 2850.460 2874.630 ;
        RECT 2849.400 2847.430 2850.460 2847.570 ;
        RECT 2849.400 2839.410 2849.540 2847.430 ;
        RECT 2848.940 2839.270 2849.540 2839.410 ;
        RECT 2848.940 2759.850 2849.080 2839.270 ;
        RECT 2848.940 2759.710 2850.460 2759.850 ;
        RECT 2850.320 2757.130 2850.460 2759.710 ;
        RECT 2848.940 2756.990 2850.460 2757.130 ;
        RECT 2848.940 2655.130 2849.080 2756.990 ;
        RECT 2848.940 2655.050 2850.000 2655.130 ;
        RECT 2848.940 2654.990 2850.060 2655.050 ;
        RECT 2849.800 2654.730 2850.060 2654.990 ;
        RECT 2849.800 2644.250 2850.060 2644.510 ;
        RECT 2848.940 2644.190 2850.060 2644.250 ;
        RECT 2848.940 2644.110 2850.000 2644.190 ;
        RECT 2848.940 2613.650 2849.080 2644.110 ;
        RECT 2848.480 2613.510 2849.080 2613.650 ;
        RECT 2848.480 2612.290 2848.620 2613.510 ;
        RECT 2849.800 2612.290 2850.060 2612.550 ;
        RECT 2848.480 2612.230 2850.060 2612.290 ;
        RECT 2848.480 2612.150 2850.000 2612.230 ;
        RECT 2849.800 2605.090 2850.060 2605.410 ;
        RECT 2849.860 2604.810 2850.000 2605.090 ;
        RECT 2848.940 2604.670 2850.000 2604.810 ;
        RECT 2848.940 2521.170 2849.080 2604.670 ;
        RECT 2848.940 2521.090 2850.000 2521.170 ;
        RECT 2848.940 2521.030 2850.060 2521.090 ;
        RECT 2849.800 2520.770 2850.060 2521.030 ;
        RECT 2849.800 2515.730 2850.060 2515.990 ;
        RECT 2848.940 2515.670 2850.060 2515.730 ;
        RECT 2848.940 2515.590 2850.000 2515.670 ;
        RECT 2848.940 2455.210 2849.080 2515.590 ;
        RECT 2848.940 2455.070 2850.000 2455.210 ;
        RECT 2849.860 2435.750 2850.000 2455.070 ;
        RECT 2849.800 2435.430 2850.060 2435.750 ;
        RECT 2899.020 2435.430 2899.280 2435.750 ;
        RECT 2899.080 2434.245 2899.220 2435.430 ;
        RECT 2899.010 2433.875 2899.290 2434.245 ;
      LAYER via2 ;
        RECT 2899.010 2433.920 2899.290 2434.200 ;
      LAYER met3 ;
        RECT 2898.985 2434.210 2899.315 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2898.985 2433.910 2924.800 2434.210 ;
        RECT 2898.985 2433.895 2899.315 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2389.845 3400.765 2390.935 3400.935 ;
        RECT 2597.765 3399.065 2597.935 3400.935 ;
        RECT 2645.605 3399.065 2645.775 3400.935 ;
        RECT 2849.845 2308.345 2850.015 2332.995 ;
        RECT 2850.305 2327.385 2850.475 2335.375 ;
        RECT 2851.225 2332.825 2851.395 2338.095 ;
        RECT 2851.685 2319.225 2851.855 2327.555 ;
        RECT 2850.305 1961.545 2850.475 1984.155 ;
        RECT 2851.225 1942.505 2851.395 1974.975 ;
        RECT 2851.685 1949.985 2851.855 1965.795 ;
        RECT 2849.385 1846.965 2850.015 1847.135 ;
        RECT 2849.385 1790.355 2849.555 1846.965 ;
        RECT 2850.305 1791.205 2850.475 1797.835 ;
        RECT 2849.385 1790.185 2850.475 1790.355 ;
        RECT 2851.685 1790.185 2851.855 1799.535 ;
        RECT 2850.305 1762.305 2850.475 1790.185 ;
        RECT 2851.225 1739.865 2851.395 1762.475 ;
        RECT 2852.145 1761.625 2852.315 1838.975 ;
        RECT 2852.605 1768.425 2852.775 1795.795 ;
        RECT 2849.385 1605.055 2849.555 1647.895 ;
        RECT 2851.225 1628.345 2851.395 1647.215 ;
        RECT 2851.685 1635.145 2851.855 1646.535 ;
        RECT 2849.385 1604.885 2850.475 1605.055 ;
        RECT 2849.385 1604.205 2850.015 1604.375 ;
        RECT 2849.385 1579.895 2849.555 1604.205 ;
        RECT 2851.225 1604.035 2851.395 1627.835 ;
        RECT 2850.305 1603.865 2851.395 1604.035 ;
        RECT 2849.385 1579.725 2850.015 1579.895 ;
        RECT 2850.305 1579.555 2850.475 1603.865 ;
        RECT 2849.385 1579.385 2850.475 1579.555 ;
        RECT 2849.385 1521.755 2849.555 1579.385 ;
        RECT 2849.845 1579.045 2850.475 1579.215 ;
        RECT 2849.845 1530.765 2850.015 1578.195 ;
        RECT 2850.305 1545.385 2850.475 1579.045 ;
        RECT 2849.385 1521.585 2850.935 1521.755 ;
        RECT 2849.845 1504.245 2850.015 1509.515 ;
        RECT 2849.845 1492.685 2850.015 1500.335 ;
        RECT 2850.765 1480.785 2850.935 1521.585 ;
        RECT 2851.225 1492.005 2851.395 1513.935 ;
        RECT 2852.145 1509.345 2852.315 1535.015 ;
        RECT 2850.765 1463.275 2850.935 1480.275 ;
        RECT 2849.385 1463.105 2850.935 1463.275 ;
        RECT 2849.385 1428.255 2849.555 1463.105 ;
        RECT 2852.145 1462.085 2852.315 1505.775 ;
        RECT 2849.385 1428.085 2850.015 1428.255 ;
        RECT 2849.845 1418.565 2850.015 1425.875 ;
        RECT 2850.305 1371.475 2850.475 1418.055 ;
        RECT 2850.765 1371.645 2850.935 1426.895 ;
        RECT 2851.225 1417.885 2851.395 1428.255 ;
        RECT 2851.685 1416.865 2851.855 1424.855 ;
        RECT 2852.605 1417.545 2852.775 1448.315 ;
        RECT 2850.305 1371.305 2850.935 1371.475 ;
        RECT 2849.845 1357.705 2850.015 1365.355 ;
        RECT 2850.765 1352.265 2850.935 1371.305 ;
        RECT 2851.685 1350.225 2851.855 1371.815 ;
        RECT 2852.605 1354.985 2852.775 1386.435 ;
        RECT 2853.065 1362.465 2853.235 1424.175 ;
        RECT 2853.525 1364.505 2853.695 1372.495 ;
        RECT 2849.385 1151.155 2849.555 1226.975 ;
        RECT 2850.765 1205.895 2850.935 1329.655 ;
        RECT 2851.225 1232.585 2851.395 1254.855 ;
        RECT 2852.605 1226.805 2852.775 1253.155 ;
        RECT 2850.765 1205.725 2851.395 1205.895 ;
        RECT 2849.385 1150.985 2850.015 1151.155 ;
        RECT 2851.225 1148.605 2851.395 1205.725 ;
        RECT 2849.385 1148.265 2850.015 1148.435 ;
        RECT 2849.385 1025.015 2849.555 1148.265 ;
        RECT 2852.145 1129.395 2852.315 1197.395 ;
        RECT 2851.225 1129.225 2852.315 1129.395 ;
        RECT 2849.385 1024.845 2850.475 1025.015 ;
        RECT 2850.305 1023.825 2850.475 1024.845 ;
        RECT 2850.765 1014.985 2850.935 1072.955 ;
        RECT 2851.225 1027.735 2851.395 1129.225 ;
        RECT 2851.685 1073.125 2851.855 1129.055 ;
        RECT 2851.225 1027.565 2851.855 1027.735 ;
        RECT 2851.685 1017.705 2851.855 1027.565 ;
        RECT 2851.225 890.035 2851.395 959.735 ;
        RECT 2851.225 889.865 2851.855 890.035 ;
        RECT 2849.845 818.465 2850.015 874.735 ;
        RECT 2849.385 793.645 2850.015 793.815 ;
        RECT 2851.685 793.645 2851.855 889.865 ;
        RECT 2852.145 810.985 2852.315 859.775 ;
        RECT 2849.385 790.075 2849.555 793.645 ;
        RECT 2849.385 789.905 2850.015 790.075 ;
        RECT 2850.765 738.225 2850.935 790.075 ;
        RECT 2851.685 778.515 2851.855 787.015 ;
        RECT 2851.685 778.345 2852.315 778.515 ;
        RECT 2852.145 766.955 2852.315 778.345 ;
        RECT 2852.605 774.945 2852.775 788.375 ;
        RECT 2851.225 766.785 2852.315 766.955 ;
        RECT 2851.225 739.585 2851.395 766.785 ;
        RECT 2849.845 284.665 2850.015 379.695 ;
        RECT 2851.225 379.525 2851.395 383.095 ;
        RECT 2851.685 379.355 2851.855 381.055 ;
        RECT 2851.225 379.185 2851.855 379.355 ;
        RECT 2851.225 299.625 2851.395 379.185 ;
        RECT 2851.685 362.185 2851.855 374.255 ;
        RECT 2852.145 364.905 2852.315 368.135 ;
        RECT 2851.685 303.705 2851.855 340.255 ;
        RECT 2852.605 330.565 2852.775 367.115 ;
        RECT 2849.845 198.305 2850.015 204.935 ;
        RECT 2850.305 196.945 2850.475 208.335 ;
        RECT 2850.765 199.325 2850.935 205.615 ;
        RECT 2849.845 115.345 2850.015 139.655 ;
        RECT 2851.225 139.485 2851.395 211.055 ;
        RECT 2852.145 200.005 2852.315 202.215 ;
        RECT 2853.065 173.825 2853.235 201.535 ;
        RECT 2850.305 73.525 2850.475 128.775 ;
        RECT 2851.225 118.745 2851.395 132.515 ;
        RECT 2852.145 120.785 2852.315 127.755 ;
        RECT 2850.765 88.145 2850.935 115.515 ;
        RECT 9.805 7.905 9.975 43.775 ;
        RECT 955.105 8.925 956.655 9.095 ;
        RECT 955.105 8.755 955.275 8.925 ;
        RECT 25.445 6.205 26.535 6.375 ;
        RECT 129.865 4.845 130.035 7.055 ;
        RECT 176.785 4.845 176.955 8.755 ;
        RECT 243.945 8.585 245.495 8.755 ;
        RECT 243.945 7.565 244.115 8.585 ;
        RECT 951.425 8.415 951.595 8.755 ;
        RECT 952.345 8.585 955.275 8.755 ;
        RECT 956.485 8.585 956.655 8.925 ;
        RECT 952.345 8.415 952.515 8.585 ;
        RECT 278.905 4.675 279.075 8.415 ;
        RECT 795.485 8.245 800.255 8.415 ;
        RECT 951.425 8.245 952.515 8.415 ;
        RECT 958.325 8.415 958.495 8.755 ;
        RECT 983.625 8.585 984.715 8.755 ;
        RECT 958.325 8.245 959.415 8.415 ;
        RECT 419.665 7.905 435.475 8.075 ;
        RECT 278.905 4.505 284.595 4.675 ;
        RECT 196.565 1.785 196.735 3.315 ;
        RECT 52.585 0.425 52.755 1.275 ;
        RECT 289.945 0.935 290.115 4.675 ;
        RECT 364.925 1.275 365.095 1.615 ;
        RECT 291.325 0.935 291.495 1.275 ;
        RECT 364.925 1.105 365.555 1.275 ;
        RECT 289.945 0.765 291.495 0.935 ;
        RECT 365.385 0.935 365.555 1.105 ;
        RECT 366.305 0.935 366.475 3.315 ;
        RECT 377.805 3.145 377.975 4.675 ;
        RECT 369.525 1.785 371.995 1.955 ;
        RECT 365.385 0.765 366.475 0.935 ;
        RECT 382.865 0.765 383.035 1.955 ;
        RECT 419.665 0.935 419.835 7.905 ;
        RECT 435.305 6.545 435.475 7.905 ;
        RECT 438.065 7.565 465.835 7.735 ;
        RECT 438.065 6.545 438.235 7.565 ;
        RECT 465.665 6.545 465.835 7.565 ;
        RECT 509.365 6.545 510.455 6.715 ;
        RECT 454.625 6.205 458.935 6.375 ;
        RECT 510.285 6.205 510.455 6.545 ;
        RECT 428.865 3.655 429.035 6.035 ;
        RECT 428.865 3.485 438.235 3.655 ;
        RECT 438.065 1.275 438.235 3.485 ;
        RECT 438.065 1.105 439.155 1.275 ;
        RECT 416.905 0.765 419.835 0.935 ;
        RECT 421.965 0.255 422.135 0.935 ;
        RECT 438.985 0.765 439.155 1.105 ;
        RECT 454.625 0.255 454.795 6.205 ;
        RECT 458.765 5.865 458.935 6.205 ;
        RECT 460.605 5.865 465.835 6.035 ;
        RECT 465.665 3.825 465.835 5.865 ;
        RECT 514.425 3.995 514.595 4.675 ;
        RECT 502.925 3.825 504.015 3.995 ;
        RECT 503.845 3.655 504.015 3.825 ;
        RECT 510.745 3.825 511.375 3.995 ;
        RECT 512.585 3.825 514.595 3.995 ;
        RECT 510.745 3.655 510.915 3.825 ;
        RECT 457.385 0.595 457.555 0.935 ;
        RECT 457.845 0.765 458.015 3.655 ;
        RECT 503.845 3.485 510.915 3.655 ;
        RECT 489.125 3.145 491.595 3.315 ;
        RECT 489.125 1.275 489.295 3.145 ;
        RECT 491.425 2.805 491.595 3.145 ;
        RECT 511.665 2.635 511.835 2.975 ;
        RECT 512.585 2.635 512.755 3.825 ;
        RECT 511.665 2.465 512.755 2.635 ;
        RECT 605.505 1.955 605.675 6.375 ;
        RECT 640.465 6.205 644.315 6.375 ;
        RECT 645.985 5.695 646.155 6.375 ;
        RECT 659.785 5.695 659.955 6.715 ;
        RECT 645.985 5.525 659.955 5.695 ;
        RECT 646.445 1.955 646.615 4.675 ;
        RECT 676.805 4.505 676.975 6.375 ;
        RECT 680.485 6.205 697.215 6.375 ;
        RECT 680.485 4.505 680.655 6.205 ;
        RECT 697.045 5.865 697.215 6.205 ;
        RECT 750.405 4.505 750.575 5.695 ;
        RECT 757.305 5.525 757.475 7.055 ;
        RECT 763.745 6.205 763.915 7.055 ;
        RECT 795.485 6.715 795.655 8.245 ;
        RECT 766.505 6.545 768.515 6.715 ;
        RECT 765.125 3.655 765.295 6.375 ;
        RECT 766.505 6.205 766.675 6.545 ;
        RECT 768.345 6.375 768.515 6.545 ;
        RECT 794.565 6.545 795.655 6.715 ;
        RECT 768.345 6.205 772.655 6.375 ;
        RECT 767.425 5.865 768.975 6.035 ;
        RECT 767.425 5.695 767.595 5.865 ;
        RECT 766.965 5.525 767.595 5.695 ;
        RECT 768.805 5.525 768.975 5.865 ;
        RECT 770.185 5.865 772.195 6.035 ;
        RECT 770.185 5.525 770.355 5.865 ;
        RECT 772.025 3.825 772.195 5.865 ;
        RECT 772.485 5.695 772.655 6.205 ;
        RECT 772.485 5.525 774.035 5.695 ;
        RECT 752.245 3.485 758.395 3.655 ;
        RECT 752.245 3.315 752.415 3.485 ;
        RECT 751.325 3.145 752.415 3.315 ;
        RECT 758.225 3.315 758.395 3.485 ;
        RECT 761.905 3.485 765.295 3.655 ;
        RECT 761.905 3.315 762.075 3.485 ;
        RECT 758.225 3.145 762.075 3.315 ;
        RECT 462.905 1.105 489.295 1.275 ;
        RECT 559.045 1.785 561.975 1.955 ;
        RECT 605.505 1.785 646.615 1.955 ;
        RECT 462.905 0.935 463.075 1.105 ;
        RECT 458.305 0.765 463.075 0.935 ;
        RECT 559.045 0.765 559.215 1.785 ;
        RECT 561.805 0.765 561.975 1.785 ;
        RECT 773.865 1.615 774.035 5.525 ;
        RECT 794.565 5.355 794.735 6.545 ;
        RECT 800.085 6.375 800.255 8.245 ;
        RECT 959.245 8.075 959.415 8.245 ;
        RECT 983.625 8.075 983.795 8.585 ;
        RECT 850.685 7.905 860.515 8.075 ;
        RECT 959.245 7.905 983.795 8.075 ;
        RECT 850.685 7.395 850.855 7.905 ;
        RECT 846.545 7.225 848.095 7.395 ;
        RECT 850.685 7.225 851.315 7.395 ;
        RECT 847.925 7.055 848.095 7.225 ;
        RECT 800.085 6.205 800.715 6.375 ;
        RECT 800.545 6.035 800.715 6.205 ;
        RECT 800.545 5.865 804.855 6.035 ;
        RECT 791.805 5.185 794.735 5.355 ;
        RECT 784.445 4.505 785.995 4.675 ;
        RECT 791.805 4.505 791.975 5.185 ;
        RECT 804.685 4.675 804.855 5.865 ;
        RECT 810.665 4.675 810.835 7.055 ;
        RECT 824.005 6.715 824.175 7.055 ;
        RECT 847.925 6.885 850.855 7.055 ;
        RECT 818.025 6.545 824.175 6.715 ;
        RECT 784.445 3.825 784.615 4.505 ;
        RECT 798.245 1.615 798.415 4.675 ;
        RECT 804.225 4.335 804.395 4.675 ;
        RECT 804.685 4.505 806.235 4.675 ;
        RECT 806.985 4.505 810.835 4.675 ;
        RECT 812.045 4.505 812.215 6.375 ;
        RECT 818.025 6.205 818.195 6.545 ;
        RECT 850.685 6.035 850.855 6.885 ;
        RECT 849.305 5.865 850.855 6.035 ;
        RECT 804.225 4.165 804.855 4.335 ;
        RECT 804.685 2.975 804.855 4.165 ;
        RECT 806.985 2.975 807.155 4.505 ;
        RECT 849.305 3.315 849.475 5.865 ;
        RECT 851.145 4.335 851.315 7.225 ;
        RECT 860.345 6.715 860.515 7.905 ;
        RECT 985.925 7.395 986.095 8.755 ;
        RECT 1596.805 8.245 1599.275 8.415 ;
        RECT 990.065 7.905 1004.495 8.075 ;
        RECT 1071.945 7.905 1072.575 8.075 ;
        RECT 990.065 7.395 990.235 7.905 ;
        RECT 869.085 6.885 880.295 7.055 ;
        RECT 869.085 6.715 869.255 6.885 ;
        RECT 860.345 6.545 869.255 6.715 ;
        RECT 878.745 6.545 879.835 6.715 ;
        RECT 880.125 6.375 880.295 6.885 ;
        RECT 884.265 6.375 884.435 7.055 ;
        RECT 880.125 6.205 884.435 6.375 ;
        RECT 953.725 6.885 955.735 7.055 ;
        RECT 953.725 6.205 953.895 6.885 ;
        RECT 955.565 6.545 955.735 6.885 ;
        RECT 956.945 6.545 957.115 7.395 ;
        RECT 957.865 6.035 958.035 7.395 ;
        RECT 985.925 7.225 990.235 7.395 ;
        RECT 1004.325 7.225 1004.495 7.905 ;
        RECT 960.625 6.885 977.355 7.055 ;
        RECT 960.625 6.035 960.795 6.885 ;
        RECT 957.865 5.865 960.795 6.035 ;
        RECT 849.765 4.165 851.315 4.335 ;
        RECT 852.065 4.165 869.715 4.335 ;
        RECT 849.765 3.485 849.935 4.165 ;
        RECT 852.065 3.655 852.235 4.165 ;
        RECT 850.685 3.485 852.235 3.655 ;
        RECT 869.545 3.655 869.715 4.165 ;
        RECT 869.545 3.485 883.055 3.655 ;
        RECT 886.565 3.485 888.115 3.655 ;
        RECT 850.685 3.315 850.855 3.485 ;
        RECT 849.305 3.145 850.855 3.315 ;
        RECT 887.945 3.145 888.115 3.485 ;
        RECT 918.765 3.145 919.855 3.315 ;
        RECT 804.685 2.805 807.155 2.975 ;
        RECT 919.685 2.295 919.855 3.145 ;
        RECT 977.185 2.635 977.355 6.885 ;
        RECT 1055.845 6.885 1056.935 7.055 ;
        RECT 1055.845 6.715 1056.015 6.885 ;
        RECT 1002.025 3.655 1002.195 6.715 ;
        RECT 1014.445 6.545 1056.015 6.715 ;
        RECT 1056.765 6.375 1056.935 6.885 ;
        RECT 1072.405 6.545 1072.575 7.905 ;
        RECT 1593.585 7.565 1595.135 7.735 ;
        RECT 1596.805 7.565 1596.975 8.245 ;
        RECT 1088.045 7.225 1089.135 7.395 ;
        RECT 1056.765 6.205 1063.835 6.375 ;
        RECT 996.045 3.485 1002.195 3.655 ;
        RECT 977.185 2.465 981.035 2.635 ;
        RECT 919.685 2.125 921.695 2.295 ;
        RECT 773.865 1.445 798.415 1.615 ;
        RECT 921.525 0.765 921.695 2.125 ;
        RECT 980.865 1.615 981.035 2.465 ;
        RECT 982.705 2.125 992.535 2.295 ;
        RECT 982.705 1.785 982.875 2.125 ;
        RECT 996.045 1.615 996.215 3.485 ;
        RECT 1063.665 3.145 1063.835 6.205 ;
        RECT 1088.045 6.035 1088.215 7.225 ;
        RECT 1088.965 6.885 1089.135 7.225 ;
        RECT 1091.725 7.225 1093.275 7.395 ;
        RECT 1483.645 7.225 1484.275 7.395 ;
        RECT 1091.725 6.885 1091.895 7.225 ;
        RECT 1093.105 6.545 1093.275 7.225 ;
        RECT 1140.945 6.885 1142.955 7.055 ;
        RECT 1140.945 6.545 1141.115 6.885 ;
        RECT 1072.865 5.865 1088.215 6.035 ;
        RECT 1141.405 5.865 1141.575 6.715 ;
        RECT 1142.785 6.035 1142.955 6.885 ;
        RECT 1484.105 6.205 1484.275 7.225 ;
        RECT 1489.625 6.035 1489.795 6.375 ;
        RECT 1142.785 5.865 1159.055 6.035 ;
        RECT 1489.625 5.865 1490.715 6.035 ;
        RECT 1072.865 3.315 1073.035 5.865 ;
        RECT 1127.605 4.675 1127.775 5.695 ;
        RECT 1158.885 5.525 1159.055 5.865 ;
        RECT 1236.625 5.525 1238.175 5.695 ;
        RECT 1593.585 5.355 1593.755 7.565 ;
        RECT 1125.305 4.505 1127.775 4.675 ;
        RECT 1574.265 5.185 1593.755 5.355 ;
        RECT 1107.365 3.315 1107.535 3.655 ;
        RECT 1125.305 3.485 1125.475 4.505 ;
        RECT 1193.845 3.655 1194.015 3.995 ;
        RECT 1197.985 3.825 1209.655 3.995 ;
        RECT 1197.985 3.655 1198.155 3.825 ;
        RECT 1193.845 3.485 1198.155 3.655 ;
        RECT 1573.345 3.655 1573.515 3.995 ;
        RECT 1574.265 3.655 1574.435 5.185 ;
        RECT 1728.825 4.845 1728.995 8.415 ;
        RECT 1951.925 6.545 1953.935 6.715 ;
        RECT 2777.165 6.205 2777.335 7.395 ;
        RECT 2801.085 6.545 2801.255 7.395 ;
        RECT 1780.805 4.505 1780.975 6.035 ;
        RECT 1863.605 5.525 1864.695 5.695 ;
        RECT 1953.305 5.525 1954.395 5.695 ;
        RECT 1863.605 4.845 1863.775 5.525 ;
        RECT 1864.525 5.015 1864.695 5.525 ;
        RECT 2469.425 5.355 2469.595 5.695 ;
        RECT 2608.345 5.525 2608.975 5.695 ;
        RECT 2469.425 5.185 2470.515 5.355 ;
        RECT 1864.525 4.845 1865.615 5.015 ;
        RECT 1862.225 4.165 1864.235 4.335 ;
        RECT 2691.145 4.165 2691.315 5.695 ;
        RECT 2715.525 4.165 2715.695 5.695 ;
        RECT 2746.345 5.525 2746.975 5.695 ;
        RECT 2797.405 4.505 2797.575 5.695 ;
        RECT 1862.225 3.825 1862.395 4.165 ;
        RECT 1573.345 3.485 1574.435 3.655 ;
        RECT 1070.105 3.145 1073.035 3.315 ;
        RECT 1105.065 3.145 1107.535 3.315 ;
        RECT 1120.705 2.975 1120.875 3.315 ;
        RECT 1127.145 2.975 1127.315 3.315 ;
        RECT 1120.705 2.805 1127.315 2.975 ;
        RECT 1931.685 2.295 1931.855 3.995 ;
        RECT 1932.605 2.295 1932.775 2.635 ;
        RECT 1931.685 2.125 1932.775 2.295 ;
        RECT 980.865 1.445 996.215 1.615 ;
        RECT 1676.845 0.765 1678.395 0.935 ;
        RECT 1737.565 0.765 1738.655 0.935 ;
        RECT 1861.765 0.765 1866.535 0.935 ;
        RECT 1883.845 0.765 1884.935 0.935 ;
        RECT 458.305 0.595 458.475 0.765 ;
        RECT 457.385 0.425 458.475 0.595 ;
        RECT 421.965 0.085 454.795 0.255 ;
        RECT 460.605 0.255 460.775 0.595 ;
        RECT 462.445 0.255 462.615 0.595 ;
        RECT 460.605 0.085 462.615 0.255 ;
        RECT 917.845 0.255 918.015 0.595 ;
        RECT 920.145 0.255 920.315 0.595 ;
        RECT 1677.765 0.425 1678.855 0.595 ;
        RECT 1737.105 0.425 1738.195 0.595 ;
        RECT 1862.225 0.425 1863.775 0.595 ;
        RECT 2153.865 0.425 2154.035 3.995 ;
        RECT 2180.545 0.425 2180.715 3.995 ;
        RECT 2367.305 0.765 2368.395 0.935 ;
        RECT 917.845 0.085 920.315 0.255 ;
        RECT 1677.305 0.085 1678.395 0.255 ;
        RECT 1736.645 0.085 1738.655 0.255 ;
        RECT 2841.565 0.085 2841.735 8.755 ;
      LAYER mcon ;
        RECT 2390.765 3400.765 2390.935 3400.935 ;
        RECT 2597.765 3400.765 2597.935 3400.935 ;
        RECT 2645.605 3400.765 2645.775 3400.935 ;
        RECT 2851.225 2337.925 2851.395 2338.095 ;
        RECT 2850.305 2335.205 2850.475 2335.375 ;
        RECT 2849.845 2332.825 2850.015 2332.995 ;
        RECT 2851.685 2327.385 2851.855 2327.555 ;
        RECT 2850.305 1983.985 2850.475 1984.155 ;
        RECT 2851.225 1974.805 2851.395 1974.975 ;
        RECT 2851.685 1965.625 2851.855 1965.795 ;
        RECT 2849.845 1846.965 2850.015 1847.135 ;
        RECT 2852.145 1838.805 2852.315 1838.975 ;
        RECT 2851.685 1799.365 2851.855 1799.535 ;
        RECT 2850.305 1797.665 2850.475 1797.835 ;
        RECT 2851.225 1762.305 2851.395 1762.475 ;
        RECT 2852.605 1795.625 2852.775 1795.795 ;
        RECT 2849.385 1647.725 2849.555 1647.895 ;
        RECT 2851.225 1647.045 2851.395 1647.215 ;
        RECT 2851.685 1646.365 2851.855 1646.535 ;
        RECT 2851.225 1627.665 2851.395 1627.835 ;
        RECT 2850.305 1604.885 2850.475 1605.055 ;
        RECT 2849.845 1604.205 2850.015 1604.375 ;
        RECT 2849.845 1579.725 2850.015 1579.895 ;
        RECT 2849.845 1578.025 2850.015 1578.195 ;
        RECT 2852.145 1534.845 2852.315 1535.015 ;
        RECT 2849.845 1509.345 2850.015 1509.515 ;
        RECT 2849.845 1500.165 2850.015 1500.335 ;
        RECT 2851.225 1513.765 2851.395 1513.935 ;
        RECT 2852.145 1505.605 2852.315 1505.775 ;
        RECT 2850.765 1480.105 2850.935 1480.275 ;
        RECT 2852.605 1448.145 2852.775 1448.315 ;
        RECT 2849.845 1428.085 2850.015 1428.255 ;
        RECT 2851.225 1428.085 2851.395 1428.255 ;
        RECT 2850.765 1426.725 2850.935 1426.895 ;
        RECT 2849.845 1425.705 2850.015 1425.875 ;
        RECT 2850.305 1417.885 2850.475 1418.055 ;
        RECT 2851.685 1424.685 2851.855 1424.855 ;
        RECT 2853.065 1424.005 2853.235 1424.175 ;
        RECT 2852.605 1386.265 2852.775 1386.435 ;
        RECT 2851.685 1371.645 2851.855 1371.815 ;
        RECT 2849.845 1365.185 2850.015 1365.355 ;
        RECT 2853.525 1372.325 2853.695 1372.495 ;
        RECT 2850.765 1329.485 2850.935 1329.655 ;
        RECT 2849.385 1226.805 2849.555 1226.975 ;
        RECT 2851.225 1254.685 2851.395 1254.855 ;
        RECT 2852.605 1252.985 2852.775 1253.155 ;
        RECT 2849.845 1150.985 2850.015 1151.155 ;
        RECT 2852.145 1197.225 2852.315 1197.395 ;
        RECT 2849.845 1148.265 2850.015 1148.435 ;
        RECT 2850.765 1072.785 2850.935 1072.955 ;
        RECT 2851.685 1128.885 2851.855 1129.055 ;
        RECT 2851.225 959.565 2851.395 959.735 ;
        RECT 2849.845 874.565 2850.015 874.735 ;
        RECT 2852.145 859.605 2852.315 859.775 ;
        RECT 2849.845 793.645 2850.015 793.815 ;
        RECT 2849.845 789.905 2850.015 790.075 ;
        RECT 2850.765 789.905 2850.935 790.075 ;
        RECT 2852.605 788.205 2852.775 788.375 ;
        RECT 2851.685 786.845 2851.855 787.015 ;
        RECT 2851.225 382.925 2851.395 383.095 ;
        RECT 2849.845 379.525 2850.015 379.695 ;
        RECT 2851.685 380.885 2851.855 381.055 ;
        RECT 2851.685 374.085 2851.855 374.255 ;
        RECT 2852.145 367.965 2852.315 368.135 ;
        RECT 2852.605 366.945 2852.775 367.115 ;
        RECT 2851.685 340.085 2851.855 340.255 ;
        RECT 2851.225 210.885 2851.395 211.055 ;
        RECT 2850.305 208.165 2850.475 208.335 ;
        RECT 2849.845 204.765 2850.015 204.935 ;
        RECT 2850.765 205.445 2850.935 205.615 ;
        RECT 2852.145 202.045 2852.315 202.215 ;
        RECT 2853.065 201.365 2853.235 201.535 ;
        RECT 2849.845 139.485 2850.015 139.655 ;
        RECT 2851.225 132.345 2851.395 132.515 ;
        RECT 2850.305 128.605 2850.475 128.775 ;
        RECT 2852.145 127.585 2852.315 127.755 ;
        RECT 2850.765 115.345 2850.935 115.515 ;
        RECT 9.805 43.605 9.975 43.775 ;
        RECT 176.785 8.585 176.955 8.755 ;
        RECT 129.865 6.885 130.035 7.055 ;
        RECT 26.365 6.205 26.535 6.375 ;
        RECT 245.325 8.585 245.495 8.755 ;
        RECT 951.425 8.585 951.595 8.755 ;
        RECT 958.325 8.585 958.495 8.755 ;
        RECT 278.905 8.245 279.075 8.415 ;
        RECT 984.545 8.585 984.715 8.755 ;
        RECT 985.925 8.585 986.095 8.755 ;
        RECT 284.425 4.505 284.595 4.675 ;
        RECT 289.945 4.505 290.115 4.675 ;
        RECT 196.565 3.145 196.735 3.315 ;
        RECT 52.585 1.105 52.755 1.275 ;
        RECT 377.805 4.505 377.975 4.675 ;
        RECT 366.305 3.145 366.475 3.315 ;
        RECT 364.925 1.445 365.095 1.615 ;
        RECT 291.325 1.105 291.495 1.275 ;
        RECT 371.825 1.785 371.995 1.955 ;
        RECT 382.865 1.785 383.035 1.955 ;
        RECT 757.305 6.885 757.475 7.055 ;
        RECT 659.785 6.545 659.955 6.715 ;
        RECT 605.505 6.205 605.675 6.375 ;
        RECT 644.145 6.205 644.315 6.375 ;
        RECT 645.985 6.205 646.155 6.375 ;
        RECT 428.865 5.865 429.035 6.035 ;
        RECT 421.965 0.765 422.135 0.935 ;
        RECT 514.425 4.505 514.595 4.675 ;
        RECT 511.205 3.825 511.375 3.995 ;
        RECT 457.845 3.485 458.015 3.655 ;
        RECT 511.665 2.805 511.835 2.975 ;
        RECT 676.805 6.205 676.975 6.375 ;
        RECT 646.445 4.505 646.615 4.675 ;
        RECT 763.745 6.885 763.915 7.055 ;
        RECT 765.125 6.205 765.295 6.375 ;
        RECT 750.405 5.525 750.575 5.695 ;
        RECT 457.385 0.765 457.555 0.935 ;
        RECT 810.665 6.885 810.835 7.055 ;
        RECT 824.005 6.885 824.175 7.055 ;
        RECT 785.825 4.505 785.995 4.675 ;
        RECT 798.245 4.505 798.415 4.675 ;
        RECT 804.225 4.505 804.395 4.675 ;
        RECT 806.065 4.505 806.235 4.675 ;
        RECT 812.045 6.205 812.215 6.375 ;
        RECT 2841.565 8.585 2841.735 8.755 ;
        RECT 1599.105 8.245 1599.275 8.415 ;
        RECT 1728.825 8.245 1728.995 8.415 ;
        RECT 956.945 7.225 957.115 7.395 ;
        RECT 879.665 6.545 879.835 6.715 ;
        RECT 884.265 6.885 884.435 7.055 ;
        RECT 957.865 7.225 958.035 7.395 ;
        RECT 882.885 3.485 883.055 3.655 ;
        RECT 1002.025 6.545 1002.195 6.715 ;
        RECT 1594.965 7.565 1595.135 7.735 ;
        RECT 992.365 2.125 992.535 2.295 ;
        RECT 1141.405 6.545 1141.575 6.715 ;
        RECT 1489.625 6.205 1489.795 6.375 ;
        RECT 1490.545 5.865 1490.715 6.035 ;
        RECT 1127.605 5.525 1127.775 5.695 ;
        RECT 1238.005 5.525 1238.175 5.695 ;
        RECT 1107.365 3.485 1107.535 3.655 ;
        RECT 1193.845 3.825 1194.015 3.995 ;
        RECT 1209.485 3.825 1209.655 3.995 ;
        RECT 1573.345 3.825 1573.515 3.995 ;
        RECT 2777.165 7.225 2777.335 7.395 ;
        RECT 1953.765 6.545 1953.935 6.715 ;
        RECT 2801.085 7.225 2801.255 7.395 ;
        RECT 1780.805 5.865 1780.975 6.035 ;
        RECT 1954.225 5.525 1954.395 5.695 ;
        RECT 2469.425 5.525 2469.595 5.695 ;
        RECT 2608.805 5.525 2608.975 5.695 ;
        RECT 2691.145 5.525 2691.315 5.695 ;
        RECT 2470.345 5.185 2470.515 5.355 ;
        RECT 1865.445 4.845 1865.615 5.015 ;
        RECT 1864.065 4.165 1864.235 4.335 ;
        RECT 2715.525 5.525 2715.695 5.695 ;
        RECT 2746.805 5.525 2746.975 5.695 ;
        RECT 2797.405 5.525 2797.575 5.695 ;
        RECT 1931.685 3.825 1931.855 3.995 ;
        RECT 1120.705 3.145 1120.875 3.315 ;
        RECT 1127.145 3.145 1127.315 3.315 ;
        RECT 2153.865 3.825 2154.035 3.995 ;
        RECT 1932.605 2.465 1932.775 2.635 ;
        RECT 1678.225 0.765 1678.395 0.935 ;
        RECT 1738.485 0.765 1738.655 0.935 ;
        RECT 1866.365 0.765 1866.535 0.935 ;
        RECT 1884.765 0.765 1884.935 0.935 ;
        RECT 460.605 0.425 460.775 0.595 ;
        RECT 462.445 0.425 462.615 0.595 ;
        RECT 917.845 0.425 918.015 0.595 ;
        RECT 920.145 0.425 920.315 0.595 ;
        RECT 1678.685 0.425 1678.855 0.595 ;
        RECT 1738.025 0.425 1738.195 0.595 ;
        RECT 1863.605 0.425 1863.775 0.595 ;
        RECT 2180.545 3.825 2180.715 3.995 ;
        RECT 2368.225 0.765 2368.395 0.935 ;
        RECT 1678.225 0.085 1678.395 0.255 ;
        RECT 1738.485 0.085 1738.655 0.255 ;
      LAYER met1 ;
        RECT 2019.470 3416.220 2019.790 3416.280 ;
        RECT 2042.010 3416.220 2042.330 3416.280 ;
        RECT 2019.470 3416.080 2042.330 3416.220 ;
        RECT 2019.470 3416.020 2019.790 3416.080 ;
        RECT 2042.010 3416.020 2042.330 3416.080 ;
        RECT 1529.570 3405.000 1529.890 3405.060 ;
        RECT 1638.130 3405.000 1638.450 3405.060 ;
        RECT 1529.570 3404.860 1638.450 3405.000 ;
        RECT 1529.570 3404.800 1529.890 3404.860 ;
        RECT 1638.130 3404.800 1638.450 3404.860 ;
        RECT 1638.130 3401.400 1638.450 3401.660 ;
        RECT 2042.010 3401.400 2042.330 3401.660 ;
        RECT 2773.870 3401.400 2774.190 3401.660 ;
        RECT 1638.220 3401.260 1638.360 3401.400 ;
        RECT 2042.100 3401.260 2042.240 3401.400 ;
        RECT 1638.220 3401.120 1652.620 3401.260 ;
        RECT 2042.100 3401.120 2042.700 3401.260 ;
        RECT 1652.480 3398.200 1652.620 3401.120 ;
        RECT 2042.560 3400.920 2042.700 3401.120 ;
        RECT 2389.785 3400.920 2390.075 3400.965 ;
        RECT 2042.560 3400.780 2390.075 3400.920 ;
        RECT 2389.785 3400.735 2390.075 3400.780 ;
        RECT 2390.705 3400.920 2390.995 3400.965 ;
        RECT 2597.705 3400.920 2597.995 3400.965 ;
        RECT 2390.705 3400.780 2597.995 3400.920 ;
        RECT 2390.705 3400.735 2390.995 3400.780 ;
        RECT 2597.705 3400.735 2597.995 3400.780 ;
        RECT 2645.545 3400.920 2645.835 3400.965 ;
        RECT 2773.960 3400.920 2774.100 3401.400 ;
        RECT 2645.545 3400.780 2774.100 3400.920 ;
        RECT 2645.545 3400.735 2645.835 3400.780 ;
        RECT 2597.705 3399.220 2597.995 3399.265 ;
        RECT 2645.545 3399.220 2645.835 3399.265 ;
        RECT 2597.705 3399.080 2645.835 3399.220 ;
        RECT 2597.705 3399.035 2597.995 3399.080 ;
        RECT 2645.545 3399.035 2645.835 3399.080 ;
        RECT 2841.950 3398.200 2842.270 3398.260 ;
        RECT 1652.480 3398.060 2842.270 3398.200 ;
        RECT 2841.950 3398.000 2842.270 3398.060 ;
        RECT 2849.770 3151.020 2850.090 3151.080 ;
        RECT 2863.570 3151.020 2863.890 3151.080 ;
        RECT 2849.770 3150.880 2863.890 3151.020 ;
        RECT 2849.770 3150.820 2850.090 3150.880 ;
        RECT 2863.570 3150.820 2863.890 3150.880 ;
        RECT 2849.770 3048.340 2850.090 3048.400 ;
        RECT 2851.610 3048.340 2851.930 3048.400 ;
        RECT 2849.770 3048.200 2851.930 3048.340 ;
        RECT 2849.770 3048.140 2850.090 3048.200 ;
        RECT 2851.610 3048.140 2851.930 3048.200 ;
        RECT 2849.770 2856.920 2850.090 2856.980 ;
        RECT 2863.570 2856.920 2863.890 2856.980 ;
        RECT 2849.770 2856.780 2863.890 2856.920 ;
        RECT 2849.770 2856.720 2850.090 2856.780 ;
        RECT 2863.570 2856.720 2863.890 2856.780 ;
        RECT 2866.790 2663.800 2867.110 2663.860 ;
        RECT 2900.830 2663.800 2901.150 2663.860 ;
        RECT 2866.790 2663.660 2901.150 2663.800 ;
        RECT 2866.790 2663.600 2867.110 2663.660 ;
        RECT 2900.830 2663.600 2901.150 2663.660 ;
        RECT 2849.770 2611.780 2850.090 2611.840 ;
        RECT 2866.790 2611.780 2867.110 2611.840 ;
        RECT 2849.770 2611.640 2867.110 2611.780 ;
        RECT 2849.770 2611.580 2850.090 2611.640 ;
        RECT 2866.790 2611.580 2867.110 2611.640 ;
        RECT 2849.770 2338.080 2850.090 2338.140 ;
        RECT 2851.165 2338.080 2851.455 2338.125 ;
        RECT 2849.770 2337.940 2851.455 2338.080 ;
        RECT 2849.770 2337.880 2850.090 2337.940 ;
        RECT 2851.165 2337.895 2851.455 2337.940 ;
        RECT 2850.230 2335.360 2850.550 2335.420 ;
        RECT 2850.035 2335.220 2850.550 2335.360 ;
        RECT 2850.230 2335.160 2850.550 2335.220 ;
        RECT 2849.785 2332.980 2850.075 2333.025 ;
        RECT 2851.165 2332.980 2851.455 2333.025 ;
        RECT 2849.785 2332.840 2851.455 2332.980 ;
        RECT 2849.785 2332.795 2850.075 2332.840 ;
        RECT 2851.165 2332.795 2851.455 2332.840 ;
        RECT 2850.245 2327.540 2850.535 2327.585 ;
        RECT 2851.625 2327.540 2851.915 2327.585 ;
        RECT 2850.245 2327.400 2851.915 2327.540 ;
        RECT 2850.245 2327.355 2850.535 2327.400 ;
        RECT 2851.625 2327.355 2851.915 2327.400 ;
        RECT 2849.310 2321.220 2849.630 2321.480 ;
        RECT 2849.400 2320.740 2849.540 2321.220 ;
        RECT 2850.230 2320.740 2850.550 2320.800 ;
        RECT 2849.400 2320.600 2850.550 2320.740 ;
        RECT 2850.230 2320.540 2850.550 2320.600 ;
        RECT 2849.770 2320.060 2850.090 2320.120 ;
        RECT 2849.400 2319.920 2850.090 2320.060 ;
        RECT 2849.400 2318.700 2849.540 2319.920 ;
        RECT 2849.770 2319.860 2850.090 2319.920 ;
        RECT 2849.770 2319.380 2850.090 2319.440 ;
        RECT 2851.625 2319.380 2851.915 2319.425 ;
        RECT 2849.770 2319.240 2851.915 2319.380 ;
        RECT 2849.770 2319.180 2850.090 2319.240 ;
        RECT 2851.625 2319.195 2851.915 2319.240 ;
        RECT 2849.770 2318.700 2850.090 2318.760 ;
        RECT 2849.400 2318.560 2850.090 2318.700 ;
        RECT 2849.770 2318.500 2850.090 2318.560 ;
        RECT 2849.770 2308.500 2850.090 2308.560 ;
        RECT 2849.575 2308.360 2850.090 2308.500 ;
        RECT 2849.770 2308.300 2850.090 2308.360 ;
        RECT 2852.990 2059.960 2853.310 2060.020 ;
        RECT 2863.570 2059.960 2863.890 2060.020 ;
        RECT 2852.990 2059.820 2863.890 2059.960 ;
        RECT 2852.990 2059.760 2853.310 2059.820 ;
        RECT 2863.570 2059.760 2863.890 2059.820 ;
        RECT 2849.770 2008.280 2850.090 2008.340 ;
        RECT 2852.990 2008.280 2853.310 2008.340 ;
        RECT 2849.770 2008.140 2853.310 2008.280 ;
        RECT 2849.770 2008.080 2850.090 2008.140 ;
        RECT 2852.990 2008.080 2853.310 2008.140 ;
        RECT 2849.770 1984.140 2850.090 1984.200 ;
        RECT 2850.245 1984.140 2850.535 1984.185 ;
        RECT 2849.770 1984.000 2850.535 1984.140 ;
        RECT 2849.770 1983.940 2850.090 1984.000 ;
        RECT 2850.245 1983.955 2850.535 1984.000 ;
        RECT 2849.770 1974.960 2850.090 1975.020 ;
        RECT 2851.165 1974.960 2851.455 1975.005 ;
        RECT 2849.770 1974.820 2851.455 1974.960 ;
        RECT 2849.770 1974.760 2850.090 1974.820 ;
        RECT 2851.165 1974.775 2851.455 1974.820 ;
        RECT 2849.770 1965.780 2850.090 1965.840 ;
        RECT 2851.625 1965.780 2851.915 1965.825 ;
        RECT 2849.770 1965.640 2851.915 1965.780 ;
        RECT 2849.770 1965.580 2850.090 1965.640 ;
        RECT 2851.625 1965.595 2851.915 1965.640 ;
        RECT 2849.770 1964.560 2850.090 1964.820 ;
        RECT 2849.860 1963.800 2850.000 1964.560 ;
        RECT 2849.770 1963.540 2850.090 1963.800 ;
        RECT 2849.770 1963.060 2850.090 1963.120 ;
        RECT 2851.610 1963.060 2851.930 1963.120 ;
        RECT 2849.770 1962.920 2851.930 1963.060 ;
        RECT 2849.770 1962.860 2850.090 1962.920 ;
        RECT 2851.610 1962.860 2851.930 1962.920 ;
        RECT 2849.770 1961.700 2850.090 1961.760 ;
        RECT 2850.245 1961.700 2850.535 1961.745 ;
        RECT 2849.770 1961.560 2850.535 1961.700 ;
        RECT 2849.770 1961.500 2850.090 1961.560 ;
        RECT 2850.245 1961.515 2850.535 1961.560 ;
        RECT 2849.770 1950.140 2850.090 1950.200 ;
        RECT 2851.625 1950.140 2851.915 1950.185 ;
        RECT 2849.770 1950.000 2851.915 1950.140 ;
        RECT 2849.770 1949.940 2850.090 1950.000 ;
        RECT 2851.625 1949.955 2851.915 1950.000 ;
        RECT 2849.770 1942.660 2850.090 1942.720 ;
        RECT 2851.165 1942.660 2851.455 1942.705 ;
        RECT 2849.770 1942.520 2851.455 1942.660 ;
        RECT 2849.770 1942.460 2850.090 1942.520 ;
        RECT 2851.165 1942.475 2851.455 1942.520 ;
        RECT 2849.770 1847.120 2850.090 1847.180 ;
        RECT 2849.575 1846.980 2850.090 1847.120 ;
        RECT 2849.770 1846.920 2850.090 1846.980 ;
        RECT 2849.770 1838.960 2850.090 1839.020 ;
        RECT 2852.085 1838.960 2852.375 1839.005 ;
        RECT 2849.770 1838.820 2852.375 1838.960 ;
        RECT 2849.770 1838.760 2850.090 1838.820 ;
        RECT 2852.085 1838.775 2852.375 1838.820 ;
        RECT 2849.770 1800.200 2850.090 1800.260 ;
        RECT 2851.610 1800.200 2851.930 1800.260 ;
        RECT 2849.770 1800.060 2851.930 1800.200 ;
        RECT 2849.770 1800.000 2850.090 1800.060 ;
        RECT 2851.610 1800.000 2851.930 1800.060 ;
        RECT 2849.770 1799.520 2850.090 1799.580 ;
        RECT 2851.625 1799.520 2851.915 1799.565 ;
        RECT 2849.770 1799.380 2851.915 1799.520 ;
        RECT 2849.770 1799.320 2850.090 1799.380 ;
        RECT 2851.625 1799.335 2851.915 1799.380 ;
        RECT 2849.770 1797.820 2850.090 1797.880 ;
        RECT 2850.245 1797.820 2850.535 1797.865 ;
        RECT 2849.770 1797.680 2850.535 1797.820 ;
        RECT 2849.770 1797.620 2850.090 1797.680 ;
        RECT 2850.245 1797.635 2850.535 1797.680 ;
        RECT 2849.770 1795.780 2850.090 1795.840 ;
        RECT 2852.545 1795.780 2852.835 1795.825 ;
        RECT 2849.770 1795.640 2852.835 1795.780 ;
        RECT 2849.770 1795.580 2850.090 1795.640 ;
        RECT 2852.545 1795.595 2852.835 1795.640 ;
        RECT 2849.770 1794.420 2850.090 1794.480 ;
        RECT 2849.400 1794.280 2850.090 1794.420 ;
        RECT 2849.400 1793.060 2849.540 1794.280 ;
        RECT 2849.770 1794.220 2850.090 1794.280 ;
        RECT 2849.770 1793.740 2850.090 1793.800 ;
        RECT 2851.150 1793.740 2851.470 1793.800 ;
        RECT 2849.770 1793.600 2851.470 1793.740 ;
        RECT 2849.770 1793.540 2850.090 1793.600 ;
        RECT 2851.150 1793.540 2851.470 1793.600 ;
        RECT 2849.770 1793.060 2850.090 1793.120 ;
        RECT 2849.400 1792.920 2850.090 1793.060 ;
        RECT 2849.770 1792.860 2850.090 1792.920 ;
        RECT 2849.770 1791.360 2850.090 1791.420 ;
        RECT 2850.245 1791.360 2850.535 1791.405 ;
        RECT 2849.770 1791.220 2850.535 1791.360 ;
        RECT 2849.770 1791.160 2850.090 1791.220 ;
        RECT 2850.245 1791.175 2850.535 1791.220 ;
        RECT 2851.150 1790.340 2851.470 1790.400 ;
        RECT 2851.625 1790.340 2851.915 1790.385 ;
        RECT 2851.150 1790.200 2851.915 1790.340 ;
        RECT 2851.150 1790.140 2851.470 1790.200 ;
        RECT 2851.625 1790.155 2851.915 1790.200 ;
        RECT 2849.770 1768.720 2850.090 1768.980 ;
        RECT 2849.860 1768.580 2850.000 1768.720 ;
        RECT 2852.545 1768.580 2852.835 1768.625 ;
        RECT 2849.860 1768.440 2852.835 1768.580 ;
        RECT 2852.545 1768.395 2852.835 1768.440 ;
        RECT 2851.610 1766.540 2851.930 1766.600 ;
        RECT 2849.400 1766.400 2851.930 1766.540 ;
        RECT 2849.400 1766.260 2849.540 1766.400 ;
        RECT 2851.610 1766.340 2851.930 1766.400 ;
        RECT 2849.310 1766.000 2849.630 1766.260 ;
        RECT 2850.245 1762.460 2850.535 1762.505 ;
        RECT 2851.165 1762.460 2851.455 1762.505 ;
        RECT 2850.245 1762.320 2851.455 1762.460 ;
        RECT 2850.245 1762.275 2850.535 1762.320 ;
        RECT 2851.165 1762.275 2851.455 1762.320 ;
        RECT 2849.770 1761.780 2850.090 1761.840 ;
        RECT 2852.085 1761.780 2852.375 1761.825 ;
        RECT 2849.770 1761.640 2852.375 1761.780 ;
        RECT 2849.770 1761.580 2850.090 1761.640 ;
        RECT 2852.085 1761.595 2852.375 1761.640 ;
        RECT 2849.770 1740.020 2850.090 1740.080 ;
        RECT 2851.165 1740.020 2851.455 1740.065 ;
        RECT 2849.770 1739.880 2851.455 1740.020 ;
        RECT 2849.770 1739.820 2850.090 1739.880 ;
        RECT 2851.165 1739.835 2851.455 1739.880 ;
        RECT 2849.325 1647.880 2849.615 1647.925 ;
        RECT 2849.770 1647.880 2850.090 1647.940 ;
        RECT 2849.325 1647.740 2850.090 1647.880 ;
        RECT 2849.325 1647.695 2849.615 1647.740 ;
        RECT 2849.770 1647.680 2850.090 1647.740 ;
        RECT 2849.770 1647.200 2850.090 1647.260 ;
        RECT 2851.165 1647.200 2851.455 1647.245 ;
        RECT 2849.770 1647.060 2851.455 1647.200 ;
        RECT 2849.770 1647.000 2850.090 1647.060 ;
        RECT 2851.165 1647.015 2851.455 1647.060 ;
        RECT 2849.770 1646.520 2850.090 1646.580 ;
        RECT 2851.625 1646.520 2851.915 1646.565 ;
        RECT 2849.770 1646.380 2851.915 1646.520 ;
        RECT 2849.770 1646.320 2850.090 1646.380 ;
        RECT 2851.625 1646.335 2851.915 1646.380 ;
        RECT 2849.770 1639.040 2850.090 1639.100 ;
        RECT 2849.400 1638.900 2850.090 1639.040 ;
        RECT 2849.400 1635.980 2849.540 1638.900 ;
        RECT 2849.770 1638.840 2850.090 1638.900 ;
        RECT 2849.770 1638.360 2850.090 1638.420 ;
        RECT 2863.570 1638.360 2863.890 1638.420 ;
        RECT 2849.770 1638.220 2863.890 1638.360 ;
        RECT 2849.770 1638.160 2850.090 1638.220 ;
        RECT 2863.570 1638.160 2863.890 1638.220 ;
        RECT 2849.770 1635.980 2850.090 1636.040 ;
        RECT 2849.400 1635.840 2850.090 1635.980 ;
        RECT 2849.770 1635.780 2850.090 1635.840 ;
        RECT 2849.770 1635.300 2850.090 1635.360 ;
        RECT 2851.625 1635.300 2851.915 1635.345 ;
        RECT 2849.770 1635.160 2851.915 1635.300 ;
        RECT 2849.770 1635.100 2850.090 1635.160 ;
        RECT 2851.625 1635.115 2851.915 1635.160 ;
        RECT 2849.770 1628.500 2850.090 1628.560 ;
        RECT 2851.165 1628.500 2851.455 1628.545 ;
        RECT 2849.770 1628.360 2851.455 1628.500 ;
        RECT 2849.770 1628.300 2850.090 1628.360 ;
        RECT 2851.165 1628.315 2851.455 1628.360 ;
        RECT 2850.690 1627.820 2851.010 1627.880 ;
        RECT 2851.165 1627.820 2851.455 1627.865 ;
        RECT 2850.690 1627.680 2851.455 1627.820 ;
        RECT 2850.690 1627.620 2851.010 1627.680 ;
        RECT 2851.165 1627.635 2851.455 1627.680 ;
        RECT 2850.245 1605.040 2850.535 1605.085 ;
        RECT 2850.690 1605.040 2851.010 1605.100 ;
        RECT 2850.245 1604.900 2851.010 1605.040 ;
        RECT 2850.245 1604.855 2850.535 1604.900 ;
        RECT 2850.690 1604.840 2851.010 1604.900 ;
        RECT 2849.770 1604.360 2850.090 1604.420 ;
        RECT 2849.770 1604.220 2850.285 1604.360 ;
        RECT 2849.770 1604.160 2850.090 1604.220 ;
        RECT 2849.785 1579.695 2850.075 1579.925 ;
        RECT 2849.860 1579.245 2850.000 1579.695 ;
        RECT 2849.785 1579.015 2850.075 1579.245 ;
        RECT 2850.230 1579.200 2850.550 1579.260 ;
        RECT 2851.610 1579.200 2851.930 1579.260 ;
        RECT 2850.230 1579.060 2851.930 1579.200 ;
        RECT 2850.230 1579.000 2850.550 1579.060 ;
        RECT 2851.610 1579.000 2851.930 1579.060 ;
        RECT 2849.770 1578.180 2850.090 1578.240 ;
        RECT 2849.770 1578.040 2850.285 1578.180 ;
        RECT 2849.770 1577.980 2850.090 1578.040 ;
        RECT 2849.770 1545.540 2850.090 1545.600 ;
        RECT 2850.245 1545.540 2850.535 1545.585 ;
        RECT 2849.770 1545.400 2850.535 1545.540 ;
        RECT 2849.770 1545.340 2850.090 1545.400 ;
        RECT 2850.245 1545.355 2850.535 1545.400 ;
        RECT 2849.770 1535.000 2850.090 1535.060 ;
        RECT 2852.085 1535.000 2852.375 1535.045 ;
        RECT 2849.770 1534.860 2852.375 1535.000 ;
        RECT 2849.770 1534.800 2850.090 1534.860 ;
        RECT 2852.085 1534.815 2852.375 1534.860 ;
        RECT 2849.770 1530.920 2850.090 1530.980 ;
        RECT 2849.575 1530.780 2850.090 1530.920 ;
        RECT 2849.770 1530.720 2850.090 1530.780 ;
        RECT 2849.770 1513.920 2850.090 1513.980 ;
        RECT 2851.165 1513.920 2851.455 1513.965 ;
        RECT 2849.770 1513.780 2851.455 1513.920 ;
        RECT 2849.770 1513.720 2850.090 1513.780 ;
        RECT 2851.165 1513.735 2851.455 1513.780 ;
        RECT 2849.785 1509.500 2850.075 1509.545 ;
        RECT 2852.085 1509.500 2852.375 1509.545 ;
        RECT 2849.785 1509.360 2852.375 1509.500 ;
        RECT 2849.785 1509.315 2850.075 1509.360 ;
        RECT 2852.085 1509.315 2852.375 1509.360 ;
        RECT 2849.770 1505.760 2850.090 1505.820 ;
        RECT 2852.085 1505.760 2852.375 1505.805 ;
        RECT 2849.770 1505.620 2852.375 1505.760 ;
        RECT 2849.770 1505.560 2850.090 1505.620 ;
        RECT 2852.085 1505.575 2852.375 1505.620 ;
        RECT 2849.770 1504.400 2850.090 1504.460 ;
        RECT 2849.770 1504.260 2850.285 1504.400 ;
        RECT 2849.770 1504.200 2850.090 1504.260 ;
        RECT 2849.770 1500.320 2850.090 1500.380 ;
        RECT 2849.575 1500.180 2850.090 1500.320 ;
        RECT 2849.770 1500.120 2850.090 1500.180 ;
        RECT 2849.770 1492.840 2850.090 1492.900 ;
        RECT 2849.575 1492.700 2850.090 1492.840 ;
        RECT 2849.770 1492.640 2850.090 1492.700 ;
        RECT 2849.770 1492.160 2850.090 1492.220 ;
        RECT 2851.165 1492.160 2851.455 1492.205 ;
        RECT 2849.770 1492.020 2851.455 1492.160 ;
        RECT 2849.770 1491.960 2850.090 1492.020 ;
        RECT 2851.165 1491.975 2851.455 1492.020 ;
        RECT 2850.230 1480.940 2850.550 1481.000 ;
        RECT 2850.705 1480.940 2850.995 1480.985 ;
        RECT 2850.230 1480.800 2850.995 1480.940 ;
        RECT 2850.230 1480.740 2850.550 1480.800 ;
        RECT 2850.705 1480.755 2850.995 1480.800 ;
        RECT 2850.705 1480.260 2850.995 1480.305 ;
        RECT 2851.150 1480.260 2851.470 1480.320 ;
        RECT 2850.705 1480.120 2851.470 1480.260 ;
        RECT 2850.705 1480.075 2850.995 1480.120 ;
        RECT 2851.150 1480.060 2851.470 1480.120 ;
        RECT 2849.770 1462.240 2850.090 1462.300 ;
        RECT 2852.085 1462.240 2852.375 1462.285 ;
        RECT 2849.770 1462.100 2852.375 1462.240 ;
        RECT 2849.770 1462.040 2850.090 1462.100 ;
        RECT 2852.085 1462.055 2852.375 1462.100 ;
        RECT 2849.770 1448.300 2850.090 1448.360 ;
        RECT 2852.545 1448.300 2852.835 1448.345 ;
        RECT 2849.770 1448.160 2852.835 1448.300 ;
        RECT 2849.770 1448.100 2850.090 1448.160 ;
        RECT 2852.545 1448.115 2852.835 1448.160 ;
        RECT 2849.785 1428.240 2850.075 1428.285 ;
        RECT 2851.165 1428.240 2851.455 1428.285 ;
        RECT 2849.785 1428.100 2851.455 1428.240 ;
        RECT 2849.785 1428.055 2850.075 1428.100 ;
        RECT 2851.165 1428.055 2851.455 1428.100 ;
        RECT 2849.770 1426.880 2850.090 1426.940 ;
        RECT 2850.705 1426.880 2850.995 1426.925 ;
        RECT 2849.770 1426.740 2850.995 1426.880 ;
        RECT 2849.770 1426.680 2850.090 1426.740 ;
        RECT 2850.705 1426.695 2850.995 1426.740 ;
        RECT 2849.770 1425.860 2850.090 1425.920 ;
        RECT 2849.575 1425.720 2850.090 1425.860 ;
        RECT 2849.770 1425.660 2850.090 1425.720 ;
        RECT 2849.770 1424.840 2850.090 1424.900 ;
        RECT 2851.625 1424.840 2851.915 1424.885 ;
        RECT 2849.770 1424.700 2851.915 1424.840 ;
        RECT 2849.770 1424.640 2850.090 1424.700 ;
        RECT 2851.625 1424.655 2851.915 1424.700 ;
        RECT 2849.770 1424.160 2850.090 1424.220 ;
        RECT 2853.005 1424.160 2853.295 1424.205 ;
        RECT 2849.770 1424.020 2853.295 1424.160 ;
        RECT 2849.770 1423.960 2850.090 1424.020 ;
        RECT 2853.005 1423.975 2853.295 1424.020 ;
        RECT 2849.770 1423.140 2850.090 1423.200 ;
        RECT 2852.530 1423.140 2852.850 1423.200 ;
        RECT 2849.770 1423.000 2852.850 1423.140 ;
        RECT 2849.770 1422.940 2850.090 1423.000 ;
        RECT 2852.530 1422.940 2852.850 1423.000 ;
        RECT 2849.770 1419.400 2850.090 1419.460 ;
        RECT 2849.770 1419.260 2850.460 1419.400 ;
        RECT 2849.770 1419.200 2850.090 1419.260 ;
        RECT 2849.770 1418.720 2850.090 1418.780 ;
        RECT 2849.575 1418.580 2850.090 1418.720 ;
        RECT 2849.770 1418.520 2850.090 1418.580 ;
        RECT 2850.320 1418.380 2850.460 1419.260 ;
        RECT 2849.400 1418.240 2850.460 1418.380 ;
        RECT 2849.400 1416.680 2849.540 1418.240 ;
        RECT 2850.245 1418.040 2850.535 1418.085 ;
        RECT 2851.165 1418.040 2851.455 1418.085 ;
        RECT 2850.245 1417.900 2851.455 1418.040 ;
        RECT 2850.245 1417.855 2850.535 1417.900 ;
        RECT 2851.165 1417.855 2851.455 1417.900 ;
        RECT 2849.770 1417.700 2850.090 1417.760 ;
        RECT 2852.545 1417.700 2852.835 1417.745 ;
        RECT 2849.770 1417.560 2852.835 1417.700 ;
        RECT 2849.770 1417.500 2850.090 1417.560 ;
        RECT 2852.545 1417.515 2852.835 1417.560 ;
        RECT 2849.770 1417.020 2850.090 1417.080 ;
        RECT 2851.625 1417.020 2851.915 1417.065 ;
        RECT 2849.770 1416.880 2851.915 1417.020 ;
        RECT 2849.770 1416.820 2850.090 1416.880 ;
        RECT 2851.625 1416.835 2851.915 1416.880 ;
        RECT 2850.230 1416.680 2850.550 1416.740 ;
        RECT 2849.400 1416.540 2850.550 1416.680 ;
        RECT 2850.230 1416.480 2850.550 1416.540 ;
        RECT 2849.770 1389.820 2850.090 1389.880 ;
        RECT 2851.610 1389.820 2851.930 1389.880 ;
        RECT 2849.770 1389.680 2851.930 1389.820 ;
        RECT 2849.770 1389.620 2850.090 1389.680 ;
        RECT 2851.610 1389.620 2851.930 1389.680 ;
        RECT 2849.770 1387.780 2850.090 1387.840 ;
        RECT 2850.690 1387.780 2851.010 1387.840 ;
        RECT 2849.770 1387.640 2851.010 1387.780 ;
        RECT 2849.770 1387.580 2850.090 1387.640 ;
        RECT 2850.690 1387.580 2851.010 1387.640 ;
        RECT 2849.770 1386.420 2850.090 1386.480 ;
        RECT 2852.545 1386.420 2852.835 1386.465 ;
        RECT 2849.770 1386.280 2852.835 1386.420 ;
        RECT 2849.770 1386.220 2850.090 1386.280 ;
        RECT 2852.545 1386.235 2852.835 1386.280 ;
        RECT 2849.770 1372.480 2850.090 1372.540 ;
        RECT 2853.465 1372.480 2853.755 1372.525 ;
        RECT 2849.770 1372.340 2853.755 1372.480 ;
        RECT 2849.770 1372.280 2850.090 1372.340 ;
        RECT 2853.465 1372.295 2853.755 1372.340 ;
        RECT 2850.705 1371.800 2850.995 1371.845 ;
        RECT 2851.625 1371.800 2851.915 1371.845 ;
        RECT 2850.705 1371.660 2851.915 1371.800 ;
        RECT 2850.705 1371.615 2850.995 1371.660 ;
        RECT 2851.625 1371.615 2851.915 1371.660 ;
        RECT 2849.770 1371.120 2850.090 1371.180 ;
        RECT 2849.400 1370.980 2850.090 1371.120 ;
        RECT 2849.400 1368.740 2849.540 1370.980 ;
        RECT 2849.770 1370.920 2850.090 1370.980 ;
        RECT 2850.230 1368.740 2850.550 1368.800 ;
        RECT 2849.400 1368.600 2850.550 1368.740 ;
        RECT 2850.230 1368.540 2850.550 1368.600 ;
        RECT 2849.770 1365.340 2850.090 1365.400 ;
        RECT 2849.575 1365.200 2850.090 1365.340 ;
        RECT 2849.770 1365.140 2850.090 1365.200 ;
        RECT 2849.770 1364.660 2850.090 1364.720 ;
        RECT 2853.465 1364.660 2853.755 1364.705 ;
        RECT 2849.770 1364.520 2853.755 1364.660 ;
        RECT 2849.770 1364.460 2850.090 1364.520 ;
        RECT 2853.465 1364.475 2853.755 1364.520 ;
        RECT 2849.770 1363.980 2850.090 1364.040 ;
        RECT 2863.570 1363.980 2863.890 1364.040 ;
        RECT 2849.770 1363.840 2863.890 1363.980 ;
        RECT 2849.770 1363.780 2850.090 1363.840 ;
        RECT 2863.570 1363.780 2863.890 1363.840 ;
        RECT 2849.770 1362.960 2850.090 1363.020 ;
        RECT 2852.070 1362.960 2852.390 1363.020 ;
        RECT 2849.770 1362.820 2852.390 1362.960 ;
        RECT 2849.770 1362.760 2850.090 1362.820 ;
        RECT 2852.070 1362.760 2852.390 1362.820 ;
        RECT 2853.005 1362.620 2853.295 1362.665 ;
        RECT 2849.400 1362.480 2853.295 1362.620 ;
        RECT 2849.400 1362.000 2849.540 1362.480 ;
        RECT 2853.005 1362.435 2853.295 1362.480 ;
        RECT 2849.310 1361.740 2849.630 1362.000 ;
        RECT 2849.770 1357.860 2850.090 1357.920 ;
        RECT 2849.575 1357.720 2850.090 1357.860 ;
        RECT 2849.770 1357.660 2850.090 1357.720 ;
        RECT 2849.770 1355.140 2850.090 1355.200 ;
        RECT 2852.545 1355.140 2852.835 1355.185 ;
        RECT 2849.770 1355.000 2852.835 1355.140 ;
        RECT 2849.770 1354.940 2850.090 1355.000 ;
        RECT 2852.545 1354.955 2852.835 1355.000 ;
        RECT 2849.770 1354.460 2850.090 1354.520 ;
        RECT 2850.690 1354.460 2851.010 1354.520 ;
        RECT 2849.770 1354.320 2851.010 1354.460 ;
        RECT 2849.770 1354.260 2850.090 1354.320 ;
        RECT 2850.690 1354.260 2851.010 1354.320 ;
        RECT 2849.770 1353.100 2850.090 1353.160 ;
        RECT 2851.610 1353.100 2851.930 1353.160 ;
        RECT 2849.770 1352.960 2851.930 1353.100 ;
        RECT 2849.770 1352.900 2850.090 1352.960 ;
        RECT 2851.610 1352.900 2851.930 1352.960 ;
        RECT 2849.770 1352.420 2850.090 1352.480 ;
        RECT 2850.705 1352.420 2850.995 1352.465 ;
        RECT 2849.770 1352.280 2850.995 1352.420 ;
        RECT 2849.770 1352.220 2850.090 1352.280 ;
        RECT 2850.705 1352.235 2850.995 1352.280 ;
        RECT 2849.770 1350.380 2850.090 1350.440 ;
        RECT 2851.625 1350.380 2851.915 1350.425 ;
        RECT 2849.770 1350.240 2851.915 1350.380 ;
        RECT 2849.770 1350.180 2850.090 1350.240 ;
        RECT 2851.625 1350.195 2851.915 1350.240 ;
        RECT 2849.770 1329.640 2850.090 1329.700 ;
        RECT 2850.705 1329.640 2850.995 1329.685 ;
        RECT 2849.770 1329.500 2850.995 1329.640 ;
        RECT 2849.770 1329.440 2850.090 1329.500 ;
        RECT 2850.705 1329.455 2850.995 1329.500 ;
        RECT 2849.770 1258.920 2850.090 1258.980 ;
        RECT 2850.690 1258.920 2851.010 1258.980 ;
        RECT 2849.770 1258.780 2851.010 1258.920 ;
        RECT 2849.770 1258.720 2850.090 1258.780 ;
        RECT 2850.690 1258.720 2851.010 1258.780 ;
        RECT 2849.770 1254.840 2850.090 1254.900 ;
        RECT 2851.165 1254.840 2851.455 1254.885 ;
        RECT 2849.770 1254.700 2851.455 1254.840 ;
        RECT 2849.770 1254.640 2850.090 1254.700 ;
        RECT 2851.165 1254.655 2851.455 1254.700 ;
        RECT 2849.770 1254.160 2850.090 1254.220 ;
        RECT 2851.610 1254.160 2851.930 1254.220 ;
        RECT 2849.770 1254.020 2851.930 1254.160 ;
        RECT 2849.770 1253.960 2850.090 1254.020 ;
        RECT 2851.610 1253.960 2851.930 1254.020 ;
        RECT 2849.770 1253.140 2850.090 1253.200 ;
        RECT 2852.545 1253.140 2852.835 1253.185 ;
        RECT 2849.770 1253.000 2852.835 1253.140 ;
        RECT 2849.770 1252.940 2850.090 1253.000 ;
        RECT 2852.545 1252.955 2852.835 1253.000 ;
        RECT 2850.230 1232.740 2850.550 1232.800 ;
        RECT 2851.165 1232.740 2851.455 1232.785 ;
        RECT 2850.230 1232.600 2851.455 1232.740 ;
        RECT 2850.230 1232.540 2850.550 1232.600 ;
        RECT 2851.165 1232.555 2851.455 1232.600 ;
        RECT 2849.325 1226.960 2849.615 1227.005 ;
        RECT 2852.545 1226.960 2852.835 1227.005 ;
        RECT 2849.325 1226.820 2852.835 1226.960 ;
        RECT 2849.325 1226.775 2849.615 1226.820 ;
        RECT 2852.545 1226.775 2852.835 1226.820 ;
        RECT 2850.690 1197.380 2851.010 1197.440 ;
        RECT 2852.085 1197.380 2852.375 1197.425 ;
        RECT 2850.690 1197.240 2852.375 1197.380 ;
        RECT 2850.690 1197.180 2851.010 1197.240 ;
        RECT 2852.085 1197.195 2852.375 1197.240 ;
        RECT 2849.770 1167.800 2850.090 1167.860 ;
        RECT 2850.690 1167.800 2851.010 1167.860 ;
        RECT 2849.770 1167.660 2851.010 1167.800 ;
        RECT 2849.770 1167.600 2850.090 1167.660 ;
        RECT 2850.690 1167.600 2851.010 1167.660 ;
        RECT 2849.770 1151.140 2850.090 1151.200 ;
        RECT 2849.575 1151.000 2850.090 1151.140 ;
        RECT 2849.770 1150.940 2850.090 1151.000 ;
        RECT 2849.770 1150.120 2850.090 1150.180 ;
        RECT 2850.690 1150.120 2851.010 1150.180 ;
        RECT 2849.770 1149.980 2851.010 1150.120 ;
        RECT 2849.770 1149.920 2850.090 1149.980 ;
        RECT 2850.690 1149.920 2851.010 1149.980 ;
        RECT 2849.770 1149.100 2850.090 1149.160 ;
        RECT 2851.610 1149.100 2851.930 1149.160 ;
        RECT 2849.770 1148.960 2851.930 1149.100 ;
        RECT 2849.770 1148.900 2850.090 1148.960 ;
        RECT 2851.610 1148.900 2851.930 1148.960 ;
        RECT 2850.690 1148.760 2851.010 1148.820 ;
        RECT 2851.165 1148.760 2851.455 1148.805 ;
        RECT 2850.690 1148.620 2851.455 1148.760 ;
        RECT 2850.690 1148.560 2851.010 1148.620 ;
        RECT 2851.165 1148.575 2851.455 1148.620 ;
        RECT 2849.785 1148.420 2850.075 1148.465 ;
        RECT 2850.230 1148.420 2850.550 1148.480 ;
        RECT 2849.785 1148.280 2850.550 1148.420 ;
        RECT 2849.785 1148.235 2850.075 1148.280 ;
        RECT 2850.230 1148.220 2850.550 1148.280 ;
        RECT 2849.770 1129.040 2850.090 1129.100 ;
        RECT 2851.625 1129.040 2851.915 1129.085 ;
        RECT 2849.770 1128.900 2851.915 1129.040 ;
        RECT 2849.770 1128.840 2850.090 1128.900 ;
        RECT 2851.625 1128.855 2851.915 1128.900 ;
        RECT 2849.770 1078.380 2850.090 1078.440 ;
        RECT 2849.400 1078.240 2850.090 1078.380 ;
        RECT 2849.400 1077.020 2849.540 1078.240 ;
        RECT 2849.770 1078.180 2850.090 1078.240 ;
        RECT 2849.770 1077.020 2850.090 1077.080 ;
        RECT 2849.400 1076.880 2850.090 1077.020 ;
        RECT 2849.770 1076.820 2850.090 1076.880 ;
        RECT 2849.770 1073.280 2850.090 1073.340 ;
        RECT 2851.625 1073.280 2851.915 1073.325 ;
        RECT 2849.770 1073.140 2851.915 1073.280 ;
        RECT 2849.770 1073.080 2850.090 1073.140 ;
        RECT 2851.625 1073.095 2851.915 1073.140 ;
        RECT 2850.690 1072.940 2851.010 1073.000 ;
        RECT 2850.495 1072.800 2851.010 1072.940 ;
        RECT 2850.690 1072.740 2851.010 1072.800 ;
        RECT 2849.770 1023.980 2850.090 1024.040 ;
        RECT 2850.245 1023.980 2850.535 1024.025 ;
        RECT 2849.770 1023.840 2850.535 1023.980 ;
        RECT 2849.770 1023.780 2850.090 1023.840 ;
        RECT 2850.245 1023.795 2850.535 1023.840 ;
        RECT 2849.770 1017.860 2850.090 1017.920 ;
        RECT 2851.625 1017.860 2851.915 1017.905 ;
        RECT 2849.770 1017.720 2851.915 1017.860 ;
        RECT 2849.770 1017.660 2850.090 1017.720 ;
        RECT 2851.625 1017.675 2851.915 1017.720 ;
        RECT 2849.770 1015.140 2850.090 1015.200 ;
        RECT 2850.705 1015.140 2850.995 1015.185 ;
        RECT 2849.770 1015.000 2850.995 1015.140 ;
        RECT 2849.770 1014.940 2850.090 1015.000 ;
        RECT 2850.705 1014.955 2850.995 1015.000 ;
        RECT 2850.230 960.060 2850.550 960.120 ;
        RECT 2849.400 959.920 2850.550 960.060 ;
        RECT 2849.400 959.380 2849.540 959.920 ;
        RECT 2850.230 959.860 2850.550 959.920 ;
        RECT 2849.770 959.720 2850.090 959.780 ;
        RECT 2851.165 959.720 2851.455 959.765 ;
        RECT 2849.770 959.580 2851.455 959.720 ;
        RECT 2849.770 959.520 2850.090 959.580 ;
        RECT 2851.165 959.535 2851.455 959.580 ;
        RECT 2849.400 959.240 2850.460 959.380 ;
        RECT 2850.320 958.760 2850.460 959.240 ;
        RECT 2849.770 958.700 2850.090 958.760 ;
        RECT 2849.400 958.560 2850.090 958.700 ;
        RECT 2849.400 957.340 2849.540 958.560 ;
        RECT 2849.770 958.500 2850.090 958.560 ;
        RECT 2850.230 958.500 2850.550 958.760 ;
        RECT 2849.770 958.020 2850.090 958.080 ;
        RECT 2851.610 958.020 2851.930 958.080 ;
        RECT 2849.770 957.880 2851.930 958.020 ;
        RECT 2849.770 957.820 2850.090 957.880 ;
        RECT 2851.610 957.820 2851.930 957.880 ;
        RECT 2849.770 957.340 2850.090 957.400 ;
        RECT 2849.400 957.200 2850.090 957.340 ;
        RECT 2849.770 957.140 2850.090 957.200 ;
        RECT 2849.770 943.060 2850.090 943.120 ;
        RECT 2851.150 943.060 2851.470 943.120 ;
        RECT 2849.770 942.920 2851.470 943.060 ;
        RECT 2849.770 942.860 2850.090 942.920 ;
        RECT 2851.150 942.860 2851.470 942.920 ;
        RECT 2849.770 874.720 2850.090 874.780 ;
        RECT 2849.575 874.580 2850.090 874.720 ;
        RECT 2849.770 874.520 2850.090 874.580 ;
        RECT 2849.770 868.260 2850.090 868.320 ;
        RECT 2850.690 868.260 2851.010 868.320 ;
        RECT 2849.770 868.120 2851.010 868.260 ;
        RECT 2849.770 868.060 2850.090 868.120 ;
        RECT 2850.690 868.060 2851.010 868.120 ;
        RECT 2850.230 859.760 2850.550 859.820 ;
        RECT 2852.085 859.760 2852.375 859.805 ;
        RECT 2850.230 859.620 2852.375 859.760 ;
        RECT 2850.230 859.560 2850.550 859.620 ;
        RECT 2852.085 859.575 2852.375 859.620 ;
        RECT 2849.770 846.640 2850.090 846.900 ;
        RECT 2849.860 845.880 2850.000 846.640 ;
        RECT 2849.770 845.620 2850.090 845.880 ;
        RECT 2849.770 845.140 2850.090 845.200 ;
        RECT 2850.690 845.140 2851.010 845.200 ;
        RECT 2849.770 845.000 2851.010 845.140 ;
        RECT 2849.770 844.940 2850.090 845.000 ;
        RECT 2850.690 844.940 2851.010 845.000 ;
        RECT 2849.770 818.620 2850.090 818.680 ;
        RECT 2849.575 818.480 2850.090 818.620 ;
        RECT 2849.770 818.420 2850.090 818.480 ;
        RECT 2852.070 811.140 2852.390 811.200 ;
        RECT 2851.875 811.000 2852.390 811.140 ;
        RECT 2852.070 810.940 2852.390 811.000 ;
        RECT 2849.785 793.800 2850.075 793.845 ;
        RECT 2851.625 793.800 2851.915 793.845 ;
        RECT 2849.785 793.660 2851.915 793.800 ;
        RECT 2849.785 793.615 2850.075 793.660 ;
        RECT 2851.625 793.615 2851.915 793.660 ;
        RECT 2849.785 790.060 2850.075 790.105 ;
        RECT 2850.705 790.060 2850.995 790.105 ;
        RECT 2849.785 789.920 2850.995 790.060 ;
        RECT 2849.785 789.875 2850.075 789.920 ;
        RECT 2850.705 789.875 2850.995 789.920 ;
        RECT 2850.690 788.360 2851.010 788.420 ;
        RECT 2852.545 788.360 2852.835 788.405 ;
        RECT 2850.690 788.220 2852.835 788.360 ;
        RECT 2850.690 788.160 2851.010 788.220 ;
        RECT 2852.545 788.175 2852.835 788.220 ;
        RECT 2849.770 787.680 2850.090 787.740 ;
        RECT 2850.690 787.680 2851.010 787.740 ;
        RECT 2849.770 787.540 2851.010 787.680 ;
        RECT 2849.770 787.480 2850.090 787.540 ;
        RECT 2850.690 787.480 2851.010 787.540 ;
        RECT 2849.770 787.000 2850.090 787.060 ;
        RECT 2851.625 787.000 2851.915 787.045 ;
        RECT 2849.770 786.860 2851.915 787.000 ;
        RECT 2849.770 786.800 2850.090 786.860 ;
        RECT 2851.625 786.815 2851.915 786.860 ;
        RECT 2849.770 779.320 2850.090 779.580 ;
        RECT 2849.860 778.840 2850.000 779.320 ;
        RECT 2851.150 778.840 2851.470 778.900 ;
        RECT 2849.860 778.700 2851.470 778.840 ;
        RECT 2851.150 778.640 2851.470 778.700 ;
        RECT 2849.770 775.920 2850.090 776.180 ;
        RECT 2849.310 775.580 2849.630 775.840 ;
        RECT 2849.400 774.420 2849.540 775.580 ;
        RECT 2849.860 775.440 2850.000 775.920 ;
        RECT 2850.230 775.440 2850.550 775.500 ;
        RECT 2849.860 775.300 2850.550 775.440 ;
        RECT 2850.230 775.240 2850.550 775.300 ;
        RECT 2849.770 775.100 2850.090 775.160 ;
        RECT 2852.545 775.100 2852.835 775.145 ;
        RECT 2849.770 774.960 2852.835 775.100 ;
        RECT 2849.770 774.900 2850.090 774.960 ;
        RECT 2852.545 774.915 2852.835 774.960 ;
        RECT 2849.770 774.420 2850.090 774.480 ;
        RECT 2849.400 774.280 2850.090 774.420 ;
        RECT 2849.770 774.220 2850.090 774.280 ;
        RECT 2849.770 769.320 2850.090 769.380 ;
        RECT 2851.150 769.320 2851.470 769.380 ;
        RECT 2849.770 769.180 2851.470 769.320 ;
        RECT 2849.770 769.120 2850.090 769.180 ;
        RECT 2851.150 769.120 2851.470 769.180 ;
        RECT 2851.150 745.520 2851.470 745.580 ;
        RECT 2852.070 745.520 2852.390 745.580 ;
        RECT 2851.150 745.380 2852.390 745.520 ;
        RECT 2851.150 745.320 2851.470 745.380 ;
        RECT 2852.070 745.320 2852.390 745.380 ;
        RECT 2849.770 739.740 2850.090 739.800 ;
        RECT 2851.165 739.740 2851.455 739.785 ;
        RECT 2849.770 739.600 2851.455 739.740 ;
        RECT 2849.770 739.540 2850.090 739.600 ;
        RECT 2851.165 739.555 2851.455 739.600 ;
        RECT 2849.770 739.060 2850.090 739.120 ;
        RECT 2850.690 739.060 2851.010 739.120 ;
        RECT 2849.770 738.920 2851.010 739.060 ;
        RECT 2849.770 738.860 2850.090 738.920 ;
        RECT 2850.690 738.860 2851.010 738.920 ;
        RECT 2849.770 738.380 2850.090 738.440 ;
        RECT 2850.705 738.380 2850.995 738.425 ;
        RECT 2849.770 738.240 2850.995 738.380 ;
        RECT 2849.770 738.180 2850.090 738.240 ;
        RECT 2850.705 738.195 2850.995 738.240 ;
        RECT 2849.770 671.740 2850.090 671.800 ;
        RECT 2851.150 671.740 2851.470 671.800 ;
        RECT 2849.770 671.600 2851.470 671.740 ;
        RECT 2849.770 671.540 2850.090 671.600 ;
        RECT 2851.150 671.540 2851.470 671.600 ;
        RECT 2849.770 383.080 2850.090 383.140 ;
        RECT 2851.165 383.080 2851.455 383.125 ;
        RECT 2849.770 382.940 2851.455 383.080 ;
        RECT 2849.770 382.880 2850.090 382.940 ;
        RECT 2851.165 382.895 2851.455 382.940 ;
        RECT 2849.770 381.040 2850.090 381.100 ;
        RECT 2851.625 381.040 2851.915 381.085 ;
        RECT 2849.770 380.900 2851.915 381.040 ;
        RECT 2849.770 380.840 2850.090 380.900 ;
        RECT 2851.625 380.855 2851.915 380.900 ;
        RECT 2849.785 379.680 2850.075 379.725 ;
        RECT 2851.165 379.680 2851.455 379.725 ;
        RECT 2849.785 379.540 2851.455 379.680 ;
        RECT 2849.785 379.495 2850.075 379.540 ;
        RECT 2851.165 379.495 2851.455 379.540 ;
        RECT 2849.770 374.240 2850.090 374.300 ;
        RECT 2851.625 374.240 2851.915 374.285 ;
        RECT 2849.770 374.100 2851.915 374.240 ;
        RECT 2849.770 374.040 2850.090 374.100 ;
        RECT 2851.625 374.055 2851.915 374.100 ;
        RECT 2849.770 373.560 2850.090 373.620 ;
        RECT 2851.150 373.560 2851.470 373.620 ;
        RECT 2849.770 373.420 2851.470 373.560 ;
        RECT 2849.770 373.360 2850.090 373.420 ;
        RECT 2851.150 373.360 2851.470 373.420 ;
        RECT 2849.770 368.800 2850.090 368.860 ;
        RECT 2849.400 368.660 2850.090 368.800 ;
        RECT 2849.400 365.740 2849.540 368.660 ;
        RECT 2849.770 368.600 2850.090 368.660 ;
        RECT 2849.770 368.120 2850.090 368.180 ;
        RECT 2852.085 368.120 2852.375 368.165 ;
        RECT 2849.770 367.980 2852.375 368.120 ;
        RECT 2849.770 367.920 2850.090 367.980 ;
        RECT 2852.085 367.935 2852.375 367.980 ;
        RECT 2849.770 367.100 2850.090 367.160 ;
        RECT 2852.545 367.100 2852.835 367.145 ;
        RECT 2849.770 366.960 2852.835 367.100 ;
        RECT 2849.770 366.900 2850.090 366.960 ;
        RECT 2852.545 366.915 2852.835 366.960 ;
        RECT 2849.770 366.420 2850.090 366.480 ;
        RECT 2851.150 366.420 2851.470 366.480 ;
        RECT 2849.770 366.280 2851.470 366.420 ;
        RECT 2849.770 366.220 2850.090 366.280 ;
        RECT 2851.150 366.220 2851.470 366.280 ;
        RECT 2849.770 365.740 2850.090 365.800 ;
        RECT 2849.400 365.600 2850.090 365.740 ;
        RECT 2849.770 365.540 2850.090 365.600 ;
        RECT 2849.770 365.060 2850.090 365.120 ;
        RECT 2852.085 365.060 2852.375 365.105 ;
        RECT 2849.770 364.920 2852.375 365.060 ;
        RECT 2849.770 364.860 2850.090 364.920 ;
        RECT 2852.085 364.875 2852.375 364.920 ;
        RECT 2849.770 362.340 2850.090 362.400 ;
        RECT 2851.625 362.340 2851.915 362.385 ;
        RECT 2849.770 362.200 2851.915 362.340 ;
        RECT 2849.770 362.140 2850.090 362.200 ;
        RECT 2851.625 362.155 2851.915 362.200 ;
        RECT 2849.770 341.940 2850.090 342.000 ;
        RECT 2851.150 341.940 2851.470 342.000 ;
        RECT 2849.770 341.800 2851.470 341.940 ;
        RECT 2849.770 341.740 2850.090 341.800 ;
        RECT 2851.150 341.740 2851.470 341.800 ;
        RECT 2849.770 340.240 2850.090 340.300 ;
        RECT 2851.625 340.240 2851.915 340.285 ;
        RECT 2849.770 340.100 2851.915 340.240 ;
        RECT 2849.770 340.040 2850.090 340.100 ;
        RECT 2851.625 340.055 2851.915 340.100 ;
        RECT 2850.690 330.720 2851.010 330.780 ;
        RECT 2852.545 330.720 2852.835 330.765 ;
        RECT 2850.690 330.580 2852.835 330.720 ;
        RECT 2850.690 330.520 2851.010 330.580 ;
        RECT 2852.545 330.535 2852.835 330.580 ;
        RECT 2849.770 308.620 2850.090 308.680 ;
        RECT 2849.400 308.480 2850.090 308.620 ;
        RECT 2849.400 306.580 2849.540 308.480 ;
        RECT 2849.770 308.420 2850.090 308.480 ;
        RECT 2849.770 307.940 2850.090 308.000 ;
        RECT 2850.690 307.940 2851.010 308.000 ;
        RECT 2849.770 307.800 2851.010 307.940 ;
        RECT 2849.770 307.740 2850.090 307.800 ;
        RECT 2850.690 307.740 2851.010 307.800 ;
        RECT 2850.230 306.580 2850.550 306.640 ;
        RECT 2849.400 306.440 2850.550 306.580 ;
        RECT 2850.230 306.380 2850.550 306.440 ;
        RECT 2849.770 303.860 2850.090 303.920 ;
        RECT 2851.625 303.860 2851.915 303.905 ;
        RECT 2849.770 303.720 2851.915 303.860 ;
        RECT 2849.770 303.660 2850.090 303.720 ;
        RECT 2851.625 303.675 2851.915 303.720 ;
        RECT 2849.770 299.780 2850.090 299.840 ;
        RECT 2851.165 299.780 2851.455 299.825 ;
        RECT 2849.770 299.640 2851.455 299.780 ;
        RECT 2849.770 299.580 2850.090 299.640 ;
        RECT 2851.165 299.595 2851.455 299.640 ;
        RECT 2849.770 284.820 2850.090 284.880 ;
        RECT 2849.575 284.680 2850.090 284.820 ;
        RECT 2849.770 284.620 2850.090 284.680 ;
        RECT 2849.770 211.040 2850.090 211.100 ;
        RECT 2851.165 211.040 2851.455 211.085 ;
        RECT 2849.770 210.900 2851.455 211.040 ;
        RECT 2849.770 210.840 2850.090 210.900 ;
        RECT 2851.165 210.855 2851.455 210.900 ;
        RECT 2849.770 208.320 2850.090 208.380 ;
        RECT 2850.245 208.320 2850.535 208.365 ;
        RECT 2849.770 208.180 2850.535 208.320 ;
        RECT 2849.770 208.120 2850.090 208.180 ;
        RECT 2850.245 208.135 2850.535 208.180 ;
        RECT 2849.770 205.600 2850.090 205.660 ;
        RECT 2850.705 205.600 2850.995 205.645 ;
        RECT 2849.770 205.460 2850.995 205.600 ;
        RECT 2849.770 205.400 2850.090 205.460 ;
        RECT 2850.705 205.415 2850.995 205.460 ;
        RECT 2849.770 204.920 2850.090 204.980 ;
        RECT 2849.575 204.780 2850.090 204.920 ;
        RECT 2849.770 204.720 2850.090 204.780 ;
        RECT 2849.770 203.560 2850.090 203.620 ;
        RECT 2849.400 203.420 2850.090 203.560 ;
        RECT 2849.400 200.840 2849.540 203.420 ;
        RECT 2849.770 203.360 2850.090 203.420 ;
        RECT 2849.770 202.200 2850.090 202.260 ;
        RECT 2852.085 202.200 2852.375 202.245 ;
        RECT 2849.770 202.060 2852.375 202.200 ;
        RECT 2849.770 202.000 2850.090 202.060 ;
        RECT 2852.085 202.015 2852.375 202.060 ;
        RECT 2849.770 201.520 2850.090 201.580 ;
        RECT 2853.005 201.520 2853.295 201.565 ;
        RECT 2849.770 201.380 2853.295 201.520 ;
        RECT 2849.770 201.320 2850.090 201.380 ;
        RECT 2853.005 201.335 2853.295 201.380 ;
        RECT 2849.770 200.840 2850.090 200.900 ;
        RECT 2849.400 200.700 2850.090 200.840 ;
        RECT 2849.770 200.640 2850.090 200.700 ;
        RECT 2849.770 200.160 2850.090 200.220 ;
        RECT 2852.085 200.160 2852.375 200.205 ;
        RECT 2849.770 200.020 2852.375 200.160 ;
        RECT 2849.770 199.960 2850.090 200.020 ;
        RECT 2852.085 199.975 2852.375 200.020 ;
        RECT 2849.770 199.480 2850.090 199.540 ;
        RECT 2850.705 199.480 2850.995 199.525 ;
        RECT 2849.770 199.340 2850.995 199.480 ;
        RECT 2849.770 199.280 2850.090 199.340 ;
        RECT 2850.705 199.295 2850.995 199.340 ;
        RECT 2849.770 198.460 2850.090 198.520 ;
        RECT 2849.575 198.320 2850.090 198.460 ;
        RECT 2849.770 198.260 2850.090 198.320 ;
        RECT 2849.770 197.100 2850.090 197.160 ;
        RECT 2850.245 197.100 2850.535 197.145 ;
        RECT 2849.770 196.960 2850.535 197.100 ;
        RECT 2849.770 196.900 2850.090 196.960 ;
        RECT 2850.245 196.915 2850.535 196.960 ;
        RECT 2851.610 173.980 2851.930 174.040 ;
        RECT 2853.005 173.980 2853.295 174.025 ;
        RECT 2851.610 173.840 2853.295 173.980 ;
        RECT 2851.610 173.780 2851.930 173.840 ;
        RECT 2853.005 173.795 2853.295 173.840 ;
        RECT 2849.785 139.640 2850.075 139.685 ;
        RECT 2851.165 139.640 2851.455 139.685 ;
        RECT 2849.785 139.500 2851.455 139.640 ;
        RECT 2849.785 139.455 2850.075 139.500 ;
        RECT 2851.165 139.455 2851.455 139.500 ;
        RECT 2849.770 132.500 2850.090 132.560 ;
        RECT 2851.165 132.500 2851.455 132.545 ;
        RECT 2849.770 132.360 2851.455 132.500 ;
        RECT 2849.770 132.300 2850.090 132.360 ;
        RECT 2851.165 132.315 2851.455 132.360 ;
        RECT 2849.770 128.760 2850.090 128.820 ;
        RECT 2850.245 128.760 2850.535 128.805 ;
        RECT 2849.770 128.620 2850.535 128.760 ;
        RECT 2849.770 128.560 2850.090 128.620 ;
        RECT 2850.245 128.575 2850.535 128.620 ;
        RECT 2849.770 127.740 2850.090 127.800 ;
        RECT 2852.085 127.740 2852.375 127.785 ;
        RECT 2849.770 127.600 2852.375 127.740 ;
        RECT 2849.770 127.540 2850.090 127.600 ;
        RECT 2852.085 127.555 2852.375 127.600 ;
        RECT 2849.770 125.700 2850.090 125.760 ;
        RECT 2851.150 125.700 2851.470 125.760 ;
        RECT 2849.770 125.560 2851.470 125.700 ;
        RECT 2849.770 125.500 2850.090 125.560 ;
        RECT 2851.150 125.500 2851.470 125.560 ;
        RECT 2849.770 121.620 2850.090 121.680 ;
        RECT 2851.610 121.620 2851.930 121.680 ;
        RECT 2849.770 121.480 2851.930 121.620 ;
        RECT 2849.770 121.420 2850.090 121.480 ;
        RECT 2851.610 121.420 2851.930 121.480 ;
        RECT 2849.770 120.940 2850.090 121.000 ;
        RECT 2852.085 120.940 2852.375 120.985 ;
        RECT 2849.770 120.800 2852.375 120.940 ;
        RECT 2849.770 120.740 2850.090 120.800 ;
        RECT 2852.085 120.755 2852.375 120.800 ;
        RECT 2849.770 118.900 2850.090 118.960 ;
        RECT 2851.165 118.900 2851.455 118.945 ;
        RECT 2849.770 118.760 2851.455 118.900 ;
        RECT 2849.770 118.700 2850.090 118.760 ;
        RECT 2851.165 118.715 2851.455 118.760 ;
        RECT 2849.770 117.880 2850.090 117.940 ;
        RECT 2851.150 117.880 2851.470 117.940 ;
        RECT 2849.770 117.740 2851.470 117.880 ;
        RECT 2849.770 117.680 2850.090 117.740 ;
        RECT 2851.150 117.680 2851.470 117.740 ;
        RECT 2849.785 115.500 2850.075 115.545 ;
        RECT 2850.705 115.500 2850.995 115.545 ;
        RECT 2849.785 115.360 2850.995 115.500 ;
        RECT 2849.785 115.315 2850.075 115.360 ;
        RECT 2850.705 115.315 2850.995 115.360 ;
        RECT 2849.770 88.300 2850.090 88.360 ;
        RECT 2850.705 88.300 2850.995 88.345 ;
        RECT 2849.770 88.160 2850.995 88.300 ;
        RECT 2849.770 88.100 2850.090 88.160 ;
        RECT 2850.705 88.115 2850.995 88.160 ;
        RECT 2850.245 73.680 2850.535 73.725 ;
        RECT 2851.610 73.680 2851.930 73.740 ;
        RECT 2850.245 73.540 2851.930 73.680 ;
        RECT 2850.245 73.495 2850.535 73.540 ;
        RECT 2851.610 73.480 2851.930 73.540 ;
        RECT 5.590 64.160 5.910 64.220 ;
        RECT 9.730 64.160 10.050 64.220 ;
        RECT 5.590 64.020 10.050 64.160 ;
        RECT 5.590 63.960 5.910 64.020 ;
        RECT 9.730 63.960 10.050 64.020 ;
        RECT 7.890 43.760 8.210 43.820 ;
        RECT 9.745 43.760 10.035 43.805 ;
        RECT 7.890 43.620 10.035 43.760 ;
        RECT 7.890 43.560 8.210 43.620 ;
        RECT 9.745 43.575 10.035 43.620 ;
        RECT 2849.770 43.080 2850.090 43.140 ;
        RECT 2851.610 43.080 2851.930 43.140 ;
        RECT 2849.770 42.940 2851.930 43.080 ;
        RECT 2849.770 42.880 2850.090 42.940 ;
        RECT 2851.610 42.880 2851.930 42.940 ;
        RECT 2845.170 9.080 2845.490 9.140 ;
        RECT 2846.090 9.080 2846.410 9.140 ;
        RECT 2845.170 8.940 2846.410 9.080 ;
        RECT 2845.170 8.880 2845.490 8.940 ;
        RECT 2846.090 8.880 2846.410 8.940 ;
        RECT 110.470 8.740 110.790 8.800 ;
        RECT 51.220 8.600 110.790 8.740 ;
        RECT 9.745 8.060 10.035 8.105 ;
        RECT 51.220 8.060 51.360 8.600 ;
        RECT 110.470 8.540 110.790 8.600 ;
        RECT 176.725 8.740 177.015 8.785 ;
        RECT 245.265 8.740 245.555 8.785 ;
        RECT 253.070 8.740 253.390 8.800 ;
        RECT 176.725 8.600 228.460 8.740 ;
        RECT 176.725 8.555 177.015 8.600 ;
        RECT 228.320 8.400 228.460 8.600 ;
        RECT 245.265 8.600 253.390 8.740 ;
        RECT 245.265 8.555 245.555 8.600 ;
        RECT 253.070 8.540 253.390 8.600 ;
        RECT 889.250 8.740 889.570 8.800 ;
        RECT 918.690 8.740 919.010 8.800 ;
        RECT 951.365 8.740 951.655 8.785 ;
        RECT 889.250 8.600 893.620 8.740 ;
        RECT 889.250 8.540 889.570 8.600 ;
        RECT 278.845 8.400 279.135 8.445 ;
        RECT 228.320 8.260 279.135 8.400 ;
        RECT 893.480 8.400 893.620 8.600 ;
        RECT 918.690 8.600 951.655 8.740 ;
        RECT 918.690 8.540 919.010 8.600 ;
        RECT 951.365 8.555 951.655 8.600 ;
        RECT 956.425 8.740 956.715 8.785 ;
        RECT 958.265 8.740 958.555 8.785 ;
        RECT 956.425 8.600 958.555 8.740 ;
        RECT 956.425 8.555 956.715 8.600 ;
        RECT 958.265 8.555 958.555 8.600 ;
        RECT 984.485 8.740 984.775 8.785 ;
        RECT 985.865 8.740 986.155 8.785 ;
        RECT 984.485 8.600 986.155 8.740 ;
        RECT 984.485 8.555 984.775 8.600 ;
        RECT 985.865 8.555 986.155 8.600 ;
        RECT 2795.490 8.740 2795.810 8.800 ;
        RECT 2836.430 8.740 2836.750 8.800 ;
        RECT 2841.490 8.740 2841.810 8.800 ;
        RECT 2795.490 8.600 2836.750 8.740 ;
        RECT 2841.295 8.600 2841.810 8.740 ;
        RECT 2795.490 8.540 2795.810 8.600 ;
        RECT 2836.430 8.540 2836.750 8.600 ;
        RECT 2841.490 8.540 2841.810 8.600 ;
        RECT 895.230 8.400 895.550 8.460 ;
        RECT 893.480 8.260 895.550 8.400 ;
        RECT 278.845 8.215 279.135 8.260 ;
        RECT 895.230 8.200 895.550 8.260 ;
        RECT 1599.045 8.400 1599.335 8.445 ;
        RECT 1728.765 8.400 1729.055 8.445 ;
        RECT 1599.045 8.260 1729.055 8.400 ;
        RECT 1599.045 8.215 1599.335 8.260 ;
        RECT 1728.765 8.215 1729.055 8.260 ;
        RECT 9.745 7.920 51.360 8.060 ;
        RECT 1070.950 8.060 1071.270 8.120 ;
        RECT 1071.885 8.060 1072.175 8.105 ;
        RECT 1070.950 7.920 1072.175 8.060 ;
        RECT 9.745 7.875 10.035 7.920 ;
        RECT 1070.950 7.860 1071.270 7.920 ;
        RECT 1071.885 7.875 1072.175 7.920 ;
        RECT 1074.630 8.060 1074.950 8.120 ;
        RECT 1082.910 8.060 1083.230 8.120 ;
        RECT 1074.630 7.920 1083.230 8.060 ;
        RECT 1074.630 7.860 1074.950 7.920 ;
        RECT 1082.910 7.860 1083.230 7.920 ;
        RECT 2841.490 8.060 2841.810 8.120 ;
        RECT 2843.330 8.060 2843.650 8.120 ;
        RECT 2841.490 7.920 2843.650 8.060 ;
        RECT 2841.490 7.860 2841.810 7.920 ;
        RECT 2843.330 7.860 2843.650 7.920 ;
        RECT 227.310 7.720 227.630 7.780 ;
        RECT 243.885 7.720 244.175 7.765 ;
        RECT 1023.110 7.720 1023.430 7.780 ;
        RECT 227.310 7.580 244.175 7.720 ;
        RECT 227.310 7.520 227.630 7.580 ;
        RECT 243.885 7.535 244.175 7.580 ;
        RECT 1014.920 7.580 1023.430 7.720 ;
        RECT 846.485 7.380 846.775 7.425 ;
        RECT 824.020 7.240 846.775 7.380 ;
        RECT 129.805 7.040 130.095 7.085 ;
        RECT 65.480 6.900 130.095 7.040 ;
        RECT 52.970 6.700 53.290 6.760 ;
        RECT 65.480 6.700 65.620 6.900 ;
        RECT 129.805 6.855 130.095 6.900 ;
        RECT 696.050 7.040 696.370 7.100 ;
        RECT 701.570 7.040 701.890 7.100 ;
        RECT 696.050 6.900 701.890 7.040 ;
        RECT 696.050 6.840 696.370 6.900 ;
        RECT 701.570 6.840 701.890 6.900 ;
        RECT 757.245 7.040 757.535 7.085 ;
        RECT 763.685 7.040 763.975 7.085 ;
        RECT 757.245 6.900 763.975 7.040 ;
        RECT 757.245 6.855 757.535 6.900 ;
        RECT 763.685 6.855 763.975 6.900 ;
        RECT 810.605 7.040 810.895 7.085 ;
        RECT 814.270 7.040 814.590 7.100 ;
        RECT 824.020 7.085 824.160 7.240 ;
        RECT 846.485 7.195 846.775 7.240 ;
        RECT 956.885 7.380 957.175 7.425 ;
        RECT 957.805 7.380 958.095 7.425 ;
        RECT 956.885 7.240 958.095 7.380 ;
        RECT 956.885 7.195 957.175 7.240 ;
        RECT 957.805 7.195 958.095 7.240 ;
        RECT 1004.265 7.380 1004.555 7.425 ;
        RECT 1014.920 7.380 1015.060 7.580 ;
        RECT 1023.110 7.520 1023.430 7.580 ;
        RECT 1594.905 7.720 1595.195 7.765 ;
        RECT 1596.745 7.720 1597.035 7.765 ;
        RECT 1594.905 7.580 1597.035 7.720 ;
        RECT 1594.905 7.535 1595.195 7.580 ;
        RECT 1596.745 7.535 1597.035 7.580 ;
        RECT 2842.410 7.720 2842.730 7.780 ;
        RECT 2843.790 7.720 2844.110 7.780 ;
        RECT 2842.410 7.580 2844.110 7.720 ;
        RECT 2842.410 7.520 2842.730 7.580 ;
        RECT 2843.790 7.520 2844.110 7.580 ;
        RECT 1004.265 7.240 1015.060 7.380 ;
        RECT 1476.670 7.380 1476.990 7.440 ;
        RECT 1483.585 7.380 1483.875 7.425 ;
        RECT 1476.670 7.240 1483.875 7.380 ;
        RECT 1004.265 7.195 1004.555 7.240 ;
        RECT 1476.670 7.180 1476.990 7.240 ;
        RECT 1483.585 7.195 1483.875 7.240 ;
        RECT 1484.030 7.380 1484.350 7.440 ;
        RECT 1499.670 7.380 1499.990 7.440 ;
        RECT 1484.030 7.240 1499.990 7.380 ;
        RECT 1484.030 7.180 1484.350 7.240 ;
        RECT 1499.670 7.180 1499.990 7.240 ;
        RECT 2777.105 7.380 2777.395 7.425 ;
        RECT 2801.025 7.380 2801.315 7.425 ;
        RECT 2777.105 7.240 2801.315 7.380 ;
        RECT 2777.105 7.195 2777.395 7.240 ;
        RECT 2801.025 7.195 2801.315 7.240 ;
        RECT 810.605 6.900 814.590 7.040 ;
        RECT 810.605 6.855 810.895 6.900 ;
        RECT 814.270 6.840 814.590 6.900 ;
        RECT 823.945 6.855 824.235 7.085 ;
        RECT 884.205 7.040 884.495 7.085 ;
        RECT 887.410 7.040 887.730 7.100 ;
        RECT 884.205 6.900 887.730 7.040 ;
        RECT 884.205 6.855 884.495 6.900 ;
        RECT 887.410 6.840 887.730 6.900 ;
        RECT 1088.905 7.040 1089.195 7.085 ;
        RECT 1090.270 7.040 1090.590 7.100 ;
        RECT 1088.905 6.900 1090.590 7.040 ;
        RECT 1088.905 6.855 1089.195 6.900 ;
        RECT 1090.270 6.840 1090.590 6.900 ;
        RECT 1091.665 7.040 1091.955 7.085 ;
        RECT 1092.110 7.040 1092.430 7.100 ;
        RECT 1091.665 6.900 1092.430 7.040 ;
        RECT 1091.665 6.855 1091.955 6.900 ;
        RECT 1092.110 6.840 1092.430 6.900 ;
        RECT 52.970 6.560 65.620 6.700 ;
        RECT 435.245 6.700 435.535 6.745 ;
        RECT 438.005 6.700 438.295 6.745 ;
        RECT 435.245 6.560 438.295 6.700 ;
        RECT 52.970 6.500 53.290 6.560 ;
        RECT 435.245 6.515 435.535 6.560 ;
        RECT 438.005 6.515 438.295 6.560 ;
        RECT 465.605 6.700 465.895 6.745 ;
        RECT 509.305 6.700 509.595 6.745 ;
        RECT 659.725 6.700 660.015 6.745 ;
        RECT 751.250 6.700 751.570 6.760 ;
        RECT 465.605 6.560 509.595 6.700 ;
        RECT 465.605 6.515 465.895 6.560 ;
        RECT 509.305 6.515 509.595 6.560 ;
        RECT 511.680 6.560 607.960 6.700 ;
        RECT 15.710 6.360 16.030 6.420 ;
        RECT 25.385 6.360 25.675 6.405 ;
        RECT 15.710 6.220 25.675 6.360 ;
        RECT 15.710 6.160 16.030 6.220 ;
        RECT 25.385 6.175 25.675 6.220 ;
        RECT 26.305 6.360 26.595 6.405 ;
        RECT 44.230 6.360 44.550 6.420 ;
        RECT 26.305 6.220 44.550 6.360 ;
        RECT 26.305 6.175 26.595 6.220 ;
        RECT 44.230 6.160 44.550 6.220 ;
        RECT 393.830 6.360 394.150 6.420 ;
        RECT 411.770 6.360 412.090 6.420 ;
        RECT 393.830 6.220 412.090 6.360 ;
        RECT 393.830 6.160 394.150 6.220 ;
        RECT 411.770 6.160 412.090 6.220 ;
        RECT 510.225 6.360 510.515 6.405 ;
        RECT 511.680 6.360 511.820 6.560 ;
        RECT 510.225 6.220 511.820 6.360 ;
        RECT 605.445 6.360 605.735 6.405 ;
        RECT 606.810 6.360 607.130 6.420 ;
        RECT 605.445 6.220 607.130 6.360 ;
        RECT 607.820 6.360 607.960 6.560 ;
        RECT 609.660 6.560 640.620 6.700 ;
        RECT 609.660 6.360 609.800 6.560 ;
        RECT 640.480 6.405 640.620 6.560 ;
        RECT 659.725 6.560 751.570 6.700 ;
        RECT 659.725 6.515 660.015 6.560 ;
        RECT 751.250 6.500 751.570 6.560 ;
        RECT 759.530 6.700 759.850 6.760 ;
        RECT 878.685 6.700 878.975 6.745 ;
        RECT 759.530 6.560 761.140 6.700 ;
        RECT 759.530 6.500 759.850 6.560 ;
        RECT 607.820 6.220 609.800 6.360 ;
        RECT 510.225 6.175 510.515 6.220 ;
        RECT 605.445 6.175 605.735 6.220 ;
        RECT 606.810 6.160 607.130 6.220 ;
        RECT 640.405 6.175 640.695 6.405 ;
        RECT 644.085 6.360 644.375 6.405 ;
        RECT 645.925 6.360 646.215 6.405 ;
        RECT 644.085 6.220 646.215 6.360 ;
        RECT 644.085 6.175 644.375 6.220 ;
        RECT 645.925 6.175 646.215 6.220 ;
        RECT 673.970 6.360 674.290 6.420 ;
        RECT 676.745 6.360 677.035 6.405 ;
        RECT 673.970 6.220 677.035 6.360 ;
        RECT 761.000 6.360 761.140 6.560 ;
        RECT 762.380 6.560 878.975 6.700 ;
        RECT 762.380 6.360 762.520 6.560 ;
        RECT 878.685 6.515 878.975 6.560 ;
        RECT 879.605 6.700 879.895 6.745 ;
        RECT 955.505 6.700 955.795 6.745 ;
        RECT 956.885 6.700 957.175 6.745 ;
        RECT 879.605 6.560 949.740 6.700 ;
        RECT 879.605 6.515 879.895 6.560 ;
        RECT 761.000 6.220 762.520 6.360 ;
        RECT 763.685 6.360 763.975 6.405 ;
        RECT 765.065 6.360 765.355 6.405 ;
        RECT 766.445 6.360 766.735 6.405 ;
        RECT 763.685 6.220 764.820 6.360 ;
        RECT 673.970 6.160 674.290 6.220 ;
        RECT 676.745 6.175 677.035 6.220 ;
        RECT 763.685 6.175 763.975 6.220 ;
        RECT 424.650 6.020 424.970 6.080 ;
        RECT 428.805 6.020 429.095 6.065 ;
        RECT 424.650 5.880 429.095 6.020 ;
        RECT 424.650 5.820 424.970 5.880 ;
        RECT 428.805 5.835 429.095 5.880 ;
        RECT 458.705 6.020 458.995 6.065 ;
        RECT 460.545 6.020 460.835 6.065 ;
        RECT 458.705 5.880 460.835 6.020 ;
        RECT 458.705 5.835 458.995 5.880 ;
        RECT 460.545 5.835 460.835 5.880 ;
        RECT 532.750 6.020 533.070 6.080 ;
        RECT 552.530 6.020 552.850 6.080 ;
        RECT 532.750 5.880 552.850 6.020 ;
        RECT 532.750 5.820 533.070 5.880 ;
        RECT 552.530 5.820 552.850 5.880 ;
        RECT 696.985 6.020 697.275 6.065 ;
        RECT 697.430 6.020 697.750 6.080 ;
        RECT 696.985 5.880 697.750 6.020 ;
        RECT 696.985 5.835 697.275 5.880 ;
        RECT 697.430 5.820 697.750 5.880 ;
        RECT 616.010 5.680 616.330 5.740 ;
        RECT 673.970 5.680 674.290 5.740 ;
        RECT 616.010 5.540 674.290 5.680 ;
        RECT 616.010 5.480 616.330 5.540 ;
        RECT 673.970 5.480 674.290 5.540 ;
        RECT 711.690 5.680 712.010 5.740 ;
        RECT 737.910 5.680 738.230 5.740 ;
        RECT 711.690 5.540 738.230 5.680 ;
        RECT 711.690 5.480 712.010 5.540 ;
        RECT 737.910 5.480 738.230 5.540 ;
        RECT 750.345 5.680 750.635 5.725 ;
        RECT 757.245 5.680 757.535 5.725 ;
        RECT 750.345 5.540 757.535 5.680 ;
        RECT 764.680 5.680 764.820 6.220 ;
        RECT 765.065 6.220 766.735 6.360 ;
        RECT 765.065 6.175 765.355 6.220 ;
        RECT 766.445 6.175 766.735 6.220 ;
        RECT 811.985 6.360 812.275 6.405 ;
        RECT 817.965 6.360 818.255 6.405 ;
        RECT 811.985 6.220 818.255 6.360 ;
        RECT 811.985 6.175 812.275 6.220 ;
        RECT 817.965 6.175 818.255 6.220 ;
        RECT 818.410 6.360 818.730 6.420 ;
        RECT 849.690 6.360 850.010 6.420 ;
        RECT 818.410 6.220 850.010 6.360 ;
        RECT 949.600 6.360 949.740 6.560 ;
        RECT 955.505 6.560 957.175 6.700 ;
        RECT 955.505 6.515 955.795 6.560 ;
        RECT 956.885 6.515 957.175 6.560 ;
        RECT 1001.965 6.700 1002.255 6.745 ;
        RECT 1014.385 6.700 1014.675 6.745 ;
        RECT 1001.965 6.560 1014.675 6.700 ;
        RECT 1001.965 6.515 1002.255 6.560 ;
        RECT 1014.385 6.515 1014.675 6.560 ;
        RECT 1072.345 6.700 1072.635 6.745 ;
        RECT 1073.710 6.700 1074.030 6.760 ;
        RECT 1072.345 6.560 1074.030 6.700 ;
        RECT 1072.345 6.515 1072.635 6.560 ;
        RECT 1073.710 6.500 1074.030 6.560 ;
        RECT 1093.045 6.700 1093.335 6.745 ;
        RECT 1127.530 6.700 1127.850 6.760 ;
        RECT 1140.885 6.700 1141.175 6.745 ;
        RECT 1093.045 6.560 1122.700 6.700 ;
        RECT 1093.045 6.515 1093.335 6.560 ;
        RECT 953.665 6.360 953.955 6.405 ;
        RECT 949.600 6.220 953.955 6.360 ;
        RECT 1122.560 6.360 1122.700 6.560 ;
        RECT 1127.530 6.560 1141.175 6.700 ;
        RECT 1127.530 6.500 1127.850 6.560 ;
        RECT 1140.885 6.515 1141.175 6.560 ;
        RECT 1141.345 6.700 1141.635 6.745 ;
        RECT 1951.865 6.700 1952.155 6.745 ;
        RECT 1141.345 6.560 1952.155 6.700 ;
        RECT 1141.345 6.515 1141.635 6.560 ;
        RECT 1951.865 6.515 1952.155 6.560 ;
        RECT 1953.705 6.700 1953.995 6.745 ;
        RECT 2801.025 6.700 2801.315 6.745 ;
        RECT 2841.490 6.700 2841.810 6.760 ;
        RECT 1953.705 6.560 2746.960 6.700 ;
        RECT 1953.705 6.515 1953.995 6.560 ;
        RECT 1162.030 6.360 1162.350 6.420 ;
        RECT 1165.250 6.360 1165.570 6.420 ;
        RECT 1122.560 6.220 1124.540 6.360 ;
        RECT 818.410 6.160 818.730 6.220 ;
        RECT 849.690 6.160 850.010 6.220 ;
        RECT 953.665 6.175 953.955 6.220 ;
        RECT 1124.400 6.020 1124.540 6.220 ;
        RECT 1162.030 6.220 1165.570 6.360 ;
        RECT 1162.030 6.160 1162.350 6.220 ;
        RECT 1165.250 6.160 1165.570 6.220 ;
        RECT 1199.290 6.360 1199.610 6.420 ;
        RECT 1206.190 6.360 1206.510 6.420 ;
        RECT 1199.290 6.220 1206.510 6.360 ;
        RECT 1199.290 6.160 1199.610 6.220 ;
        RECT 1206.190 6.160 1206.510 6.220 ;
        RECT 1283.010 6.360 1283.330 6.420 ;
        RECT 1301.870 6.360 1302.190 6.420 ;
        RECT 1283.010 6.220 1302.190 6.360 ;
        RECT 1283.010 6.160 1283.330 6.220 ;
        RECT 1301.870 6.160 1302.190 6.220 ;
        RECT 1484.045 6.360 1484.335 6.405 ;
        RECT 1489.565 6.360 1489.855 6.405 ;
        RECT 1484.045 6.220 1489.855 6.360 ;
        RECT 1484.045 6.175 1484.335 6.220 ;
        RECT 1489.565 6.175 1489.855 6.220 ;
        RECT 1637.670 6.360 1637.990 6.420 ;
        RECT 1648.250 6.360 1648.570 6.420 ;
        RECT 1637.670 6.220 1648.570 6.360 ;
        RECT 2746.820 6.360 2746.960 6.560 ;
        RECT 2801.025 6.560 2841.810 6.700 ;
        RECT 2801.025 6.515 2801.315 6.560 ;
        RECT 2841.490 6.500 2841.810 6.560 ;
        RECT 2777.105 6.360 2777.395 6.405 ;
        RECT 2746.820 6.220 2777.395 6.360 ;
        RECT 1637.670 6.160 1637.990 6.220 ;
        RECT 1648.250 6.160 1648.570 6.220 ;
        RECT 2777.105 6.175 2777.395 6.220 ;
        RECT 1141.345 6.020 1141.635 6.065 ;
        RECT 1124.400 5.880 1141.635 6.020 ;
        RECT 1141.345 5.835 1141.635 5.880 ;
        RECT 1490.485 6.020 1490.775 6.065 ;
        RECT 1503.350 6.020 1503.670 6.080 ;
        RECT 1490.485 5.880 1503.670 6.020 ;
        RECT 1490.485 5.835 1490.775 5.880 ;
        RECT 1503.350 5.820 1503.670 5.880 ;
        RECT 1780.745 6.020 1781.035 6.065 ;
        RECT 1784.870 6.020 1785.190 6.080 ;
        RECT 1780.745 5.880 1785.190 6.020 ;
        RECT 1780.745 5.835 1781.035 5.880 ;
        RECT 1784.870 5.820 1785.190 5.880 ;
        RECT 766.905 5.680 767.195 5.725 ;
        RECT 764.680 5.540 767.195 5.680 ;
        RECT 750.345 5.495 750.635 5.540 ;
        RECT 757.245 5.495 757.535 5.540 ;
        RECT 766.905 5.495 767.195 5.540 ;
        RECT 768.745 5.680 769.035 5.725 ;
        RECT 770.125 5.680 770.415 5.725 ;
        RECT 1127.530 5.680 1127.850 5.740 ;
        RECT 768.745 5.540 770.415 5.680 ;
        RECT 1127.335 5.540 1127.850 5.680 ;
        RECT 768.745 5.495 769.035 5.540 ;
        RECT 770.125 5.495 770.415 5.540 ;
        RECT 1127.530 5.480 1127.850 5.540 ;
        RECT 1158.825 5.680 1159.115 5.725 ;
        RECT 1236.565 5.680 1236.855 5.725 ;
        RECT 1158.825 5.540 1236.855 5.680 ;
        RECT 1158.825 5.495 1159.115 5.540 ;
        RECT 1236.565 5.495 1236.855 5.540 ;
        RECT 1237.945 5.680 1238.235 5.725 ;
        RECT 1953.245 5.680 1953.535 5.725 ;
        RECT 1237.945 5.540 1953.535 5.680 ;
        RECT 1237.945 5.495 1238.235 5.540 ;
        RECT 1953.245 5.495 1953.535 5.540 ;
        RECT 1954.165 5.680 1954.455 5.725 ;
        RECT 2469.365 5.680 2469.655 5.725 ;
        RECT 2608.285 5.680 2608.575 5.725 ;
        RECT 1954.165 5.540 2469.655 5.680 ;
        RECT 1954.165 5.495 1954.455 5.540 ;
        RECT 2469.365 5.495 2469.655 5.540 ;
        RECT 2471.280 5.540 2608.575 5.680 ;
        RECT 2470.285 5.340 2470.575 5.385 ;
        RECT 2471.280 5.340 2471.420 5.540 ;
        RECT 2608.285 5.495 2608.575 5.540 ;
        RECT 2608.745 5.680 2609.035 5.725 ;
        RECT 2691.085 5.680 2691.375 5.725 ;
        RECT 2608.745 5.540 2691.375 5.680 ;
        RECT 2608.745 5.495 2609.035 5.540 ;
        RECT 2691.085 5.495 2691.375 5.540 ;
        RECT 2715.465 5.680 2715.755 5.725 ;
        RECT 2746.285 5.680 2746.575 5.725 ;
        RECT 2715.465 5.540 2746.575 5.680 ;
        RECT 2715.465 5.495 2715.755 5.540 ;
        RECT 2746.285 5.495 2746.575 5.540 ;
        RECT 2746.745 5.680 2747.035 5.725 ;
        RECT 2797.345 5.680 2797.635 5.725 ;
        RECT 2746.745 5.540 2797.635 5.680 ;
        RECT 2746.745 5.495 2747.035 5.540 ;
        RECT 2797.345 5.495 2797.635 5.540 ;
        RECT 2470.285 5.200 2471.420 5.340 ;
        RECT 2470.285 5.155 2470.575 5.200 ;
        RECT 129.805 5.000 130.095 5.045 ;
        RECT 176.725 5.000 177.015 5.045 ;
        RECT 658.330 5.000 658.650 5.060 ;
        RECT 129.805 4.860 177.015 5.000 ;
        RECT 129.805 4.815 130.095 4.860 ;
        RECT 176.725 4.815 177.015 4.860 ;
        RECT 645.080 4.860 658.650 5.000 ;
        RECT 284.365 4.660 284.655 4.705 ;
        RECT 289.885 4.660 290.175 4.705 ;
        RECT 284.365 4.520 290.175 4.660 ;
        RECT 284.365 4.475 284.655 4.520 ;
        RECT 289.885 4.475 290.175 4.520 ;
        RECT 377.745 4.660 378.035 4.705 ;
        RECT 382.330 4.660 382.650 4.720 ;
        RECT 377.745 4.520 382.650 4.660 ;
        RECT 377.745 4.475 378.035 4.520 ;
        RECT 382.330 4.460 382.650 4.520 ;
        RECT 514.365 4.660 514.655 4.705 ;
        RECT 582.890 4.660 583.210 4.720 ;
        RECT 514.365 4.520 583.210 4.660 ;
        RECT 514.365 4.475 514.655 4.520 ;
        RECT 582.890 4.460 583.210 4.520 ;
        RECT 617.850 4.660 618.170 4.720 ;
        RECT 645.080 4.660 645.220 4.860 ;
        RECT 658.330 4.800 658.650 4.860 ;
        RECT 1534.630 5.000 1534.950 5.060 ;
        RECT 1593.050 5.000 1593.370 5.060 ;
        RECT 1534.630 4.860 1593.370 5.000 ;
        RECT 1534.630 4.800 1534.950 4.860 ;
        RECT 1593.050 4.800 1593.370 4.860 ;
        RECT 1658.830 5.000 1659.150 5.060 ;
        RECT 1678.610 5.000 1678.930 5.060 ;
        RECT 1658.830 4.860 1678.930 5.000 ;
        RECT 1658.830 4.800 1659.150 4.860 ;
        RECT 1678.610 4.800 1678.930 4.860 ;
        RECT 1728.765 5.000 1729.055 5.045 ;
        RECT 1863.545 5.000 1863.835 5.045 ;
        RECT 1728.765 4.860 1863.835 5.000 ;
        RECT 1728.765 4.815 1729.055 4.860 ;
        RECT 1863.545 4.815 1863.835 4.860 ;
        RECT 1865.385 5.000 1865.675 5.045 ;
        RECT 2841.030 5.000 2841.350 5.060 ;
        RECT 1865.385 4.860 2841.350 5.000 ;
        RECT 1865.385 4.815 1865.675 4.860 ;
        RECT 2841.030 4.800 2841.350 4.860 ;
        RECT 617.850 4.520 645.220 4.660 ;
        RECT 646.385 4.660 646.675 4.705 ;
        RECT 647.290 4.660 647.610 4.720 ;
        RECT 646.385 4.520 647.610 4.660 ;
        RECT 617.850 4.460 618.170 4.520 ;
        RECT 646.385 4.475 646.675 4.520 ;
        RECT 647.290 4.460 647.610 4.520 ;
        RECT 676.745 4.660 677.035 4.705 ;
        RECT 680.425 4.660 680.715 4.705 ;
        RECT 676.745 4.520 680.715 4.660 ;
        RECT 676.745 4.475 677.035 4.520 ;
        RECT 680.425 4.475 680.715 4.520 ;
        RECT 747.570 4.660 747.890 4.720 ;
        RECT 750.345 4.660 750.635 4.705 ;
        RECT 747.570 4.520 750.635 4.660 ;
        RECT 747.570 4.460 747.890 4.520 ;
        RECT 750.345 4.475 750.635 4.520 ;
        RECT 785.765 4.660 786.055 4.705 ;
        RECT 791.745 4.660 792.035 4.705 ;
        RECT 785.765 4.520 792.035 4.660 ;
        RECT 785.765 4.475 786.055 4.520 ;
        RECT 791.745 4.475 792.035 4.520 ;
        RECT 798.185 4.660 798.475 4.705 ;
        RECT 804.165 4.660 804.455 4.705 ;
        RECT 798.185 4.520 804.455 4.660 ;
        RECT 798.185 4.475 798.475 4.520 ;
        RECT 804.165 4.475 804.455 4.520 ;
        RECT 806.005 4.660 806.295 4.705 ;
        RECT 811.985 4.660 812.275 4.705 ;
        RECT 806.005 4.520 812.275 4.660 ;
        RECT 806.005 4.475 806.295 4.520 ;
        RECT 811.985 4.475 812.275 4.520 ;
        RECT 1648.710 4.660 1649.030 4.720 ;
        RECT 1715.410 4.660 1715.730 4.720 ;
        RECT 1648.710 4.520 1715.730 4.660 ;
        RECT 1648.710 4.460 1649.030 4.520 ;
        RECT 1715.410 4.460 1715.730 4.520 ;
        RECT 1747.610 4.660 1747.930 4.720 ;
        RECT 1780.745 4.660 1781.035 4.705 ;
        RECT 1869.510 4.660 1869.830 4.720 ;
        RECT 1747.610 4.520 1781.035 4.660 ;
        RECT 1747.610 4.460 1747.930 4.520 ;
        RECT 1780.745 4.475 1781.035 4.520 ;
        RECT 1864.540 4.520 1869.830 4.660 ;
        RECT 888.790 4.320 889.110 4.380 ;
        RECT 897.990 4.320 898.310 4.380 ;
        RECT 888.790 4.180 898.310 4.320 ;
        RECT 888.790 4.120 889.110 4.180 ;
        RECT 897.990 4.120 898.310 4.180 ;
        RECT 1437.570 4.320 1437.890 4.380 ;
        RECT 1448.150 4.320 1448.470 4.380 ;
        RECT 1437.570 4.180 1448.470 4.320 ;
        RECT 1437.570 4.120 1437.890 4.180 ;
        RECT 1448.150 4.120 1448.470 4.180 ;
        RECT 1864.005 4.320 1864.295 4.365 ;
        RECT 1864.540 4.320 1864.680 4.520 ;
        RECT 1869.510 4.460 1869.830 4.520 ;
        RECT 1900.790 4.660 1901.110 4.720 ;
        RECT 1946.790 4.660 1947.110 4.720 ;
        RECT 1900.790 4.520 1947.110 4.660 ;
        RECT 1900.790 4.460 1901.110 4.520 ;
        RECT 1946.790 4.460 1947.110 4.520 ;
        RECT 2797.345 4.660 2797.635 4.705 ;
        RECT 2847.010 4.660 2847.330 4.720 ;
        RECT 2797.345 4.520 2847.330 4.660 ;
        RECT 2797.345 4.475 2797.635 4.520 ;
        RECT 2847.010 4.460 2847.330 4.520 ;
        RECT 1864.005 4.180 1864.680 4.320 ;
        RECT 2691.085 4.320 2691.375 4.365 ;
        RECT 2715.465 4.320 2715.755 4.365 ;
        RECT 2691.085 4.180 2715.755 4.320 ;
        RECT 1864.005 4.135 1864.295 4.180 ;
        RECT 2691.085 4.135 2691.375 4.180 ;
        RECT 2715.465 4.135 2715.755 4.180 ;
        RECT 465.605 3.980 465.895 4.025 ;
        RECT 502.865 3.980 503.155 4.025 ;
        RECT 465.605 3.840 503.155 3.980 ;
        RECT 465.605 3.795 465.895 3.840 ;
        RECT 502.865 3.795 503.155 3.840 ;
        RECT 511.145 3.980 511.435 4.025 ;
        RECT 534.590 3.980 534.910 4.040 ;
        RECT 511.145 3.840 534.910 3.980 ;
        RECT 511.145 3.795 511.435 3.840 ;
        RECT 534.590 3.780 534.910 3.840 ;
        RECT 771.965 3.980 772.255 4.025 ;
        RECT 784.385 3.980 784.675 4.025 ;
        RECT 771.965 3.840 784.675 3.980 ;
        RECT 771.965 3.795 772.255 3.840 ;
        RECT 784.385 3.795 784.675 3.840 ;
        RECT 1192.390 3.980 1192.710 4.040 ;
        RECT 1193.785 3.980 1194.075 4.025 ;
        RECT 1192.390 3.840 1194.075 3.980 ;
        RECT 1192.390 3.780 1192.710 3.840 ;
        RECT 1193.785 3.795 1194.075 3.840 ;
        RECT 1209.425 3.980 1209.715 4.025 ;
        RECT 1573.285 3.980 1573.575 4.025 ;
        RECT 1209.425 3.840 1573.575 3.980 ;
        RECT 1209.425 3.795 1209.715 3.840 ;
        RECT 1573.285 3.795 1573.575 3.840 ;
        RECT 1782.570 3.980 1782.890 4.040 ;
        RECT 1862.165 3.980 1862.455 4.025 ;
        RECT 1782.570 3.840 1862.455 3.980 ;
        RECT 1782.570 3.780 1782.890 3.840 ;
        RECT 1862.165 3.795 1862.455 3.840 ;
        RECT 1862.610 3.980 1862.930 4.040 ;
        RECT 1931.625 3.980 1931.915 4.025 ;
        RECT 1862.610 3.840 1931.915 3.980 ;
        RECT 1862.610 3.780 1862.930 3.840 ;
        RECT 1931.625 3.795 1931.915 3.840 ;
        RECT 2056.270 3.980 2056.590 4.040 ;
        RECT 2128.490 3.980 2128.810 4.040 ;
        RECT 2056.270 3.840 2128.810 3.980 ;
        RECT 2056.270 3.780 2056.590 3.840 ;
        RECT 2128.490 3.780 2128.810 3.840 ;
        RECT 2153.805 3.980 2154.095 4.025 ;
        RECT 2180.485 3.980 2180.775 4.025 ;
        RECT 2153.805 3.840 2180.775 3.980 ;
        RECT 2153.805 3.795 2154.095 3.840 ;
        RECT 2180.485 3.795 2180.775 3.840 ;
        RECT 2383.790 3.980 2384.110 4.040 ;
        RECT 2430.710 3.980 2431.030 4.040 ;
        RECT 2383.790 3.840 2431.030 3.980 ;
        RECT 2383.790 3.780 2384.110 3.840 ;
        RECT 2430.710 3.780 2431.030 3.840 ;
        RECT 419.130 3.640 419.450 3.700 ;
        RECT 457.785 3.640 458.075 3.685 ;
        RECT 419.130 3.500 458.075 3.640 ;
        RECT 419.130 3.440 419.450 3.500 ;
        RECT 457.785 3.455 458.075 3.500 ;
        RECT 848.310 3.640 848.630 3.700 ;
        RECT 849.705 3.640 849.995 3.685 ;
        RECT 848.310 3.500 849.995 3.640 ;
        RECT 848.310 3.440 848.630 3.500 ;
        RECT 849.705 3.455 849.995 3.500 ;
        RECT 882.825 3.640 883.115 3.685 ;
        RECT 886.505 3.640 886.795 3.685 ;
        RECT 882.825 3.500 886.795 3.640 ;
        RECT 882.825 3.455 883.115 3.500 ;
        RECT 886.505 3.455 886.795 3.500 ;
        RECT 1107.305 3.640 1107.595 3.685 ;
        RECT 1125.245 3.640 1125.535 3.685 ;
        RECT 1107.305 3.500 1125.535 3.640 ;
        RECT 1107.305 3.455 1107.595 3.500 ;
        RECT 1125.245 3.455 1125.535 3.500 ;
        RECT 2174.950 3.640 2175.270 3.700 ;
        RECT 2214.050 3.640 2214.370 3.700 ;
        RECT 2174.950 3.500 2214.370 3.640 ;
        RECT 2174.950 3.440 2175.270 3.500 ;
        RECT 2214.050 3.440 2214.370 3.500 ;
        RECT 133.470 3.300 133.790 3.360 ;
        RECT 196.505 3.300 196.795 3.345 ;
        RECT 133.470 3.160 196.795 3.300 ;
        RECT 133.470 3.100 133.790 3.160 ;
        RECT 196.505 3.115 196.795 3.160 ;
        RECT 366.245 3.300 366.535 3.345 ;
        RECT 377.745 3.300 378.035 3.345 ;
        RECT 751.250 3.300 751.570 3.360 ;
        RECT 366.245 3.160 378.035 3.300 ;
        RECT 751.055 3.160 751.570 3.300 ;
        RECT 366.245 3.115 366.535 3.160 ;
        RECT 377.745 3.115 378.035 3.160 ;
        RECT 751.250 3.100 751.570 3.160 ;
        RECT 887.885 3.300 888.175 3.345 ;
        RECT 889.710 3.300 890.030 3.360 ;
        RECT 887.885 3.160 890.030 3.300 ;
        RECT 887.885 3.115 888.175 3.160 ;
        RECT 889.710 3.100 890.030 3.160 ;
        RECT 917.770 3.300 918.090 3.360 ;
        RECT 918.705 3.300 918.995 3.345 ;
        RECT 917.770 3.160 918.995 3.300 ;
        RECT 917.770 3.100 918.090 3.160 ;
        RECT 918.705 3.115 918.995 3.160 ;
        RECT 1063.605 3.300 1063.895 3.345 ;
        RECT 1070.045 3.300 1070.335 3.345 ;
        RECT 1063.605 3.160 1070.335 3.300 ;
        RECT 1063.605 3.115 1063.895 3.160 ;
        RECT 1070.045 3.115 1070.335 3.160 ;
        RECT 1075.090 3.300 1075.410 3.360 ;
        RECT 1087.970 3.300 1088.290 3.360 ;
        RECT 1075.090 3.160 1088.290 3.300 ;
        RECT 1075.090 3.100 1075.410 3.160 ;
        RECT 1087.970 3.100 1088.290 3.160 ;
        RECT 1098.090 3.300 1098.410 3.360 ;
        RECT 1105.005 3.300 1105.295 3.345 ;
        RECT 1098.090 3.160 1105.295 3.300 ;
        RECT 1098.090 3.100 1098.410 3.160 ;
        RECT 1105.005 3.115 1105.295 3.160 ;
        RECT 1105.450 3.300 1105.770 3.360 ;
        RECT 1120.645 3.300 1120.935 3.345 ;
        RECT 1105.450 3.160 1120.935 3.300 ;
        RECT 1105.450 3.100 1105.770 3.160 ;
        RECT 1120.645 3.115 1120.935 3.160 ;
        RECT 1127.085 3.300 1127.375 3.345 ;
        RECT 1157.430 3.300 1157.750 3.360 ;
        RECT 1127.085 3.160 1157.750 3.300 ;
        RECT 1127.085 3.115 1127.375 3.160 ;
        RECT 1157.430 3.100 1157.750 3.160 ;
        RECT 1158.350 3.300 1158.670 3.360 ;
        RECT 1165.710 3.300 1166.030 3.360 ;
        RECT 1158.350 3.160 1166.030 3.300 ;
        RECT 1158.350 3.100 1158.670 3.160 ;
        RECT 1165.710 3.100 1166.030 3.160 ;
        RECT 1307.850 3.300 1308.170 3.360 ;
        RECT 1334.990 3.300 1335.310 3.360 ;
        RECT 1307.850 3.160 1335.310 3.300 ;
        RECT 1307.850 3.100 1308.170 3.160 ;
        RECT 1334.990 3.100 1335.310 3.160 ;
        RECT 1484.950 3.300 1485.270 3.360 ;
        RECT 1503.350 3.300 1503.670 3.360 ;
        RECT 1484.950 3.160 1503.670 3.300 ;
        RECT 1484.950 3.100 1485.270 3.160 ;
        RECT 1503.350 3.100 1503.670 3.160 ;
        RECT 491.365 2.960 491.655 3.005 ;
        RECT 511.605 2.960 511.895 3.005 ;
        RECT 491.365 2.820 511.895 2.960 ;
        RECT 491.365 2.775 491.655 2.820 ;
        RECT 511.605 2.775 511.895 2.820 ;
        RECT 2549.390 2.960 2549.710 3.020 ;
        RECT 2584.350 2.960 2584.670 3.020 ;
        RECT 2549.390 2.820 2584.670 2.960 ;
        RECT 2549.390 2.760 2549.710 2.820 ;
        RECT 2584.350 2.760 2584.670 2.820 ;
        RECT 1359.370 2.620 1359.690 2.680 ;
        RECT 1396.630 2.620 1396.950 2.680 ;
        RECT 1359.370 2.480 1396.950 2.620 ;
        RECT 1359.370 2.420 1359.690 2.480 ;
        RECT 1396.630 2.420 1396.950 2.480 ;
        RECT 1450.450 2.620 1450.770 2.680 ;
        RECT 1469.310 2.620 1469.630 2.680 ;
        RECT 1450.450 2.480 1469.630 2.620 ;
        RECT 1450.450 2.420 1450.770 2.480 ;
        RECT 1469.310 2.420 1469.630 2.480 ;
        RECT 1932.545 2.620 1932.835 2.665 ;
        RECT 1967.030 2.620 1967.350 2.680 ;
        RECT 1932.545 2.480 1967.350 2.620 ;
        RECT 1932.545 2.435 1932.835 2.480 ;
        RECT 1967.030 2.420 1967.350 2.480 ;
        RECT 711.690 2.280 712.010 2.340 ;
        RECT 723.650 2.280 723.970 2.340 ;
        RECT 711.690 2.140 723.970 2.280 ;
        RECT 711.690 2.080 712.010 2.140 ;
        RECT 723.650 2.080 723.970 2.140 ;
        RECT 992.290 2.280 992.610 2.340 ;
        RECT 1594.890 2.280 1595.210 2.340 ;
        RECT 1615.130 2.280 1615.450 2.340 ;
        RECT 992.290 2.140 992.805 2.280 ;
        RECT 1594.890 2.140 1615.450 2.280 ;
        RECT 992.290 2.080 992.610 2.140 ;
        RECT 1594.890 2.080 1595.210 2.140 ;
        RECT 1615.130 2.080 1615.450 2.140 ;
        RECT 196.505 1.940 196.795 1.985 ;
        RECT 369.465 1.940 369.755 1.985 ;
        RECT 196.505 1.800 369.755 1.940 ;
        RECT 196.505 1.755 196.795 1.800 ;
        RECT 369.465 1.755 369.755 1.800 ;
        RECT 371.765 1.940 372.055 1.985 ;
        RECT 382.805 1.940 383.095 1.985 ;
        RECT 371.765 1.800 383.095 1.940 ;
        RECT 371.765 1.755 372.055 1.800 ;
        RECT 382.805 1.755 383.095 1.800 ;
        RECT 967.910 1.940 968.230 2.000 ;
        RECT 982.645 1.940 982.935 1.985 ;
        RECT 967.910 1.800 982.935 1.940 ;
        RECT 967.910 1.740 968.230 1.800 ;
        RECT 982.645 1.755 982.935 1.800 ;
        RECT 984.930 1.940 985.250 2.000 ;
        RECT 990.910 1.940 991.230 2.000 ;
        RECT 984.930 1.800 991.230 1.940 ;
        RECT 984.930 1.740 985.250 1.800 ;
        RECT 990.910 1.740 991.230 1.800 ;
        RECT 364.865 1.600 365.155 1.645 ;
        RECT 304.680 1.460 365.155 1.600 ;
        RECT 52.525 1.260 52.815 1.305 ;
        RECT 126.570 1.260 126.890 1.320 ;
        RECT 52.525 1.120 126.890 1.260 ;
        RECT 52.525 1.075 52.815 1.120 ;
        RECT 126.570 1.060 126.890 1.120 ;
        RECT 291.265 1.260 291.555 1.305 ;
        RECT 304.680 1.260 304.820 1.460 ;
        RECT 364.865 1.415 365.155 1.460 ;
        RECT 291.265 1.120 304.820 1.260 ;
        RECT 291.265 1.075 291.555 1.120 ;
        RECT 382.805 0.920 383.095 0.965 ;
        RECT 416.845 0.920 417.135 0.965 ;
        RECT 382.805 0.780 417.135 0.920 ;
        RECT 382.805 0.735 383.095 0.780 ;
        RECT 416.845 0.735 417.135 0.780 ;
        RECT 417.290 0.920 417.610 0.980 ;
        RECT 421.905 0.920 422.195 0.965 ;
        RECT 417.290 0.780 422.195 0.920 ;
        RECT 417.290 0.720 417.610 0.780 ;
        RECT 421.905 0.735 422.195 0.780 ;
        RECT 438.925 0.920 439.215 0.965 ;
        RECT 457.325 0.920 457.615 0.965 ;
        RECT 438.925 0.780 457.615 0.920 ;
        RECT 438.925 0.735 439.215 0.780 ;
        RECT 457.325 0.735 457.615 0.780 ;
        RECT 457.785 0.920 458.075 0.965 ;
        RECT 558.985 0.920 559.275 0.965 ;
        RECT 457.785 0.780 559.275 0.920 ;
        RECT 457.785 0.735 458.075 0.780 ;
        RECT 558.985 0.735 559.275 0.780 ;
        RECT 561.745 0.920 562.035 0.965 ;
        RECT 917.310 0.920 917.630 0.980 ;
        RECT 561.745 0.780 917.630 0.920 ;
        RECT 561.745 0.735 562.035 0.780 ;
        RECT 917.310 0.720 917.630 0.780 ;
        RECT 921.465 0.920 921.755 0.965 ;
        RECT 1676.785 0.920 1677.075 0.965 ;
        RECT 921.465 0.780 1677.075 0.920 ;
        RECT 921.465 0.735 921.755 0.780 ;
        RECT 1676.785 0.735 1677.075 0.780 ;
        RECT 1678.165 0.920 1678.455 0.965 ;
        RECT 1737.505 0.920 1737.795 0.965 ;
        RECT 1678.165 0.780 1737.795 0.920 ;
        RECT 1678.165 0.735 1678.455 0.780 ;
        RECT 1737.505 0.735 1737.795 0.780 ;
        RECT 1738.425 0.920 1738.715 0.965 ;
        RECT 1861.705 0.920 1861.995 0.965 ;
        RECT 1738.425 0.780 1861.995 0.920 ;
        RECT 1738.425 0.735 1738.715 0.780 ;
        RECT 1861.705 0.735 1861.995 0.780 ;
        RECT 1866.305 0.920 1866.595 0.965 ;
        RECT 1883.785 0.920 1884.075 0.965 ;
        RECT 1866.305 0.780 1884.075 0.920 ;
        RECT 1866.305 0.735 1866.595 0.780 ;
        RECT 1883.785 0.735 1884.075 0.780 ;
        RECT 1884.705 0.920 1884.995 0.965 ;
        RECT 2367.245 0.920 2367.535 0.965 ;
        RECT 1884.705 0.780 2367.535 0.920 ;
        RECT 1884.705 0.735 1884.995 0.780 ;
        RECT 2367.245 0.735 2367.535 0.780 ;
        RECT 2368.165 0.920 2368.455 0.965 ;
        RECT 2846.090 0.920 2846.410 0.980 ;
        RECT 2368.165 0.780 2846.410 0.920 ;
        RECT 2368.165 0.735 2368.455 0.780 ;
        RECT 2846.090 0.720 2846.410 0.780 ;
        RECT 49.290 0.580 49.610 0.640 ;
        RECT 52.525 0.580 52.815 0.625 ;
        RECT 49.290 0.440 52.815 0.580 ;
        RECT 49.290 0.380 49.610 0.440 ;
        RECT 52.525 0.395 52.815 0.440 ;
        RECT 276.990 0.580 277.310 0.640 ;
        RECT 460.545 0.580 460.835 0.625 ;
        RECT 276.990 0.440 460.835 0.580 ;
        RECT 276.990 0.380 277.310 0.440 ;
        RECT 460.545 0.395 460.835 0.440 ;
        RECT 462.385 0.580 462.675 0.625 ;
        RECT 917.785 0.580 918.075 0.625 ;
        RECT 920.085 0.580 920.375 0.625 ;
        RECT 1677.705 0.580 1677.995 0.625 ;
        RECT 462.385 0.440 918.075 0.580 ;
        RECT 462.385 0.395 462.675 0.440 ;
        RECT 917.785 0.395 918.075 0.440 ;
        RECT 918.320 0.440 919.380 0.580 ;
        RECT 87.010 0.240 87.330 0.300 ;
        RECT 918.320 0.240 918.460 0.440 ;
        RECT 87.010 0.100 918.460 0.240 ;
        RECT 919.240 0.240 919.380 0.440 ;
        RECT 920.085 0.440 1677.995 0.580 ;
        RECT 920.085 0.395 920.375 0.440 ;
        RECT 1677.705 0.395 1677.995 0.440 ;
        RECT 1678.625 0.580 1678.915 0.625 ;
        RECT 1737.045 0.580 1737.335 0.625 ;
        RECT 1678.625 0.440 1737.335 0.580 ;
        RECT 1678.625 0.395 1678.915 0.440 ;
        RECT 1737.045 0.395 1737.335 0.440 ;
        RECT 1737.965 0.580 1738.255 0.625 ;
        RECT 1862.165 0.580 1862.455 0.625 ;
        RECT 1737.965 0.440 1862.455 0.580 ;
        RECT 1737.965 0.395 1738.255 0.440 ;
        RECT 1862.165 0.395 1862.455 0.440 ;
        RECT 1863.545 0.580 1863.835 0.625 ;
        RECT 2153.805 0.580 2154.095 0.625 ;
        RECT 1863.545 0.440 2154.095 0.580 ;
        RECT 1863.545 0.395 1863.835 0.440 ;
        RECT 2153.805 0.395 2154.095 0.440 ;
        RECT 2180.485 0.580 2180.775 0.625 ;
        RECT 2844.250 0.580 2844.570 0.640 ;
        RECT 2180.485 0.440 2844.570 0.580 ;
        RECT 2180.485 0.395 2180.775 0.440 ;
        RECT 2844.250 0.380 2844.570 0.440 ;
        RECT 1677.245 0.240 1677.535 0.285 ;
        RECT 919.240 0.100 1677.535 0.240 ;
        RECT 87.010 0.040 87.330 0.100 ;
        RECT 1677.245 0.055 1677.535 0.100 ;
        RECT 1678.165 0.240 1678.455 0.285 ;
        RECT 1736.585 0.240 1736.875 0.285 ;
        RECT 1678.165 0.100 1736.875 0.240 ;
        RECT 1678.165 0.055 1678.455 0.100 ;
        RECT 1736.585 0.055 1736.875 0.100 ;
        RECT 1738.425 0.240 1738.715 0.285 ;
        RECT 2366.770 0.240 2367.090 0.300 ;
        RECT 1738.425 0.100 2367.090 0.240 ;
        RECT 1738.425 0.055 1738.715 0.100 ;
        RECT 2366.770 0.040 2367.090 0.100 ;
        RECT 2368.610 0.240 2368.930 0.300 ;
        RECT 2841.505 0.240 2841.795 0.285 ;
        RECT 2368.610 0.100 2841.795 0.240 ;
        RECT 2368.610 0.040 2368.930 0.100 ;
        RECT 2841.505 0.055 2841.795 0.100 ;
      LAYER via ;
        RECT 2019.500 3416.020 2019.760 3416.280 ;
        RECT 2042.040 3416.020 2042.300 3416.280 ;
        RECT 1529.600 3404.800 1529.860 3405.060 ;
        RECT 1638.160 3404.800 1638.420 3405.060 ;
        RECT 1638.160 3401.400 1638.420 3401.660 ;
        RECT 2042.040 3401.400 2042.300 3401.660 ;
        RECT 2773.900 3401.400 2774.160 3401.660 ;
        RECT 2841.980 3398.000 2842.240 3398.260 ;
        RECT 2849.800 3150.820 2850.060 3151.080 ;
        RECT 2863.600 3150.820 2863.860 3151.080 ;
        RECT 2849.800 3048.140 2850.060 3048.400 ;
        RECT 2851.640 3048.140 2851.900 3048.400 ;
        RECT 2849.800 2856.720 2850.060 2856.980 ;
        RECT 2863.600 2856.720 2863.860 2856.980 ;
        RECT 2866.820 2663.600 2867.080 2663.860 ;
        RECT 2900.860 2663.600 2901.120 2663.860 ;
        RECT 2849.800 2611.580 2850.060 2611.840 ;
        RECT 2866.820 2611.580 2867.080 2611.840 ;
        RECT 2849.800 2337.880 2850.060 2338.140 ;
        RECT 2850.260 2335.160 2850.520 2335.420 ;
        RECT 2849.340 2321.220 2849.600 2321.480 ;
        RECT 2850.260 2320.540 2850.520 2320.800 ;
        RECT 2849.800 2319.860 2850.060 2320.120 ;
        RECT 2849.800 2319.180 2850.060 2319.440 ;
        RECT 2849.800 2318.500 2850.060 2318.760 ;
        RECT 2849.800 2308.300 2850.060 2308.560 ;
        RECT 2853.020 2059.760 2853.280 2060.020 ;
        RECT 2863.600 2059.760 2863.860 2060.020 ;
        RECT 2849.800 2008.080 2850.060 2008.340 ;
        RECT 2853.020 2008.080 2853.280 2008.340 ;
        RECT 2849.800 1983.940 2850.060 1984.200 ;
        RECT 2849.800 1974.760 2850.060 1975.020 ;
        RECT 2849.800 1965.580 2850.060 1965.840 ;
        RECT 2849.800 1964.560 2850.060 1964.820 ;
        RECT 2849.800 1963.540 2850.060 1963.800 ;
        RECT 2849.800 1962.860 2850.060 1963.120 ;
        RECT 2851.640 1962.860 2851.900 1963.120 ;
        RECT 2849.800 1961.500 2850.060 1961.760 ;
        RECT 2849.800 1949.940 2850.060 1950.200 ;
        RECT 2849.800 1942.460 2850.060 1942.720 ;
        RECT 2849.800 1846.920 2850.060 1847.180 ;
        RECT 2849.800 1838.760 2850.060 1839.020 ;
        RECT 2849.800 1800.000 2850.060 1800.260 ;
        RECT 2851.640 1800.000 2851.900 1800.260 ;
        RECT 2849.800 1799.320 2850.060 1799.580 ;
        RECT 2849.800 1797.620 2850.060 1797.880 ;
        RECT 2849.800 1795.580 2850.060 1795.840 ;
        RECT 2849.800 1794.220 2850.060 1794.480 ;
        RECT 2849.800 1793.540 2850.060 1793.800 ;
        RECT 2851.180 1793.540 2851.440 1793.800 ;
        RECT 2849.800 1792.860 2850.060 1793.120 ;
        RECT 2849.800 1791.160 2850.060 1791.420 ;
        RECT 2851.180 1790.140 2851.440 1790.400 ;
        RECT 2849.800 1768.720 2850.060 1768.980 ;
        RECT 2851.640 1766.340 2851.900 1766.600 ;
        RECT 2849.340 1766.000 2849.600 1766.260 ;
        RECT 2849.800 1761.580 2850.060 1761.840 ;
        RECT 2849.800 1739.820 2850.060 1740.080 ;
        RECT 2849.800 1647.680 2850.060 1647.940 ;
        RECT 2849.800 1647.000 2850.060 1647.260 ;
        RECT 2849.800 1646.320 2850.060 1646.580 ;
        RECT 2849.800 1638.840 2850.060 1639.100 ;
        RECT 2849.800 1638.160 2850.060 1638.420 ;
        RECT 2863.600 1638.160 2863.860 1638.420 ;
        RECT 2849.800 1635.780 2850.060 1636.040 ;
        RECT 2849.800 1635.100 2850.060 1635.360 ;
        RECT 2849.800 1628.300 2850.060 1628.560 ;
        RECT 2850.720 1627.620 2850.980 1627.880 ;
        RECT 2850.720 1604.840 2850.980 1605.100 ;
        RECT 2849.800 1604.160 2850.060 1604.420 ;
        RECT 2850.260 1579.000 2850.520 1579.260 ;
        RECT 2851.640 1579.000 2851.900 1579.260 ;
        RECT 2849.800 1577.980 2850.060 1578.240 ;
        RECT 2849.800 1545.340 2850.060 1545.600 ;
        RECT 2849.800 1534.800 2850.060 1535.060 ;
        RECT 2849.800 1530.720 2850.060 1530.980 ;
        RECT 2849.800 1513.720 2850.060 1513.980 ;
        RECT 2849.800 1505.560 2850.060 1505.820 ;
        RECT 2849.800 1504.200 2850.060 1504.460 ;
        RECT 2849.800 1500.120 2850.060 1500.380 ;
        RECT 2849.800 1492.640 2850.060 1492.900 ;
        RECT 2849.800 1491.960 2850.060 1492.220 ;
        RECT 2850.260 1480.740 2850.520 1481.000 ;
        RECT 2851.180 1480.060 2851.440 1480.320 ;
        RECT 2849.800 1462.040 2850.060 1462.300 ;
        RECT 2849.800 1448.100 2850.060 1448.360 ;
        RECT 2849.800 1426.680 2850.060 1426.940 ;
        RECT 2849.800 1425.660 2850.060 1425.920 ;
        RECT 2849.800 1424.640 2850.060 1424.900 ;
        RECT 2849.800 1423.960 2850.060 1424.220 ;
        RECT 2849.800 1422.940 2850.060 1423.200 ;
        RECT 2852.560 1422.940 2852.820 1423.200 ;
        RECT 2849.800 1419.200 2850.060 1419.460 ;
        RECT 2849.800 1418.520 2850.060 1418.780 ;
        RECT 2849.800 1417.500 2850.060 1417.760 ;
        RECT 2849.800 1416.820 2850.060 1417.080 ;
        RECT 2850.260 1416.480 2850.520 1416.740 ;
        RECT 2849.800 1389.620 2850.060 1389.880 ;
        RECT 2851.640 1389.620 2851.900 1389.880 ;
        RECT 2849.800 1387.580 2850.060 1387.840 ;
        RECT 2850.720 1387.580 2850.980 1387.840 ;
        RECT 2849.800 1386.220 2850.060 1386.480 ;
        RECT 2849.800 1372.280 2850.060 1372.540 ;
        RECT 2849.800 1370.920 2850.060 1371.180 ;
        RECT 2850.260 1368.540 2850.520 1368.800 ;
        RECT 2849.800 1365.140 2850.060 1365.400 ;
        RECT 2849.800 1364.460 2850.060 1364.720 ;
        RECT 2849.800 1363.780 2850.060 1364.040 ;
        RECT 2863.600 1363.780 2863.860 1364.040 ;
        RECT 2849.800 1362.760 2850.060 1363.020 ;
        RECT 2852.100 1362.760 2852.360 1363.020 ;
        RECT 2849.340 1361.740 2849.600 1362.000 ;
        RECT 2849.800 1357.660 2850.060 1357.920 ;
        RECT 2849.800 1354.940 2850.060 1355.200 ;
        RECT 2849.800 1354.260 2850.060 1354.520 ;
        RECT 2850.720 1354.260 2850.980 1354.520 ;
        RECT 2849.800 1352.900 2850.060 1353.160 ;
        RECT 2851.640 1352.900 2851.900 1353.160 ;
        RECT 2849.800 1352.220 2850.060 1352.480 ;
        RECT 2849.800 1350.180 2850.060 1350.440 ;
        RECT 2849.800 1329.440 2850.060 1329.700 ;
        RECT 2849.800 1258.720 2850.060 1258.980 ;
        RECT 2850.720 1258.720 2850.980 1258.980 ;
        RECT 2849.800 1254.640 2850.060 1254.900 ;
        RECT 2849.800 1253.960 2850.060 1254.220 ;
        RECT 2851.640 1253.960 2851.900 1254.220 ;
        RECT 2849.800 1252.940 2850.060 1253.200 ;
        RECT 2850.260 1232.540 2850.520 1232.800 ;
        RECT 2850.720 1197.180 2850.980 1197.440 ;
        RECT 2849.800 1167.600 2850.060 1167.860 ;
        RECT 2850.720 1167.600 2850.980 1167.860 ;
        RECT 2849.800 1150.940 2850.060 1151.200 ;
        RECT 2849.800 1149.920 2850.060 1150.180 ;
        RECT 2850.720 1149.920 2850.980 1150.180 ;
        RECT 2849.800 1148.900 2850.060 1149.160 ;
        RECT 2851.640 1148.900 2851.900 1149.160 ;
        RECT 2850.720 1148.560 2850.980 1148.820 ;
        RECT 2850.260 1148.220 2850.520 1148.480 ;
        RECT 2849.800 1128.840 2850.060 1129.100 ;
        RECT 2849.800 1078.180 2850.060 1078.440 ;
        RECT 2849.800 1076.820 2850.060 1077.080 ;
        RECT 2849.800 1073.080 2850.060 1073.340 ;
        RECT 2850.720 1072.740 2850.980 1073.000 ;
        RECT 2849.800 1023.780 2850.060 1024.040 ;
        RECT 2849.800 1017.660 2850.060 1017.920 ;
        RECT 2849.800 1014.940 2850.060 1015.200 ;
        RECT 2850.260 959.860 2850.520 960.120 ;
        RECT 2849.800 959.520 2850.060 959.780 ;
        RECT 2849.800 958.500 2850.060 958.760 ;
        RECT 2850.260 958.500 2850.520 958.760 ;
        RECT 2849.800 957.820 2850.060 958.080 ;
        RECT 2851.640 957.820 2851.900 958.080 ;
        RECT 2849.800 957.140 2850.060 957.400 ;
        RECT 2849.800 942.860 2850.060 943.120 ;
        RECT 2851.180 942.860 2851.440 943.120 ;
        RECT 2849.800 874.520 2850.060 874.780 ;
        RECT 2849.800 868.060 2850.060 868.320 ;
        RECT 2850.720 868.060 2850.980 868.320 ;
        RECT 2850.260 859.560 2850.520 859.820 ;
        RECT 2849.800 846.640 2850.060 846.900 ;
        RECT 2849.800 845.620 2850.060 845.880 ;
        RECT 2849.800 844.940 2850.060 845.200 ;
        RECT 2850.720 844.940 2850.980 845.200 ;
        RECT 2849.800 818.420 2850.060 818.680 ;
        RECT 2852.100 810.940 2852.360 811.200 ;
        RECT 2850.720 788.160 2850.980 788.420 ;
        RECT 2849.800 787.480 2850.060 787.740 ;
        RECT 2850.720 787.480 2850.980 787.740 ;
        RECT 2849.800 786.800 2850.060 787.060 ;
        RECT 2849.800 779.320 2850.060 779.580 ;
        RECT 2851.180 778.640 2851.440 778.900 ;
        RECT 2849.800 775.920 2850.060 776.180 ;
        RECT 2849.340 775.580 2849.600 775.840 ;
        RECT 2850.260 775.240 2850.520 775.500 ;
        RECT 2849.800 774.900 2850.060 775.160 ;
        RECT 2849.800 774.220 2850.060 774.480 ;
        RECT 2849.800 769.120 2850.060 769.380 ;
        RECT 2851.180 769.120 2851.440 769.380 ;
        RECT 2851.180 745.320 2851.440 745.580 ;
        RECT 2852.100 745.320 2852.360 745.580 ;
        RECT 2849.800 739.540 2850.060 739.800 ;
        RECT 2849.800 738.860 2850.060 739.120 ;
        RECT 2850.720 738.860 2850.980 739.120 ;
        RECT 2849.800 738.180 2850.060 738.440 ;
        RECT 2849.800 671.540 2850.060 671.800 ;
        RECT 2851.180 671.540 2851.440 671.800 ;
        RECT 2849.800 382.880 2850.060 383.140 ;
        RECT 2849.800 380.840 2850.060 381.100 ;
        RECT 2849.800 374.040 2850.060 374.300 ;
        RECT 2849.800 373.360 2850.060 373.620 ;
        RECT 2851.180 373.360 2851.440 373.620 ;
        RECT 2849.800 368.600 2850.060 368.860 ;
        RECT 2849.800 367.920 2850.060 368.180 ;
        RECT 2849.800 366.900 2850.060 367.160 ;
        RECT 2849.800 366.220 2850.060 366.480 ;
        RECT 2851.180 366.220 2851.440 366.480 ;
        RECT 2849.800 365.540 2850.060 365.800 ;
        RECT 2849.800 364.860 2850.060 365.120 ;
        RECT 2849.800 362.140 2850.060 362.400 ;
        RECT 2849.800 341.740 2850.060 342.000 ;
        RECT 2851.180 341.740 2851.440 342.000 ;
        RECT 2849.800 340.040 2850.060 340.300 ;
        RECT 2850.720 330.520 2850.980 330.780 ;
        RECT 2849.800 308.420 2850.060 308.680 ;
        RECT 2849.800 307.740 2850.060 308.000 ;
        RECT 2850.720 307.740 2850.980 308.000 ;
        RECT 2850.260 306.380 2850.520 306.640 ;
        RECT 2849.800 303.660 2850.060 303.920 ;
        RECT 2849.800 299.580 2850.060 299.840 ;
        RECT 2849.800 284.620 2850.060 284.880 ;
        RECT 2849.800 210.840 2850.060 211.100 ;
        RECT 2849.800 208.120 2850.060 208.380 ;
        RECT 2849.800 205.400 2850.060 205.660 ;
        RECT 2849.800 204.720 2850.060 204.980 ;
        RECT 2849.800 203.360 2850.060 203.620 ;
        RECT 2849.800 202.000 2850.060 202.260 ;
        RECT 2849.800 201.320 2850.060 201.580 ;
        RECT 2849.800 200.640 2850.060 200.900 ;
        RECT 2849.800 199.960 2850.060 200.220 ;
        RECT 2849.800 199.280 2850.060 199.540 ;
        RECT 2849.800 198.260 2850.060 198.520 ;
        RECT 2849.800 196.900 2850.060 197.160 ;
        RECT 2851.640 173.780 2851.900 174.040 ;
        RECT 2849.800 132.300 2850.060 132.560 ;
        RECT 2849.800 128.560 2850.060 128.820 ;
        RECT 2849.800 127.540 2850.060 127.800 ;
        RECT 2849.800 125.500 2850.060 125.760 ;
        RECT 2851.180 125.500 2851.440 125.760 ;
        RECT 2849.800 121.420 2850.060 121.680 ;
        RECT 2851.640 121.420 2851.900 121.680 ;
        RECT 2849.800 120.740 2850.060 121.000 ;
        RECT 2849.800 118.700 2850.060 118.960 ;
        RECT 2849.800 117.680 2850.060 117.940 ;
        RECT 2851.180 117.680 2851.440 117.940 ;
        RECT 2849.800 88.100 2850.060 88.360 ;
        RECT 2851.640 73.480 2851.900 73.740 ;
        RECT 5.620 63.960 5.880 64.220 ;
        RECT 9.760 63.960 10.020 64.220 ;
        RECT 7.920 43.560 8.180 43.820 ;
        RECT 2849.800 42.880 2850.060 43.140 ;
        RECT 2851.640 42.880 2851.900 43.140 ;
        RECT 2845.200 8.880 2845.460 9.140 ;
        RECT 2846.120 8.880 2846.380 9.140 ;
        RECT 110.500 8.540 110.760 8.800 ;
        RECT 253.100 8.540 253.360 8.800 ;
        RECT 889.280 8.540 889.540 8.800 ;
        RECT 918.720 8.540 918.980 8.800 ;
        RECT 2795.520 8.540 2795.780 8.800 ;
        RECT 2836.460 8.540 2836.720 8.800 ;
        RECT 2841.520 8.540 2841.780 8.800 ;
        RECT 895.260 8.200 895.520 8.460 ;
        RECT 1070.980 7.860 1071.240 8.120 ;
        RECT 1074.660 7.860 1074.920 8.120 ;
        RECT 1082.940 7.860 1083.200 8.120 ;
        RECT 2841.520 7.860 2841.780 8.120 ;
        RECT 2843.360 7.860 2843.620 8.120 ;
        RECT 227.340 7.520 227.600 7.780 ;
        RECT 53.000 6.500 53.260 6.760 ;
        RECT 696.080 6.840 696.340 7.100 ;
        RECT 701.600 6.840 701.860 7.100 ;
        RECT 814.300 6.840 814.560 7.100 ;
        RECT 1023.140 7.520 1023.400 7.780 ;
        RECT 2842.440 7.520 2842.700 7.780 ;
        RECT 2843.820 7.520 2844.080 7.780 ;
        RECT 1476.700 7.180 1476.960 7.440 ;
        RECT 1484.060 7.180 1484.320 7.440 ;
        RECT 1499.700 7.180 1499.960 7.440 ;
        RECT 887.440 6.840 887.700 7.100 ;
        RECT 1090.300 6.840 1090.560 7.100 ;
        RECT 1092.140 6.840 1092.400 7.100 ;
        RECT 15.740 6.160 16.000 6.420 ;
        RECT 44.260 6.160 44.520 6.420 ;
        RECT 393.860 6.160 394.120 6.420 ;
        RECT 411.800 6.160 412.060 6.420 ;
        RECT 606.840 6.160 607.100 6.420 ;
        RECT 751.280 6.500 751.540 6.760 ;
        RECT 759.560 6.500 759.820 6.760 ;
        RECT 674.000 6.160 674.260 6.420 ;
        RECT 424.680 5.820 424.940 6.080 ;
        RECT 532.780 5.820 533.040 6.080 ;
        RECT 552.560 5.820 552.820 6.080 ;
        RECT 697.460 5.820 697.720 6.080 ;
        RECT 616.040 5.480 616.300 5.740 ;
        RECT 674.000 5.480 674.260 5.740 ;
        RECT 711.720 5.480 711.980 5.740 ;
        RECT 737.940 5.480 738.200 5.740 ;
        RECT 818.440 6.160 818.700 6.420 ;
        RECT 849.720 6.160 849.980 6.420 ;
        RECT 1073.740 6.500 1074.000 6.760 ;
        RECT 1127.560 6.500 1127.820 6.760 ;
        RECT 1162.060 6.160 1162.320 6.420 ;
        RECT 1165.280 6.160 1165.540 6.420 ;
        RECT 1199.320 6.160 1199.580 6.420 ;
        RECT 1206.220 6.160 1206.480 6.420 ;
        RECT 1283.040 6.160 1283.300 6.420 ;
        RECT 1301.900 6.160 1302.160 6.420 ;
        RECT 1637.700 6.160 1637.960 6.420 ;
        RECT 1648.280 6.160 1648.540 6.420 ;
        RECT 2841.520 6.500 2841.780 6.760 ;
        RECT 1503.380 5.820 1503.640 6.080 ;
        RECT 1784.900 5.820 1785.160 6.080 ;
        RECT 1127.560 5.480 1127.820 5.740 ;
        RECT 382.360 4.460 382.620 4.720 ;
        RECT 582.920 4.460 583.180 4.720 ;
        RECT 617.880 4.460 618.140 4.720 ;
        RECT 658.360 4.800 658.620 5.060 ;
        RECT 1534.660 4.800 1534.920 5.060 ;
        RECT 1593.080 4.800 1593.340 5.060 ;
        RECT 1658.860 4.800 1659.120 5.060 ;
        RECT 1678.640 4.800 1678.900 5.060 ;
        RECT 2841.060 4.800 2841.320 5.060 ;
        RECT 647.320 4.460 647.580 4.720 ;
        RECT 747.600 4.460 747.860 4.720 ;
        RECT 1648.740 4.460 1649.000 4.720 ;
        RECT 1715.440 4.460 1715.700 4.720 ;
        RECT 1747.640 4.460 1747.900 4.720 ;
        RECT 888.820 4.120 889.080 4.380 ;
        RECT 898.020 4.120 898.280 4.380 ;
        RECT 1437.600 4.120 1437.860 4.380 ;
        RECT 1448.180 4.120 1448.440 4.380 ;
        RECT 1869.540 4.460 1869.800 4.720 ;
        RECT 1900.820 4.460 1901.080 4.720 ;
        RECT 1946.820 4.460 1947.080 4.720 ;
        RECT 2847.040 4.460 2847.300 4.720 ;
        RECT 534.620 3.780 534.880 4.040 ;
        RECT 1192.420 3.780 1192.680 4.040 ;
        RECT 1782.600 3.780 1782.860 4.040 ;
        RECT 1862.640 3.780 1862.900 4.040 ;
        RECT 2056.300 3.780 2056.560 4.040 ;
        RECT 2128.520 3.780 2128.780 4.040 ;
        RECT 2383.820 3.780 2384.080 4.040 ;
        RECT 2430.740 3.780 2431.000 4.040 ;
        RECT 419.160 3.440 419.420 3.700 ;
        RECT 848.340 3.440 848.600 3.700 ;
        RECT 2174.980 3.440 2175.240 3.700 ;
        RECT 2214.080 3.440 2214.340 3.700 ;
        RECT 133.500 3.100 133.760 3.360 ;
        RECT 751.280 3.100 751.540 3.360 ;
        RECT 889.740 3.100 890.000 3.360 ;
        RECT 917.800 3.100 918.060 3.360 ;
        RECT 1075.120 3.100 1075.380 3.360 ;
        RECT 1088.000 3.100 1088.260 3.360 ;
        RECT 1098.120 3.100 1098.380 3.360 ;
        RECT 1105.480 3.100 1105.740 3.360 ;
        RECT 1157.460 3.100 1157.720 3.360 ;
        RECT 1158.380 3.100 1158.640 3.360 ;
        RECT 1165.740 3.100 1166.000 3.360 ;
        RECT 1307.880 3.100 1308.140 3.360 ;
        RECT 1335.020 3.100 1335.280 3.360 ;
        RECT 1484.980 3.100 1485.240 3.360 ;
        RECT 1503.380 3.100 1503.640 3.360 ;
        RECT 2549.420 2.760 2549.680 3.020 ;
        RECT 2584.380 2.760 2584.640 3.020 ;
        RECT 1359.400 2.420 1359.660 2.680 ;
        RECT 1396.660 2.420 1396.920 2.680 ;
        RECT 1450.480 2.420 1450.740 2.680 ;
        RECT 1469.340 2.420 1469.600 2.680 ;
        RECT 1967.060 2.420 1967.320 2.680 ;
        RECT 711.720 2.080 711.980 2.340 ;
        RECT 723.680 2.080 723.940 2.340 ;
        RECT 992.320 2.080 992.580 2.340 ;
        RECT 1594.920 2.080 1595.180 2.340 ;
        RECT 1615.160 2.080 1615.420 2.340 ;
        RECT 967.940 1.740 968.200 2.000 ;
        RECT 984.960 1.740 985.220 2.000 ;
        RECT 990.940 1.740 991.200 2.000 ;
        RECT 126.600 1.060 126.860 1.320 ;
        RECT 417.320 0.720 417.580 0.980 ;
        RECT 917.340 0.720 917.600 0.980 ;
        RECT 2846.120 0.720 2846.380 0.980 ;
        RECT 49.320 0.380 49.580 0.640 ;
        RECT 277.020 0.380 277.280 0.640 ;
        RECT 87.040 0.040 87.300 0.300 ;
        RECT 2844.280 0.380 2844.540 0.640 ;
        RECT 2366.800 0.040 2367.060 0.300 ;
        RECT 2368.640 0.040 2368.900 0.300 ;
      LAYER met2 ;
        RECT 2019.500 3415.990 2019.760 3416.310 ;
        RECT 2042.040 3415.990 2042.300 3416.310 ;
        RECT 1527.690 3404.490 1527.970 3405.000 ;
        RECT 1529.600 3404.770 1529.860 3405.090 ;
        RECT 1638.160 3404.770 1638.420 3405.090 ;
        RECT 2019.560 3405.000 2019.700 3415.990 ;
        RECT 1529.660 3404.490 1529.800 3404.770 ;
        RECT 1527.690 3404.350 1529.800 3404.490 ;
        RECT 1527.690 3401.000 1527.970 3404.350 ;
        RECT 1638.220 3401.690 1638.360 3404.770 ;
        RECT 1638.160 3401.370 1638.420 3401.690 ;
        RECT 2019.430 3401.000 2019.710 3405.000 ;
        RECT 2042.100 3401.690 2042.240 3415.990 ;
        RECT 2773.890 3402.195 2774.170 3402.565 ;
        RECT 2773.960 3401.690 2774.100 3402.195 ;
        RECT 2042.040 3401.370 2042.300 3401.690 ;
        RECT 2773.900 3401.370 2774.160 3401.690 ;
        RECT 2841.120 3398.290 2842.180 3398.370 ;
        RECT 2841.120 3398.230 2842.240 3398.290 ;
        RECT 2841.120 3367.090 2841.260 3398.230 ;
        RECT 2841.980 3397.970 2842.240 3398.230 ;
        RECT 2841.120 3366.950 2841.720 3367.090 ;
        RECT 2841.580 3319.490 2841.720 3366.950 ;
        RECT 2841.580 3319.350 2842.640 3319.490 ;
        RECT 2842.500 3295.010 2842.640 3319.350 ;
        RECT 2841.580 3294.870 2842.640 3295.010 ;
        RECT 2841.580 3201.850 2841.720 3294.870 ;
        RECT 2841.580 3201.710 2842.180 3201.850 ;
        RECT 2842.040 3105.290 2842.180 3201.710 ;
        RECT 2863.590 3200.915 2863.870 3201.285 ;
        RECT 2863.660 3151.110 2863.800 3200.915 ;
        RECT 2849.800 3150.850 2850.060 3151.110 ;
        RECT 2841.120 3105.150 2842.180 3105.290 ;
        RECT 2844.340 3150.790 2850.060 3150.850 ;
        RECT 2863.600 3150.790 2863.860 3151.110 ;
        RECT 2844.340 3150.710 2850.000 3150.790 ;
        RECT 2841.120 3067.210 2841.260 3105.150 ;
        RECT 2844.340 3104.610 2844.480 3150.710 ;
        RECT 2843.880 3104.470 2844.480 3104.610 ;
        RECT 2841.120 3067.070 2841.720 3067.210 ;
        RECT 2841.580 3021.650 2841.720 3067.070 ;
        RECT 2843.880 3054.970 2844.020 3104.470 ;
        RECT 2851.630 3062.195 2851.910 3062.565 ;
        RECT 2843.880 3054.830 2844.480 3054.970 ;
        RECT 2844.340 3053.610 2844.480 3054.830 ;
        RECT 2843.880 3053.470 2844.480 3053.610 ;
        RECT 2841.580 3021.510 2843.100 3021.650 ;
        RECT 2842.960 2975.410 2843.100 3021.510 ;
        RECT 2841.580 2975.270 2843.100 2975.410 ;
        RECT 2841.580 2974.730 2841.720 2975.270 ;
        RECT 2841.120 2974.590 2841.720 2974.730 ;
        RECT 2841.120 2944.810 2841.260 2974.590 ;
        RECT 2843.880 2974.050 2844.020 3053.470 ;
        RECT 2851.700 3048.430 2851.840 3062.195 ;
        RECT 2849.800 3048.170 2850.060 3048.430 ;
        RECT 2842.960 2973.910 2844.020 2974.050 ;
        RECT 2847.100 3048.110 2850.060 3048.170 ;
        RECT 2851.640 3048.110 2851.900 3048.430 ;
        RECT 2847.100 3048.030 2850.000 3048.110 ;
        RECT 2842.960 2963.850 2843.100 2973.910 ;
        RECT 2847.100 2963.850 2847.240 3048.030 ;
        RECT 2842.960 2963.710 2844.020 2963.850 ;
        RECT 2847.100 2963.710 2847.700 2963.850 ;
        RECT 2843.880 2945.490 2844.020 2963.710 ;
        RECT 2843.420 2945.350 2844.020 2945.490 ;
        RECT 2841.120 2944.670 2842.180 2944.810 ;
        RECT 2842.040 2922.370 2842.180 2944.670 ;
        RECT 2841.580 2922.230 2842.180 2922.370 ;
        RECT 2841.580 2897.890 2841.720 2922.230 ;
        RECT 2841.120 2897.750 2841.720 2897.890 ;
        RECT 2841.120 2883.610 2841.260 2897.750 ;
        RECT 2841.120 2883.470 2841.720 2883.610 ;
        RECT 2841.580 2770.730 2841.720 2883.470 ;
        RECT 2843.420 2842.130 2843.560 2945.350 ;
        RECT 2847.560 2873.410 2847.700 2963.710 ;
        RECT 2863.590 2928.915 2863.870 2929.285 ;
        RECT 2846.180 2873.270 2847.700 2873.410 ;
        RECT 2843.420 2841.990 2844.020 2842.130 ;
        RECT 2841.580 2770.590 2842.640 2770.730 ;
        RECT 2842.500 2766.650 2842.640 2770.590 ;
        RECT 2842.040 2766.510 2842.640 2766.650 ;
        RECT 2842.040 2746.250 2842.180 2766.510 ;
        RECT 2842.040 2746.110 2842.640 2746.250 ;
        RECT 2842.500 2704.090 2842.640 2746.110 ;
        RECT 2843.880 2717.690 2844.020 2841.990 ;
        RECT 2842.960 2717.550 2844.020 2717.690 ;
        RECT 2842.960 2704.770 2843.100 2717.550 ;
        RECT 2846.180 2716.330 2846.320 2873.270 ;
        RECT 2863.660 2857.010 2863.800 2928.915 ;
        RECT 2849.800 2856.920 2850.060 2857.010 ;
        RECT 2845.260 2716.190 2846.320 2716.330 ;
        RECT 2846.640 2856.780 2850.060 2856.920 ;
        RECT 2845.260 2704.770 2845.400 2716.190 ;
        RECT 2842.960 2704.630 2843.560 2704.770 ;
        RECT 2845.260 2704.630 2846.320 2704.770 ;
        RECT 2841.580 2703.950 2842.640 2704.090 ;
        RECT 2841.580 2679.610 2841.720 2703.950 ;
        RECT 2841.580 2679.470 2842.180 2679.610 ;
        RECT 2842.040 2622.490 2842.180 2679.470 ;
        RECT 2843.420 2642.890 2843.560 2704.630 ;
        RECT 2841.580 2622.350 2842.180 2622.490 ;
        RECT 2842.960 2642.750 2843.560 2642.890 ;
        RECT 2841.580 2428.690 2841.720 2622.350 ;
        RECT 2842.960 2574.210 2843.100 2642.750 ;
        RECT 2842.960 2574.070 2843.560 2574.210 ;
        RECT 2843.420 2538.850 2843.560 2574.070 ;
        RECT 2846.180 2573.530 2846.320 2704.630 ;
        RECT 2844.800 2573.390 2846.320 2573.530 ;
        RECT 2843.420 2538.710 2844.020 2538.850 ;
        RECT 2843.880 2518.450 2844.020 2538.710 ;
        RECT 2842.960 2518.310 2844.020 2518.450 ;
        RECT 2842.960 2470.850 2843.100 2518.310 ;
        RECT 2844.800 2494.650 2844.940 2573.390 ;
        RECT 2846.640 2572.850 2846.780 2856.780 ;
        RECT 2849.800 2856.690 2850.060 2856.780 ;
        RECT 2863.600 2856.690 2863.860 2857.010 ;
        RECT 2900.850 2669.155 2901.130 2669.525 ;
        RECT 2900.920 2663.890 2901.060 2669.155 ;
        RECT 2866.820 2663.570 2867.080 2663.890 ;
        RECT 2900.860 2663.570 2901.120 2663.890 ;
        RECT 2866.880 2611.870 2867.020 2663.570 ;
        RECT 2849.800 2611.610 2850.060 2611.870 ;
        RECT 2846.180 2572.710 2846.780 2572.850 ;
        RECT 2848.020 2611.550 2850.060 2611.610 ;
        RECT 2866.820 2611.550 2867.080 2611.870 ;
        RECT 2848.020 2611.470 2850.000 2611.550 ;
        RECT 2844.800 2494.510 2845.400 2494.650 ;
        RECT 2842.960 2470.710 2844.020 2470.850 ;
        RECT 2843.880 2428.690 2844.020 2470.710 ;
        RECT 2841.580 2428.550 2842.640 2428.690 ;
        RECT 2842.500 2407.610 2842.640 2428.550 ;
        RECT 2841.580 2407.470 2842.640 2407.610 ;
        RECT 2843.420 2428.550 2844.020 2428.690 ;
        RECT 2841.580 2092.090 2841.720 2407.470 ;
        RECT 2843.420 2332.130 2843.560 2428.550 ;
        RECT 2845.260 2404.890 2845.400 2494.510 ;
        RECT 2846.180 2453.170 2846.320 2572.710 ;
        RECT 2845.720 2453.030 2846.320 2453.170 ;
        RECT 2845.720 2428.690 2845.860 2453.030 ;
        RECT 2845.720 2428.550 2846.320 2428.690 ;
        RECT 2846.180 2428.010 2846.320 2428.550 ;
        RECT 2846.180 2427.870 2846.780 2428.010 ;
        RECT 2845.260 2404.750 2845.860 2404.890 ;
        RECT 2845.720 2373.610 2845.860 2404.750 ;
        RECT 2842.960 2331.990 2843.560 2332.130 ;
        RECT 2845.260 2373.470 2845.860 2373.610 ;
        RECT 2842.960 2277.050 2843.100 2331.990 ;
        RECT 2845.260 2324.650 2845.400 2373.470 ;
        RECT 2846.640 2325.160 2846.780 2427.870 ;
        RECT 2848.020 2340.290 2848.160 2611.470 ;
        RECT 2851.630 2382.450 2851.910 2382.565 ;
        RECT 2850.320 2382.310 2851.910 2382.450 ;
        RECT 2848.020 2340.150 2850.000 2340.290 ;
        RECT 2849.860 2338.170 2850.000 2340.150 ;
        RECT 2849.800 2337.850 2850.060 2338.170 ;
        RECT 2850.320 2335.450 2850.460 2382.310 ;
        RECT 2851.630 2382.195 2851.910 2382.310 ;
        RECT 2850.260 2335.130 2850.520 2335.450 ;
        RECT 2846.640 2325.020 2850.460 2325.160 ;
        RECT 2845.260 2324.510 2850.000 2324.650 ;
        RECT 2849.340 2321.190 2849.600 2321.510 ;
        RECT 2849.400 2319.890 2849.540 2321.190 ;
        RECT 2849.860 2320.150 2850.000 2324.510 ;
        RECT 2850.320 2320.830 2850.460 2325.020 ;
        RECT 2850.260 2320.510 2850.520 2320.830 ;
        RECT 2843.880 2319.750 2849.540 2319.890 ;
        RECT 2849.800 2319.830 2850.060 2320.150 ;
        RECT 2842.960 2276.910 2843.560 2277.050 ;
        RECT 2843.420 2260.050 2843.560 2276.910 ;
        RECT 2842.960 2259.910 2843.560 2260.050 ;
        RECT 2842.960 2245.090 2843.100 2259.910 ;
        RECT 2843.880 2255.290 2844.020 2319.750 ;
        RECT 2849.800 2319.210 2850.060 2319.470 ;
        RECT 2844.800 2319.150 2850.060 2319.210 ;
        RECT 2844.800 2319.070 2850.000 2319.150 ;
        RECT 2844.800 2277.050 2844.940 2319.070 ;
        RECT 2849.800 2318.530 2850.060 2318.790 ;
        RECT 2846.640 2318.470 2850.060 2318.530 ;
        RECT 2846.640 2318.390 2850.000 2318.470 ;
        RECT 2844.800 2276.910 2846.320 2277.050 ;
        RECT 2843.420 2255.150 2844.020 2255.290 ;
        RECT 2843.420 2248.490 2843.560 2255.150 ;
        RECT 2843.420 2248.350 2845.860 2248.490 ;
        RECT 2845.720 2247.130 2845.860 2248.350 ;
        RECT 2846.180 2247.130 2846.320 2276.910 ;
        RECT 2845.260 2246.990 2846.320 2247.130 ;
        RECT 2842.960 2244.950 2844.480 2245.090 ;
        RECT 2844.340 2216.530 2844.480 2244.950 ;
        RECT 2842.040 2216.390 2844.480 2216.530 ;
        RECT 2842.040 2170.290 2842.180 2216.390 ;
        RECT 2845.260 2213.810 2845.400 2246.990 ;
        RECT 2842.960 2213.670 2845.400 2213.810 ;
        RECT 2842.040 2170.150 2842.640 2170.290 ;
        RECT 2842.500 2097.530 2842.640 2170.150 ;
        RECT 2842.960 2103.650 2843.100 2213.670 ;
        RECT 2845.720 2212.450 2845.860 2246.990 ;
        RECT 2846.640 2212.450 2846.780 2318.390 ;
        RECT 2849.800 2308.500 2850.060 2308.590 ;
        RECT 2848.480 2308.360 2850.060 2308.500 ;
        RECT 2848.480 2287.930 2848.620 2308.360 ;
        RECT 2849.800 2308.270 2850.060 2308.360 ;
        RECT 2843.420 2212.310 2846.780 2212.450 ;
        RECT 2848.020 2287.790 2848.620 2287.930 ;
        RECT 2843.420 2204.290 2843.560 2212.310 ;
        RECT 2845.720 2211.770 2845.860 2212.310 ;
        RECT 2845.720 2211.630 2846.320 2211.770 ;
        RECT 2846.180 2210.410 2846.320 2211.630 ;
        RECT 2846.180 2210.270 2846.780 2210.410 ;
        RECT 2843.420 2204.150 2844.480 2204.290 ;
        RECT 2844.340 2170.290 2844.480 2204.150 ;
        RECT 2844.340 2170.150 2845.860 2170.290 ;
        RECT 2845.720 2111.130 2845.860 2170.150 ;
        RECT 2844.340 2110.990 2845.860 2111.130 ;
        RECT 2844.340 2109.770 2844.480 2110.990 ;
        RECT 2844.340 2109.630 2844.940 2109.770 ;
        RECT 2844.800 2108.410 2844.940 2109.630 ;
        RECT 2844.340 2108.270 2844.940 2108.410 ;
        RECT 2844.340 2105.690 2844.480 2108.270 ;
        RECT 2843.880 2105.550 2844.480 2105.690 ;
        RECT 2843.880 2104.330 2844.020 2105.550 ;
        RECT 2843.880 2104.190 2844.480 2104.330 ;
        RECT 2844.340 2103.650 2844.480 2104.190 ;
        RECT 2842.960 2103.510 2845.860 2103.650 ;
        RECT 2844.340 2102.970 2844.480 2103.510 ;
        RECT 2844.340 2102.830 2844.940 2102.970 ;
        RECT 2842.500 2097.390 2844.480 2097.530 ;
        RECT 2841.580 2091.950 2842.180 2092.090 ;
        RECT 2842.040 2090.900 2842.180 2091.950 ;
        RECT 2841.580 2090.760 2842.180 2090.900 ;
        RECT 2841.580 2056.730 2841.720 2090.760 ;
        RECT 2841.120 2056.590 2841.720 2056.730 ;
        RECT 2841.120 1997.740 2841.260 2056.590 ;
        RECT 2844.340 2034.290 2844.480 2097.390 ;
        RECT 2842.960 2034.150 2844.480 2034.290 ;
        RECT 2842.960 2032.930 2843.100 2034.150 ;
        RECT 2842.040 2032.790 2843.100 2032.930 ;
        RECT 2842.040 2028.170 2842.180 2032.790 ;
        RECT 2844.800 2029.530 2844.940 2102.830 ;
        RECT 2845.720 2066.930 2845.860 2103.510 ;
        RECT 2843.420 2029.390 2844.940 2029.530 ;
        RECT 2845.260 2066.790 2845.860 2066.930 ;
        RECT 2842.040 2028.030 2842.640 2028.170 ;
        RECT 2842.500 2003.690 2842.640 2028.030 ;
        RECT 2843.420 2004.370 2843.560 2029.390 ;
        RECT 2845.260 2027.490 2845.400 2066.790 ;
        RECT 2845.260 2027.350 2846.320 2027.490 ;
        RECT 2843.420 2004.230 2844.480 2004.370 ;
        RECT 2842.500 2003.550 2844.020 2003.690 ;
        RECT 2841.120 1997.600 2842.180 1997.740 ;
        RECT 2842.040 1970.370 2842.180 1997.600 ;
        RECT 2841.580 1970.230 2842.180 1970.370 ;
        RECT 2841.580 1952.010 2841.720 1970.230 ;
        RECT 2843.880 1969.690 2844.020 2003.550 ;
        RECT 2841.120 1951.870 2841.720 1952.010 ;
        RECT 2842.040 1969.550 2844.020 1969.690 ;
        RECT 2841.120 1872.450 2841.260 1951.870 ;
        RECT 2842.040 1945.380 2842.180 1969.550 ;
        RECT 2844.340 1969.180 2844.480 2004.230 ;
        RECT 2843.420 1969.040 2844.480 1969.180 ;
        RECT 2843.420 1964.250 2843.560 1969.040 ;
        RECT 2846.180 1965.610 2846.320 2027.350 ;
        RECT 2846.640 1968.330 2846.780 2210.270 ;
        RECT 2848.020 1996.890 2848.160 2287.790 ;
        RECT 2863.590 2112.915 2863.870 2113.285 ;
        RECT 2863.660 2060.050 2863.800 2112.915 ;
        RECT 2853.020 2059.730 2853.280 2060.050 ;
        RECT 2863.600 2059.730 2863.860 2060.050 ;
        RECT 2853.080 2008.370 2853.220 2059.730 ;
        RECT 2849.800 2008.050 2850.060 2008.370 ;
        RECT 2853.020 2008.050 2853.280 2008.370 ;
        RECT 2848.020 1996.750 2848.620 1996.890 ;
        RECT 2848.480 1974.960 2848.620 1996.750 ;
        RECT 2849.860 1984.230 2850.000 2008.050 ;
        RECT 2849.800 1983.910 2850.060 1984.230 ;
        RECT 2849.800 1974.960 2850.060 1975.050 ;
        RECT 2848.480 1974.820 2850.060 1974.960 ;
        RECT 2849.800 1974.730 2850.060 1974.820 ;
        RECT 2851.630 1974.195 2851.910 1974.565 ;
        RECT 2846.640 1968.190 2849.080 1968.330 ;
        RECT 2848.940 1966.290 2849.080 1968.190 ;
        RECT 2848.940 1966.150 2850.000 1966.290 ;
        RECT 2849.860 1965.870 2850.000 1966.150 ;
        RECT 2846.180 1965.470 2849.540 1965.610 ;
        RECT 2849.800 1965.550 2850.060 1965.870 ;
        RECT 2849.400 1964.930 2849.540 1965.470 ;
        RECT 2849.400 1964.850 2850.000 1964.930 ;
        RECT 2849.400 1964.790 2850.060 1964.850 ;
        RECT 2849.800 1964.530 2850.060 1964.790 ;
        RECT 2843.420 1964.110 2850.460 1964.250 ;
        RECT 2849.800 1963.740 2850.060 1963.830 ;
        RECT 2842.960 1963.600 2850.060 1963.740 ;
        RECT 2842.960 1945.380 2843.100 1963.600 ;
        RECT 2849.800 1963.510 2850.060 1963.600 ;
        RECT 2849.800 1962.830 2850.060 1963.150 ;
        RECT 2849.860 1962.210 2850.000 1962.830 ;
        RECT 2845.720 1962.070 2850.000 1962.210 ;
        RECT 2845.720 1949.290 2845.860 1962.070 ;
        RECT 2849.800 1961.700 2850.060 1961.790 ;
        RECT 2847.100 1961.560 2850.060 1961.700 ;
        RECT 2847.100 1961.530 2847.240 1961.560 ;
        RECT 2843.880 1949.150 2845.860 1949.290 ;
        RECT 2846.180 1961.390 2847.240 1961.530 ;
        RECT 2849.800 1961.470 2850.060 1961.560 ;
        RECT 2842.040 1945.240 2842.640 1945.380 ;
        RECT 2842.960 1945.240 2843.560 1945.380 ;
        RECT 2842.500 1943.850 2842.640 1945.240 ;
        RECT 2842.500 1943.710 2843.100 1943.850 ;
        RECT 2842.960 1873.130 2843.100 1943.710 ;
        RECT 2843.420 1883.330 2843.560 1945.240 ;
        RECT 2843.880 1886.050 2844.020 1949.150 ;
        RECT 2846.180 1948.610 2846.320 1961.390 ;
        RECT 2850.320 1960.850 2850.460 1964.110 ;
        RECT 2851.700 1963.150 2851.840 1974.195 ;
        RECT 2851.640 1962.830 2851.900 1963.150 ;
        RECT 2845.260 1948.470 2846.320 1948.610 ;
        RECT 2847.560 1960.710 2850.460 1960.850 ;
        RECT 2845.260 1905.770 2845.400 1948.470 ;
        RECT 2847.560 1947.930 2847.700 1960.710 ;
        RECT 2849.800 1949.970 2850.060 1950.230 ;
        RECT 2844.800 1905.630 2845.400 1905.770 ;
        RECT 2846.180 1947.790 2847.700 1947.930 ;
        RECT 2848.020 1949.910 2850.060 1949.970 ;
        RECT 2848.020 1949.830 2850.000 1949.910 ;
        RECT 2844.800 1904.410 2844.940 1905.630 ;
        RECT 2844.800 1904.270 2845.400 1904.410 ;
        RECT 2843.880 1885.910 2844.940 1886.050 ;
        RECT 2843.420 1883.190 2844.480 1883.330 ;
        RECT 2841.580 1872.990 2843.100 1873.130 ;
        RECT 2841.580 1872.450 2841.720 1872.990 ;
        RECT 2841.120 1872.310 2844.020 1872.450 ;
        RECT 2841.580 1870.410 2841.720 1872.310 ;
        RECT 2841.120 1870.270 2841.720 1870.410 ;
        RECT 2841.120 1814.650 2841.260 1870.270 ;
        RECT 2843.880 1865.650 2844.020 1872.310 ;
        RECT 2841.580 1865.510 2844.020 1865.650 ;
        RECT 2841.580 1857.490 2841.720 1865.510 ;
        RECT 2841.580 1857.350 2842.640 1857.490 ;
        RECT 2842.500 1820.770 2842.640 1857.350 ;
        RECT 2842.500 1820.630 2843.100 1820.770 ;
        RECT 2842.960 1816.010 2843.100 1820.630 ;
        RECT 2844.340 1819.410 2844.480 1883.190 ;
        RECT 2844.800 1820.090 2844.940 1885.910 ;
        RECT 2845.260 1837.770 2845.400 1904.270 ;
        RECT 2846.180 1890.810 2846.320 1947.790 ;
        RECT 2848.020 1946.570 2848.160 1949.830 ;
        RECT 2845.720 1890.670 2846.320 1890.810 ;
        RECT 2846.640 1946.430 2848.160 1946.570 ;
        RECT 2845.720 1838.450 2845.860 1890.670 ;
        RECT 2846.640 1890.130 2846.780 1946.430 ;
        RECT 2849.800 1942.490 2850.060 1942.750 ;
        RECT 2848.020 1942.430 2850.060 1942.490 ;
        RECT 2848.020 1942.350 2850.000 1942.430 ;
        RECT 2848.020 1892.170 2848.160 1942.350 ;
        RECT 2848.020 1892.030 2849.540 1892.170 ;
        RECT 2846.180 1889.990 2846.780 1890.130 ;
        RECT 2846.180 1839.810 2846.320 1889.990 ;
        RECT 2849.400 1885.370 2849.540 1892.030 ;
        RECT 2848.020 1885.230 2849.540 1885.370 ;
        RECT 2848.020 1847.290 2848.160 1885.230 ;
        RECT 2848.020 1847.210 2850.000 1847.290 ;
        RECT 2848.020 1847.150 2850.060 1847.210 ;
        RECT 2849.800 1846.890 2850.060 1847.150 ;
        RECT 2846.180 1839.670 2847.240 1839.810 ;
        RECT 2847.100 1838.960 2847.240 1839.670 ;
        RECT 2849.800 1838.960 2850.060 1839.050 ;
        RECT 2847.100 1838.820 2850.060 1838.960 ;
        RECT 2849.800 1838.730 2850.060 1838.820 ;
        RECT 2845.720 1838.310 2850.000 1838.450 ;
        RECT 2845.260 1837.630 2848.160 1837.770 ;
        RECT 2844.800 1819.950 2847.240 1820.090 ;
        RECT 2844.340 1819.270 2844.940 1819.410 ;
        RECT 2844.800 1818.050 2844.940 1819.270 ;
        RECT 2844.800 1817.910 2846.780 1818.050 ;
        RECT 2842.960 1815.870 2844.020 1816.010 ;
        RECT 2843.880 1814.650 2844.020 1815.870 ;
        RECT 2841.120 1814.510 2845.400 1814.650 ;
        RECT 2843.880 1813.970 2844.020 1814.510 ;
        RECT 2842.960 1813.830 2844.020 1813.970 ;
        RECT 2842.960 1793.570 2843.100 1813.830 ;
        RECT 2845.260 1794.420 2845.400 1814.510 ;
        RECT 2846.640 1813.970 2846.780 1817.910 ;
        RECT 2845.720 1813.830 2846.780 1813.970 ;
        RECT 2845.720 1795.780 2845.860 1813.830 ;
        RECT 2847.100 1797.820 2847.240 1819.950 ;
        RECT 2848.020 1799.520 2848.160 1837.630 ;
        RECT 2849.860 1800.290 2850.000 1838.310 ;
        RECT 2851.630 1838.195 2851.910 1838.565 ;
        RECT 2851.700 1800.880 2851.840 1838.195 ;
        RECT 2851.240 1800.740 2851.840 1800.880 ;
        RECT 2849.800 1799.970 2850.060 1800.290 ;
        RECT 2849.800 1799.520 2850.060 1799.610 ;
        RECT 2848.020 1799.380 2850.060 1799.520 ;
        RECT 2849.800 1799.290 2850.060 1799.380 ;
        RECT 2849.800 1797.820 2850.060 1797.910 ;
        RECT 2847.100 1797.680 2850.060 1797.820 ;
        RECT 2849.800 1797.590 2850.060 1797.680 ;
        RECT 2849.800 1795.780 2850.060 1795.870 ;
        RECT 2845.720 1795.640 2850.060 1795.780 ;
        RECT 2849.800 1795.550 2850.060 1795.640 ;
        RECT 2849.800 1794.420 2850.060 1794.510 ;
        RECT 2845.260 1794.280 2850.060 1794.420 ;
        RECT 2849.800 1794.190 2850.060 1794.280 ;
        RECT 2851.240 1793.830 2851.380 1800.740 ;
        RECT 2851.640 1799.970 2851.900 1800.290 ;
        RECT 2849.800 1793.740 2850.060 1793.830 ;
        RECT 2841.120 1793.430 2843.100 1793.570 ;
        RECT 2843.420 1793.600 2850.060 1793.740 ;
        RECT 2841.120 1695.650 2841.260 1793.430 ;
        RECT 2842.040 1792.750 2843.100 1792.890 ;
        RECT 2842.040 1792.210 2842.180 1792.750 ;
        RECT 2841.580 1792.070 2842.180 1792.210 ;
        RECT 2842.960 1792.210 2843.100 1792.750 ;
        RECT 2843.420 1792.210 2843.560 1793.600 ;
        RECT 2849.800 1793.510 2850.060 1793.600 ;
        RECT 2851.180 1793.510 2851.440 1793.830 ;
        RECT 2849.800 1793.060 2850.060 1793.150 ;
        RECT 2842.960 1792.070 2843.560 1792.210 ;
        RECT 2849.400 1792.920 2850.060 1793.060 ;
        RECT 2841.580 1697.010 2841.720 1792.070 ;
        RECT 2849.400 1791.360 2849.540 1792.920 ;
        RECT 2849.800 1792.830 2850.060 1792.920 ;
        RECT 2842.960 1791.220 2849.540 1791.360 ;
        RECT 2842.960 1718.770 2843.100 1791.220 ;
        RECT 2849.800 1791.130 2850.060 1791.450 ;
        RECT 2849.860 1790.680 2850.000 1791.130 ;
        RECT 2844.340 1790.540 2850.000 1790.680 ;
        RECT 2844.340 1784.730 2844.480 1790.540 ;
        RECT 2851.180 1790.170 2851.440 1790.430 ;
        RECT 2843.420 1784.590 2844.480 1784.730 ;
        RECT 2846.180 1790.110 2851.440 1790.170 ;
        RECT 2846.180 1790.030 2851.380 1790.110 ;
        RECT 2843.420 1720.130 2843.560 1784.590 ;
        RECT 2846.180 1783.370 2846.320 1790.030 ;
        RECT 2844.800 1783.230 2846.320 1783.370 ;
        RECT 2844.800 1748.010 2844.940 1783.230 ;
        RECT 2844.340 1747.870 2844.940 1748.010 ;
        RECT 2845.260 1771.670 2848.160 1771.810 ;
        RECT 2844.340 1724.210 2844.480 1747.870 ;
        RECT 2845.260 1747.330 2845.400 1771.670 ;
        RECT 2848.020 1768.920 2848.160 1771.670 ;
        RECT 2849.800 1768.920 2850.060 1769.010 ;
        RECT 2848.020 1768.780 2850.060 1768.920 ;
        RECT 2849.800 1768.690 2850.060 1768.780 ;
        RECT 2851.700 1766.630 2851.840 1799.970 ;
        RECT 2851.640 1766.310 2851.900 1766.630 ;
        RECT 2849.340 1765.970 2849.600 1766.290 ;
        RECT 2844.800 1747.190 2845.400 1747.330 ;
        RECT 2844.800 1724.210 2844.940 1747.190 ;
        RECT 2849.400 1745.970 2849.540 1765.970 ;
        RECT 2849.800 1761.550 2850.060 1761.870 ;
        RECT 2843.880 1724.070 2844.940 1724.210 ;
        RECT 2846.180 1745.830 2849.540 1745.970 ;
        RECT 2843.880 1720.810 2844.020 1724.070 ;
        RECT 2844.340 1721.490 2844.480 1724.070 ;
        RECT 2844.340 1721.350 2845.400 1721.490 ;
        RECT 2843.880 1720.670 2844.480 1720.810 ;
        RECT 2843.420 1719.990 2844.020 1720.130 ;
        RECT 2842.960 1718.630 2843.560 1718.770 ;
        RECT 2841.580 1696.870 2843.100 1697.010 ;
        RECT 2841.120 1695.510 2842.640 1695.650 ;
        RECT 2842.500 1687.490 2842.640 1695.510 ;
        RECT 2841.580 1687.350 2842.640 1687.490 ;
        RECT 2841.580 1686.810 2841.720 1687.350 ;
        RECT 2842.960 1686.810 2843.100 1696.870 ;
        RECT 2841.120 1686.670 2843.100 1686.810 ;
        RECT 2841.120 1577.840 2841.260 1686.670 ;
        RECT 2841.580 1601.130 2841.720 1686.670 ;
        RECT 2843.420 1663.690 2843.560 1718.630 ;
        RECT 2842.960 1663.550 2843.560 1663.690 ;
        RECT 2842.960 1663.010 2843.100 1663.550 ;
        RECT 2843.880 1663.010 2844.020 1719.990 ;
        RECT 2842.500 1662.870 2843.100 1663.010 ;
        RECT 2843.420 1662.870 2844.020 1663.010 ;
        RECT 2842.500 1639.040 2842.640 1662.870 ;
        RECT 2843.420 1639.890 2843.560 1662.870 ;
        RECT 2844.340 1644.650 2844.480 1720.670 ;
        RECT 2845.260 1688.170 2845.400 1721.350 ;
        RECT 2846.180 1698.370 2846.320 1745.830 ;
        RECT 2849.860 1745.290 2850.000 1761.550 ;
        RECT 2847.100 1745.150 2850.000 1745.290 ;
        RECT 2847.100 1741.890 2847.240 1745.150 ;
        RECT 2846.640 1741.750 2847.240 1741.890 ;
        RECT 2846.640 1699.050 2846.780 1741.750 ;
        RECT 2849.800 1740.020 2850.060 1740.110 ;
        RECT 2848.020 1739.880 2850.060 1740.020 ;
        RECT 2848.020 1701.090 2848.160 1739.880 ;
        RECT 2849.800 1739.790 2850.060 1739.880 ;
        RECT 2863.590 1704.915 2863.870 1705.285 ;
        RECT 2848.020 1700.950 2849.080 1701.090 ;
        RECT 2846.640 1698.910 2847.700 1699.050 ;
        RECT 2846.180 1698.230 2847.240 1698.370 ;
        RECT 2847.100 1688.170 2847.240 1698.230 ;
        RECT 2844.800 1688.030 2845.400 1688.170 ;
        RECT 2845.720 1688.030 2847.240 1688.170 ;
        RECT 2844.800 1646.690 2844.940 1688.030 ;
        RECT 2844.800 1646.550 2845.400 1646.690 ;
        RECT 2845.260 1645.330 2845.400 1646.550 ;
        RECT 2845.720 1646.010 2845.860 1688.030 ;
        RECT 2847.560 1686.810 2847.700 1698.910 ;
        RECT 2846.640 1686.670 2847.700 1686.810 ;
        RECT 2846.640 1648.050 2846.780 1686.670 ;
        RECT 2848.940 1680.010 2849.080 1700.950 ;
        RECT 2848.020 1679.870 2849.080 1680.010 ;
        RECT 2848.020 1652.130 2848.160 1679.870 ;
        RECT 2848.020 1651.990 2850.920 1652.130 ;
        RECT 2846.640 1647.970 2850.000 1648.050 ;
        RECT 2846.640 1647.910 2850.060 1647.970 ;
        RECT 2849.800 1647.650 2850.060 1647.910 ;
        RECT 2847.100 1647.290 2850.000 1647.370 ;
        RECT 2847.100 1647.230 2850.060 1647.290 ;
        RECT 2847.100 1646.010 2847.240 1647.230 ;
        RECT 2849.800 1646.970 2850.060 1647.230 ;
        RECT 2845.720 1645.870 2847.240 1646.010 ;
        RECT 2847.560 1646.610 2850.000 1646.690 ;
        RECT 2847.560 1646.550 2850.060 1646.610 ;
        RECT 2847.560 1645.330 2847.700 1646.550 ;
        RECT 2849.800 1646.290 2850.060 1646.550 ;
        RECT 2845.260 1645.190 2847.700 1645.330 ;
        RECT 2844.340 1644.510 2845.400 1644.650 ;
        RECT 2843.420 1639.750 2844.480 1639.890 ;
        RECT 2842.040 1638.900 2842.640 1639.040 ;
        RECT 2842.040 1622.210 2842.180 1638.900 ;
        RECT 2842.040 1622.070 2843.100 1622.210 ;
        RECT 2841.580 1600.990 2842.180 1601.130 ;
        RECT 2842.040 1579.200 2842.180 1600.990 ;
        RECT 2842.960 1589.740 2843.100 1622.070 ;
        RECT 2844.340 1620.850 2844.480 1639.750 ;
        RECT 2845.260 1639.040 2845.400 1644.510 ;
        RECT 2849.800 1639.040 2850.060 1639.130 ;
        RECT 2845.260 1638.900 2850.060 1639.040 ;
        RECT 2849.800 1638.810 2850.060 1638.900 ;
        RECT 2846.180 1638.390 2848.160 1638.530 ;
        RECT 2844.340 1620.710 2844.940 1620.850 ;
        RECT 2844.800 1614.730 2844.940 1620.710 ;
        RECT 2846.180 1614.730 2846.320 1638.390 ;
        RECT 2848.020 1638.360 2848.160 1638.390 ;
        RECT 2849.800 1638.360 2850.060 1638.450 ;
        RECT 2848.020 1638.220 2850.060 1638.360 ;
        RECT 2849.800 1638.130 2850.060 1638.220 ;
        RECT 2849.800 1635.980 2850.060 1636.070 ;
        RECT 2843.420 1614.590 2844.940 1614.730 ;
        RECT 2845.260 1614.590 2846.320 1614.730 ;
        RECT 2847.560 1635.840 2850.060 1635.980 ;
        RECT 2843.420 1600.450 2843.560 1614.590 ;
        RECT 2845.260 1607.930 2845.400 1614.590 ;
        RECT 2845.260 1607.790 2846.320 1607.930 ;
        RECT 2843.420 1600.310 2845.860 1600.450 ;
        RECT 2842.960 1589.600 2844.020 1589.740 ;
        RECT 2842.040 1579.060 2843.560 1579.200 ;
        RECT 2841.120 1577.700 2841.720 1577.840 ;
        RECT 2841.580 1577.500 2841.720 1577.700 ;
        RECT 2841.120 1577.360 2841.720 1577.500 ;
        RECT 2841.120 1575.970 2841.260 1577.360 ;
        RECT 2841.120 1575.830 2841.720 1575.970 ;
        RECT 2841.580 1573.930 2841.720 1575.830 ;
        RECT 2843.420 1573.930 2843.560 1579.060 ;
        RECT 2841.120 1573.790 2843.560 1573.930 ;
        RECT 2843.880 1573.930 2844.020 1589.600 ;
        RECT 2845.720 1575.970 2845.860 1600.310 ;
        RECT 2846.180 1577.500 2846.320 1607.790 ;
        RECT 2847.560 1600.450 2847.700 1635.840 ;
        RECT 2849.800 1635.750 2850.060 1635.840 ;
        RECT 2849.800 1635.300 2850.060 1635.390 ;
        RECT 2848.940 1635.160 2850.060 1635.300 ;
        RECT 2848.940 1603.680 2849.080 1635.160 ;
        RECT 2849.800 1635.070 2850.060 1635.160 ;
        RECT 2849.800 1628.500 2850.060 1628.590 ;
        RECT 2849.400 1628.360 2850.060 1628.500 ;
        RECT 2849.400 1604.530 2849.540 1628.360 ;
        RECT 2849.800 1628.270 2850.060 1628.360 ;
        RECT 2850.780 1627.910 2850.920 1651.990 ;
        RECT 2863.660 1638.450 2863.800 1704.915 ;
        RECT 2863.600 1638.130 2863.860 1638.450 ;
        RECT 2850.720 1627.590 2850.980 1627.910 ;
        RECT 2850.720 1604.810 2850.980 1605.130 ;
        RECT 2849.400 1604.450 2850.000 1604.530 ;
        RECT 2849.400 1604.390 2850.060 1604.450 ;
        RECT 2849.800 1604.130 2850.060 1604.390 ;
        RECT 2848.940 1603.540 2849.540 1603.680 ;
        RECT 2849.400 1602.490 2849.540 1603.540 ;
        RECT 2850.780 1603.170 2850.920 1604.810 ;
        RECT 2848.940 1602.350 2849.540 1602.490 ;
        RECT 2850.320 1603.030 2850.920 1603.170 ;
        RECT 2847.560 1600.310 2848.160 1600.450 ;
        RECT 2846.180 1577.360 2847.700 1577.500 ;
        RECT 2845.720 1575.830 2846.320 1575.970 ;
        RECT 2843.880 1573.790 2844.480 1573.930 ;
        RECT 2841.120 1501.850 2841.260 1573.790 ;
        RECT 2841.580 1549.280 2841.720 1573.790 ;
        RECT 2844.340 1573.270 2844.480 1573.790 ;
        RECT 2844.340 1573.130 2844.940 1573.270 ;
        RECT 2844.800 1552.850 2844.940 1573.130 ;
        RECT 2842.040 1552.710 2844.940 1552.850 ;
        RECT 2842.040 1549.280 2842.180 1552.710 ;
        RECT 2841.580 1549.140 2842.640 1549.280 ;
        RECT 2842.040 1548.770 2842.180 1549.140 ;
        RECT 2841.580 1548.630 2842.180 1548.770 ;
        RECT 2841.580 1541.970 2841.720 1548.630 ;
        RECT 2842.500 1546.730 2842.640 1549.140 ;
        RECT 2842.040 1546.590 2842.640 1546.730 ;
        RECT 2842.960 1546.590 2844.940 1546.730 ;
        RECT 2842.040 1542.650 2842.180 1546.590 ;
        RECT 2842.960 1545.540 2843.100 1546.590 ;
        RECT 2844.800 1545.540 2844.940 1546.590 ;
        RECT 2842.500 1545.400 2843.100 1545.540 ;
        RECT 2844.340 1545.400 2844.940 1545.540 ;
        RECT 2842.500 1542.650 2842.640 1545.400 ;
        RECT 2844.340 1543.330 2844.480 1545.400 ;
        RECT 2844.340 1543.190 2845.400 1543.330 ;
        RECT 2842.040 1542.510 2844.940 1542.650 ;
        RECT 2842.500 1541.970 2842.640 1542.510 ;
        RECT 2841.580 1541.830 2843.560 1541.970 ;
        RECT 2842.500 1503.210 2842.640 1541.830 ;
        RECT 2843.420 1505.250 2843.560 1541.830 ;
        RECT 2844.800 1514.090 2844.940 1542.510 ;
        RECT 2845.260 1524.970 2845.400 1543.190 ;
        RECT 2846.180 1524.970 2846.320 1575.830 ;
        RECT 2847.560 1573.250 2847.700 1577.360 ;
        RECT 2848.020 1576.650 2848.160 1600.310 ;
        RECT 2848.940 1578.180 2849.080 1602.350 ;
        RECT 2850.320 1579.290 2850.460 1603.030 ;
        RECT 2850.260 1578.970 2850.520 1579.290 ;
        RECT 2851.640 1578.970 2851.900 1579.290 ;
        RECT 2849.800 1578.180 2850.060 1578.270 ;
        RECT 2848.940 1578.040 2850.060 1578.180 ;
        RECT 2849.800 1577.950 2850.060 1578.040 ;
        RECT 2848.020 1576.510 2850.000 1576.650 ;
        RECT 2847.100 1573.110 2847.700 1573.250 ;
        RECT 2847.100 1549.280 2847.240 1573.110 ;
        RECT 2845.260 1524.830 2846.320 1524.970 ;
        RECT 2846.640 1549.140 2847.240 1549.280 ;
        RECT 2844.800 1513.950 2845.860 1514.090 ;
        RECT 2845.720 1505.250 2845.860 1513.950 ;
        RECT 2843.420 1505.110 2846.320 1505.250 ;
        RECT 2845.720 1504.400 2845.860 1505.110 ;
        RECT 2845.260 1504.260 2845.860 1504.400 ;
        RECT 2842.500 1503.070 2843.560 1503.210 ;
        RECT 2841.120 1501.710 2842.640 1501.850 ;
        RECT 2842.500 1500.660 2842.640 1501.710 ;
        RECT 2843.420 1501.170 2843.560 1503.070 ;
        RECT 2842.960 1501.030 2843.560 1501.170 ;
        RECT 2842.960 1500.660 2843.100 1501.030 ;
        RECT 2841.120 1500.520 2843.100 1500.660 ;
        RECT 2841.120 1371.120 2841.260 1500.520 ;
        RECT 2842.500 1420.250 2842.640 1500.520 ;
        RECT 2845.260 1500.490 2845.400 1504.260 ;
        RECT 2843.420 1500.350 2845.400 1500.490 ;
        RECT 2843.420 1500.320 2843.560 1500.350 ;
        RECT 2842.960 1500.180 2843.560 1500.320 ;
        RECT 2842.960 1421.610 2843.100 1500.180 ;
        RECT 2846.180 1475.840 2846.320 1505.110 ;
        RECT 2845.720 1475.700 2846.320 1475.840 ;
        RECT 2845.720 1423.140 2845.860 1475.700 ;
        RECT 2846.640 1475.330 2846.780 1549.140 ;
        RECT 2849.860 1546.050 2850.000 1576.510 ;
        RECT 2848.940 1545.910 2850.000 1546.050 ;
        RECT 2848.940 1545.370 2849.080 1545.910 ;
        RECT 2847.560 1545.230 2849.080 1545.370 ;
        RECT 2849.800 1545.310 2850.060 1545.630 ;
        RECT 2847.560 1505.930 2847.700 1545.230 ;
        RECT 2849.860 1539.250 2850.000 1545.310 ;
        RECT 2849.400 1539.110 2850.000 1539.250 ;
        RECT 2849.400 1537.890 2849.540 1539.110 ;
        RECT 2849.400 1537.750 2850.000 1537.890 ;
        RECT 2849.860 1535.090 2850.000 1537.750 ;
        RECT 2849.800 1534.770 2850.060 1535.090 ;
        RECT 2849.800 1530.920 2850.060 1531.010 ;
        RECT 2848.020 1530.780 2850.060 1530.920 ;
        RECT 2848.020 1513.920 2848.160 1530.780 ;
        RECT 2849.800 1530.690 2850.060 1530.780 ;
        RECT 2851.700 1514.770 2851.840 1578.970 ;
        RECT 2863.590 1568.915 2863.870 1569.285 ;
        RECT 2851.240 1514.630 2851.840 1514.770 ;
        RECT 2849.800 1513.920 2850.060 1514.010 ;
        RECT 2848.020 1513.780 2850.060 1513.920 ;
        RECT 2849.800 1513.690 2850.060 1513.780 ;
        RECT 2847.560 1505.850 2850.000 1505.930 ;
        RECT 2847.560 1505.790 2850.060 1505.850 ;
        RECT 2849.800 1505.530 2850.060 1505.790 ;
        RECT 2849.800 1504.170 2850.060 1504.490 ;
        RECT 2849.860 1500.410 2850.000 1504.170 ;
        RECT 2849.800 1500.090 2850.060 1500.410 ;
        RECT 2849.800 1492.840 2850.060 1492.930 ;
        RECT 2848.020 1492.700 2850.060 1492.840 ;
        RECT 2848.020 1482.130 2848.160 1492.700 ;
        RECT 2849.800 1492.610 2850.060 1492.700 ;
        RECT 2849.800 1491.930 2850.060 1492.250 ;
        RECT 2846.180 1475.190 2846.780 1475.330 ;
        RECT 2847.560 1481.990 2848.160 1482.130 ;
        RECT 2846.180 1457.650 2846.320 1475.190 ;
        RECT 2847.560 1471.250 2847.700 1481.990 ;
        RECT 2849.860 1481.450 2850.000 1491.930 ;
        RECT 2847.100 1471.110 2847.700 1471.250 ;
        RECT 2848.020 1481.310 2850.000 1481.450 ;
        RECT 2846.180 1457.510 2846.780 1457.650 ;
        RECT 2846.640 1424.330 2846.780 1457.510 ;
        RECT 2847.100 1425.010 2847.240 1471.110 ;
        RECT 2848.020 1468.530 2848.160 1481.310 ;
        RECT 2850.260 1480.710 2850.520 1481.030 ;
        RECT 2847.560 1468.390 2848.160 1468.530 ;
        RECT 2847.560 1425.860 2847.700 1468.390 ;
        RECT 2850.320 1466.490 2850.460 1480.710 ;
        RECT 2851.240 1480.350 2851.380 1514.630 ;
        RECT 2851.180 1480.030 2851.440 1480.350 ;
        RECT 2848.940 1466.350 2850.460 1466.490 ;
        RECT 2848.940 1439.290 2849.080 1466.350 ;
        RECT 2849.800 1462.010 2850.060 1462.330 ;
        RECT 2849.860 1448.390 2850.000 1462.010 ;
        RECT 2849.800 1448.070 2850.060 1448.390 ;
        RECT 2848.940 1439.150 2850.000 1439.290 ;
        RECT 2849.860 1426.970 2850.000 1439.150 ;
        RECT 2852.090 1430.195 2852.370 1430.565 ;
        RECT 2849.800 1426.650 2850.060 1426.970 ;
        RECT 2849.800 1425.860 2850.060 1425.950 ;
        RECT 2847.560 1425.720 2850.060 1425.860 ;
        RECT 2849.800 1425.630 2850.060 1425.720 ;
        RECT 2847.100 1424.930 2850.000 1425.010 ;
        RECT 2847.100 1424.870 2850.060 1424.930 ;
        RECT 2849.800 1424.610 2850.060 1424.870 ;
        RECT 2846.640 1424.250 2850.000 1424.330 ;
        RECT 2846.640 1424.190 2850.060 1424.250 ;
        RECT 2849.800 1423.930 2850.060 1424.190 ;
        RECT 2849.800 1423.140 2850.060 1423.230 ;
        RECT 2845.720 1423.000 2850.060 1423.140 ;
        RECT 2849.800 1422.910 2850.060 1423.000 ;
        RECT 2842.960 1421.470 2850.000 1421.610 ;
        RECT 2842.500 1420.110 2843.560 1420.250 ;
        RECT 2843.420 1418.210 2843.560 1420.110 ;
        RECT 2849.860 1419.490 2850.000 1421.470 ;
        RECT 2849.800 1419.170 2850.060 1419.490 ;
        RECT 2849.800 1418.490 2850.060 1418.810 ;
        RECT 2849.860 1418.210 2850.000 1418.490 ;
        RECT 2842.500 1418.070 2843.560 1418.210 ;
        RECT 2845.260 1418.070 2850.000 1418.210 ;
        RECT 2842.500 1384.210 2842.640 1418.070 ;
        RECT 2845.260 1386.930 2845.400 1418.070 ;
        RECT 2849.800 1417.530 2850.060 1417.790 ;
        RECT 2845.720 1417.470 2850.060 1417.530 ;
        RECT 2845.720 1417.390 2850.000 1417.470 ;
        RECT 2845.720 1387.780 2845.860 1417.390 ;
        RECT 2849.800 1417.020 2850.060 1417.110 ;
        RECT 2846.180 1416.880 2850.060 1417.020 ;
        RECT 2846.180 1389.820 2846.320 1416.880 ;
        RECT 2849.800 1416.790 2850.060 1416.880 ;
        RECT 2850.260 1416.450 2850.520 1416.770 ;
        RECT 2849.800 1389.820 2850.060 1389.910 ;
        RECT 2846.180 1389.680 2850.060 1389.820 ;
        RECT 2849.800 1389.590 2850.060 1389.680 ;
        RECT 2849.800 1387.780 2850.060 1387.870 ;
        RECT 2845.720 1387.640 2850.060 1387.780 ;
        RECT 2849.800 1387.550 2850.060 1387.640 ;
        RECT 2845.260 1386.790 2846.320 1386.930 ;
        RECT 2846.180 1386.420 2846.320 1386.790 ;
        RECT 2849.800 1386.420 2850.060 1386.510 ;
        RECT 2846.180 1386.280 2850.060 1386.420 ;
        RECT 2849.800 1386.190 2850.060 1386.280 ;
        RECT 2842.500 1384.070 2850.000 1384.210 ;
        RECT 2849.860 1372.570 2850.000 1384.070 ;
        RECT 2849.800 1372.250 2850.060 1372.570 ;
        RECT 2849.800 1371.120 2850.060 1371.210 ;
        RECT 2841.120 1370.980 2850.060 1371.120 ;
        RECT 2849.800 1370.890 2850.060 1370.980 ;
        RECT 2850.320 1370.610 2850.460 1416.450 ;
        RECT 2851.640 1389.590 2851.900 1389.910 ;
        RECT 2850.720 1387.550 2850.980 1387.870 ;
        RECT 2849.860 1370.470 2850.460 1370.610 ;
        RECT 2849.860 1365.430 2850.000 1370.470 ;
        RECT 2850.260 1368.510 2850.520 1368.830 ;
        RECT 2849.800 1365.110 2850.060 1365.430 ;
        RECT 2849.800 1364.490 2850.060 1364.750 ;
        RECT 2841.120 1364.430 2850.060 1364.490 ;
        RECT 2841.120 1364.350 2850.000 1364.430 ;
        RECT 2841.120 1184.290 2841.260 1364.350 ;
        RECT 2849.800 1363.980 2850.060 1364.070 ;
        RECT 2842.500 1363.840 2850.060 1363.980 ;
        RECT 2841.970 1242.090 2842.250 1242.205 ;
        RECT 2841.580 1241.950 2842.250 1242.090 ;
        RECT 2841.580 1184.970 2841.720 1241.950 ;
        RECT 2841.970 1241.835 2842.250 1241.950 ;
        RECT 2842.500 1218.970 2842.640 1363.840 ;
        RECT 2849.800 1363.750 2850.060 1363.840 ;
        RECT 2849.800 1362.730 2850.060 1363.050 ;
        RECT 2849.340 1361.710 2849.600 1362.030 ;
        RECT 2849.400 1359.050 2849.540 1361.710 ;
        RECT 2843.420 1358.910 2849.540 1359.050 ;
        RECT 2843.420 1269.290 2843.560 1358.910 ;
        RECT 2849.860 1358.370 2850.000 1362.730 ;
        RECT 2844.340 1358.230 2850.000 1358.370 ;
        RECT 2844.340 1357.010 2844.480 1358.230 ;
        RECT 2849.800 1357.630 2850.060 1357.950 ;
        RECT 2843.880 1356.870 2844.480 1357.010 ;
        RECT 2843.880 1314.170 2844.020 1356.870 ;
        RECT 2849.860 1356.330 2850.000 1357.630 ;
        RECT 2844.340 1356.190 2850.000 1356.330 ;
        RECT 2844.340 1314.850 2844.480 1356.190 ;
        RECT 2850.320 1355.820 2850.460 1368.510 ;
        RECT 2844.800 1355.680 2850.460 1355.820 ;
        RECT 2844.800 1315.530 2844.940 1355.680 ;
        RECT 2849.800 1354.970 2850.060 1355.230 ;
        RECT 2845.260 1354.910 2850.060 1354.970 ;
        RECT 2845.260 1354.830 2850.000 1354.910 ;
        RECT 2845.260 1316.210 2845.400 1354.830 ;
        RECT 2850.780 1354.550 2850.920 1387.550 ;
        RECT 2849.800 1354.290 2850.060 1354.550 ;
        RECT 2845.720 1354.230 2850.060 1354.290 ;
        RECT 2850.720 1354.230 2850.980 1354.550 ;
        RECT 2845.720 1354.150 2850.000 1354.230 ;
        RECT 2845.720 1316.890 2845.860 1354.150 ;
        RECT 2851.700 1353.190 2851.840 1389.590 ;
        RECT 2852.160 1363.050 2852.300 1430.195 ;
        RECT 2852.560 1423.085 2852.820 1423.230 ;
        RECT 2852.550 1422.715 2852.830 1423.085 ;
        RECT 2863.660 1364.070 2863.800 1568.915 ;
        RECT 2863.600 1363.750 2863.860 1364.070 ;
        RECT 2852.100 1362.730 2852.360 1363.050 ;
        RECT 2849.800 1352.930 2850.060 1353.190 ;
        RECT 2846.180 1352.870 2850.060 1352.930 ;
        RECT 2851.640 1352.870 2851.900 1353.190 ;
        RECT 2846.180 1352.790 2850.000 1352.870 ;
        RECT 2846.180 1317.570 2846.320 1352.790 ;
        RECT 2849.800 1352.250 2850.060 1352.510 ;
        RECT 2846.640 1352.190 2850.060 1352.250 ;
        RECT 2846.640 1352.110 2850.000 1352.190 ;
        RECT 2846.640 1318.250 2846.780 1352.110 ;
        RECT 2849.800 1350.210 2850.060 1350.470 ;
        RECT 2848.020 1350.150 2850.060 1350.210 ;
        RECT 2848.020 1350.070 2850.000 1350.150 ;
        RECT 2848.020 1331.680 2848.160 1350.070 ;
        RECT 2848.020 1331.540 2849.080 1331.680 ;
        RECT 2848.940 1331.170 2849.080 1331.540 ;
        RECT 2848.940 1331.030 2849.540 1331.170 ;
        RECT 2849.400 1329.640 2849.540 1331.030 ;
        RECT 2849.800 1329.640 2850.060 1329.730 ;
        RECT 2849.400 1329.500 2850.060 1329.640 ;
        RECT 2849.800 1329.410 2850.060 1329.500 ;
        RECT 2846.640 1318.110 2848.620 1318.250 ;
        RECT 2846.180 1317.430 2847.700 1317.570 ;
        RECT 2845.720 1316.750 2847.240 1316.890 ;
        RECT 2845.260 1316.070 2846.780 1316.210 ;
        RECT 2844.800 1315.390 2846.320 1315.530 ;
        RECT 2844.340 1314.710 2845.860 1314.850 ;
        RECT 2843.880 1314.030 2844.480 1314.170 ;
        RECT 2842.960 1269.150 2843.560 1269.290 ;
        RECT 2842.960 1250.930 2843.100 1269.150 ;
        RECT 2844.340 1252.460 2844.480 1314.030 ;
        RECT 2845.720 1280.170 2845.860 1314.710 ;
        RECT 2846.180 1300.685 2846.320 1315.390 ;
        RECT 2846.110 1300.315 2846.390 1300.685 ;
        RECT 2844.800 1280.030 2845.860 1280.170 ;
        RECT 2844.800 1253.140 2844.940 1280.030 ;
        RECT 2846.640 1273.370 2846.780 1316.070 ;
        RECT 2845.260 1273.230 2846.780 1273.370 ;
        RECT 2845.260 1253.650 2845.400 1273.230 ;
        RECT 2847.100 1272.690 2847.240 1316.750 ;
        RECT 2845.720 1272.550 2847.240 1272.690 ;
        RECT 2845.720 1254.330 2845.860 1272.550 ;
        RECT 2847.560 1258.410 2847.700 1317.430 ;
        RECT 2848.480 1262.490 2848.620 1318.110 ;
        RECT 2848.480 1262.350 2850.000 1262.490 ;
        RECT 2849.860 1259.010 2850.000 1262.350 ;
        RECT 2849.800 1258.690 2850.060 1259.010 ;
        RECT 2850.720 1258.690 2850.980 1259.010 ;
        RECT 2847.560 1258.270 2850.000 1258.410 ;
        RECT 2849.860 1254.930 2850.000 1258.270 ;
        RECT 2849.800 1254.610 2850.060 1254.930 ;
        RECT 2845.720 1254.250 2850.000 1254.330 ;
        RECT 2845.720 1254.190 2850.060 1254.250 ;
        RECT 2849.800 1253.930 2850.060 1254.190 ;
        RECT 2845.260 1253.510 2847.240 1253.650 ;
        RECT 2847.100 1253.140 2847.240 1253.510 ;
        RECT 2849.800 1253.140 2850.060 1253.230 ;
        RECT 2844.800 1253.000 2846.780 1253.140 ;
        RECT 2847.100 1253.000 2850.060 1253.140 ;
        RECT 2844.340 1252.320 2846.320 1252.460 ;
        RECT 2842.960 1250.790 2845.860 1250.930 ;
        RECT 2842.040 1218.830 2842.640 1218.970 ;
        RECT 2842.040 1214.890 2842.180 1218.830 ;
        RECT 2845.720 1217.780 2845.860 1250.790 ;
        RECT 2845.260 1217.640 2845.860 1217.780 ;
        RECT 2842.040 1214.750 2843.560 1214.890 ;
        RECT 2843.420 1214.210 2843.560 1214.750 ;
        RECT 2843.420 1214.070 2844.940 1214.210 ;
        RECT 2844.800 1203.330 2844.940 1214.070 ;
        RECT 2845.260 1203.330 2845.400 1217.640 ;
        RECT 2846.180 1204.010 2846.320 1252.320 ;
        RECT 2846.640 1204.690 2846.780 1253.000 ;
        RECT 2849.800 1252.910 2850.060 1253.000 ;
        RECT 2850.260 1232.510 2850.520 1232.830 ;
        RECT 2846.640 1204.550 2848.160 1204.690 ;
        RECT 2846.180 1203.870 2847.700 1204.010 ;
        RECT 2844.800 1203.190 2846.320 1203.330 ;
        RECT 2845.260 1201.970 2845.400 1203.190 ;
        RECT 2846.180 1202.650 2846.320 1203.190 ;
        RECT 2846.180 1202.510 2847.240 1202.650 ;
        RECT 2845.260 1201.830 2846.320 1201.970 ;
        RECT 2846.180 1188.370 2846.320 1201.830 ;
        RECT 2842.960 1188.230 2846.320 1188.370 ;
        RECT 2842.960 1184.970 2843.100 1188.230 ;
        RECT 2841.580 1184.830 2843.560 1184.970 ;
        RECT 2841.120 1184.150 2842.640 1184.290 ;
        RECT 2842.500 1182.930 2842.640 1184.150 ;
        RECT 2842.040 1182.790 2842.640 1182.930 ;
        RECT 2842.040 1180.890 2842.180 1182.790 ;
        RECT 2842.040 1180.750 2842.640 1180.890 ;
        RECT 2842.500 1176.810 2842.640 1180.750 ;
        RECT 2841.580 1176.670 2842.640 1176.810 ;
        RECT 2841.580 1176.130 2841.720 1176.670 ;
        RECT 2842.960 1176.130 2843.100 1184.830 ;
        RECT 2843.420 1182.250 2843.560 1184.830 ;
        RECT 2843.420 1182.110 2844.020 1182.250 ;
        RECT 2841.120 1175.990 2843.100 1176.130 ;
        RECT 2841.120 1044.890 2841.260 1175.990 ;
        RECT 2841.580 1170.690 2841.720 1175.990 ;
        RECT 2841.580 1170.550 2843.100 1170.690 ;
        RECT 2842.960 1155.730 2843.100 1170.550 ;
        RECT 2843.880 1160.490 2844.020 1182.110 ;
        RECT 2843.880 1160.350 2845.400 1160.490 ;
        RECT 2842.500 1155.590 2843.100 1155.730 ;
        RECT 2842.500 1118.330 2842.640 1155.590 ;
        RECT 2845.260 1128.530 2845.400 1160.350 ;
        RECT 2847.100 1158.450 2847.240 1202.510 ;
        RECT 2844.800 1128.390 2845.400 1128.530 ;
        RECT 2846.180 1158.310 2847.240 1158.450 ;
        RECT 2842.500 1118.190 2843.560 1118.330 ;
        RECT 2841.120 1044.750 2841.720 1044.890 ;
        RECT 2841.580 1042.000 2841.720 1044.750 ;
        RECT 2843.420 1042.000 2843.560 1118.190 ;
        RECT 2844.270 1111.530 2844.550 1111.645 ;
        RECT 2844.800 1111.530 2844.940 1128.390 ;
        RECT 2846.180 1127.850 2846.320 1158.310 ;
        RECT 2847.560 1157.770 2847.700 1203.870 ;
        RECT 2848.020 1167.970 2848.160 1204.550 ;
        RECT 2848.020 1167.890 2850.000 1167.970 ;
        RECT 2848.020 1167.830 2850.060 1167.890 ;
        RECT 2849.800 1167.570 2850.060 1167.830 ;
        RECT 2844.270 1111.390 2844.940 1111.530 ;
        RECT 2845.260 1127.710 2846.320 1127.850 ;
        RECT 2846.640 1157.630 2847.700 1157.770 ;
        RECT 2844.270 1111.275 2844.550 1111.390 ;
        RECT 2845.260 1102.690 2845.400 1127.710 ;
        RECT 2844.340 1102.550 2845.400 1102.690 ;
        RECT 2844.340 1047.610 2844.480 1102.550 ;
        RECT 2846.640 1093.850 2846.780 1157.630 ;
        RECT 2849.800 1150.970 2850.060 1151.230 ;
        RECT 2847.560 1150.910 2850.060 1150.970 ;
        RECT 2847.560 1150.830 2850.000 1150.910 ;
        RECT 2847.560 1119.690 2847.700 1150.830 ;
        RECT 2849.800 1149.890 2850.060 1150.210 ;
        RECT 2849.860 1149.610 2850.000 1149.890 ;
        RECT 2848.480 1149.470 2850.000 1149.610 ;
        RECT 2848.480 1121.730 2848.620 1149.470 ;
        RECT 2849.800 1148.930 2850.060 1149.190 ;
        RECT 2848.940 1148.870 2850.060 1148.930 ;
        RECT 2848.940 1148.790 2850.000 1148.870 ;
        RECT 2848.940 1129.040 2849.080 1148.790 ;
        RECT 2850.320 1148.510 2850.460 1232.510 ;
        RECT 2850.780 1197.470 2850.920 1258.690 ;
        RECT 2851.640 1253.930 2851.900 1254.250 ;
        RECT 2850.720 1197.150 2850.980 1197.470 ;
        RECT 2850.720 1167.570 2850.980 1167.890 ;
        RECT 2850.780 1150.210 2850.920 1167.570 ;
        RECT 2850.720 1149.890 2850.980 1150.210 ;
        RECT 2851.700 1149.190 2851.840 1253.930 ;
        RECT 2851.640 1148.870 2851.900 1149.190 ;
        RECT 2850.720 1148.530 2850.980 1148.850 ;
        RECT 2850.260 1148.190 2850.520 1148.510 ;
        RECT 2849.800 1129.040 2850.060 1129.130 ;
        RECT 2848.940 1128.900 2850.060 1129.040 ;
        RECT 2849.800 1128.810 2850.060 1128.900 ;
        RECT 2848.020 1121.590 2848.620 1121.730 ;
        RECT 2848.020 1120.370 2848.160 1121.590 ;
        RECT 2848.020 1120.230 2850.000 1120.370 ;
        RECT 2847.560 1119.550 2849.540 1119.690 ;
        RECT 2844.800 1093.710 2846.780 1093.850 ;
        RECT 2844.800 1048.290 2844.940 1093.710 ;
        RECT 2849.400 1080.250 2849.540 1119.550 ;
        RECT 2845.720 1080.110 2849.540 1080.250 ;
        RECT 2845.720 1048.970 2845.860 1080.110 ;
        RECT 2849.860 1078.470 2850.000 1120.230 ;
        RECT 2849.800 1078.150 2850.060 1078.470 ;
        RECT 2849.800 1077.020 2850.060 1077.110 ;
        RECT 2847.560 1076.880 2850.060 1077.020 ;
        RECT 2845.720 1048.830 2847.240 1048.970 ;
        RECT 2844.800 1048.150 2845.860 1048.290 ;
        RECT 2844.340 1047.470 2844.940 1047.610 ;
        RECT 2844.800 1046.930 2844.940 1047.470 ;
        RECT 2844.800 1046.790 2845.400 1046.930 ;
        RECT 2845.260 1042.850 2845.400 1046.790 ;
        RECT 2843.880 1042.710 2845.400 1042.850 ;
        RECT 2843.880 1042.000 2844.020 1042.710 ;
        RECT 2841.120 1041.860 2844.020 1042.000 ;
        RECT 2841.120 967.370 2841.260 1041.860 ;
        RECT 2841.580 1015.140 2841.720 1041.860 ;
        RECT 2843.420 1041.490 2843.560 1041.860 ;
        RECT 2843.420 1041.350 2844.020 1041.490 ;
        RECT 2843.880 1040.130 2844.020 1041.350 ;
        RECT 2843.420 1039.990 2844.020 1040.130 ;
        RECT 2843.420 1027.890 2843.560 1039.990 ;
        RECT 2845.720 1027.890 2845.860 1048.150 ;
        RECT 2842.500 1027.750 2845.860 1027.890 ;
        RECT 2842.500 1017.010 2842.640 1027.750 ;
        RECT 2843.420 1027.210 2843.560 1027.750 ;
        RECT 2842.960 1027.070 2843.560 1027.210 ;
        RECT 2842.960 1025.850 2843.100 1027.070 ;
        RECT 2847.100 1026.530 2847.240 1048.830 ;
        RECT 2844.800 1026.390 2847.240 1026.530 ;
        RECT 2842.960 1025.710 2843.560 1025.850 ;
        RECT 2843.420 1017.010 2843.560 1025.710 ;
        RECT 2844.800 1019.730 2844.940 1026.390 ;
        RECT 2847.560 1025.170 2847.700 1076.880 ;
        RECT 2849.800 1076.790 2850.060 1076.880 ;
        RECT 2849.800 1073.050 2850.060 1073.370 ;
        RECT 2849.860 1070.730 2850.000 1073.050 ;
        RECT 2850.780 1073.030 2850.920 1148.530 ;
        RECT 2850.720 1072.710 2850.980 1073.030 ;
        RECT 2848.480 1070.590 2850.000 1070.730 ;
        RECT 2848.480 1051.010 2848.620 1070.590 ;
        RECT 2844.340 1019.590 2844.940 1019.730 ;
        RECT 2845.260 1025.030 2847.700 1025.170 ;
        RECT 2848.020 1050.870 2848.620 1051.010 ;
        RECT 2844.340 1017.010 2844.480 1019.590 ;
        RECT 2845.260 1018.370 2845.400 1025.030 ;
        RECT 2848.020 1024.490 2848.160 1050.870 ;
        RECT 2846.180 1024.350 2848.160 1024.490 ;
        RECT 2846.180 1021.600 2846.320 1024.350 ;
        RECT 2849.800 1023.980 2850.060 1024.070 ;
        RECT 2844.800 1018.230 2845.400 1018.370 ;
        RECT 2845.720 1021.460 2846.320 1021.600 ;
        RECT 2846.640 1023.840 2850.060 1023.980 ;
        RECT 2844.800 1017.010 2844.940 1018.230 ;
        RECT 2842.500 1016.870 2843.100 1017.010 ;
        RECT 2843.420 1016.870 2844.020 1017.010 ;
        RECT 2844.340 1016.870 2845.400 1017.010 ;
        RECT 2842.960 1015.140 2843.100 1016.870 ;
        RECT 2843.880 1015.650 2844.020 1016.870 ;
        RECT 2843.880 1015.510 2844.480 1015.650 ;
        RECT 2841.580 1015.000 2844.020 1015.140 ;
        RECT 2842.960 968.165 2843.100 1015.000 ;
        RECT 2842.890 967.795 2843.170 968.165 ;
        RECT 2841.510 967.370 2841.790 967.485 ;
        RECT 2841.120 967.230 2841.790 967.370 ;
        RECT 2841.510 967.115 2841.790 967.230 ;
        RECT 2843.880 959.210 2844.020 1015.000 ;
        RECT 2843.420 959.070 2844.020 959.210 ;
        RECT 2843.420 941.530 2843.560 959.070 ;
        RECT 2844.340 942.040 2844.480 1015.510 ;
        RECT 2842.960 941.390 2843.560 941.530 ;
        RECT 2843.880 941.900 2844.480 942.040 ;
        RECT 2842.960 940.170 2843.100 941.390 ;
        RECT 2843.880 940.170 2844.020 941.900 ;
        RECT 2844.800 941.530 2844.940 1016.870 ;
        RECT 2845.260 942.040 2845.400 1016.870 ;
        RECT 2845.720 958.700 2845.860 1021.460 ;
        RECT 2846.640 1018.540 2846.780 1023.840 ;
        RECT 2849.800 1023.750 2850.060 1023.840 ;
        RECT 2846.180 1018.400 2846.780 1018.540 ;
        RECT 2846.180 959.210 2846.320 1018.400 ;
        RECT 2849.800 1017.860 2850.060 1017.950 ;
        RECT 2846.640 1017.720 2850.060 1017.860 ;
        RECT 2846.640 960.570 2846.780 1017.720 ;
        RECT 2849.800 1017.630 2850.060 1017.720 ;
        RECT 2849.800 1014.970 2850.060 1015.230 ;
        RECT 2848.020 1014.910 2850.060 1014.970 ;
        RECT 2848.020 1014.830 2850.000 1014.910 ;
        RECT 2848.020 962.440 2848.160 1014.830 ;
        RECT 2851.630 967.795 2851.910 968.165 ;
        RECT 2848.020 962.300 2849.540 962.440 ;
        RECT 2849.400 961.930 2849.540 962.300 ;
        RECT 2849.400 961.790 2850.460 961.930 ;
        RECT 2846.640 960.430 2847.240 960.570 ;
        RECT 2847.100 959.890 2847.240 960.430 ;
        RECT 2850.320 960.150 2850.460 961.790 ;
        RECT 2847.100 959.810 2850.000 959.890 ;
        RECT 2850.260 959.830 2850.520 960.150 ;
        RECT 2847.100 959.750 2850.060 959.810 ;
        RECT 2849.800 959.490 2850.060 959.750 ;
        RECT 2846.180 959.070 2851.380 959.210 ;
        RECT 2849.800 958.700 2850.060 958.790 ;
        RECT 2845.720 958.560 2850.060 958.700 ;
        RECT 2849.800 958.470 2850.060 958.560 ;
        RECT 2850.260 958.470 2850.520 958.790 ;
        RECT 2849.800 957.850 2850.060 958.110 ;
        RECT 2846.640 957.790 2850.060 957.850 ;
        RECT 2846.640 957.710 2850.000 957.790 ;
        RECT 2846.640 942.040 2846.780 957.710 ;
        RECT 2849.800 957.110 2850.060 957.430 ;
        RECT 2849.860 956.490 2850.000 957.110 ;
        RECT 2849.400 956.350 2850.000 956.490 ;
        RECT 2849.400 943.570 2849.540 956.350 ;
        RECT 2848.480 943.430 2849.540 943.570 ;
        RECT 2845.260 941.900 2848.160 942.040 ;
        RECT 2844.800 941.390 2845.860 941.530 ;
        RECT 2841.120 940.030 2844.020 940.170 ;
        RECT 2841.120 679.050 2841.260 940.030 ;
        RECT 2842.960 938.810 2843.100 940.030 ;
        RECT 2842.040 938.670 2843.100 938.810 ;
        RECT 2842.040 899.370 2842.180 938.670 ;
        RECT 2845.720 937.450 2845.860 941.390 ;
        RECT 2842.500 937.310 2845.860 937.450 ;
        RECT 2842.500 900.050 2842.640 937.310 ;
        RECT 2846.640 936.090 2846.780 941.900 ;
        RECT 2845.260 935.950 2846.780 936.090 ;
        RECT 2845.260 900.730 2845.400 935.950 ;
        RECT 2845.260 900.590 2845.860 900.730 ;
        RECT 2842.500 899.910 2843.100 900.050 ;
        RECT 2842.960 899.370 2843.100 899.910 ;
        RECT 2842.040 899.230 2842.640 899.370 ;
        RECT 2842.960 899.230 2843.560 899.370 ;
        RECT 2842.500 893.930 2842.640 899.230 ;
        RECT 2841.580 893.790 2842.640 893.930 ;
        RECT 2841.580 816.410 2841.720 893.790 ;
        RECT 2842.500 892.430 2843.100 892.570 ;
        RECT 2842.500 872.965 2842.640 892.430 ;
        RECT 2842.430 872.595 2842.710 872.965 ;
        RECT 2842.960 816.410 2843.100 892.430 ;
        RECT 2843.420 870.130 2843.560 899.230 ;
        RECT 2843.420 869.990 2845.400 870.130 ;
        RECT 2845.260 831.370 2845.400 869.990 ;
        RECT 2845.720 859.930 2845.860 900.590 ;
        RECT 2846.110 892.315 2846.390 892.685 ;
        RECT 2846.180 860.610 2846.320 892.315 ;
        RECT 2848.020 867.410 2848.160 941.900 ;
        RECT 2848.480 935.410 2848.620 943.430 ;
        RECT 2849.800 942.890 2850.060 943.150 ;
        RECT 2848.940 942.830 2850.060 942.890 ;
        RECT 2848.940 942.750 2850.000 942.830 ;
        RECT 2848.940 936.090 2849.080 942.750 ;
        RECT 2848.940 935.950 2849.540 936.090 ;
        RECT 2848.480 935.270 2849.080 935.410 ;
        RECT 2848.940 872.850 2849.080 935.270 ;
        RECT 2849.400 874.890 2849.540 935.950 ;
        RECT 2849.400 874.810 2850.000 874.890 ;
        RECT 2849.400 874.750 2850.060 874.810 ;
        RECT 2849.800 874.490 2850.060 874.750 ;
        RECT 2848.940 872.710 2850.000 872.850 ;
        RECT 2849.860 868.350 2850.000 872.710 ;
        RECT 2849.800 868.030 2850.060 868.350 ;
        RECT 2848.020 867.270 2848.620 867.410 ;
        RECT 2848.480 860.610 2848.620 867.270 ;
        RECT 2849.400 861.150 2850.000 861.290 ;
        RECT 2849.400 860.610 2849.540 861.150 ;
        RECT 2846.180 860.470 2847.700 860.610 ;
        RECT 2848.480 860.470 2849.540 860.610 ;
        RECT 2845.720 859.790 2846.780 859.930 ;
        RECT 2846.640 859.250 2846.780 859.790 ;
        RECT 2846.640 859.110 2847.240 859.250 ;
        RECT 2847.100 851.770 2847.240 859.110 ;
        RECT 2845.720 851.630 2847.240 851.770 ;
        RECT 2845.720 847.690 2845.860 851.630 ;
        RECT 2845.720 847.550 2847.240 847.690 ;
        RECT 2845.260 831.230 2846.780 831.370 ;
        RECT 2841.580 816.270 2843.560 816.410 ;
        RECT 2842.960 815.730 2843.100 816.270 ;
        RECT 2841.580 815.590 2843.100 815.730 ;
        RECT 2841.580 769.490 2841.720 815.590 ;
        RECT 2843.420 811.650 2843.560 816.270 ;
        RECT 2842.960 811.510 2843.560 811.650 ;
        RECT 2842.960 810.290 2843.100 811.510 ;
        RECT 2842.960 810.150 2844.480 810.290 ;
        RECT 2844.340 804.850 2844.480 810.150 ;
        RECT 2843.880 804.710 2844.480 804.850 ;
        RECT 2841.580 769.350 2842.180 769.490 ;
        RECT 2842.040 738.380 2842.180 769.350 ;
        RECT 2843.880 758.610 2844.020 804.710 ;
        RECT 2846.640 776.120 2846.780 831.230 ;
        RECT 2847.100 779.010 2847.240 847.550 ;
        RECT 2847.560 846.330 2847.700 860.470 ;
        RECT 2849.860 846.930 2850.000 861.150 ;
        RECT 2850.320 859.850 2850.460 958.470 ;
        RECT 2851.240 943.150 2851.380 959.070 ;
        RECT 2851.700 958.110 2851.840 967.795 ;
        RECT 2851.640 957.790 2851.900 958.110 ;
        RECT 2851.180 942.830 2851.440 943.150 ;
        RECT 2850.720 868.030 2850.980 868.350 ;
        RECT 2850.260 859.530 2850.520 859.850 ;
        RECT 2849.800 846.610 2850.060 846.930 ;
        RECT 2847.560 846.190 2850.460 846.330 ;
        RECT 2849.800 845.820 2850.060 845.910 ;
        RECT 2847.560 845.680 2850.060 845.820 ;
        RECT 2847.560 781.050 2847.700 845.680 ;
        RECT 2849.800 845.590 2850.060 845.680 ;
        RECT 2849.800 844.910 2850.060 845.230 ;
        RECT 2849.860 819.810 2850.000 844.910 ;
        RECT 2850.320 844.290 2850.460 846.190 ;
        RECT 2850.780 845.230 2850.920 868.030 ;
        RECT 2850.720 844.910 2850.980 845.230 ;
        RECT 2850.320 844.150 2850.920 844.290 ;
        RECT 2848.940 819.670 2850.000 819.810 ;
        RECT 2848.940 787.000 2849.080 819.670 ;
        RECT 2849.800 818.450 2850.060 818.710 ;
        RECT 2849.400 818.390 2850.060 818.450 ;
        RECT 2849.400 818.310 2850.000 818.390 ;
        RECT 2849.400 787.680 2849.540 818.310 ;
        RECT 2850.780 788.450 2850.920 844.150 ;
        RECT 2852.100 810.910 2852.360 811.230 ;
        RECT 2850.720 788.130 2850.980 788.450 ;
        RECT 2849.800 787.680 2850.060 787.770 ;
        RECT 2849.400 787.540 2850.060 787.680 ;
        RECT 2849.800 787.450 2850.060 787.540 ;
        RECT 2850.720 787.450 2850.980 787.770 ;
        RECT 2849.800 787.000 2850.060 787.090 ;
        RECT 2848.940 786.860 2850.060 787.000 ;
        RECT 2849.800 786.770 2850.060 786.860 ;
        RECT 2847.560 780.910 2850.000 781.050 ;
        RECT 2849.860 779.610 2850.000 780.910 ;
        RECT 2849.800 779.290 2850.060 779.610 ;
        RECT 2847.100 778.870 2850.000 779.010 ;
        RECT 2849.860 776.210 2850.000 778.870 ;
        RECT 2846.640 775.980 2849.080 776.120 ;
        RECT 2848.940 775.780 2849.080 775.980 ;
        RECT 2849.800 775.890 2850.060 776.210 ;
        RECT 2849.340 775.780 2849.600 775.870 ;
        RECT 2848.940 775.640 2849.600 775.780 ;
        RECT 2847.100 775.470 2848.160 775.610 ;
        RECT 2849.340 775.550 2849.600 775.640 ;
        RECT 2847.100 758.610 2847.240 775.470 ;
        RECT 2848.020 775.100 2848.160 775.470 ;
        RECT 2850.260 775.210 2850.520 775.530 ;
        RECT 2849.800 775.100 2850.060 775.190 ;
        RECT 2848.020 774.960 2850.060 775.100 ;
        RECT 2849.800 774.870 2850.060 774.960 ;
        RECT 2849.800 774.420 2850.060 774.510 ;
        RECT 2843.420 758.470 2844.020 758.610 ;
        RECT 2844.340 758.470 2847.240 758.610 ;
        RECT 2847.560 774.280 2850.060 774.420 ;
        RECT 2842.040 738.240 2843.100 738.380 ;
        RECT 2842.960 732.770 2843.100 738.240 ;
        RECT 2842.500 732.630 2843.100 732.770 ;
        RECT 2842.500 717.130 2842.640 732.630 ;
        RECT 2843.420 719.850 2843.560 758.470 ;
        RECT 2844.340 757.930 2844.480 758.470 ;
        RECT 2842.040 716.990 2842.640 717.130 ;
        RECT 2842.960 719.710 2843.560 719.850 ;
        RECT 2843.880 757.790 2844.480 757.930 ;
        RECT 2842.040 697.410 2842.180 716.990 ;
        RECT 2842.960 698.090 2843.100 719.710 ;
        RECT 2842.960 697.950 2843.560 698.090 ;
        RECT 2842.040 697.270 2843.100 697.410 ;
        RECT 2841.120 678.910 2842.180 679.050 ;
        RECT 2842.040 607.650 2842.180 678.910 ;
        RECT 2841.580 607.510 2842.180 607.650 ;
        RECT 2841.580 493.410 2841.720 607.510 ;
        RECT 2841.120 493.270 2841.720 493.410 ;
        RECT 2841.120 481.850 2841.260 493.270 ;
        RECT 2842.960 485.250 2843.100 697.270 ;
        RECT 2842.040 485.110 2843.100 485.250 ;
        RECT 2841.120 481.710 2841.720 481.850 ;
        RECT 2841.580 385.970 2841.720 481.710 ;
        RECT 2842.040 469.610 2842.180 485.110 ;
        RECT 2843.420 483.210 2843.560 697.950 ;
        RECT 2842.960 483.070 2843.560 483.210 ;
        RECT 2842.960 480.490 2843.100 483.070 ;
        RECT 2843.880 482.700 2844.020 757.790 ;
        RECT 2847.560 756.570 2847.700 774.280 ;
        RECT 2849.800 774.190 2850.060 774.280 ;
        RECT 2850.320 771.020 2850.460 775.210 ;
        RECT 2842.500 480.350 2843.100 480.490 ;
        RECT 2843.420 482.560 2844.020 482.700 ;
        RECT 2844.340 756.430 2847.700 756.570 ;
        RECT 2849.400 770.880 2850.460 771.020 ;
        RECT 2842.500 475.730 2842.640 480.350 ;
        RECT 2842.500 475.590 2843.100 475.730 ;
        RECT 2842.040 469.470 2842.640 469.610 ;
        RECT 2842.500 428.130 2842.640 469.470 ;
        RECT 2842.960 437.650 2843.100 475.590 ;
        RECT 2843.420 439.010 2843.560 482.560 ;
        RECT 2843.420 438.870 2844.020 439.010 ;
        RECT 2842.960 437.510 2843.560 437.650 ;
        RECT 2842.500 427.990 2843.100 428.130 ;
        RECT 2841.580 385.830 2842.640 385.970 ;
        RECT 2842.500 365.740 2842.640 385.830 ;
        RECT 2841.580 365.600 2842.640 365.740 ;
        RECT 2841.580 200.160 2841.720 365.600 ;
        RECT 2842.960 276.490 2843.100 427.990 ;
        RECT 2843.420 322.050 2843.560 437.510 ;
        RECT 2843.880 322.730 2844.020 438.870 ;
        RECT 2844.340 367.610 2844.480 756.430 ;
        RECT 2849.400 755.890 2849.540 770.880 ;
        RECT 2849.800 769.090 2850.060 769.410 ;
        RECT 2845.720 755.750 2849.540 755.890 ;
        RECT 2845.720 734.980 2845.860 755.750 ;
        RECT 2849.860 747.220 2850.000 769.090 ;
        RECT 2844.800 734.840 2845.860 734.980 ;
        RECT 2846.180 747.080 2850.000 747.220 ;
        RECT 2844.800 368.290 2844.940 734.840 ;
        RECT 2846.180 710.500 2846.320 747.080 ;
        RECT 2849.800 739.740 2850.060 739.830 ;
        RECT 2847.560 739.600 2850.060 739.740 ;
        RECT 2847.560 713.730 2847.700 739.600 ;
        RECT 2849.800 739.510 2850.060 739.600 ;
        RECT 2850.780 739.150 2850.920 787.450 ;
        RECT 2851.180 778.610 2851.440 778.930 ;
        RECT 2851.240 769.410 2851.380 778.610 ;
        RECT 2851.180 769.090 2851.440 769.410 ;
        RECT 2852.160 745.610 2852.300 810.910 ;
        RECT 2851.180 745.290 2851.440 745.610 ;
        RECT 2852.100 745.290 2852.360 745.610 ;
        RECT 2849.800 739.060 2850.060 739.150 ;
        RECT 2847.100 713.590 2847.700 713.730 ;
        RECT 2848.020 738.920 2850.060 739.060 ;
        RECT 2847.100 711.690 2847.240 713.590 ;
        RECT 2845.260 710.360 2846.320 710.500 ;
        RECT 2846.640 711.550 2847.240 711.690 ;
        RECT 2845.260 370.330 2845.400 710.360 ;
        RECT 2846.640 694.010 2846.780 711.550 ;
        RECT 2848.020 711.180 2848.160 738.920 ;
        RECT 2849.800 738.830 2850.060 738.920 ;
        RECT 2850.720 738.830 2850.980 739.150 ;
        RECT 2849.800 738.380 2850.060 738.470 ;
        RECT 2845.720 693.870 2846.780 694.010 ;
        RECT 2847.100 711.040 2848.160 711.180 ;
        RECT 2848.480 738.240 2850.060 738.380 ;
        RECT 2845.720 380.530 2845.860 693.870 ;
        RECT 2847.100 693.330 2847.240 711.040 ;
        RECT 2848.480 710.500 2848.620 738.240 ;
        RECT 2849.800 738.150 2850.060 738.240 ;
        RECT 2846.180 693.190 2847.240 693.330 ;
        RECT 2848.020 710.360 2848.620 710.500 ;
        RECT 2846.180 381.210 2846.320 693.190 ;
        RECT 2848.020 691.290 2848.160 710.360 ;
        RECT 2846.640 691.150 2848.160 691.290 ;
        RECT 2846.640 381.720 2846.780 691.150 ;
        RECT 2851.240 671.830 2851.380 745.290 ;
        RECT 2849.800 671.570 2850.060 671.830 ;
        RECT 2848.020 671.510 2850.060 671.570 ;
        RECT 2851.180 671.510 2851.440 671.830 ;
        RECT 2848.020 671.430 2850.000 671.510 ;
        RECT 2848.020 383.760 2848.160 671.430 ;
        RECT 2851.630 496.555 2851.910 496.925 ;
        RECT 2851.700 450.685 2851.840 496.555 ;
        RECT 2851.630 450.315 2851.910 450.685 ;
        RECT 2848.020 383.620 2848.620 383.760 ;
        RECT 2848.480 383.080 2848.620 383.620 ;
        RECT 2849.400 383.170 2850.000 383.250 ;
        RECT 2849.400 383.110 2850.060 383.170 ;
        RECT 2849.400 383.080 2849.540 383.110 ;
        RECT 2848.480 382.940 2849.540 383.080 ;
        RECT 2849.800 382.850 2850.060 383.110 ;
        RECT 2846.640 381.580 2847.240 381.720 ;
        RECT 2847.100 381.210 2847.240 381.580 ;
        RECT 2846.180 381.070 2846.780 381.210 ;
        RECT 2847.100 381.130 2850.000 381.210 ;
        RECT 2847.100 381.070 2850.060 381.130 ;
        RECT 2846.640 380.530 2846.780 381.070 ;
        RECT 2849.800 380.810 2850.060 381.070 ;
        RECT 2845.720 380.390 2846.320 380.530 ;
        RECT 2846.640 380.390 2847.240 380.530 ;
        RECT 2846.180 379.850 2846.320 380.390 ;
        RECT 2846.180 379.710 2846.780 379.850 ;
        RECT 2846.640 373.560 2846.780 379.710 ;
        RECT 2847.100 374.240 2847.240 380.390 ;
        RECT 2849.800 374.240 2850.060 374.330 ;
        RECT 2847.100 374.100 2850.060 374.240 ;
        RECT 2849.800 374.010 2850.060 374.100 ;
        RECT 2849.800 373.560 2850.060 373.650 ;
        RECT 2846.640 373.420 2850.060 373.560 ;
        RECT 2849.800 373.330 2850.060 373.420 ;
        RECT 2851.180 373.330 2851.440 373.650 ;
        RECT 2845.260 370.190 2850.000 370.330 ;
        RECT 2849.860 368.890 2850.000 370.190 ;
        RECT 2849.800 368.570 2850.060 368.890 ;
        RECT 2844.800 368.210 2850.000 368.290 ;
        RECT 2844.800 368.150 2850.060 368.210 ;
        RECT 2849.800 367.890 2850.060 368.150 ;
        RECT 2844.340 367.470 2850.000 367.610 ;
        RECT 2849.860 367.190 2850.000 367.470 ;
        RECT 2844.800 366.790 2848.620 366.930 ;
        RECT 2849.800 366.870 2850.060 367.190 ;
        RECT 2844.800 323.410 2844.940 366.790 ;
        RECT 2848.480 366.420 2848.620 366.790 ;
        RECT 2851.240 366.510 2851.380 373.330 ;
        RECT 2849.800 366.420 2850.060 366.510 ;
        RECT 2848.480 366.280 2850.060 366.420 ;
        RECT 2845.260 366.110 2847.240 366.250 ;
        RECT 2849.800 366.190 2850.060 366.280 ;
        RECT 2851.180 366.190 2851.440 366.510 ;
        RECT 2845.260 324.090 2845.400 366.110 ;
        RECT 2847.100 365.740 2847.240 366.110 ;
        RECT 2849.800 365.740 2850.060 365.830 ;
        RECT 2847.100 365.600 2850.060 365.740 ;
        RECT 2849.800 365.510 2850.060 365.600 ;
        RECT 2849.800 365.060 2850.060 365.150 ;
        RECT 2848.020 364.920 2850.060 365.060 ;
        RECT 2848.020 340.410 2848.160 364.920 ;
        RECT 2849.800 364.830 2850.060 364.920 ;
        RECT 2849.800 362.340 2850.060 362.430 ;
        RECT 2848.480 362.200 2850.060 362.340 ;
        RECT 2848.480 341.940 2848.620 362.200 ;
        RECT 2849.800 362.110 2850.060 362.200 ;
        RECT 2849.800 341.940 2850.060 342.030 ;
        RECT 2848.480 341.800 2850.060 341.940 ;
        RECT 2849.800 341.710 2850.060 341.800 ;
        RECT 2851.180 341.710 2851.440 342.030 ;
        RECT 2848.020 340.330 2850.000 340.410 ;
        RECT 2848.020 340.270 2850.060 340.330 ;
        RECT 2849.800 340.010 2850.060 340.270 ;
        RECT 2850.720 330.490 2850.980 330.810 ;
        RECT 2845.260 323.950 2850.000 324.090 ;
        RECT 2844.800 323.270 2847.240 323.410 ;
        RECT 2843.880 322.590 2846.780 322.730 ;
        RECT 2843.420 321.910 2844.940 322.050 ;
        RECT 2844.800 320.010 2844.940 321.910 ;
        RECT 2844.800 319.870 2845.860 320.010 ;
        RECT 2845.720 315.930 2845.860 319.870 ;
        RECT 2842.040 276.350 2843.100 276.490 ;
        RECT 2843.420 315.790 2845.860 315.930 ;
        RECT 2842.040 271.730 2842.180 276.350 ;
        RECT 2842.040 271.590 2842.640 271.730 ;
        RECT 2842.500 245.210 2842.640 271.590 ;
        RECT 2843.420 248.610 2843.560 315.790 ;
        RECT 2846.640 315.250 2846.780 322.590 ;
        RECT 2841.120 200.020 2841.720 200.160 ;
        RECT 2842.040 245.070 2842.640 245.210 ;
        RECT 2842.960 248.470 2843.560 248.610 ;
        RECT 2843.880 315.110 2846.780 315.250 ;
        RECT 2.390 89.915 2.670 90.285 ;
        RECT 2.460 51.410 2.600 89.915 ;
        RECT 5.610 64.075 5.890 64.445 ;
        RECT 9.760 64.160 10.020 64.250 ;
        RECT 5.620 63.930 5.880 64.075 ;
        RECT 9.760 64.020 15.940 64.160 ;
        RECT 9.760 63.930 10.020 64.020 ;
        RECT 2.460 51.270 3.520 51.410 ;
        RECT 3.380 3.925 3.520 51.270 ;
        RECT 7.910 43.675 8.190 44.045 ;
        RECT 7.920 43.530 8.180 43.675 ;
        RECT 15.800 6.450 15.940 64.020 ;
        RECT 110.500 8.510 110.760 8.830 ;
        RECT 53.000 6.700 53.260 6.790 ;
        RECT 52.600 6.560 53.260 6.700 ;
        RECT 15.740 6.130 16.000 6.450 ;
        RECT 44.260 6.130 44.520 6.450 ;
        RECT 3.310 3.555 3.590 3.925 ;
        RECT 44.320 2.400 44.460 6.130 ;
        RECT 52.600 4.490 52.740 6.560 ;
        RECT 53.000 6.470 53.260 6.560 ;
        RECT 110.560 4.605 110.700 8.510 ;
        RECT 218.530 7.210 218.810 9.000 ;
        RECT 253.100 8.510 253.360 8.830 ;
        RECT 889.280 8.740 889.540 8.830 ;
        RECT 918.720 8.740 918.980 8.830 ;
        RECT 413.170 8.570 413.450 8.685 ;
        RECT 227.340 7.490 227.600 7.810 ;
        RECT 227.400 7.325 227.540 7.490 ;
        RECT 253.160 7.380 253.300 8.510 ;
        RECT 411.860 8.430 413.450 8.570 ;
        RECT 254.930 7.890 255.210 8.005 ;
        RECT 254.540 7.750 255.210 7.890 ;
        RECT 254.540 7.380 254.680 7.750 ;
        RECT 254.930 7.635 255.210 7.750 ;
        RECT 380.970 7.635 381.250 8.005 ;
        RECT 220.430 7.210 220.710 7.325 ;
        RECT 218.530 7.070 220.710 7.210 ;
        RECT 218.530 5.000 218.810 7.070 ;
        RECT 220.430 6.955 220.710 7.070 ;
        RECT 227.330 6.955 227.610 7.325 ;
        RECT 253.160 7.240 254.680 7.380 ;
        RECT 366.320 5.710 368.300 5.850 ;
        RECT 51.220 4.350 52.740 4.490 ;
        RECT 51.220 3.925 51.360 4.350 ;
        RECT 110.490 4.235 110.770 4.605 ;
        RECT 139.470 4.235 139.750 4.605 ;
        RECT 51.150 3.555 51.430 3.925 ;
        RECT 86.180 2.990 87.240 3.130 ;
        RECT 86.180 2.400 86.320 2.990 ;
        RECT 44.110 -4.800 44.670 2.400 ;
        RECT 49.320 0.525 49.580 0.670 ;
        RECT 49.310 0.155 49.590 0.525 ;
        RECT 85.970 -4.800 86.530 2.400 ;
        RECT 87.100 0.330 87.240 2.990 ;
        RECT 126.660 2.990 127.720 3.130 ;
        RECT 133.500 3.070 133.760 3.390 ;
        RECT 126.660 1.350 126.800 2.990 ;
        RECT 127.580 2.400 127.720 2.990 ;
        RECT 133.560 2.400 133.700 3.070 ;
        RECT 139.540 2.400 139.680 4.235 ;
        RECT 366.320 3.130 366.460 5.710 ;
        RECT 368.160 4.660 368.300 5.710 ;
        RECT 368.160 4.520 372.900 4.660 ;
        RECT 276.160 2.990 277.220 3.130 ;
        RECT 276.160 2.400 276.300 2.990 ;
        RECT 126.600 1.030 126.860 1.350 ;
        RECT 87.040 0.010 87.300 0.330 ;
        RECT 127.370 -4.800 127.930 2.400 ;
        RECT 133.350 -4.800 133.910 2.400 ;
        RECT 139.330 -4.800 139.890 2.400 ;
        RECT 275.950 -4.800 276.510 2.400 ;
        RECT 277.080 0.670 277.220 2.990 ;
        RECT 365.400 2.990 366.460 3.130 ;
        RECT 365.400 2.400 365.540 2.990 ;
        RECT 277.020 0.350 277.280 0.670 ;
        RECT 365.190 -4.800 365.750 2.400 ;
        RECT 372.760 0.525 372.900 4.520 ;
        RECT 381.040 2.565 381.180 7.635 ;
        RECT 411.860 6.450 412.000 8.430 ;
        RECT 413.170 8.315 413.450 8.430 ;
        RECT 603.150 8.570 603.430 8.685 ;
        RECT 603.150 8.430 607.040 8.570 ;
        RECT 603.150 8.315 603.430 8.430 ;
        RECT 512.990 6.530 513.270 6.645 ;
        RECT 393.860 6.360 394.120 6.450 ;
        RECT 392.540 6.220 394.120 6.360 ;
        RECT 382.360 4.430 382.620 4.750 ;
        RECT 382.420 3.810 382.560 4.430 ;
        RECT 382.420 3.670 383.480 3.810 ;
        RECT 380.970 2.195 381.250 2.565 ;
        RECT 383.340 2.400 383.480 3.670 ;
        RECT 392.540 2.565 392.680 6.220 ;
        RECT 393.860 6.130 394.120 6.220 ;
        RECT 411.800 6.130 412.060 6.450 ;
        RECT 512.140 6.390 513.270 6.530 ;
        RECT 424.680 5.790 424.940 6.110 ;
        RECT 419.160 3.410 419.420 3.730 ;
        RECT 407.260 2.990 408.320 3.130 ;
        RECT 372.690 0.155 372.970 0.525 ;
        RECT 383.130 -4.800 383.690 2.400 ;
        RECT 392.470 2.195 392.750 2.565 ;
        RECT 407.260 2.400 407.400 2.990 ;
        RECT 407.050 -4.800 407.610 2.400 ;
        RECT 408.180 0.525 408.320 2.990 ;
        RECT 419.220 2.400 419.360 3.410 ;
        RECT 424.740 2.400 424.880 5.790 ;
        RECT 512.140 5.170 512.280 6.390 ;
        RECT 512.990 6.275 513.270 6.390 ;
        RECT 519.040 6.390 531.600 6.530 ;
        RECT 606.900 6.450 607.040 8.430 ;
        RECT 678.130 8.315 678.410 8.685 ;
        RECT 887.500 8.600 889.540 8.740 ;
        RECT 678.200 8.060 678.340 8.315 ;
        RECT 678.200 7.920 682.480 8.060 ;
        RECT 647.380 7.240 659.940 7.380 ;
        RECT 504.780 5.030 512.280 5.170 ;
        RECT 504.780 4.320 504.920 5.030 ;
        RECT 496.500 4.180 504.920 4.320 ;
        RECT 496.500 2.400 496.640 4.180 ;
        RECT 519.040 3.925 519.180 6.390 ;
        RECT 531.460 6.020 531.600 6.390 ;
        RECT 536.520 6.220 537.580 6.360 ;
        RECT 532.780 6.020 533.040 6.110 ;
        RECT 531.460 5.880 533.040 6.020 ;
        RECT 532.780 5.790 533.040 5.880 ;
        RECT 518.970 3.555 519.250 3.925 ;
        RECT 534.620 3.750 534.880 4.070 ;
        RECT 534.680 2.960 534.820 3.750 ;
        RECT 536.520 2.960 536.660 6.220 ;
        RECT 537.440 6.020 537.580 6.220 ;
        RECT 606.840 6.130 607.100 6.450 ;
        RECT 537.440 5.880 546.320 6.020 ;
        RECT 552.560 5.965 552.820 6.110 ;
        RECT 546.180 5.285 546.320 5.880 ;
        RECT 552.550 5.595 552.830 5.965 ;
        RECT 616.040 5.680 616.300 5.770 ;
        RECT 614.720 5.540 616.300 5.680 ;
        RECT 546.110 4.915 546.390 5.285 ;
        RECT 614.720 5.170 614.860 5.540 ;
        RECT 616.040 5.450 616.300 5.540 ;
        RECT 613.800 5.030 614.860 5.170 ;
        RECT 582.920 4.430 583.180 4.750 ;
        RECT 582.980 3.925 583.120 4.430 ;
        RECT 613.800 3.925 613.940 5.030 ;
        RECT 617.870 4.915 618.150 5.285 ;
        RECT 617.940 4.750 618.080 4.915 ;
        RECT 647.380 4.750 647.520 7.240 ;
        RECT 659.800 7.040 659.940 7.240 ;
        RECT 659.800 6.900 673.740 7.040 ;
        RECT 673.600 6.645 673.740 6.900 ;
        RECT 673.530 6.275 673.810 6.645 ;
        RECT 682.340 6.530 682.480 7.920 ;
        RECT 696.070 6.955 696.350 7.325 ;
        RECT 697.910 6.955 698.190 7.325 ;
        RECT 700.210 6.955 700.490 7.325 ;
        RECT 887.500 7.130 887.640 8.600 ;
        RECT 889.280 8.510 889.540 8.600 ;
        RECT 895.250 8.315 895.530 8.685 ;
        RECT 898.080 8.600 918.980 8.740 ;
        RECT 895.260 8.170 895.520 8.315 ;
        RECT 696.080 6.810 696.340 6.955 ;
        RECT 684.570 6.530 684.850 6.645 ;
        RECT 674.000 6.130 674.260 6.450 ;
        RECT 682.340 6.390 684.850 6.530 ;
        RECT 684.570 6.275 684.850 6.390 ;
        RECT 674.060 5.770 674.200 6.130 ;
        RECT 697.460 6.020 697.720 6.110 ;
        RECT 697.980 6.020 698.120 6.955 ;
        RECT 697.460 5.880 698.120 6.020 ;
        RECT 697.460 5.790 697.720 5.880 ;
        RECT 674.000 5.450 674.260 5.770 ;
        RECT 658.350 4.915 658.630 5.285 ;
        RECT 658.360 4.770 658.620 4.915 ;
        RECT 617.880 4.430 618.140 4.750 ;
        RECT 647.320 4.430 647.580 4.750 ;
        RECT 582.910 3.555 583.190 3.925 ;
        RECT 613.730 3.555 614.010 3.925 ;
        RECT 648.230 3.555 648.510 3.925 ;
        RECT 696.990 3.640 697.270 3.925 ;
        RECT 697.910 3.640 698.190 3.925 ;
        RECT 696.990 3.555 698.190 3.640 ;
        RECT 648.300 3.300 648.440 3.555 ;
        RECT 697.060 3.500 698.120 3.555 ;
        RECT 648.300 3.160 675.580 3.300 ;
        RECT 700.280 3.245 700.420 6.955 ;
        RECT 701.600 6.810 701.860 7.130 ;
        RECT 814.300 6.810 814.560 7.130 ;
        RECT 887.440 6.810 887.700 7.130 ;
        RECT 701.660 5.170 701.800 6.810 ;
        RECT 751.280 6.700 751.540 6.790 ;
        RECT 759.560 6.700 759.820 6.790 ;
        RECT 751.280 6.560 759.820 6.700 ;
        RECT 751.280 6.470 751.540 6.560 ;
        RECT 759.560 6.470 759.820 6.560 ;
        RECT 814.360 6.360 814.500 6.810 ;
        RECT 818.440 6.360 818.700 6.450 ;
        RECT 814.360 6.220 818.700 6.360 ;
        RECT 818.440 6.130 818.700 6.220 ;
        RECT 849.720 6.360 849.980 6.450 ;
        RECT 849.720 6.220 852.220 6.360 ;
        RECT 888.810 6.275 889.090 6.645 ;
        RECT 849.720 6.130 849.980 6.220 ;
        RECT 711.720 5.680 711.980 5.770 ;
        RECT 710.400 5.540 711.980 5.680 ;
        RECT 727.350 5.595 727.630 5.965 ;
        RECT 710.400 5.170 710.540 5.540 ;
        RECT 711.720 5.450 711.980 5.540 ;
        RECT 701.660 5.030 710.540 5.170 ;
        RECT 703.040 4.180 711.920 4.320 ;
        RECT 534.680 2.820 536.660 2.960 ;
        RECT 417.320 0.690 417.580 1.010 ;
        RECT 408.110 0.155 408.390 0.525 ;
        RECT 414.550 0.410 414.830 0.525 ;
        RECT 417.380 0.410 417.520 0.690 ;
        RECT 414.550 0.270 417.520 0.410 ;
        RECT 414.550 0.155 414.830 0.270 ;
        RECT 419.010 -4.800 419.570 2.400 ;
        RECT 421.910 0.835 422.190 1.205 ;
        RECT 420.990 0.410 421.270 0.525 ;
        RECT 421.980 0.410 422.120 0.835 ;
        RECT 420.990 0.270 422.120 0.410 ;
        RECT 420.990 0.155 421.270 0.270 ;
        RECT 424.530 -4.800 425.090 2.400 ;
        RECT 496.290 -4.800 496.850 2.400 ;
        RECT 675.440 1.770 675.580 3.160 ;
        RECT 677.740 2.820 699.500 2.960 ;
        RECT 700.210 2.875 700.490 3.245 ;
        RECT 677.740 1.770 677.880 2.820 ;
        RECT 675.440 1.630 677.880 1.770 ;
        RECT 699.360 1.770 699.500 2.820 ;
        RECT 703.040 1.770 703.180 4.180 ;
        RECT 711.250 3.555 711.530 3.925 ;
        RECT 711.780 3.810 711.920 4.180 ;
        RECT 712.170 3.810 712.450 3.925 ;
        RECT 711.780 3.670 712.450 3.810 ;
        RECT 712.170 3.555 712.450 3.670 ;
        RECT 720.910 3.810 721.190 3.925 ;
        RECT 727.420 3.810 727.560 5.595 ;
        RECT 737.940 5.450 738.200 5.770 ;
        RECT 746.210 5.595 746.490 5.965 ;
        RECT 738.000 3.980 738.140 5.450 ;
        RECT 746.280 3.980 746.420 5.595 ;
        RECT 747.600 4.430 747.860 4.750 ;
        RECT 852.080 4.490 852.220 6.220 ;
        RECT 738.000 3.840 746.420 3.980 ;
        RECT 720.910 3.670 727.560 3.810 ;
        RECT 720.910 3.555 721.190 3.670 ;
        RECT 711.320 3.300 711.460 3.555 ;
        RECT 747.660 3.300 747.800 4.430 ;
        RECT 852.080 4.350 880.740 4.490 ;
        RECT 888.880 4.410 889.020 6.275 ;
        RECT 898.080 4.410 898.220 8.600 ;
        RECT 918.720 8.510 918.980 8.600 ;
        RECT 982.190 8.315 982.470 8.685 ;
        RECT 1238.410 8.570 1238.690 8.685 ;
        RECT 1228.360 8.430 1238.690 8.570 ;
        RECT 982.260 4.490 982.400 8.315 ;
        RECT 1084.380 8.260 1093.260 8.400 ;
        RECT 1070.980 8.060 1071.240 8.150 ;
        RECT 1074.660 8.060 1074.920 8.150 ;
        RECT 1027.270 7.890 1027.550 8.005 ;
        RECT 1023.140 7.490 1023.400 7.810 ;
        RECT 1026.420 7.750 1027.550 7.890 ;
        RECT 1023.200 6.530 1023.340 7.490 ;
        RECT 1021.360 6.390 1023.340 6.530 ;
        RECT 880.600 3.810 880.740 4.350 ;
        RECT 888.820 4.090 889.080 4.410 ;
        RECT 898.020 4.090 898.280 4.410 ;
        RECT 982.260 4.350 985.160 4.490 ;
        RECT 880.990 3.810 881.270 3.925 ;
        RECT 848.340 3.410 848.600 3.730 ;
        RECT 880.600 3.670 881.270 3.810 ;
        RECT 880.990 3.555 881.270 3.670 ;
        RECT 921.010 3.555 921.290 3.925 ;
        RECT 711.320 3.160 711.920 3.300 ;
        RECT 711.780 2.370 711.920 3.160 ;
        RECT 723.740 3.160 747.800 3.300 ;
        RECT 751.280 3.245 751.540 3.390 ;
        RECT 848.400 3.245 848.540 3.410 ;
        RECT 889.740 3.245 890.000 3.390 ;
        RECT 917.800 3.300 918.060 3.390 ;
        RECT 723.740 2.370 723.880 3.160 ;
        RECT 751.270 2.875 751.550 3.245 ;
        RECT 848.330 2.875 848.610 3.245 ;
        RECT 889.730 2.875 890.010 3.245 ;
        RECT 917.400 3.160 918.060 3.300 ;
        RECT 711.720 2.050 711.980 2.370 ;
        RECT 723.680 2.050 723.940 2.370 ;
        RECT 699.360 1.630 703.180 1.770 ;
        RECT 917.400 1.010 917.540 3.160 ;
        RECT 917.800 3.070 918.060 3.160 ;
        RECT 921.080 3.130 921.220 3.555 ;
        RECT 952.820 3.500 955.720 3.640 ;
        RECT 952.820 3.300 952.960 3.500 ;
        RECT 939.020 3.160 952.960 3.300 ;
        RECT 939.020 3.130 939.160 3.160 ;
        RECT 921.080 2.990 939.160 3.130 ;
        RECT 955.580 1.940 955.720 3.500 ;
        RECT 958.340 3.500 968.140 3.640 ;
        RECT 958.340 3.130 958.480 3.500 ;
        RECT 956.960 2.990 958.480 3.130 ;
        RECT 956.960 1.940 957.100 2.990 ;
        RECT 968.000 2.030 968.140 3.500 ;
        RECT 985.020 2.030 985.160 4.350 ;
        RECT 993.230 3.555 993.510 3.925 ;
        RECT 986.790 2.875 987.070 3.245 ;
        RECT 992.310 3.130 992.590 3.245 ;
        RECT 988.700 2.990 992.590 3.130 ;
        RECT 955.580 1.800 957.100 1.940 ;
        RECT 967.940 1.710 968.200 2.030 ;
        RECT 984.960 1.710 985.220 2.030 ;
        RECT 986.860 1.940 987.000 2.875 ;
        RECT 988.700 1.940 988.840 2.990 ;
        RECT 992.310 2.875 992.590 2.990 ;
        RECT 990.930 2.195 991.210 2.565 ;
        RECT 991.000 2.030 991.140 2.195 ;
        RECT 992.320 2.050 992.580 2.370 ;
        RECT 986.860 1.800 988.840 1.940 ;
        RECT 990.940 1.710 991.200 2.030 ;
        RECT 992.380 1.770 992.520 2.050 ;
        RECT 993.300 1.770 993.440 3.555 ;
        RECT 1021.360 3.245 1021.500 6.390 ;
        RECT 1026.420 4.490 1026.560 7.750 ;
        RECT 1027.270 7.635 1027.550 7.750 ;
        RECT 1036.470 7.635 1036.750 8.005 ;
        RECT 1062.760 7.920 1071.240 8.060 ;
        RECT 1036.540 7.210 1036.680 7.635 ;
        RECT 1038.770 7.210 1039.050 7.325 ;
        RECT 1036.540 7.070 1039.050 7.210 ;
        RECT 1038.770 6.955 1039.050 7.070 ;
        RECT 1049.420 7.070 1056.460 7.210 ;
        RECT 1049.420 6.645 1049.560 7.070 ;
        RECT 1049.350 6.275 1049.630 6.645 ;
        RECT 1056.320 6.530 1056.460 7.070 ;
        RECT 1062.760 6.530 1062.900 7.920 ;
        RECT 1070.980 7.830 1071.240 7.920 ;
        RECT 1074.260 7.920 1074.920 8.060 ;
        RECT 1056.320 6.390 1062.900 6.530 ;
        RECT 1073.740 6.470 1074.000 6.790 ;
        RECT 1074.260 6.645 1074.400 7.920 ;
        RECT 1074.660 7.830 1074.920 7.920 ;
        RECT 1082.940 7.890 1083.200 8.150 ;
        RECT 1084.380 7.890 1084.520 8.260 ;
        RECT 1082.940 7.830 1084.520 7.890 ;
        RECT 1083.000 7.750 1084.520 7.830 ;
        RECT 1093.120 7.720 1093.260 8.260 ;
        RECT 1194.710 7.890 1194.990 8.005 ;
        RECT 1125.320 7.750 1128.220 7.890 ;
        RECT 1090.360 7.580 1092.340 7.720 ;
        RECT 1093.120 7.580 1108.440 7.720 ;
        RECT 1090.360 7.130 1090.500 7.580 ;
        RECT 1092.200 7.130 1092.340 7.580 ;
        RECT 1090.300 6.810 1090.560 7.130 ;
        RECT 1092.140 6.810 1092.400 7.130 ;
        RECT 1108.300 6.645 1108.440 7.580 ;
        RECT 1125.320 6.645 1125.460 7.750 ;
        RECT 1073.800 5.850 1073.940 6.470 ;
        RECT 1074.190 6.275 1074.470 6.645 ;
        RECT 1075.110 6.530 1075.390 6.645 ;
        RECT 1074.720 6.390 1075.390 6.530 ;
        RECT 1074.720 5.850 1074.860 6.390 ;
        RECT 1075.110 6.275 1075.390 6.390 ;
        RECT 1087.070 6.275 1087.350 6.645 ;
        RECT 1108.230 6.275 1108.510 6.645 ;
        RECT 1125.250 6.275 1125.530 6.645 ;
        RECT 1127.560 6.470 1127.820 6.790 ;
        RECT 1073.800 5.710 1074.860 5.850 ;
        RECT 1087.140 5.850 1087.280 6.275 ;
        RECT 1089.370 5.850 1089.650 5.965 ;
        RECT 1087.140 5.710 1089.650 5.850 ;
        RECT 1089.370 5.595 1089.650 5.710 ;
        RECT 1124.790 5.595 1125.070 5.965 ;
        RECT 1126.630 5.595 1126.910 5.965 ;
        RECT 1127.620 5.770 1127.760 6.470 ;
        RECT 1128.080 5.850 1128.220 7.750 ;
        RECT 1194.710 7.750 1199.520 7.890 ;
        RECT 1194.710 7.635 1194.990 7.750 ;
        RECT 1152.460 7.070 1158.580 7.210 ;
        RECT 1129.920 6.645 1137.420 6.700 ;
        RECT 1129.920 6.560 1137.490 6.645 ;
        RECT 1129.920 5.850 1130.060 6.560 ;
        RECT 1137.210 6.275 1137.490 6.560 ;
        RECT 1124.860 5.170 1125.000 5.595 ;
        RECT 1126.700 5.170 1126.840 5.595 ;
        RECT 1127.560 5.450 1127.820 5.770 ;
        RECT 1128.080 5.710 1130.060 5.850 ;
        RECT 1133.070 5.850 1133.350 5.965 ;
        RECT 1152.460 5.850 1152.600 7.070 ;
        RECT 1133.070 5.710 1152.600 5.850 ;
        RECT 1133.070 5.595 1133.350 5.710 ;
        RECT 1158.440 5.340 1158.580 7.070 ;
        RECT 1199.380 6.450 1199.520 7.750 ;
        RECT 1162.060 6.130 1162.320 6.450 ;
        RECT 1165.280 6.130 1165.540 6.450 ;
        RECT 1199.320 6.130 1199.580 6.450 ;
        RECT 1206.220 6.130 1206.480 6.450 ;
        RECT 1162.120 5.340 1162.260 6.130 ;
        RECT 1158.440 5.200 1160.420 5.340 ;
        RECT 1124.860 5.030 1126.840 5.170 ;
        RECT 1160.280 5.170 1160.420 5.200 ;
        RECT 1160.740 5.200 1162.260 5.340 ;
        RECT 1160.740 5.170 1160.880 5.200 ;
        RECT 1160.280 5.030 1160.880 5.170 ;
        RECT 1022.740 4.350 1026.560 4.490 ;
        RECT 1088.060 4.350 1098.320 4.490 ;
        RECT 1022.740 3.245 1022.880 4.350 ;
        RECT 1042.980 3.670 1046.800 3.810 ;
        RECT 1021.290 2.875 1021.570 3.245 ;
        RECT 1022.670 2.875 1022.950 3.245 ;
        RECT 1025.430 3.130 1025.710 3.245 ;
        RECT 1042.980 3.130 1043.120 3.670 ;
        RECT 1025.430 2.990 1038.520 3.130 ;
        RECT 1025.430 2.875 1025.710 2.990 ;
        RECT 992.380 1.630 993.440 1.770 ;
        RECT 1038.380 1.770 1038.520 2.990 ;
        RECT 1042.520 2.990 1043.120 3.130 ;
        RECT 1046.660 3.130 1046.800 3.670 ;
        RECT 1088.060 3.390 1088.200 4.350 ;
        RECT 1098.180 3.390 1098.320 4.350 ;
        RECT 1165.340 3.980 1165.480 6.130 ;
        RECT 1206.280 5.850 1206.420 6.130 ;
        RECT 1206.280 5.710 1209.180 5.850 ;
        RECT 1169.020 5.030 1170.080 5.170 ;
        RECT 1169.020 3.980 1169.160 5.030 ;
        RECT 1105.470 3.555 1105.750 3.925 ;
        RECT 1165.340 3.840 1169.160 3.980 ;
        RECT 1105.540 3.390 1105.680 3.555 ;
        RECT 1075.120 3.245 1075.380 3.390 ;
        RECT 1057.170 3.130 1057.450 3.245 ;
        RECT 1046.660 2.990 1057.450 3.130 ;
        RECT 1042.520 1.770 1042.660 2.990 ;
        RECT 1057.170 2.875 1057.450 2.990 ;
        RECT 1075.110 2.875 1075.390 3.245 ;
        RECT 1088.000 3.070 1088.260 3.390 ;
        RECT 1098.120 3.070 1098.380 3.390 ;
        RECT 1105.480 3.070 1105.740 3.390 ;
        RECT 1157.460 3.300 1157.720 3.390 ;
        RECT 1158.380 3.300 1158.640 3.390 ;
        RECT 1157.460 3.160 1158.640 3.300 ;
        RECT 1165.740 3.245 1166.000 3.390 ;
        RECT 1169.940 3.300 1170.080 5.030 ;
        RECT 1192.420 3.750 1192.680 4.070 ;
        RECT 1192.480 3.300 1192.620 3.750 ;
        RECT 1157.460 3.070 1157.720 3.160 ;
        RECT 1158.380 3.070 1158.640 3.160 ;
        RECT 1165.730 2.875 1166.010 3.245 ;
        RECT 1169.940 3.160 1192.620 3.300 ;
        RECT 1209.040 3.300 1209.180 5.710 ;
        RECT 1228.360 3.300 1228.500 8.430 ;
        RECT 1238.410 8.315 1238.690 8.430 ;
        RECT 1396.650 8.315 1396.930 8.685 ;
        RECT 1869.530 8.315 1869.810 8.685 ;
        RECT 1900.810 8.315 1901.090 8.685 ;
        RECT 1283.030 7.635 1283.310 8.005 ;
        RECT 1301.960 7.750 1303.020 7.890 ;
        RECT 1283.100 6.450 1283.240 7.635 ;
        RECT 1301.960 6.450 1302.100 7.750 ;
        RECT 1302.880 7.210 1303.020 7.750 ;
        RECT 1359.390 7.635 1359.670 8.005 ;
        RECT 1303.270 7.210 1303.550 7.325 ;
        RECT 1302.880 7.070 1303.550 7.210 ;
        RECT 1303.270 6.955 1303.550 7.070 ;
        RECT 1340.070 6.955 1340.350 7.325 ;
        RECT 1345.130 7.210 1345.410 7.325 ;
        RECT 1344.740 7.070 1345.410 7.210 ;
        RECT 1283.040 6.130 1283.300 6.450 ;
        RECT 1301.900 6.130 1302.160 6.450 ;
        RECT 1263.710 5.850 1263.990 5.965 ;
        RECT 1265.090 5.850 1265.370 5.965 ;
        RECT 1263.710 5.710 1265.370 5.850 ;
        RECT 1340.140 5.850 1340.280 6.955 ;
        RECT 1344.740 5.850 1344.880 7.070 ;
        RECT 1345.130 6.955 1345.410 7.070 ;
        RECT 1340.140 5.710 1344.880 5.850 ;
        RECT 1263.710 5.595 1263.990 5.710 ;
        RECT 1265.090 5.595 1265.370 5.710 ;
        RECT 1209.040 3.160 1228.500 3.300 ;
        RECT 1238.020 3.245 1242.300 3.300 ;
        RECT 1307.880 3.245 1308.140 3.390 ;
        RECT 1335.020 3.245 1335.280 3.390 ;
        RECT 1237.950 3.160 1242.370 3.245 ;
        RECT 1237.950 2.875 1238.230 3.160 ;
        RECT 1242.090 2.875 1242.370 3.160 ;
        RECT 1307.870 2.875 1308.150 3.245 ;
        RECT 1335.010 2.875 1335.290 3.245 ;
        RECT 1359.460 2.710 1359.600 7.635 ;
        RECT 1396.720 2.710 1396.860 8.315 ;
        RECT 1476.700 7.380 1476.960 7.470 ;
        RECT 1474.920 7.240 1476.960 7.380 ;
        RECT 1474.920 6.645 1475.060 7.240 ;
        RECT 1476.700 7.150 1476.960 7.240 ;
        RECT 1484.060 7.150 1484.320 7.470 ;
        RECT 1499.700 7.150 1499.960 7.470 ;
        RECT 1474.850 6.275 1475.130 6.645 ;
        RECT 1437.590 5.595 1437.870 5.965 ;
        RECT 1483.590 5.850 1483.870 5.965 ;
        RECT 1484.120 5.850 1484.260 7.150 ;
        RECT 1483.590 5.710 1484.260 5.850 ;
        RECT 1483.590 5.595 1483.870 5.710 ;
        RECT 1437.660 4.410 1437.800 5.595 ;
        RECT 1499.760 5.285 1499.900 7.150 ;
        RECT 1614.760 7.070 1624.560 7.210 ;
        RECT 1614.760 6.645 1614.900 7.070 ;
        RECT 1591.690 6.275 1591.970 6.645 ;
        RECT 1593.070 6.275 1593.350 6.645 ;
        RECT 1614.690 6.275 1614.970 6.645 ;
        RECT 1615.610 6.530 1615.890 6.645 ;
        RECT 1615.220 6.390 1615.890 6.530 ;
        RECT 1624.420 6.530 1624.560 7.070 ;
        RECT 1624.810 6.530 1625.090 6.645 ;
        RECT 1624.420 6.390 1625.090 6.530 ;
        RECT 1503.380 5.790 1503.640 6.110 ;
        RECT 1544.770 5.850 1545.050 5.965 ;
        RECT 1499.690 4.915 1499.970 5.285 ;
        RECT 1503.440 5.170 1503.580 5.790 ;
        RECT 1536.560 5.710 1545.050 5.850 ;
        RECT 1517.170 5.170 1517.450 5.285 ;
        RECT 1503.440 5.030 1517.450 5.170 ;
        RECT 1517.170 4.915 1517.450 5.030 ;
        RECT 1534.650 4.915 1534.930 5.285 ;
        RECT 1534.660 4.770 1534.920 4.915 ;
        RECT 1448.240 4.410 1449.300 4.490 ;
        RECT 1437.600 4.090 1437.860 4.410 ;
        RECT 1448.180 4.350 1449.300 4.410 ;
        RECT 1448.180 4.090 1448.440 4.350 ;
        RECT 1449.160 4.320 1449.300 4.350 ;
        RECT 1449.160 4.180 1450.680 4.320 ;
        RECT 1450.540 2.710 1450.680 4.180 ;
        RECT 1536.560 3.810 1536.700 5.710 ;
        RECT 1544.770 5.595 1545.050 5.710 ;
        RECT 1476.760 3.670 1485.180 3.810 ;
        RECT 1469.400 2.990 1472.760 3.130 ;
        RECT 1469.400 2.710 1469.540 2.990 ;
        RECT 1359.400 2.390 1359.660 2.710 ;
        RECT 1396.660 2.390 1396.920 2.710 ;
        RECT 1450.480 2.390 1450.740 2.710 ;
        RECT 1469.340 2.390 1469.600 2.710 ;
        RECT 1472.620 2.450 1472.760 2.990 ;
        RECT 1476.760 2.450 1476.900 3.670 ;
        RECT 1485.040 3.390 1485.180 3.670 ;
        RECT 1503.440 3.670 1536.700 3.810 ;
        RECT 1503.440 3.390 1503.580 3.670 ;
        RECT 1484.980 3.070 1485.240 3.390 ;
        RECT 1503.380 3.070 1503.640 3.390 ;
        RECT 1472.620 2.310 1476.900 2.450 ;
        RECT 1038.380 1.630 1042.660 1.770 ;
        RECT 1591.760 1.770 1591.900 6.275 ;
        RECT 1593.140 5.090 1593.280 6.275 ;
        RECT 1593.080 4.770 1593.340 5.090 ;
        RECT 1615.220 2.370 1615.360 6.390 ;
        RECT 1615.610 6.275 1615.890 6.390 ;
        RECT 1624.810 6.275 1625.090 6.390 ;
        RECT 1637.690 6.275 1637.970 6.645 ;
        RECT 1637.700 6.130 1637.960 6.275 ;
        RECT 1648.280 6.130 1648.540 6.450 ;
        RECT 1648.340 5.850 1648.480 6.130 ;
        RECT 1648.730 5.850 1649.010 5.965 ;
        RECT 1634.540 5.710 1636.060 5.850 ;
        RECT 1648.340 5.710 1649.010 5.850 ;
        RECT 1634.540 5.285 1634.680 5.710 ;
        RECT 1634.470 4.915 1634.750 5.285 ;
        RECT 1635.920 5.170 1636.060 5.710 ;
        RECT 1648.730 5.595 1649.010 5.710 ;
        RECT 1658.850 5.595 1659.130 5.965 ;
        RECT 1784.900 5.790 1785.160 6.110 ;
        RECT 1636.310 5.170 1636.590 5.285 ;
        RECT 1635.920 5.030 1636.590 5.170 ;
        RECT 1658.920 5.090 1659.060 5.595 ;
        RECT 1636.310 4.915 1636.590 5.030 ;
        RECT 1658.860 4.770 1659.120 5.090 ;
        RECT 1678.640 4.770 1678.900 5.090 ;
        RECT 1648.270 4.490 1648.550 4.605 ;
        RECT 1648.740 4.490 1649.000 4.750 ;
        RECT 1648.270 4.430 1649.000 4.490 ;
        RECT 1648.270 4.350 1648.940 4.430 ;
        RECT 1648.270 4.235 1648.550 4.350 ;
        RECT 1678.700 3.810 1678.840 4.770 ;
        RECT 1680.930 4.235 1681.210 4.605 ;
        RECT 1715.440 4.430 1715.700 4.750 ;
        RECT 1747.640 4.605 1747.900 4.750 ;
        RECT 1678.700 3.670 1680.680 3.810 ;
        RECT 1680.540 2.620 1680.680 3.670 ;
        RECT 1681.000 3.245 1681.140 4.235 ;
        RECT 1715.500 3.245 1715.640 4.430 ;
        RECT 1747.630 4.235 1747.910 4.605 ;
        RECT 1782.600 3.750 1782.860 4.070 ;
        RECT 1782.660 3.245 1782.800 3.750 ;
        RECT 1784.960 3.245 1785.100 5.790 ;
        RECT 1862.630 5.595 1862.910 5.965 ;
        RECT 1862.700 4.070 1862.840 5.595 ;
        RECT 1869.600 4.750 1869.740 8.315 ;
        RECT 1900.880 4.750 1901.020 8.315 ;
        RECT 2356.150 7.890 2356.430 9.000 ;
        RECT 2612.890 8.315 2613.170 8.685 ;
        RECT 2357.590 7.890 2357.870 8.005 ;
        RECT 2356.150 7.750 2357.870 7.890 ;
        RECT 2215.910 6.275 2216.190 6.645 ;
        RECT 1946.810 5.595 1947.090 5.965 ;
        RECT 1946.880 4.750 1947.020 5.595 ;
        RECT 1869.540 4.430 1869.800 4.750 ;
        RECT 1900.820 4.430 1901.080 4.750 ;
        RECT 1946.820 4.430 1947.080 4.750 ;
        RECT 1862.640 3.750 1862.900 4.070 ;
        RECT 2031.910 3.555 2032.190 3.925 ;
        RECT 2056.300 3.750 2056.560 4.070 ;
        RECT 2128.520 3.750 2128.780 4.070 ;
        RECT 1680.930 2.875 1681.210 3.245 ;
        RECT 1681.850 3.130 1682.130 3.245 ;
        RECT 1681.460 2.990 1682.130 3.130 ;
        RECT 1681.460 2.620 1681.600 2.990 ;
        RECT 1681.850 2.875 1682.130 2.990 ;
        RECT 1715.430 2.875 1715.710 3.245 ;
        RECT 1782.590 2.875 1782.870 3.245 ;
        RECT 1784.890 2.875 1785.170 3.245 ;
        RECT 1825.370 2.875 1825.650 3.245 ;
        RECT 1930.250 2.875 1930.530 3.245 ;
        RECT 1967.050 2.875 1967.330 3.245 ;
        RECT 1680.540 2.480 1681.600 2.620 ;
        RECT 1594.920 2.050 1595.180 2.370 ;
        RECT 1615.160 2.050 1615.420 2.370 ;
        RECT 1594.980 1.770 1595.120 2.050 ;
        RECT 1825.440 1.885 1825.580 2.875 ;
        RECT 1930.320 1.885 1930.460 2.875 ;
        RECT 1967.120 2.710 1967.260 2.875 ;
        RECT 1967.060 2.390 1967.320 2.710 ;
        RECT 2031.980 1.885 2032.120 3.555 ;
        RECT 2056.360 3.245 2056.500 3.750 ;
        RECT 2056.290 2.875 2056.570 3.245 ;
        RECT 2128.580 1.885 2128.720 3.750 ;
        RECT 2174.970 3.555 2175.250 3.925 ;
        RECT 2174.980 3.410 2175.240 3.555 ;
        RECT 2214.080 3.410 2214.340 3.730 ;
        RECT 2214.140 3.245 2214.280 3.410 ;
        RECT 2214.070 2.875 2214.350 3.245 ;
        RECT 2215.980 1.885 2216.120 6.275 ;
        RECT 2356.150 5.000 2356.430 7.750 ;
        RECT 2357.590 7.635 2357.870 7.750 ;
        RECT 2584.370 6.275 2584.650 6.645 ;
        RECT 2383.820 3.750 2384.080 4.070 ;
        RECT 2430.740 3.750 2431.000 4.070 ;
        RECT 2383.880 3.245 2384.020 3.750 ;
        RECT 2383.810 2.875 2384.090 3.245 ;
        RECT 1591.760 1.630 1595.120 1.770 ;
        RECT 1825.370 1.515 1825.650 1.885 ;
        RECT 1930.250 1.515 1930.530 1.885 ;
        RECT 2031.910 1.515 2032.190 1.885 ;
        RECT 2128.510 1.515 2128.790 1.885 ;
        RECT 2215.910 1.515 2216.190 1.885 ;
        RECT 2430.800 1.205 2430.940 3.750 ;
        RECT 2584.440 3.050 2584.580 6.275 ;
        RECT 2612.960 3.245 2613.100 8.315 ;
        RECT 2688.270 7.210 2688.550 9.000 ;
        RECT 2795.520 8.510 2795.780 8.830 ;
        RECT 2836.460 8.685 2836.720 8.830 ;
        RECT 2795.580 8.005 2795.720 8.510 ;
        RECT 2836.450 8.315 2836.730 8.685 ;
        RECT 2795.510 7.635 2795.790 8.005 ;
        RECT 2686.560 7.070 2688.550 7.210 ;
        RECT 2686.560 6.645 2686.700 7.070 ;
        RECT 2686.490 6.275 2686.770 6.645 ;
        RECT 2688.270 5.000 2688.550 7.070 ;
        RECT 2841.120 5.090 2841.260 200.020 ;
        RECT 2842.040 192.850 2842.180 245.070 ;
        RECT 2842.960 201.010 2843.100 248.470 ;
        RECT 2843.880 202.200 2844.020 315.110 ;
        RECT 2847.100 307.940 2847.240 323.270 ;
        RECT 2849.860 308.710 2850.000 323.950 ;
        RECT 2849.800 308.390 2850.060 308.710 ;
        RECT 2850.780 308.450 2850.920 330.490 ;
        RECT 2850.320 308.310 2850.920 308.450 ;
        RECT 2849.800 307.940 2850.060 308.030 ;
        RECT 2847.100 307.800 2850.060 307.940 ;
        RECT 2849.800 307.710 2850.060 307.800 ;
        RECT 2850.320 307.090 2850.460 308.310 ;
        RECT 2850.720 307.710 2850.980 308.030 ;
        RECT 2844.340 306.950 2850.460 307.090 ;
        RECT 2844.340 205.090 2844.480 306.950 ;
        RECT 2850.260 306.350 2850.520 306.670 ;
        RECT 2849.800 303.690 2850.060 303.950 ;
        RECT 2844.800 303.630 2850.060 303.690 ;
        RECT 2844.800 303.550 2850.000 303.630 ;
        RECT 2844.800 205.600 2844.940 303.550 ;
        RECT 2850.320 303.180 2850.460 306.350 ;
        RECT 2845.260 303.040 2850.460 303.180 ;
        RECT 2845.260 206.450 2845.400 303.040 ;
        RECT 2850.780 301.140 2850.920 307.710 ;
        RECT 2845.720 301.000 2850.920 301.140 ;
        RECT 2845.720 207.130 2845.860 301.000 ;
        RECT 2851.240 300.460 2851.380 341.710 ;
        RECT 2846.180 300.320 2851.380 300.460 ;
        RECT 2846.180 207.810 2846.320 300.320 ;
        RECT 2849.800 299.610 2850.060 299.870 ;
        RECT 2846.640 299.550 2850.060 299.610 ;
        RECT 2846.640 299.470 2850.000 299.550 ;
        RECT 2846.640 208.490 2846.780 299.470 ;
        RECT 2849.800 284.650 2850.060 284.910 ;
        RECT 2848.020 284.590 2850.060 284.650 ;
        RECT 2848.020 284.510 2850.000 284.590 ;
        RECT 2848.020 215.290 2848.160 284.510 ;
        RECT 2848.020 215.150 2849.540 215.290 ;
        RECT 2849.400 211.040 2849.540 215.150 ;
        RECT 2849.800 211.040 2850.060 211.130 ;
        RECT 2849.400 210.900 2850.060 211.040 ;
        RECT 2849.800 210.810 2850.060 210.900 ;
        RECT 2846.640 208.410 2850.000 208.490 ;
        RECT 2846.640 208.350 2850.060 208.410 ;
        RECT 2849.800 208.090 2850.060 208.350 ;
        RECT 2846.180 207.670 2850.000 207.810 ;
        RECT 2845.720 206.990 2847.700 207.130 ;
        RECT 2845.260 206.310 2847.240 206.450 ;
        RECT 2844.800 205.460 2845.860 205.600 ;
        RECT 2844.340 204.950 2844.940 205.090 ;
        RECT 2844.800 203.560 2844.940 204.950 ;
        RECT 2845.720 203.560 2845.860 205.460 ;
        RECT 2847.100 204.410 2847.240 206.310 ;
        RECT 2847.560 204.920 2847.700 206.990 ;
        RECT 2849.860 205.690 2850.000 207.670 ;
        RECT 2849.800 205.370 2850.060 205.690 ;
        RECT 2849.800 204.920 2850.060 205.010 ;
        RECT 2847.560 204.780 2850.060 204.920 ;
        RECT 2849.800 204.690 2850.060 204.780 ;
        RECT 2847.100 204.270 2850.920 204.410 ;
        RECT 2849.800 203.560 2850.060 203.650 ;
        RECT 2844.800 203.420 2845.400 203.560 ;
        RECT 2845.720 203.420 2850.060 203.560 ;
        RECT 2845.260 203.050 2845.400 203.420 ;
        RECT 2849.800 203.330 2850.060 203.420 ;
        RECT 2845.260 202.910 2850.460 203.050 ;
        RECT 2849.800 202.200 2850.060 202.290 ;
        RECT 2843.880 202.060 2850.060 202.200 ;
        RECT 2849.800 201.970 2850.060 202.060 ;
        RECT 2849.800 201.520 2850.060 201.610 ;
        RECT 2844.340 201.380 2850.060 201.520 ;
        RECT 2844.340 201.010 2844.480 201.380 ;
        RECT 2849.800 201.290 2850.060 201.380 ;
        RECT 2842.960 200.870 2844.480 201.010 ;
        RECT 2849.800 200.840 2850.060 200.930 ;
        RECT 2846.180 200.700 2850.060 200.840 ;
        RECT 2846.180 198.290 2846.320 200.700 ;
        RECT 2849.800 200.610 2850.060 200.700 ;
        RECT 2849.800 200.160 2850.060 200.250 ;
        RECT 2844.340 198.150 2846.320 198.290 ;
        RECT 2847.100 200.020 2850.060 200.160 ;
        RECT 2844.340 197.100 2844.480 198.150 ;
        RECT 2844.340 196.960 2845.400 197.100 ;
        RECT 2842.040 192.710 2842.640 192.850 ;
        RECT 2842.500 33.050 2842.640 192.710 ;
        RECT 2845.260 156.810 2845.400 196.960 ;
        RECT 2847.100 196.250 2847.240 200.020 ;
        RECT 2849.800 199.930 2850.060 200.020 ;
        RECT 2849.800 199.480 2850.060 199.570 ;
        RECT 2844.340 156.670 2845.400 156.810 ;
        RECT 2845.720 196.110 2847.240 196.250 ;
        RECT 2847.560 199.340 2850.060 199.480 ;
        RECT 2844.340 156.130 2844.480 156.670 ;
        RECT 2843.880 155.990 2844.480 156.130 ;
        RECT 2843.880 154.090 2844.020 155.990 ;
        RECT 2843.880 153.950 2845.400 154.090 ;
        RECT 2845.260 150.690 2845.400 153.950 ;
        RECT 2842.960 150.550 2845.400 150.690 ;
        RECT 2842.960 123.490 2843.100 150.550 ;
        RECT 2845.720 150.010 2845.860 196.110 ;
        RECT 2847.560 177.210 2847.700 199.340 ;
        RECT 2849.800 199.250 2850.060 199.340 ;
        RECT 2850.320 198.970 2850.460 202.910 ;
        RECT 2848.480 198.830 2850.460 198.970 ;
        RECT 2848.480 198.290 2848.620 198.830 ;
        RECT 2849.800 198.460 2850.060 198.550 ;
        RECT 2849.400 198.320 2850.060 198.460 ;
        RECT 2849.400 198.290 2849.540 198.320 ;
        RECT 2843.420 149.870 2845.860 150.010 ;
        RECT 2846.640 177.070 2847.700 177.210 ;
        RECT 2848.020 198.150 2848.620 198.290 ;
        RECT 2848.940 198.150 2849.540 198.290 ;
        RECT 2849.800 198.230 2850.060 198.320 ;
        RECT 2843.420 124.340 2843.560 149.870 ;
        RECT 2846.640 148.650 2846.780 177.070 ;
        RECT 2848.020 176.530 2848.160 198.150 ;
        RECT 2843.880 148.510 2846.780 148.650 ;
        RECT 2847.100 176.390 2848.160 176.530 ;
        RECT 2843.880 125.700 2844.020 148.510 ;
        RECT 2847.100 128.250 2847.240 176.390 ;
        RECT 2848.940 175.850 2849.080 198.150 ;
        RECT 2850.780 197.610 2850.920 204.270 ;
        RECT 2847.560 175.710 2849.080 175.850 ;
        RECT 2849.400 197.470 2850.920 197.610 ;
        RECT 2847.560 131.650 2847.700 175.710 ;
        RECT 2849.400 132.500 2849.540 197.470 ;
        RECT 2849.800 196.870 2850.060 197.190 ;
        RECT 2849.860 141.850 2850.000 196.870 ;
        RECT 2851.640 173.750 2851.900 174.070 ;
        RECT 2849.860 141.710 2850.460 141.850 ;
        RECT 2849.800 132.500 2850.060 132.590 ;
        RECT 2849.400 132.360 2850.060 132.500 ;
        RECT 2849.800 132.270 2850.060 132.360 ;
        RECT 2847.560 131.510 2850.000 131.650 ;
        RECT 2849.860 128.850 2850.000 131.510 ;
        RECT 2849.800 128.530 2850.060 128.850 ;
        RECT 2847.100 128.110 2850.000 128.250 ;
        RECT 2849.860 127.830 2850.000 128.110 ;
        RECT 2849.800 127.510 2850.060 127.830 ;
        RECT 2849.800 125.700 2850.060 125.790 ;
        RECT 2843.880 125.560 2850.060 125.700 ;
        RECT 2849.800 125.470 2850.060 125.560 ;
        RECT 2843.420 124.200 2844.940 124.340 ;
        RECT 2842.960 123.350 2844.480 123.490 ;
        RECT 2844.340 93.570 2844.480 123.350 ;
        RECT 2841.580 32.910 2842.640 33.050 ;
        RECT 2843.420 93.430 2844.480 93.570 ;
        RECT 2841.580 8.830 2841.720 32.910 ;
        RECT 2843.420 24.890 2843.560 93.430 ;
        RECT 2844.800 92.210 2844.940 124.200 ;
        RECT 2849.800 121.620 2850.060 121.710 ;
        RECT 2842.040 24.750 2843.560 24.890 ;
        RECT 2843.880 92.070 2844.940 92.210 ;
        RECT 2845.260 121.480 2850.060 121.620 ;
        RECT 2841.520 8.510 2841.780 8.830 ;
        RECT 2841.520 7.830 2841.780 8.150 ;
        RECT 2841.580 6.790 2841.720 7.830 ;
        RECT 2841.520 6.470 2841.780 6.790 ;
        RECT 2842.040 5.965 2842.180 24.750 ;
        RECT 2843.880 24.210 2844.020 92.070 ;
        RECT 2845.260 80.650 2845.400 121.480 ;
        RECT 2849.800 121.390 2850.060 121.480 ;
        RECT 2849.800 120.770 2850.060 121.030 ;
        RECT 2842.960 24.070 2844.020 24.210 ;
        RECT 2844.340 80.510 2845.400 80.650 ;
        RECT 2845.720 120.710 2850.060 120.770 ;
        RECT 2845.720 120.630 2850.000 120.710 ;
        RECT 2842.960 11.290 2843.100 24.070 ;
        RECT 2842.500 11.150 2843.100 11.290 ;
        RECT 2842.500 7.810 2842.640 11.150 ;
        RECT 2844.340 9.930 2844.480 80.510 ;
        RECT 2845.720 79.970 2845.860 120.630 ;
        RECT 2849.800 118.730 2850.060 118.990 ;
        RECT 2843.420 9.790 2844.480 9.930 ;
        RECT 2844.800 79.830 2845.860 79.970 ;
        RECT 2846.180 118.670 2850.060 118.730 ;
        RECT 2846.180 118.590 2850.000 118.670 ;
        RECT 2843.420 8.150 2843.560 9.790 ;
        RECT 2844.800 8.570 2844.940 79.830 ;
        RECT 2846.180 79.290 2846.320 118.590 ;
        RECT 2845.260 79.150 2846.320 79.290 ;
        RECT 2847.100 117.970 2850.000 118.050 ;
        RECT 2847.100 117.910 2850.060 117.970 ;
        RECT 2845.260 9.170 2845.400 79.150 ;
        RECT 2847.100 78.610 2847.240 117.910 ;
        RECT 2849.800 117.650 2850.060 117.910 ;
        RECT 2850.320 116.690 2850.460 141.710 ;
        RECT 2851.180 125.470 2851.440 125.790 ;
        RECT 2851.240 117.970 2851.380 125.470 ;
        RECT 2851.700 121.710 2851.840 173.750 ;
        RECT 2851.640 121.390 2851.900 121.710 ;
        RECT 2851.180 117.650 2851.440 117.970 ;
        RECT 2848.940 116.550 2850.460 116.690 ;
        RECT 2848.940 90.170 2849.080 116.550 ;
        RECT 2848.020 90.030 2849.080 90.170 ;
        RECT 2848.020 89.660 2848.160 90.030 ;
        RECT 2846.180 78.470 2847.240 78.610 ;
        RECT 2847.560 89.520 2848.160 89.660 ;
        RECT 2846.180 77.930 2846.320 78.470 ;
        RECT 2845.720 77.790 2846.320 77.930 ;
        RECT 2845.200 8.850 2845.460 9.170 ;
        RECT 2844.800 8.430 2845.400 8.570 ;
        RECT 2843.360 7.830 2843.620 8.150 ;
        RECT 2842.440 7.490 2842.700 7.810 ;
        RECT 2843.820 7.490 2844.080 7.810 ;
        RECT 2843.880 6.530 2844.020 7.490 ;
        RECT 2843.420 6.390 2844.020 6.530 ;
        RECT 2841.970 5.595 2842.250 5.965 ;
        RECT 2843.420 5.285 2843.560 6.390 ;
        RECT 2841.060 4.770 2841.320 5.090 ;
        RECT 2843.350 4.915 2843.630 5.285 ;
        RECT 2684.650 3.810 2684.930 3.925 ;
        RECT 2683.800 3.670 2684.930 3.810 ;
        RECT 2683.800 3.245 2683.940 3.670 ;
        RECT 2684.650 3.555 2684.930 3.670 ;
        RECT 2549.420 2.730 2549.680 3.050 ;
        RECT 2584.380 2.730 2584.640 3.050 ;
        RECT 2612.890 2.875 2613.170 3.245 ;
        RECT 2683.730 2.875 2684.010 3.245 ;
        RECT 2845.260 3.130 2845.400 8.430 ;
        RECT 2845.720 3.925 2845.860 77.790 ;
        RECT 2847.560 77.250 2847.700 89.520 ;
        RECT 2849.800 88.300 2850.060 88.390 ;
        RECT 2846.180 77.110 2847.700 77.250 ;
        RECT 2848.480 88.160 2850.060 88.300 ;
        RECT 2846.180 34.410 2846.320 77.110 ;
        RECT 2848.480 61.610 2848.620 88.160 ;
        RECT 2849.800 88.070 2850.060 88.160 ;
        RECT 2851.640 73.450 2851.900 73.770 ;
        RECT 2851.700 61.725 2851.840 73.450 ;
        RECT 2848.020 61.470 2848.620 61.610 ;
        RECT 2848.020 48.010 2848.160 61.470 ;
        RECT 2851.630 61.355 2851.910 61.725 ;
        RECT 2848.020 47.870 2848.620 48.010 ;
        RECT 2848.480 43.250 2848.620 47.870 ;
        RECT 2848.480 43.170 2850.000 43.250 ;
        RECT 2848.480 43.110 2850.060 43.170 ;
        RECT 2849.800 42.850 2850.060 43.110 ;
        RECT 2851.640 42.850 2851.900 43.170 ;
        RECT 2846.180 34.270 2847.240 34.410 ;
        RECT 2846.120 8.850 2846.380 9.170 ;
        RECT 2845.650 3.555 2845.930 3.925 ;
        RECT 2844.340 2.990 2845.400 3.130 ;
        RECT 2549.480 2.565 2549.620 2.730 ;
        RECT 2549.410 2.195 2549.690 2.565 ;
        RECT 2728.350 2.195 2728.630 2.565 ;
        RECT 2728.420 1.205 2728.560 2.195 ;
        RECT 917.340 0.690 917.600 1.010 ;
        RECT 2366.790 0.835 2367.070 1.205 ;
        RECT 2368.630 0.835 2368.910 1.205 ;
        RECT 2430.730 0.835 2431.010 1.205 ;
        RECT 2728.350 0.835 2728.630 1.205 ;
        RECT 2366.860 0.330 2367.000 0.835 ;
        RECT 2368.700 0.330 2368.840 0.835 ;
        RECT 2844.340 0.670 2844.480 2.990 ;
        RECT 2846.180 1.010 2846.320 8.850 ;
        RECT 2847.100 4.750 2847.240 34.270 ;
        RECT 2851.700 22.285 2851.840 42.850 ;
        RECT 2851.630 21.915 2851.910 22.285 ;
        RECT 2847.040 4.430 2847.300 4.750 ;
        RECT 2846.120 0.690 2846.380 1.010 ;
        RECT 2844.280 0.350 2844.540 0.670 ;
        RECT 2366.800 0.010 2367.060 0.330 ;
        RECT 2368.640 0.010 2368.900 0.330 ;
      LAYER via2 ;
        RECT 2773.890 3402.240 2774.170 3402.520 ;
        RECT 2863.590 3200.960 2863.870 3201.240 ;
        RECT 2851.630 3062.240 2851.910 3062.520 ;
        RECT 2863.590 2928.960 2863.870 2929.240 ;
        RECT 2900.850 2669.200 2901.130 2669.480 ;
        RECT 2851.630 2382.240 2851.910 2382.520 ;
        RECT 2863.590 2112.960 2863.870 2113.240 ;
        RECT 2851.630 1974.240 2851.910 1974.520 ;
        RECT 2851.630 1838.240 2851.910 1838.520 ;
        RECT 2863.590 1704.960 2863.870 1705.240 ;
        RECT 2863.590 1568.960 2863.870 1569.240 ;
        RECT 2852.090 1430.240 2852.370 1430.520 ;
        RECT 2841.970 1241.880 2842.250 1242.160 ;
        RECT 2852.550 1422.760 2852.830 1423.040 ;
        RECT 2846.110 1300.360 2846.390 1300.640 ;
        RECT 2844.270 1111.320 2844.550 1111.600 ;
        RECT 2842.890 967.840 2843.170 968.120 ;
        RECT 2841.510 967.160 2841.790 967.440 ;
        RECT 2851.630 967.840 2851.910 968.120 ;
        RECT 2842.430 872.640 2842.710 872.920 ;
        RECT 2846.110 892.360 2846.390 892.640 ;
        RECT 2851.630 496.600 2851.910 496.880 ;
        RECT 2851.630 450.360 2851.910 450.640 ;
        RECT 2.390 89.960 2.670 90.240 ;
        RECT 5.610 64.120 5.890 64.400 ;
        RECT 7.910 43.720 8.190 44.000 ;
        RECT 3.310 3.600 3.590 3.880 ;
        RECT 254.930 7.680 255.210 7.960 ;
        RECT 380.970 7.680 381.250 7.960 ;
        RECT 220.430 7.000 220.710 7.280 ;
        RECT 227.330 7.000 227.610 7.280 ;
        RECT 110.490 4.280 110.770 4.560 ;
        RECT 139.470 4.280 139.750 4.560 ;
        RECT 51.150 3.600 51.430 3.880 ;
        RECT 49.310 0.200 49.590 0.480 ;
        RECT 413.170 8.360 413.450 8.640 ;
        RECT 603.150 8.360 603.430 8.640 ;
        RECT 380.970 2.240 381.250 2.520 ;
        RECT 372.690 0.200 372.970 0.480 ;
        RECT 392.470 2.240 392.750 2.520 ;
        RECT 512.990 6.320 513.270 6.600 ;
        RECT 678.130 8.360 678.410 8.640 ;
        RECT 518.970 3.600 519.250 3.880 ;
        RECT 552.550 5.640 552.830 5.920 ;
        RECT 546.110 4.960 546.390 5.240 ;
        RECT 617.870 4.960 618.150 5.240 ;
        RECT 673.530 6.320 673.810 6.600 ;
        RECT 696.070 7.000 696.350 7.280 ;
        RECT 697.910 7.000 698.190 7.280 ;
        RECT 700.210 7.000 700.490 7.280 ;
        RECT 895.250 8.360 895.530 8.640 ;
        RECT 684.570 6.320 684.850 6.600 ;
        RECT 658.350 4.960 658.630 5.240 ;
        RECT 582.910 3.600 583.190 3.880 ;
        RECT 613.730 3.600 614.010 3.880 ;
        RECT 648.230 3.600 648.510 3.880 ;
        RECT 696.990 3.600 697.270 3.880 ;
        RECT 697.910 3.600 698.190 3.880 ;
        RECT 888.810 6.320 889.090 6.600 ;
        RECT 727.350 5.640 727.630 5.920 ;
        RECT 408.110 0.200 408.390 0.480 ;
        RECT 414.550 0.200 414.830 0.480 ;
        RECT 421.910 0.880 422.190 1.160 ;
        RECT 420.990 0.200 421.270 0.480 ;
        RECT 700.210 2.920 700.490 3.200 ;
        RECT 711.250 3.600 711.530 3.880 ;
        RECT 712.170 3.600 712.450 3.880 ;
        RECT 720.910 3.600 721.190 3.880 ;
        RECT 746.210 5.640 746.490 5.920 ;
        RECT 982.190 8.360 982.470 8.640 ;
        RECT 880.990 3.600 881.270 3.880 ;
        RECT 921.010 3.600 921.290 3.880 ;
        RECT 751.270 2.920 751.550 3.200 ;
        RECT 848.330 2.920 848.610 3.200 ;
        RECT 889.730 2.920 890.010 3.200 ;
        RECT 993.230 3.600 993.510 3.880 ;
        RECT 986.790 2.920 987.070 3.200 ;
        RECT 992.310 2.920 992.590 3.200 ;
        RECT 990.930 2.240 991.210 2.520 ;
        RECT 1027.270 7.680 1027.550 7.960 ;
        RECT 1036.470 7.680 1036.750 7.960 ;
        RECT 1038.770 7.000 1039.050 7.280 ;
        RECT 1049.350 6.320 1049.630 6.600 ;
        RECT 1074.190 6.320 1074.470 6.600 ;
        RECT 1075.110 6.320 1075.390 6.600 ;
        RECT 1087.070 6.320 1087.350 6.600 ;
        RECT 1108.230 6.320 1108.510 6.600 ;
        RECT 1125.250 6.320 1125.530 6.600 ;
        RECT 1089.370 5.640 1089.650 5.920 ;
        RECT 1124.790 5.640 1125.070 5.920 ;
        RECT 1126.630 5.640 1126.910 5.920 ;
        RECT 1194.710 7.680 1194.990 7.960 ;
        RECT 1137.210 6.320 1137.490 6.600 ;
        RECT 1133.070 5.640 1133.350 5.920 ;
        RECT 1021.290 2.920 1021.570 3.200 ;
        RECT 1022.670 2.920 1022.950 3.200 ;
        RECT 1025.430 2.920 1025.710 3.200 ;
        RECT 1105.470 3.600 1105.750 3.880 ;
        RECT 1057.170 2.920 1057.450 3.200 ;
        RECT 1075.110 2.920 1075.390 3.200 ;
        RECT 1165.730 2.920 1166.010 3.200 ;
        RECT 1238.410 8.360 1238.690 8.640 ;
        RECT 1396.650 8.360 1396.930 8.640 ;
        RECT 1869.530 8.360 1869.810 8.640 ;
        RECT 1900.810 8.360 1901.090 8.640 ;
        RECT 1283.030 7.680 1283.310 7.960 ;
        RECT 1359.390 7.680 1359.670 7.960 ;
        RECT 1303.270 7.000 1303.550 7.280 ;
        RECT 1340.070 7.000 1340.350 7.280 ;
        RECT 1263.710 5.640 1263.990 5.920 ;
        RECT 1265.090 5.640 1265.370 5.920 ;
        RECT 1345.130 7.000 1345.410 7.280 ;
        RECT 1237.950 2.920 1238.230 3.200 ;
        RECT 1242.090 2.920 1242.370 3.200 ;
        RECT 1307.870 2.920 1308.150 3.200 ;
        RECT 1335.010 2.920 1335.290 3.200 ;
        RECT 1474.850 6.320 1475.130 6.600 ;
        RECT 1437.590 5.640 1437.870 5.920 ;
        RECT 1483.590 5.640 1483.870 5.920 ;
        RECT 1591.690 6.320 1591.970 6.600 ;
        RECT 1593.070 6.320 1593.350 6.600 ;
        RECT 1614.690 6.320 1614.970 6.600 ;
        RECT 1499.690 4.960 1499.970 5.240 ;
        RECT 1517.170 4.960 1517.450 5.240 ;
        RECT 1534.650 4.960 1534.930 5.240 ;
        RECT 1544.770 5.640 1545.050 5.920 ;
        RECT 1615.610 6.320 1615.890 6.600 ;
        RECT 1624.810 6.320 1625.090 6.600 ;
        RECT 1637.690 6.320 1637.970 6.600 ;
        RECT 1634.470 4.960 1634.750 5.240 ;
        RECT 1648.730 5.640 1649.010 5.920 ;
        RECT 1658.850 5.640 1659.130 5.920 ;
        RECT 1636.310 4.960 1636.590 5.240 ;
        RECT 1648.270 4.280 1648.550 4.560 ;
        RECT 1680.930 4.280 1681.210 4.560 ;
        RECT 1747.630 4.280 1747.910 4.560 ;
        RECT 1862.630 5.640 1862.910 5.920 ;
        RECT 2612.890 8.360 2613.170 8.640 ;
        RECT 2215.910 6.320 2216.190 6.600 ;
        RECT 1946.810 5.640 1947.090 5.920 ;
        RECT 2031.910 3.600 2032.190 3.880 ;
        RECT 1680.930 2.920 1681.210 3.200 ;
        RECT 1681.850 2.920 1682.130 3.200 ;
        RECT 1715.430 2.920 1715.710 3.200 ;
        RECT 1782.590 2.920 1782.870 3.200 ;
        RECT 1784.890 2.920 1785.170 3.200 ;
        RECT 1825.370 2.920 1825.650 3.200 ;
        RECT 1930.250 2.920 1930.530 3.200 ;
        RECT 1967.050 2.920 1967.330 3.200 ;
        RECT 2056.290 2.920 2056.570 3.200 ;
        RECT 2174.970 3.600 2175.250 3.880 ;
        RECT 2214.070 2.920 2214.350 3.200 ;
        RECT 2357.590 7.680 2357.870 7.960 ;
        RECT 2584.370 6.320 2584.650 6.600 ;
        RECT 2383.810 2.920 2384.090 3.200 ;
        RECT 1825.370 1.560 1825.650 1.840 ;
        RECT 1930.250 1.560 1930.530 1.840 ;
        RECT 2031.910 1.560 2032.190 1.840 ;
        RECT 2128.510 1.560 2128.790 1.840 ;
        RECT 2215.910 1.560 2216.190 1.840 ;
        RECT 2836.450 8.360 2836.730 8.640 ;
        RECT 2795.510 7.680 2795.790 7.960 ;
        RECT 2686.490 6.320 2686.770 6.600 ;
        RECT 2841.970 5.640 2842.250 5.920 ;
        RECT 2843.350 4.960 2843.630 5.240 ;
        RECT 2684.650 3.600 2684.930 3.880 ;
        RECT 2612.890 2.920 2613.170 3.200 ;
        RECT 2683.730 2.920 2684.010 3.200 ;
        RECT 2851.630 61.400 2851.910 61.680 ;
        RECT 2845.650 3.600 2845.930 3.880 ;
        RECT 2549.410 2.240 2549.690 2.520 ;
        RECT 2728.350 2.240 2728.630 2.520 ;
        RECT 2366.790 0.880 2367.070 1.160 ;
        RECT 2368.630 0.880 2368.910 1.160 ;
        RECT 2430.730 0.880 2431.010 1.160 ;
        RECT 2728.350 0.880 2728.630 1.160 ;
        RECT 2851.630 21.960 2851.910 22.240 ;
      LAYER met3 ;
        RECT 2798.910 3403.890 2799.290 3403.900 ;
        RECT 2787.910 3403.590 2799.290 3403.890 ;
        RECT 2773.865 3402.530 2774.195 3402.545 ;
        RECT 2787.910 3402.530 2788.210 3403.590 ;
        RECT 2798.910 3403.580 2799.290 3403.590 ;
        RECT 2773.865 3402.230 2788.210 3402.530 ;
        RECT 2773.865 3402.215 2774.195 3402.230 ;
        RECT 2851.000 3201.250 2855.000 3201.640 ;
        RECT 2863.565 3201.250 2863.895 3201.265 ;
        RECT 2851.000 3201.040 2863.895 3201.250 ;
        RECT 2854.300 3200.950 2863.895 3201.040 ;
        RECT 2863.565 3200.935 2863.895 3200.950 ;
        RECT 2851.000 3065.040 2855.000 3065.640 ;
        RECT 2851.390 3062.545 2851.690 3065.040 ;
        RECT 2851.390 3062.230 2851.935 3062.545 ;
        RECT 2851.605 3062.215 2851.935 3062.230 ;
        RECT 2851.000 2929.250 2855.000 2929.640 ;
        RECT 2863.565 2929.250 2863.895 2929.265 ;
        RECT 2851.000 2929.040 2863.895 2929.250 ;
        RECT 2854.300 2928.950 2863.895 2929.040 ;
        RECT 2863.565 2928.935 2863.895 2928.950 ;
        RECT 2900.825 2669.490 2901.155 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2900.825 2669.190 2924.800 2669.490 ;
        RECT 2900.825 2669.175 2901.155 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
        RECT 2851.000 2385.040 2855.000 2385.640 ;
        RECT 2851.390 2382.545 2851.690 2385.040 ;
        RECT 2851.390 2382.230 2851.935 2382.545 ;
        RECT 2851.605 2382.215 2851.935 2382.230 ;
        RECT 2851.000 2113.250 2855.000 2113.640 ;
        RECT 2863.565 2113.250 2863.895 2113.265 ;
        RECT 2851.000 2113.040 2863.895 2113.250 ;
        RECT 2854.300 2112.950 2863.895 2113.040 ;
        RECT 2863.565 2112.935 2863.895 2112.950 ;
        RECT 2851.000 1977.040 2855.000 1977.640 ;
        RECT 2851.390 1974.545 2851.690 1977.040 ;
        RECT 2851.390 1974.230 2851.935 1974.545 ;
        RECT 2851.605 1974.215 2851.935 1974.230 ;
        RECT 2851.000 1841.040 2855.000 1841.640 ;
        RECT 2851.390 1838.545 2851.690 1841.040 ;
        RECT 2851.390 1838.230 2851.935 1838.545 ;
        RECT 2851.605 1838.215 2851.935 1838.230 ;
        RECT 2851.000 1705.250 2855.000 1705.640 ;
        RECT 2863.565 1705.250 2863.895 1705.265 ;
        RECT 2851.000 1705.040 2863.895 1705.250 ;
        RECT 2854.300 1704.950 2863.895 1705.040 ;
        RECT 2863.565 1704.935 2863.895 1704.950 ;
        RECT 2851.000 1569.250 2855.000 1569.640 ;
        RECT 2863.565 1569.250 2863.895 1569.265 ;
        RECT 2851.000 1569.040 2863.895 1569.250 ;
        RECT 2854.300 1568.950 2863.895 1569.040 ;
        RECT 2863.565 1568.935 2863.895 1568.950 ;
        RECT 2851.000 1433.040 2855.000 1433.640 ;
        RECT 2852.310 1430.545 2852.610 1433.040 ;
        RECT 2852.065 1430.230 2852.610 1430.545 ;
        RECT 2852.065 1430.215 2852.395 1430.230 ;
        RECT 2852.525 1423.060 2852.855 1423.065 ;
        RECT 2852.270 1423.050 2852.855 1423.060 ;
        RECT 2852.270 1422.750 2853.080 1423.050 ;
        RECT 2852.270 1422.740 2852.855 1422.750 ;
        RECT 2852.525 1422.735 2852.855 1422.740 ;
        RECT 2851.605 968.140 2851.935 968.145 ;
        RECT 2851.350 968.130 2851.935 968.140 ;
        RECT 2851.350 967.830 2852.160 968.130 ;
        RECT 2851.350 967.820 2851.935 967.830 ;
        RECT 2851.605 967.815 2851.935 967.820 ;
        RECT 2852.270 967.450 2852.650 967.460 ;
        RECT 2853.190 967.450 2853.570 967.460 ;
        RECT 2852.270 967.150 2853.570 967.450 ;
        RECT 2852.270 967.140 2852.650 967.150 ;
        RECT 2853.190 967.140 2853.570 967.150 ;
        RECT 2846.180 892.360 2846.390 892.640 ;
        RECT 2851.605 496.900 2851.935 496.905 ;
        RECT 2851.350 496.890 2851.935 496.900 ;
        RECT 2851.350 496.590 2852.160 496.890 ;
        RECT 2851.350 496.580 2851.935 496.590 ;
        RECT 2851.605 496.575 2851.935 496.580 ;
        RECT 2851.605 450.650 2851.935 450.665 ;
        RECT 2852.270 450.650 2852.650 450.660 ;
        RECT 2851.605 450.350 2852.650 450.650 ;
        RECT 2851.605 450.335 2851.935 450.350 ;
        RECT 2852.270 450.340 2852.650 450.350 ;
        RECT 2.365 90.250 2.695 90.265 ;
        RECT 7.630 90.250 8.010 90.260 ;
        RECT 2.365 89.950 8.010 90.250 ;
        RECT 2.365 89.935 2.695 89.950 ;
        RECT 7.630 89.940 8.010 89.950 ;
        RECT 4.870 64.410 5.250 64.420 ;
        RECT 5.585 64.410 5.915 64.425 ;
        RECT 4.870 64.110 5.915 64.410 ;
        RECT 4.870 64.100 5.250 64.110 ;
        RECT 5.585 64.095 5.915 64.110 ;
        RECT 2851.605 61.700 2851.935 61.705 ;
        RECT 2851.350 61.690 2851.935 61.700 ;
        RECT 2851.350 61.390 2852.160 61.690 ;
        RECT 2851.350 61.380 2851.935 61.390 ;
        RECT 2851.605 61.375 2851.935 61.380 ;
        RECT 7.885 44.020 8.215 44.025 ;
        RECT 7.630 44.010 8.215 44.020 ;
        RECT 7.630 43.710 8.440 44.010 ;
        RECT 7.630 43.700 8.215 43.710 ;
        RECT 7.885 43.695 8.215 43.700 ;
        RECT 2851.605 22.250 2851.935 22.265 ;
        RECT 2852.270 22.250 2852.650 22.260 ;
        RECT 2851.605 21.950 2852.650 22.250 ;
        RECT 2851.605 21.935 2851.935 21.950 ;
        RECT 2852.270 21.940 2852.650 21.950 ;
        RECT 413.145 8.650 413.475 8.665 ;
        RECT 417.950 8.650 418.330 8.660 ;
        RECT 413.145 8.350 418.330 8.650 ;
        RECT 413.145 8.335 413.475 8.350 ;
        RECT 417.950 8.340 418.330 8.350 ;
        RECT 428.990 8.650 429.370 8.660 ;
        RECT 440.030 8.650 440.410 8.660 ;
        RECT 428.990 8.350 440.410 8.650 ;
        RECT 428.990 8.340 429.370 8.350 ;
        RECT 440.030 8.340 440.410 8.350 ;
        RECT 557.790 8.650 558.170 8.660 ;
        RECT 603.125 8.650 603.455 8.665 ;
        RECT 678.105 8.660 678.435 8.665 ;
        RECT 557.790 8.350 603.455 8.650 ;
        RECT 557.790 8.340 558.170 8.350 ;
        RECT 603.125 8.335 603.455 8.350 ;
        RECT 629.550 8.650 629.930 8.660 ;
        RECT 639.670 8.650 640.050 8.660 ;
        RECT 629.550 8.350 640.050 8.650 ;
        RECT 629.550 8.340 629.930 8.350 ;
        RECT 639.670 8.340 640.050 8.350 ;
        RECT 678.105 8.650 678.690 8.660 ;
        RECT 895.225 8.650 895.555 8.665 ;
        RECT 974.550 8.650 974.930 8.660 ;
        RECT 982.165 8.650 982.495 8.665 ;
        RECT 678.105 8.350 678.890 8.650 ;
        RECT 895.225 8.350 924.290 8.650 ;
        RECT 678.105 8.340 678.690 8.350 ;
        RECT 678.105 8.335 678.435 8.340 ;
        RECT 895.225 8.335 895.555 8.350 ;
        RECT 254.905 7.970 255.235 7.985 ;
        RECT 261.550 7.970 261.930 7.980 ;
        RECT 254.905 7.670 261.930 7.970 ;
        RECT 254.905 7.655 255.235 7.670 ;
        RECT 261.550 7.660 261.930 7.670 ;
        RECT 377.470 7.970 377.850 7.980 ;
        RECT 380.945 7.970 381.275 7.985 ;
        RECT 377.470 7.670 381.275 7.970 ;
        RECT 377.470 7.660 377.850 7.670 ;
        RECT 380.945 7.655 381.275 7.670 ;
        RECT 509.030 7.970 509.410 7.980 ;
        RECT 516.390 7.970 516.770 7.980 ;
        RECT 509.030 7.670 516.770 7.970 ;
        RECT 923.990 7.970 924.290 8.350 ;
        RECT 974.550 8.350 982.495 8.650 ;
        RECT 974.550 8.340 974.930 8.350 ;
        RECT 982.165 8.335 982.495 8.350 ;
        RECT 1084.030 8.650 1084.410 8.660 ;
        RECT 1101.510 8.650 1101.890 8.660 ;
        RECT 1084.030 8.350 1101.890 8.650 ;
        RECT 1084.030 8.340 1084.410 8.350 ;
        RECT 1101.510 8.340 1101.890 8.350 ;
        RECT 1171.430 8.650 1171.810 8.660 ;
        RECT 1189.830 8.650 1190.210 8.660 ;
        RECT 1171.430 8.350 1190.210 8.650 ;
        RECT 1171.430 8.340 1171.810 8.350 ;
        RECT 1189.830 8.340 1190.210 8.350 ;
        RECT 1238.385 8.650 1238.715 8.665 ;
        RECT 1396.625 8.650 1396.955 8.665 ;
        RECT 1428.110 8.650 1428.490 8.660 ;
        RECT 1238.385 8.350 1249.970 8.650 ;
        RECT 1238.385 8.335 1238.715 8.350 ;
        RECT 952.470 7.970 952.850 7.980 ;
        RECT 992.030 7.970 992.410 7.980 ;
        RECT 923.990 7.670 952.850 7.970 ;
        RECT 509.030 7.660 509.410 7.670 ;
        RECT 516.390 7.660 516.770 7.670 ;
        RECT 952.470 7.660 952.850 7.670 ;
        RECT 986.550 7.670 992.410 7.970 ;
        RECT 220.405 7.290 220.735 7.305 ;
        RECT 227.305 7.290 227.635 7.305 ;
        RECT 220.405 6.990 227.635 7.290 ;
        RECT 220.405 6.975 220.735 6.990 ;
        RECT 227.305 6.975 227.635 6.990 ;
        RECT 514.550 6.980 514.930 7.300 ;
        RECT 675.550 7.290 675.930 7.300 ;
        RECT 674.670 6.990 675.930 7.290 ;
        RECT 512.965 6.610 513.295 6.625 ;
        RECT 514.590 6.610 514.890 6.980 ;
        RECT 512.965 6.310 514.890 6.610 ;
        RECT 673.505 6.610 673.835 6.625 ;
        RECT 674.670 6.610 674.970 6.990 ;
        RECT 675.550 6.980 675.930 6.990 ;
        RECT 693.950 7.290 694.330 7.300 ;
        RECT 696.045 7.290 696.375 7.305 ;
        RECT 693.950 6.990 696.375 7.290 ;
        RECT 693.950 6.980 694.330 6.990 ;
        RECT 696.045 6.975 696.375 6.990 ;
        RECT 697.885 7.290 698.215 7.305 ;
        RECT 700.185 7.290 700.515 7.305 ;
        RECT 697.885 6.990 700.515 7.290 ;
        RECT 697.885 6.975 698.215 6.990 ;
        RECT 700.185 6.975 700.515 6.990 ;
        RECT 808.030 7.290 808.410 7.300 ;
        RECT 819.990 7.290 820.370 7.300 ;
        RECT 808.030 6.990 820.370 7.290 ;
        RECT 808.030 6.980 808.410 6.990 ;
        RECT 819.990 6.980 820.370 6.990 ;
        RECT 955.230 7.290 955.610 7.300 ;
        RECT 986.550 7.290 986.850 7.670 ;
        RECT 992.030 7.660 992.410 7.670 ;
        RECT 1027.245 7.970 1027.575 7.985 ;
        RECT 1036.445 7.970 1036.775 7.985 ;
        RECT 1193.510 7.970 1193.890 7.980 ;
        RECT 1194.685 7.970 1195.015 7.985 ;
        RECT 1027.245 7.670 1036.775 7.970 ;
        RECT 1027.245 7.655 1027.575 7.670 ;
        RECT 1036.445 7.655 1036.775 7.670 ;
        RECT 1038.070 7.670 1050.330 7.970 ;
        RECT 955.230 6.990 986.850 7.290 ;
        RECT 1002.150 7.290 1002.530 7.300 ;
        RECT 1038.070 7.290 1038.370 7.670 ;
        RECT 1002.150 6.990 1038.370 7.290 ;
        RECT 1038.745 7.290 1039.075 7.305 ;
        RECT 1050.030 7.290 1050.330 7.670 ;
        RECT 1193.510 7.670 1195.015 7.970 ;
        RECT 1249.670 7.970 1249.970 8.350 ;
        RECT 1396.625 8.350 1428.490 8.650 ;
        RECT 1396.625 8.335 1396.955 8.350 ;
        RECT 1428.110 8.340 1428.490 8.350 ;
        RECT 1869.505 8.650 1869.835 8.665 ;
        RECT 1900.785 8.650 1901.115 8.665 ;
        RECT 1869.505 8.350 1901.115 8.650 ;
        RECT 1869.505 8.335 1869.835 8.350 ;
        RECT 1900.785 8.335 1901.115 8.350 ;
        RECT 2566.150 8.650 2566.530 8.660 ;
        RECT 2612.865 8.650 2613.195 8.665 ;
        RECT 2566.150 8.350 2613.195 8.650 ;
        RECT 2566.150 8.340 2566.530 8.350 ;
        RECT 2612.865 8.335 2613.195 8.350 ;
        RECT 2836.425 8.650 2836.755 8.665 ;
        RECT 2845.830 8.650 2846.210 8.660 ;
        RECT 2836.425 8.350 2846.210 8.650 ;
        RECT 2836.425 8.335 2836.755 8.350 ;
        RECT 2845.830 8.340 2846.210 8.350 ;
        RECT 1268.950 7.970 1269.330 7.980 ;
        RECT 1283.005 7.970 1283.335 7.985 ;
        RECT 1359.365 7.970 1359.695 7.985 ;
        RECT 1249.670 7.670 1265.610 7.970 ;
        RECT 1193.510 7.660 1193.890 7.670 ;
        RECT 1194.685 7.655 1195.015 7.670 ;
        RECT 1054.590 7.290 1054.970 7.300 ;
        RECT 1038.745 6.990 1041.130 7.290 ;
        RECT 1050.030 6.990 1054.970 7.290 ;
        RECT 1265.310 7.290 1265.610 7.670 ;
        RECT 1268.950 7.670 1283.335 7.970 ;
        RECT 1268.950 7.660 1269.330 7.670 ;
        RECT 1283.005 7.655 1283.335 7.670 ;
        RECT 1355.470 7.670 1359.695 7.970 ;
        RECT 1303.245 7.300 1303.575 7.305 ;
        RECT 1267.110 7.290 1267.490 7.300 ;
        RECT 1265.310 6.990 1267.490 7.290 ;
        RECT 955.230 6.980 955.610 6.990 ;
        RECT 1002.150 6.980 1002.530 6.990 ;
        RECT 1038.745 6.975 1039.075 6.990 ;
        RECT 684.545 6.620 684.875 6.625 ;
        RECT 684.545 6.610 685.130 6.620 ;
        RECT 673.505 6.310 674.970 6.610 ;
        RECT 684.320 6.310 685.130 6.610 ;
        RECT 512.965 6.295 513.295 6.310 ;
        RECT 673.505 6.295 673.835 6.310 ;
        RECT 684.545 6.300 685.130 6.310 ;
        RECT 881.630 6.610 882.010 6.620 ;
        RECT 888.785 6.610 889.115 6.625 ;
        RECT 881.630 6.310 889.115 6.610 ;
        RECT 1040.830 6.610 1041.130 6.990 ;
        RECT 1054.590 6.980 1054.970 6.990 ;
        RECT 1267.110 6.980 1267.490 6.990 ;
        RECT 1302.990 7.290 1303.575 7.300 ;
        RECT 1304.830 7.290 1305.210 7.300 ;
        RECT 1340.045 7.290 1340.375 7.305 ;
        RECT 1302.990 6.990 1303.800 7.290 ;
        RECT 1304.830 6.990 1340.375 7.290 ;
        RECT 1302.990 6.980 1303.575 6.990 ;
        RECT 1304.830 6.980 1305.210 6.990 ;
        RECT 1303.245 6.975 1303.575 6.980 ;
        RECT 1340.045 6.975 1340.375 6.990 ;
        RECT 1345.105 7.290 1345.435 7.305 ;
        RECT 1355.470 7.290 1355.770 7.670 ;
        RECT 1359.365 7.655 1359.695 7.670 ;
        RECT 2357.565 7.970 2357.895 7.985 ;
        RECT 2795.485 7.980 2795.815 7.985 ;
        RECT 2794.310 7.970 2794.690 7.980 ;
        RECT 2795.230 7.970 2795.815 7.980 ;
        RECT 2357.565 7.670 2794.690 7.970 ;
        RECT 2795.030 7.670 2795.815 7.970 ;
        RECT 2357.565 7.655 2357.895 7.670 ;
        RECT 2794.310 7.660 2794.690 7.670 ;
        RECT 2795.230 7.660 2795.815 7.670 ;
        RECT 2795.485 7.655 2795.815 7.660 ;
        RECT 1345.105 6.990 1355.770 7.290 ;
        RECT 1402.350 7.290 1402.730 7.300 ;
        RECT 1402.350 6.990 1406.370 7.290 ;
        RECT 1345.105 6.975 1345.435 6.990 ;
        RECT 1402.350 6.980 1402.730 6.990 ;
        RECT 1049.325 6.610 1049.655 6.625 ;
        RECT 1074.165 6.620 1074.495 6.625 ;
        RECT 1073.910 6.610 1074.495 6.620 ;
        RECT 1040.830 6.310 1049.655 6.610 ;
        RECT 1073.710 6.310 1074.495 6.610 ;
        RECT 881.630 6.300 882.010 6.310 ;
        RECT 684.545 6.295 684.875 6.300 ;
        RECT 888.785 6.295 889.115 6.310 ;
        RECT 1049.325 6.295 1049.655 6.310 ;
        RECT 1073.910 6.300 1074.495 6.310 ;
        RECT 1074.165 6.295 1074.495 6.300 ;
        RECT 1075.085 6.610 1075.415 6.625 ;
        RECT 1087.045 6.610 1087.375 6.625 ;
        RECT 1075.085 6.310 1087.375 6.610 ;
        RECT 1075.085 6.295 1075.415 6.310 ;
        RECT 1087.045 6.295 1087.375 6.310 ;
        RECT 1108.205 6.610 1108.535 6.625 ;
        RECT 1125.225 6.610 1125.555 6.625 ;
        RECT 1137.185 6.620 1137.515 6.625 ;
        RECT 1137.185 6.610 1137.770 6.620 ;
        RECT 1108.205 6.310 1125.555 6.610 ;
        RECT 1136.960 6.310 1137.770 6.610 ;
        RECT 1108.205 6.295 1108.535 6.310 ;
        RECT 1125.225 6.295 1125.555 6.310 ;
        RECT 1137.185 6.300 1137.770 6.310 ;
        RECT 1138.310 6.610 1138.690 6.620 ;
        RECT 1145.670 6.610 1146.050 6.620 ;
        RECT 1138.310 6.310 1146.050 6.610 ;
        RECT 1138.310 6.300 1138.690 6.310 ;
        RECT 1145.670 6.300 1146.050 6.310 ;
        RECT 1314.030 6.610 1314.410 6.620 ;
        RECT 1324.150 6.610 1324.530 6.620 ;
        RECT 1314.030 6.310 1324.530 6.610 ;
        RECT 1406.070 6.610 1406.370 6.990 ;
        RECT 1474.110 6.610 1474.490 6.620 ;
        RECT 1474.825 6.610 1475.155 6.625 ;
        RECT 1406.070 6.310 1438.570 6.610 ;
        RECT 1314.030 6.300 1314.410 6.310 ;
        RECT 1324.150 6.300 1324.530 6.310 ;
        RECT 1137.185 6.295 1137.515 6.300 ;
        RECT 462.110 5.930 462.490 5.940 ;
        RECT 506.270 5.930 506.650 5.940 ;
        RECT 462.110 5.630 506.650 5.930 ;
        RECT 462.110 5.620 462.490 5.630 ;
        RECT 506.270 5.620 506.650 5.630 ;
        RECT 552.525 5.930 552.855 5.945 ;
        RECT 556.870 5.930 557.250 5.940 ;
        RECT 552.525 5.630 557.250 5.930 ;
        RECT 552.525 5.615 552.855 5.630 ;
        RECT 556.870 5.620 557.250 5.630 ;
        RECT 634.150 5.930 634.530 5.940 ;
        RECT 641.510 5.930 641.890 5.940 ;
        RECT 634.150 5.630 641.890 5.930 ;
        RECT 634.150 5.620 634.530 5.630 ;
        RECT 641.510 5.620 641.890 5.630 ;
        RECT 727.325 5.930 727.655 5.945 ;
        RECT 737.190 5.930 737.570 5.940 ;
        RECT 727.325 5.630 737.570 5.930 ;
        RECT 727.325 5.615 727.655 5.630 ;
        RECT 737.190 5.620 737.570 5.630 ;
        RECT 746.185 5.930 746.515 5.945 ;
        RECT 753.750 5.930 754.130 5.940 ;
        RECT 746.185 5.630 754.130 5.930 ;
        RECT 746.185 5.615 746.515 5.630 ;
        RECT 753.750 5.620 754.130 5.630 ;
        RECT 1089.345 5.930 1089.675 5.945 ;
        RECT 1124.765 5.930 1125.095 5.945 ;
        RECT 1089.345 5.630 1125.095 5.930 ;
        RECT 1089.345 5.615 1089.675 5.630 ;
        RECT 1124.765 5.615 1125.095 5.630 ;
        RECT 1126.605 5.930 1126.935 5.945 ;
        RECT 1133.045 5.930 1133.375 5.945 ;
        RECT 1126.605 5.630 1133.375 5.930 ;
        RECT 1126.605 5.615 1126.935 5.630 ;
        RECT 1133.045 5.615 1133.375 5.630 ;
        RECT 1133.710 5.930 1134.090 5.940 ;
        RECT 1263.685 5.930 1264.015 5.945 ;
        RECT 1133.710 5.630 1264.015 5.930 ;
        RECT 1133.710 5.620 1134.090 5.630 ;
        RECT 1263.685 5.615 1264.015 5.630 ;
        RECT 1265.065 5.930 1265.395 5.945 ;
        RECT 1344.390 5.930 1344.770 5.940 ;
        RECT 1265.065 5.630 1344.770 5.930 ;
        RECT 1265.065 5.615 1265.395 5.630 ;
        RECT 1344.390 5.620 1344.770 5.630 ;
        RECT 1397.750 5.930 1398.130 5.940 ;
        RECT 1437.565 5.930 1437.895 5.945 ;
        RECT 1397.750 5.630 1437.895 5.930 ;
        RECT 1397.750 5.620 1398.130 5.630 ;
        RECT 1437.565 5.615 1437.895 5.630 ;
        RECT 546.085 5.250 546.415 5.265 ;
        RECT 617.845 5.250 618.175 5.265 ;
        RECT 546.085 4.950 618.175 5.250 ;
        RECT 546.085 4.935 546.415 4.950 ;
        RECT 617.845 4.935 618.175 4.950 ;
        RECT 658.325 5.250 658.655 5.265 ;
        RECT 677.390 5.250 677.770 5.260 ;
        RECT 658.325 4.950 677.770 5.250 ;
        RECT 1438.270 5.250 1438.570 6.310 ;
        RECT 1474.110 6.310 1475.155 6.610 ;
        RECT 1474.110 6.300 1474.490 6.310 ;
        RECT 1474.825 6.295 1475.155 6.310 ;
        RECT 1589.110 6.610 1589.490 6.620 ;
        RECT 1591.665 6.610 1591.995 6.625 ;
        RECT 1589.110 6.310 1591.995 6.610 ;
        RECT 1589.110 6.300 1589.490 6.310 ;
        RECT 1591.665 6.295 1591.995 6.310 ;
        RECT 1593.045 6.610 1593.375 6.625 ;
        RECT 1614.665 6.610 1614.995 6.625 ;
        RECT 1593.045 6.310 1614.995 6.610 ;
        RECT 1593.045 6.295 1593.375 6.310 ;
        RECT 1614.665 6.295 1614.995 6.310 ;
        RECT 1615.585 6.610 1615.915 6.625 ;
        RECT 1624.070 6.610 1624.450 6.620 ;
        RECT 1615.585 6.310 1624.450 6.610 ;
        RECT 1615.585 6.295 1615.915 6.310 ;
        RECT 1624.070 6.300 1624.450 6.310 ;
        RECT 1624.785 6.610 1625.115 6.625 ;
        RECT 1637.665 6.610 1637.995 6.625 ;
        RECT 2215.885 6.610 2216.215 6.625 ;
        RECT 1624.785 6.310 1637.995 6.610 ;
        RECT 1624.785 6.295 1625.115 6.310 ;
        RECT 1637.665 6.295 1637.995 6.310 ;
        RECT 2197.270 6.310 2216.215 6.610 ;
        RECT 1448.350 5.930 1448.730 5.940 ;
        RECT 1450.190 5.930 1450.570 5.940 ;
        RECT 1483.565 5.930 1483.895 5.945 ;
        RECT 1448.350 5.630 1450.570 5.930 ;
        RECT 1448.350 5.620 1448.730 5.630 ;
        RECT 1450.190 5.620 1450.570 5.630 ;
        RECT 1452.990 5.630 1483.895 5.930 ;
        RECT 1452.990 5.250 1453.290 5.630 ;
        RECT 1483.565 5.615 1483.895 5.630 ;
        RECT 1544.745 5.930 1545.075 5.945 ;
        RECT 1648.705 5.930 1649.035 5.945 ;
        RECT 1658.825 5.930 1659.155 5.945 ;
        RECT 1544.745 5.630 1548.970 5.930 ;
        RECT 1544.745 5.615 1545.075 5.630 ;
        RECT 1438.270 4.950 1453.290 5.250 ;
        RECT 1499.665 5.250 1499.995 5.265 ;
        RECT 1516.430 5.250 1516.810 5.260 ;
        RECT 1499.665 4.950 1516.810 5.250 ;
        RECT 658.325 4.935 658.655 4.950 ;
        RECT 677.390 4.940 677.770 4.950 ;
        RECT 1499.665 4.935 1499.995 4.950 ;
        RECT 1516.430 4.940 1516.810 4.950 ;
        RECT 1517.145 5.250 1517.475 5.265 ;
        RECT 1534.625 5.250 1534.955 5.265 ;
        RECT 1517.145 4.950 1534.955 5.250 ;
        RECT 1548.670 5.250 1548.970 5.630 ;
        RECT 1648.705 5.630 1659.155 5.930 ;
        RECT 1648.705 5.615 1649.035 5.630 ;
        RECT 1658.825 5.615 1659.155 5.630 ;
        RECT 1852.230 5.930 1852.610 5.940 ;
        RECT 1862.605 5.930 1862.935 5.945 ;
        RECT 1852.230 5.630 1862.935 5.930 ;
        RECT 1852.230 5.620 1852.610 5.630 ;
        RECT 1862.605 5.615 1862.935 5.630 ;
        RECT 1946.785 5.930 1947.115 5.945 ;
        RECT 2197.270 5.930 2197.570 6.310 ;
        RECT 2215.885 6.295 2216.215 6.310 ;
        RECT 2584.345 6.610 2584.675 6.625 ;
        RECT 2686.465 6.610 2686.795 6.625 ;
        RECT 2584.345 6.310 2686.795 6.610 ;
        RECT 2584.345 6.295 2584.675 6.310 ;
        RECT 2686.465 6.295 2686.795 6.310 ;
        RECT 1946.785 5.630 2197.570 5.930 ;
        RECT 2807.190 5.930 2807.570 5.940 ;
        RECT 2841.945 5.930 2842.275 5.945 ;
        RECT 2807.190 5.630 2842.275 5.930 ;
        RECT 1946.785 5.615 1947.115 5.630 ;
        RECT 2807.190 5.620 2807.570 5.630 ;
        RECT 2841.945 5.615 2842.275 5.630 ;
        RECT 1634.445 5.250 1634.775 5.265 ;
        RECT 1548.670 4.950 1634.775 5.250 ;
        RECT 1517.145 4.935 1517.475 4.950 ;
        RECT 1534.625 4.935 1534.955 4.950 ;
        RECT 1634.445 4.935 1634.775 4.950 ;
        RECT 1636.285 5.250 1636.615 5.265 ;
        RECT 2843.325 5.250 2843.655 5.265 ;
        RECT 1636.285 4.950 2843.655 5.250 ;
        RECT 1636.285 4.935 1636.615 4.950 ;
        RECT 2843.325 4.935 2843.655 4.950 ;
        RECT 110.465 4.570 110.795 4.585 ;
        RECT 139.445 4.570 139.775 4.585 ;
        RECT 110.465 4.270 139.775 4.570 ;
        RECT 110.465 4.255 110.795 4.270 ;
        RECT 139.445 4.255 139.775 4.270 ;
        RECT 679.230 4.570 679.610 4.580 ;
        RECT 1645.230 4.570 1645.610 4.580 ;
        RECT 1648.245 4.570 1648.575 4.585 ;
        RECT 679.230 4.270 689.690 4.570 ;
        RECT 679.230 4.260 679.610 4.270 ;
        RECT 3.285 3.890 3.615 3.905 ;
        RECT 51.125 3.890 51.455 3.905 ;
        RECT 3.285 3.590 51.455 3.890 ;
        RECT 3.285 3.575 3.615 3.590 ;
        RECT 51.125 3.575 51.455 3.590 ;
        RECT 514.550 3.890 514.930 3.900 ;
        RECT 518.945 3.890 519.275 3.905 ;
        RECT 514.550 3.590 519.275 3.890 ;
        RECT 514.550 3.580 514.930 3.590 ;
        RECT 518.945 3.575 519.275 3.590 ;
        RECT 582.885 3.890 583.215 3.905 ;
        RECT 613.705 3.890 614.035 3.905 ;
        RECT 582.885 3.590 614.035 3.890 ;
        RECT 582.885 3.575 583.215 3.590 ;
        RECT 613.705 3.575 614.035 3.590 ;
        RECT 646.110 3.890 646.490 3.900 ;
        RECT 648.205 3.890 648.535 3.905 ;
        RECT 646.110 3.590 648.535 3.890 ;
        RECT 689.390 3.890 689.690 4.270 ;
        RECT 1645.230 4.270 1648.575 4.570 ;
        RECT 1645.230 4.260 1645.610 4.270 ;
        RECT 1648.245 4.255 1648.575 4.270 ;
        RECT 1680.905 4.570 1681.235 4.585 ;
        RECT 1747.605 4.570 1747.935 4.585 ;
        RECT 1680.905 4.270 1747.935 4.570 ;
        RECT 1680.905 4.255 1681.235 4.270 ;
        RECT 1747.605 4.255 1747.935 4.270 ;
        RECT 696.965 3.890 697.295 3.905 ;
        RECT 689.390 3.590 697.295 3.890 ;
        RECT 646.110 3.580 646.490 3.590 ;
        RECT 648.205 3.575 648.535 3.590 ;
        RECT 696.965 3.575 697.295 3.590 ;
        RECT 697.885 3.890 698.215 3.905 ;
        RECT 711.225 3.890 711.555 3.905 ;
        RECT 697.885 3.590 711.555 3.890 ;
        RECT 697.885 3.575 698.215 3.590 ;
        RECT 711.225 3.575 711.555 3.590 ;
        RECT 712.145 3.890 712.475 3.905 ;
        RECT 720.885 3.890 721.215 3.905 ;
        RECT 712.145 3.590 721.215 3.890 ;
        RECT 712.145 3.575 712.475 3.590 ;
        RECT 720.885 3.575 721.215 3.590 ;
        RECT 880.965 3.890 881.295 3.905 ;
        RECT 920.985 3.890 921.315 3.905 ;
        RECT 880.965 3.590 921.315 3.890 ;
        RECT 880.965 3.575 881.295 3.590 ;
        RECT 920.985 3.575 921.315 3.590 ;
        RECT 993.205 3.890 993.535 3.905 ;
        RECT 1105.445 3.890 1105.775 3.905 ;
        RECT 1769.430 3.890 1769.810 3.900 ;
        RECT 993.205 3.590 1105.775 3.890 ;
        RECT 993.205 3.575 993.535 3.590 ;
        RECT 1105.445 3.575 1105.775 3.590 ;
        RECT 1749.230 3.590 1769.810 3.890 ;
        RECT 700.185 3.210 700.515 3.225 ;
        RECT 751.245 3.210 751.575 3.225 ;
        RECT 700.185 2.910 751.575 3.210 ;
        RECT 700.185 2.895 700.515 2.910 ;
        RECT 751.245 2.895 751.575 2.910 ;
        RECT 818.150 3.210 818.530 3.220 ;
        RECT 848.305 3.210 848.635 3.225 ;
        RECT 818.150 2.910 848.635 3.210 ;
        RECT 818.150 2.900 818.530 2.910 ;
        RECT 848.305 2.895 848.635 2.910 ;
        RECT 889.705 3.210 890.035 3.225 ;
        RECT 986.765 3.210 987.095 3.225 ;
        RECT 889.705 2.910 987.095 3.210 ;
        RECT 889.705 2.895 890.035 2.910 ;
        RECT 986.765 2.895 987.095 2.910 ;
        RECT 992.285 3.210 992.615 3.225 ;
        RECT 1020.550 3.210 1020.930 3.220 ;
        RECT 992.285 2.910 1020.930 3.210 ;
        RECT 992.285 2.895 992.615 2.910 ;
        RECT 1020.550 2.900 1020.930 2.910 ;
        RECT 1021.265 3.210 1021.595 3.225 ;
        RECT 1022.645 3.210 1022.975 3.225 ;
        RECT 1021.265 2.910 1022.975 3.210 ;
        RECT 1021.265 2.895 1021.595 2.910 ;
        RECT 1022.645 2.895 1022.975 2.910 ;
        RECT 1023.310 3.210 1023.690 3.220 ;
        RECT 1025.405 3.210 1025.735 3.225 ;
        RECT 1023.310 2.910 1025.735 3.210 ;
        RECT 1023.310 2.900 1023.690 2.910 ;
        RECT 1025.405 2.895 1025.735 2.910 ;
        RECT 1057.145 3.210 1057.475 3.225 ;
        RECT 1075.085 3.210 1075.415 3.225 ;
        RECT 1057.145 2.910 1075.415 3.210 ;
        RECT 1057.145 2.895 1057.475 2.910 ;
        RECT 1075.085 2.895 1075.415 2.910 ;
        RECT 1165.705 3.210 1166.035 3.225 ;
        RECT 1237.925 3.210 1238.255 3.225 ;
        RECT 1165.705 2.910 1238.255 3.210 ;
        RECT 1165.705 2.895 1166.035 2.910 ;
        RECT 1237.925 2.895 1238.255 2.910 ;
        RECT 1242.065 3.210 1242.395 3.225 ;
        RECT 1307.845 3.210 1308.175 3.225 ;
        RECT 1242.065 2.910 1308.175 3.210 ;
        RECT 1242.065 2.895 1242.395 2.910 ;
        RECT 1307.845 2.895 1308.175 2.910 ;
        RECT 1334.985 3.210 1335.315 3.225 ;
        RECT 1680.905 3.210 1681.235 3.225 ;
        RECT 1334.985 2.910 1681.235 3.210 ;
        RECT 1334.985 2.895 1335.315 2.910 ;
        RECT 1680.905 2.895 1681.235 2.910 ;
        RECT 1681.825 3.210 1682.155 3.225 ;
        RECT 1693.070 3.210 1693.450 3.220 ;
        RECT 1681.825 2.910 1693.450 3.210 ;
        RECT 1681.825 2.895 1682.155 2.910 ;
        RECT 1693.070 2.900 1693.450 2.910 ;
        RECT 1715.405 3.210 1715.735 3.225 ;
        RECT 1749.230 3.210 1749.530 3.590 ;
        RECT 1769.430 3.580 1769.810 3.590 ;
        RECT 2031.885 3.890 2032.215 3.905 ;
        RECT 2174.945 3.890 2175.275 3.905 ;
        RECT 2031.885 3.590 2175.275 3.890 ;
        RECT 2031.885 3.575 2032.215 3.590 ;
        RECT 2174.945 3.575 2175.275 3.590 ;
        RECT 2684.625 3.890 2684.955 3.905 ;
        RECT 2697.710 3.890 2698.090 3.900 ;
        RECT 2684.625 3.590 2698.090 3.890 ;
        RECT 2684.625 3.575 2684.955 3.590 ;
        RECT 2697.710 3.580 2698.090 3.590 ;
        RECT 2845.625 3.890 2845.955 3.905 ;
        RECT 2845.625 3.575 2846.170 3.890 ;
        RECT 1715.405 2.910 1749.530 3.210 ;
        RECT 1750.110 3.210 1750.490 3.220 ;
        RECT 1782.565 3.210 1782.895 3.225 ;
        RECT 1750.110 2.910 1782.895 3.210 ;
        RECT 1715.405 2.895 1715.735 2.910 ;
        RECT 1750.110 2.900 1750.490 2.910 ;
        RECT 1782.565 2.895 1782.895 2.910 ;
        RECT 1784.865 3.210 1785.195 3.225 ;
        RECT 1825.345 3.210 1825.675 3.225 ;
        RECT 1784.865 2.910 1825.675 3.210 ;
        RECT 1784.865 2.895 1785.195 2.910 ;
        RECT 1825.345 2.895 1825.675 2.910 ;
        RECT 1930.225 3.210 1930.555 3.225 ;
        RECT 1952.510 3.210 1952.890 3.220 ;
        RECT 1930.225 2.910 1952.890 3.210 ;
        RECT 1930.225 2.895 1930.555 2.910 ;
        RECT 1952.510 2.900 1952.890 2.910 ;
        RECT 1967.025 3.210 1967.355 3.225 ;
        RECT 2056.265 3.210 2056.595 3.225 ;
        RECT 1967.025 2.910 2056.595 3.210 ;
        RECT 1967.025 2.895 1967.355 2.910 ;
        RECT 2056.265 2.895 2056.595 2.910 ;
        RECT 2214.045 3.210 2214.375 3.225 ;
        RECT 2383.785 3.210 2384.115 3.225 ;
        RECT 2612.865 3.210 2613.195 3.225 ;
        RECT 2683.705 3.210 2684.035 3.225 ;
        RECT 2798.910 3.210 2799.290 3.220 ;
        RECT 2214.045 2.910 2384.115 3.210 ;
        RECT 2214.045 2.895 2214.375 2.910 ;
        RECT 2383.785 2.895 2384.115 2.910 ;
        RECT 2563.430 2.910 2612.490 3.210 ;
        RECT 380.945 2.530 381.275 2.545 ;
        RECT 392.445 2.530 392.775 2.545 ;
        RECT 990.905 2.540 991.235 2.545 ;
        RECT 380.945 2.230 392.775 2.530 ;
        RECT 380.945 2.215 381.275 2.230 ;
        RECT 392.445 2.215 392.775 2.230 ;
        RECT 396.790 2.530 397.170 2.540 ;
        RECT 401.390 2.530 401.770 2.540 ;
        RECT 990.905 2.530 991.490 2.540 ;
        RECT 396.790 2.230 401.770 2.530 ;
        RECT 990.680 2.230 991.490 2.530 ;
        RECT 396.790 2.220 397.170 2.230 ;
        RECT 401.390 2.220 401.770 2.230 ;
        RECT 990.905 2.220 991.490 2.230 ;
        RECT 2367.430 2.530 2367.810 2.540 ;
        RECT 2549.385 2.530 2549.715 2.545 ;
        RECT 2367.430 2.230 2549.715 2.530 ;
        RECT 2367.430 2.220 2367.810 2.230 ;
        RECT 990.905 2.215 991.235 2.220 ;
        RECT 2549.385 2.215 2549.715 2.230 ;
        RECT 789.630 1.850 790.010 1.860 ;
        RECT 806.190 1.850 806.570 1.860 ;
        RECT 789.630 1.550 806.570 1.850 ;
        RECT 789.630 1.540 790.010 1.550 ;
        RECT 806.190 1.540 806.570 1.550 ;
        RECT 1825.345 1.850 1825.675 1.865 ;
        RECT 1930.225 1.850 1930.555 1.865 ;
        RECT 1825.345 1.550 1930.555 1.850 ;
        RECT 1825.345 1.535 1825.675 1.550 ;
        RECT 1930.225 1.535 1930.555 1.550 ;
        RECT 1952.510 1.850 1952.890 1.860 ;
        RECT 2031.885 1.850 2032.215 1.865 ;
        RECT 1952.510 1.550 2032.215 1.850 ;
        RECT 1952.510 1.540 1952.890 1.550 ;
        RECT 2031.885 1.535 2032.215 1.550 ;
        RECT 2128.485 1.850 2128.815 1.865 ;
        RECT 2134.670 1.850 2135.050 1.860 ;
        RECT 2128.485 1.550 2135.050 1.850 ;
        RECT 2128.485 1.535 2128.815 1.550 ;
        RECT 2134.670 1.540 2135.050 1.550 ;
        RECT 2215.885 1.850 2216.215 1.865 ;
        RECT 2365.590 1.850 2365.970 1.860 ;
        RECT 2563.430 1.850 2563.730 2.910 ;
        RECT 2612.190 2.530 2612.490 2.910 ;
        RECT 2612.865 2.910 2684.035 3.210 ;
        RECT 2612.865 2.895 2613.195 2.910 ;
        RECT 2683.705 2.895 2684.035 2.910 ;
        RECT 2727.190 2.910 2799.290 3.210 ;
        RECT 2697.710 2.530 2698.090 2.540 ;
        RECT 2727.190 2.530 2727.490 2.910 ;
        RECT 2798.910 2.900 2799.290 2.910 ;
        RECT 2612.190 2.230 2643.770 2.530 ;
        RECT 2215.885 1.550 2365.970 1.850 ;
        RECT 2215.885 1.535 2216.215 1.550 ;
        RECT 2365.590 1.540 2365.970 1.550 ;
        RECT 2521.110 1.550 2563.730 1.850 ;
        RECT 421.885 1.170 422.215 1.185 ;
        RECT 427.150 1.170 427.530 1.180 ;
        RECT 421.885 0.870 427.530 1.170 ;
        RECT 421.885 0.855 422.215 0.870 ;
        RECT 427.150 0.860 427.530 0.870 ;
        RECT 2366.765 1.170 2367.095 1.185 ;
        RECT 2368.605 1.170 2368.935 1.185 ;
        RECT 2366.765 0.870 2368.935 1.170 ;
        RECT 2366.765 0.855 2367.095 0.870 ;
        RECT 2368.605 0.855 2368.935 0.870 ;
        RECT 2430.705 1.170 2431.035 1.185 ;
        RECT 2521.110 1.170 2521.410 1.550 ;
        RECT 2430.705 0.870 2521.410 1.170 ;
        RECT 2643.470 1.170 2643.770 2.230 ;
        RECT 2697.710 2.230 2727.490 2.530 ;
        RECT 2728.325 2.530 2728.655 2.545 ;
        RECT 2845.870 2.530 2846.170 3.575 ;
        RECT 2728.325 2.230 2846.170 2.530 ;
        RECT 2697.710 2.220 2698.090 2.230 ;
        RECT 2728.325 2.215 2728.655 2.230 ;
        RECT 2728.325 1.170 2728.655 1.185 ;
        RECT 2643.470 0.870 2728.655 1.170 ;
        RECT 2430.705 0.855 2431.035 0.870 ;
        RECT 2728.325 0.855 2728.655 0.870 ;
        RECT 9.470 0.490 9.850 0.500 ;
        RECT 49.285 0.490 49.615 0.505 ;
        RECT 9.470 0.190 49.615 0.490 ;
        RECT 9.470 0.180 9.850 0.190 ;
        RECT 49.285 0.175 49.615 0.190 ;
        RECT 372.665 0.490 372.995 0.505 ;
        RECT 393.110 0.490 393.490 0.500 ;
        RECT 372.665 0.190 393.490 0.490 ;
        RECT 372.665 0.175 372.995 0.190 ;
        RECT 393.110 0.180 393.490 0.190 ;
        RECT 408.085 0.490 408.415 0.505 ;
        RECT 414.525 0.490 414.855 0.505 ;
        RECT 408.085 0.190 414.855 0.490 ;
        RECT 408.085 0.175 408.415 0.190 ;
        RECT 414.525 0.175 414.855 0.190 ;
        RECT 415.190 0.490 415.570 0.500 ;
        RECT 420.965 0.490 421.295 0.505 ;
        RECT 415.190 0.190 421.295 0.490 ;
        RECT 415.190 0.180 415.570 0.190 ;
        RECT 420.965 0.175 421.295 0.190 ;
      LAYER via3 ;
        RECT 2798.940 3403.580 2799.260 3403.900 ;
        RECT 2852.300 1422.740 2852.620 1423.060 ;
        RECT 2851.380 967.820 2851.700 968.140 ;
        RECT 2852.300 967.140 2852.620 967.460 ;
        RECT 2853.220 967.140 2853.540 967.460 ;
        RECT 2851.380 496.580 2851.700 496.900 ;
        RECT 2852.300 450.340 2852.620 450.660 ;
        RECT 7.660 89.940 7.980 90.260 ;
        RECT 4.900 64.100 5.220 64.420 ;
        RECT 2851.380 61.380 2851.700 61.700 ;
        RECT 7.660 43.700 7.980 44.020 ;
        RECT 2852.300 21.940 2852.620 22.260 ;
        RECT 417.980 8.340 418.300 8.660 ;
        RECT 429.020 8.340 429.340 8.660 ;
        RECT 440.060 8.340 440.380 8.660 ;
        RECT 557.820 8.340 558.140 8.660 ;
        RECT 629.580 8.340 629.900 8.660 ;
        RECT 639.700 8.340 640.020 8.660 ;
        RECT 678.340 8.340 678.660 8.660 ;
        RECT 261.580 7.660 261.900 7.980 ;
        RECT 377.500 7.660 377.820 7.980 ;
        RECT 509.060 7.660 509.380 7.980 ;
        RECT 516.420 7.660 516.740 7.980 ;
        RECT 974.580 8.340 974.900 8.660 ;
        RECT 1084.060 8.340 1084.380 8.660 ;
        RECT 1101.540 8.340 1101.860 8.660 ;
        RECT 1171.460 8.340 1171.780 8.660 ;
        RECT 1189.860 8.340 1190.180 8.660 ;
        RECT 952.500 7.660 952.820 7.980 ;
        RECT 514.580 6.980 514.900 7.300 ;
        RECT 675.580 6.980 675.900 7.300 ;
        RECT 693.980 6.980 694.300 7.300 ;
        RECT 808.060 6.980 808.380 7.300 ;
        RECT 820.020 6.980 820.340 7.300 ;
        RECT 955.260 6.980 955.580 7.300 ;
        RECT 992.060 7.660 992.380 7.980 ;
        RECT 1002.180 6.980 1002.500 7.300 ;
        RECT 1193.540 7.660 1193.860 7.980 ;
        RECT 1428.140 8.340 1428.460 8.660 ;
        RECT 2566.180 8.340 2566.500 8.660 ;
        RECT 2845.860 8.340 2846.180 8.660 ;
        RECT 684.780 6.300 685.100 6.620 ;
        RECT 881.660 6.300 881.980 6.620 ;
        RECT 1054.620 6.980 1054.940 7.300 ;
        RECT 1268.980 7.660 1269.300 7.980 ;
        RECT 1267.140 6.980 1267.460 7.300 ;
        RECT 1303.020 6.980 1303.340 7.300 ;
        RECT 1304.860 6.980 1305.180 7.300 ;
        RECT 2794.340 7.660 2794.660 7.980 ;
        RECT 2795.260 7.660 2795.580 7.980 ;
        RECT 1402.380 6.980 1402.700 7.300 ;
        RECT 1073.940 6.300 1074.260 6.620 ;
        RECT 1137.420 6.300 1137.740 6.620 ;
        RECT 1138.340 6.300 1138.660 6.620 ;
        RECT 1145.700 6.300 1146.020 6.620 ;
        RECT 1314.060 6.300 1314.380 6.620 ;
        RECT 1324.180 6.300 1324.500 6.620 ;
        RECT 462.140 5.620 462.460 5.940 ;
        RECT 506.300 5.620 506.620 5.940 ;
        RECT 556.900 5.620 557.220 5.940 ;
        RECT 634.180 5.620 634.500 5.940 ;
        RECT 641.540 5.620 641.860 5.940 ;
        RECT 737.220 5.620 737.540 5.940 ;
        RECT 753.780 5.620 754.100 5.940 ;
        RECT 1133.740 5.620 1134.060 5.940 ;
        RECT 1344.420 5.620 1344.740 5.940 ;
        RECT 1397.780 5.620 1398.100 5.940 ;
        RECT 677.420 4.940 677.740 5.260 ;
        RECT 1474.140 6.300 1474.460 6.620 ;
        RECT 1589.140 6.300 1589.460 6.620 ;
        RECT 1624.100 6.300 1624.420 6.620 ;
        RECT 1448.380 5.620 1448.700 5.940 ;
        RECT 1450.220 5.620 1450.540 5.940 ;
        RECT 1516.460 4.940 1516.780 5.260 ;
        RECT 1852.260 5.620 1852.580 5.940 ;
        RECT 2807.220 5.620 2807.540 5.940 ;
        RECT 679.260 4.260 679.580 4.580 ;
        RECT 514.580 3.580 514.900 3.900 ;
        RECT 646.140 3.580 646.460 3.900 ;
        RECT 1645.260 4.260 1645.580 4.580 ;
        RECT 818.180 2.900 818.500 3.220 ;
        RECT 1020.580 2.900 1020.900 3.220 ;
        RECT 1023.340 2.900 1023.660 3.220 ;
        RECT 1693.100 2.900 1693.420 3.220 ;
        RECT 1769.460 3.580 1769.780 3.900 ;
        RECT 2697.740 3.580 2698.060 3.900 ;
        RECT 1750.140 2.900 1750.460 3.220 ;
        RECT 1952.540 2.900 1952.860 3.220 ;
        RECT 396.820 2.220 397.140 2.540 ;
        RECT 401.420 2.220 401.740 2.540 ;
        RECT 991.140 2.220 991.460 2.540 ;
        RECT 2367.460 2.220 2367.780 2.540 ;
        RECT 789.660 1.540 789.980 1.860 ;
        RECT 806.220 1.540 806.540 1.860 ;
        RECT 1952.540 1.540 1952.860 1.860 ;
        RECT 2134.700 1.540 2135.020 1.860 ;
        RECT 2365.620 1.540 2365.940 1.860 ;
        RECT 427.180 0.860 427.500 1.180 ;
        RECT 2697.740 2.220 2698.060 2.540 ;
        RECT 2798.940 2.900 2799.260 3.220 ;
        RECT 9.500 0.180 9.820 0.500 ;
        RECT 393.140 0.180 393.460 0.500 ;
        RECT 415.220 0.180 415.540 0.500 ;
      LAYER met4 ;
        RECT -37.580 -32.220 -34.580 3551.900 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 2798.935 3403.575 2799.265 3403.905 ;
        RECT 2798.950 3381.890 2799.250 3403.575 ;
        RECT 2793.910 3380.710 2795.090 3381.890 ;
        RECT 2798.510 3380.710 2799.690 3381.890 ;
        RECT 2794.350 3225.050 2794.650 3380.710 ;
        RECT 2793.430 3224.750 2794.650 3225.050 ;
        RECT 2793.430 3201.250 2793.730 3224.750 ;
        RECT 2793.430 3200.950 2794.650 3201.250 ;
        RECT 2794.350 3123.050 2794.650 3200.950 ;
        RECT 2794.350 3122.750 2795.570 3123.050 ;
        RECT 2795.270 3116.250 2795.570 3122.750 ;
        RECT 2794.350 3115.950 2795.570 3116.250 ;
        RECT 2794.350 1545.450 2794.650 3115.950 ;
        RECT 2794.350 1545.150 2795.570 1545.450 ;
        RECT 2795.270 1477.450 2795.570 1545.150 ;
        RECT 2794.350 1477.150 2795.570 1477.450 ;
        RECT 9.070 130.310 10.250 131.490 ;
        RECT 7.655 90.250 7.985 90.265 ;
        RECT 9.510 90.250 9.810 130.310 ;
        RECT 7.655 89.950 9.810 90.250 ;
        RECT 7.655 89.935 7.985 89.950 ;
        RECT 2794.350 80.490 2794.650 1477.150 ;
        RECT 2852.295 1423.050 2852.625 1423.065 ;
        RECT 2849.550 1422.750 2852.625 1423.050 ;
        RECT 2849.550 1419.650 2849.850 1422.750 ;
        RECT 2852.295 1422.735 2852.625 1422.750 ;
        RECT 2846.790 1419.350 2849.850 1419.650 ;
        RECT 2846.790 1368.650 2847.090 1419.350 ;
        RECT 2846.790 1368.350 2848.930 1368.650 ;
        RECT 2848.630 1338.050 2848.930 1368.350 ;
        RECT 2848.630 1337.750 2851.690 1338.050 ;
        RECT 2846.085 1300.650 2846.415 1300.665 ;
        RECT 2844.030 1300.350 2846.415 1300.650 ;
        RECT 2844.030 1263.250 2844.330 1300.350 ;
        RECT 2846.085 1300.335 2846.415 1300.350 ;
        RECT 2851.390 1290.450 2851.690 1337.750 ;
        RECT 2849.550 1290.150 2851.690 1290.450 ;
        RECT 2849.550 1283.650 2849.850 1290.150 ;
        RECT 2843.110 1262.950 2844.330 1263.250 ;
        RECT 2846.790 1283.350 2849.850 1283.650 ;
        RECT 2843.110 1242.850 2843.410 1262.950 ;
        RECT 2841.960 1242.550 2843.410 1242.850 ;
        RECT 2841.960 1242.185 2842.260 1242.550 ;
        RECT 2841.945 1241.855 2842.275 1242.185 ;
        RECT 2844.245 1111.295 2844.575 1111.625 ;
        RECT 2844.260 1110.250 2844.560 1111.295 ;
        RECT 2841.270 1109.950 2844.560 1110.250 ;
        RECT 2841.270 1049.050 2841.570 1109.950 ;
        RECT 2841.270 1048.750 2842.490 1049.050 ;
        RECT 2842.190 974.250 2842.490 1048.750 ;
        RECT 2846.790 974.250 2847.090 1283.350 ;
        RECT 2842.190 973.950 2844.330 974.250 ;
        RECT 2846.790 973.950 2853.530 974.250 ;
        RECT 2842.865 968.130 2843.195 968.145 ;
        RECT 2842.865 967.815 2843.410 968.130 ;
        RECT 2841.485 967.450 2841.815 967.465 ;
        RECT 2841.270 967.135 2841.815 967.450 ;
        RECT 2841.270 872.250 2841.570 967.135 ;
        RECT 2843.110 964.050 2843.410 967.815 ;
        RECT 2844.030 967.450 2844.330 973.950 ;
        RECT 2851.375 968.130 2851.705 968.145 ;
        RECT 2845.870 967.830 2851.705 968.130 ;
        RECT 2845.870 967.450 2846.170 967.830 ;
        RECT 2851.375 967.815 2851.705 967.830 ;
        RECT 2853.230 967.465 2853.530 973.950 ;
        RECT 2852.295 967.450 2852.625 967.465 ;
        RECT 2844.030 967.150 2846.170 967.450 ;
        RECT 2846.790 967.150 2852.625 967.450 ;
        RECT 2843.110 963.750 2844.330 964.050 ;
        RECT 2844.030 892.650 2844.330 963.750 ;
        RECT 2845.855 892.650 2846.185 892.665 ;
        RECT 2844.030 892.350 2846.185 892.650 ;
        RECT 2845.855 892.335 2846.185 892.350 ;
        RECT 2842.405 872.615 2842.735 872.945 ;
        RECT 2842.420 872.250 2842.720 872.615 ;
        RECT 2841.270 871.950 2842.720 872.250 ;
        RECT 2846.790 831.450 2847.090 967.150 ;
        RECT 2852.295 967.135 2852.625 967.150 ;
        RECT 2853.215 967.135 2853.545 967.465 ;
        RECT 2846.790 831.150 2848.930 831.450 ;
        RECT 2848.630 624.050 2848.930 831.150 ;
        RECT 2846.790 623.750 2848.930 624.050 ;
        RECT 2846.790 501.650 2847.090 623.750 ;
        RECT 2846.790 501.350 2851.690 501.650 ;
        RECT 2851.390 496.905 2851.690 501.350 ;
        RECT 2851.375 496.575 2851.705 496.905 ;
        RECT 2852.295 450.650 2852.625 450.665 ;
        RECT 2847.710 450.350 2852.625 450.650 ;
        RECT 2847.710 253.450 2848.010 450.350 ;
        RECT 2852.295 450.335 2852.625 450.350 ;
        RECT 2846.790 253.150 2848.010 253.450 ;
        RECT 2846.790 216.050 2847.090 253.150 ;
        RECT 2846.790 215.750 2852.610 216.050 ;
        RECT 2852.310 182.050 2852.610 215.750 ;
        RECT 2845.870 181.750 2852.610 182.050 ;
        RECT 2806.790 130.310 2807.970 131.490 ;
        RECT 2798.510 92.910 2799.690 94.090 ;
        RECT 2793.910 79.310 2795.090 80.490 ;
        RECT 4.470 75.910 5.650 77.090 ;
        RECT 4.910 64.425 5.210 75.910 ;
        RECT 9.070 69.110 10.250 70.290 ;
        RECT 23.790 69.110 24.970 70.290 ;
        RECT 4.895 64.095 5.225 64.425 ;
        RECT 7.230 52.110 8.410 53.290 ;
        RECT 7.670 44.025 7.970 52.110 ;
        RECT 7.655 43.695 7.985 44.025 ;
        RECT 9.510 0.505 9.810 69.110 ;
        RECT 24.230 60.090 24.530 69.110 ;
        RECT 100.150 65.710 101.330 66.890 ;
        RECT 23.790 58.910 24.970 60.090 ;
        RECT 2792.990 58.910 2794.170 60.090 ;
        RECT 2793.430 49.450 2793.730 58.910 ;
        RECT 2798.950 56.690 2799.250 92.910 ;
        RECT 2794.830 55.510 2796.010 56.690 ;
        RECT 2798.510 55.510 2799.690 56.690 ;
        RECT 2793.430 49.150 2794.650 49.450 ;
        RECT 1128.710 24.910 1129.890 26.090 ;
        RECT 261.150 14.710 262.330 15.890 ;
        RECT 374.310 14.710 375.490 15.890 ;
        RECT 513.230 14.710 514.410 15.890 ;
        RECT 626.390 15.450 627.570 15.890 ;
        RECT 626.390 15.150 628.050 15.450 ;
        RECT 626.390 14.710 627.570 15.150 ;
        RECT 261.590 7.985 261.890 14.710 ;
        RECT 261.575 7.655 261.905 7.985 ;
        RECT 374.750 7.970 375.050 14.710 ;
        RECT 460.310 11.750 466.130 12.050 ;
        RECT 460.310 9.330 460.610 11.750 ;
        RECT 440.070 9.030 442.210 9.330 ;
        RECT 440.070 8.665 440.370 9.030 ;
        RECT 417.975 8.650 418.305 8.665 ;
        RECT 429.015 8.650 429.345 8.665 ;
        RECT 417.975 8.350 429.345 8.650 ;
        RECT 417.975 8.335 418.305 8.350 ;
        RECT 429.015 8.335 429.345 8.350 ;
        RECT 440.055 8.335 440.385 8.665 ;
        RECT 441.910 8.650 442.210 9.030 ;
        RECT 459.620 9.030 460.610 9.330 ;
        RECT 465.830 9.330 466.130 11.750 ;
        RECT 465.830 9.030 475.330 9.330 ;
        RECT 459.620 8.650 459.920 9.030 ;
        RECT 441.910 8.350 459.920 8.650 ;
        RECT 377.495 7.970 377.825 7.985 ;
        RECT 374.750 7.670 377.825 7.970 ;
        RECT 377.495 7.655 377.825 7.670 ;
        RECT 475.030 7.290 475.330 9.030 ;
        RECT 509.055 7.970 509.385 7.985 ;
        RECT 479.630 7.670 509.385 7.970 ;
        RECT 479.630 7.290 479.930 7.670 ;
        RECT 509.055 7.655 509.385 7.670 ;
        RECT 475.030 6.990 479.930 7.290 ;
        RECT 513.670 7.290 513.970 14.710 ;
        RECT 518.270 11.750 580.210 12.050 ;
        RECT 516.415 7.970 516.745 7.985 ;
        RECT 518.270 7.970 518.570 11.750 ;
        RECT 579.910 9.330 580.210 11.750 ;
        RECT 627.750 9.330 628.050 15.150 ;
        RECT 678.830 14.710 680.010 15.890 ;
        RECT 768.070 14.710 769.250 15.890 ;
        RECT 776.350 14.710 777.530 15.890 ;
        RECT 1138.830 14.710 1140.010 15.890 ;
        RECT 1300.750 14.710 1301.930 15.890 ;
        RECT 2134.270 14.710 2135.450 15.890 ;
        RECT 2565.750 14.710 2566.930 15.890 ;
        RECT 639.710 11.750 671.290 12.050 ;
        RECT 579.910 9.030 623.450 9.330 ;
        RECT 627.750 9.030 630.810 9.330 ;
        RECT 557.815 8.650 558.145 8.665 ;
        RECT 516.415 7.670 518.570 7.970 ;
        RECT 556.910 8.350 558.145 8.650 ;
        RECT 623.150 8.650 623.450 9.030 ;
        RECT 629.575 8.650 629.905 8.665 ;
        RECT 623.150 8.350 629.905 8.650 ;
        RECT 516.415 7.655 516.745 7.670 ;
        RECT 514.575 7.290 514.905 7.305 ;
        RECT 513.670 6.990 514.905 7.290 ;
        RECT 514.575 6.975 514.905 6.990 ;
        RECT 401.430 6.310 414.610 6.610 ;
        RECT 401.430 2.545 401.730 6.310 ;
        RECT 396.815 2.215 397.145 2.545 ;
        RECT 401.415 2.215 401.745 2.545 ;
        RECT 396.830 1.850 397.130 2.215 ;
        RECT 395.910 1.550 397.130 1.850 ;
        RECT 9.495 0.175 9.825 0.505 ;
        RECT 393.135 0.490 393.465 0.505 ;
        RECT 395.910 0.490 396.210 1.550 ;
        RECT 393.135 0.190 396.210 0.490 ;
        RECT 414.310 0.490 414.610 6.310 ;
        RECT 556.910 5.945 557.210 8.350 ;
        RECT 557.815 8.335 558.145 8.350 ;
        RECT 629.575 8.335 629.905 8.350 ;
        RECT 462.135 5.615 462.465 5.945 ;
        RECT 506.295 5.615 506.625 5.945 ;
        RECT 556.895 5.615 557.225 5.945 ;
        RECT 630.510 5.930 630.810 9.030 ;
        RECT 639.710 8.665 640.010 11.750 ;
        RECT 670.990 9.330 671.290 11.750 ;
        RECT 670.990 9.030 677.730 9.330 ;
        RECT 639.695 8.335 640.025 8.665 ;
        RECT 677.430 8.650 677.730 9.030 ;
        RECT 678.335 8.650 678.665 8.665 ;
        RECT 677.430 8.350 678.665 8.650 ;
        RECT 678.335 8.335 678.665 8.350 ;
        RECT 679.270 7.970 679.570 14.710 ;
        RECT 768.510 9.330 768.810 14.710 ;
        RECT 770.140 9.330 771.320 9.770 ;
        RECT 675.590 7.670 679.570 7.970 ;
        RECT 735.390 9.030 763.290 9.330 ;
        RECT 768.510 9.030 771.320 9.330 ;
        RECT 675.590 7.305 675.890 7.670 ;
        RECT 675.575 6.975 675.905 7.305 ;
        RECT 693.975 6.975 694.305 7.305 ;
        RECT 684.775 6.610 685.105 6.625 ;
        RECT 693.990 6.610 694.290 6.975 ;
        RECT 684.775 6.310 694.290 6.610 ;
        RECT 735.390 6.610 735.690 9.030 ;
        RECT 762.990 7.970 763.290 9.030 ;
        RECT 770.140 8.590 771.320 9.030 ;
        RECT 776.790 8.650 777.090 14.710 ;
        RECT 1128.710 13.210 1129.890 14.390 ;
        RECT 974.150 11.310 975.330 12.490 ;
        RECT 1056.470 11.750 1077.010 12.050 ;
        RECT 774.030 8.350 777.090 8.650 ;
        RECT 794.750 8.650 795.930 9.770 ;
        RECT 974.590 8.665 974.890 11.310 ;
        RECT 794.750 8.590 800.090 8.650 ;
        RECT 795.190 8.350 800.090 8.590 ;
        RECT 774.030 7.970 774.330 8.350 ;
        RECT 762.990 7.670 774.330 7.970 ;
        RECT 799.790 7.290 800.090 8.350 ;
        RECT 859.590 8.350 866.330 8.650 ;
        RECT 799.790 6.990 801.010 7.290 ;
        RECT 808.055 7.050 808.385 7.305 ;
        RECT 820.015 7.290 820.345 7.305 ;
        RECT 735.390 6.310 737.530 6.610 ;
        RECT 684.775 6.295 685.105 6.310 ;
        RECT 737.230 5.945 737.530 6.310 ;
        RECT 753.790 6.310 759.610 6.610 ;
        RECT 753.790 5.945 754.090 6.310 ;
        RECT 634.175 5.930 634.505 5.945 ;
        RECT 630.510 5.630 634.505 5.930 ;
        RECT 634.175 5.615 634.505 5.630 ;
        RECT 641.535 5.615 641.865 5.945 ;
        RECT 737.215 5.615 737.545 5.945 ;
        RECT 753.775 5.615 754.105 5.945 ;
        RECT 462.150 3.210 462.450 5.615 ;
        RECT 506.310 5.250 506.610 5.615 ;
        RECT 506.310 4.950 514.890 5.250 ;
        RECT 514.590 3.905 514.890 4.950 ;
        RECT 514.575 3.575 514.905 3.905 ;
        RECT 641.550 3.890 641.850 5.615 ;
        RECT 677.415 4.935 677.745 5.265 ;
        RECT 677.430 4.570 677.730 4.935 ;
        RECT 679.255 4.570 679.585 4.585 ;
        RECT 677.430 4.270 679.585 4.570 ;
        RECT 679.255 4.255 679.585 4.270 ;
        RECT 646.135 3.890 646.465 3.905 ;
        RECT 641.550 3.590 646.465 3.890 ;
        RECT 646.135 3.575 646.465 3.590 ;
        RECT 437.310 2.910 462.450 3.210 ;
        RECT 427.175 0.855 427.505 1.185 ;
        RECT 415.215 0.490 415.545 0.505 ;
        RECT 414.310 0.190 415.545 0.490 ;
        RECT 427.190 0.490 427.490 0.855 ;
        RECT 437.310 0.490 437.610 2.910 ;
        RECT 759.310 1.850 759.610 6.310 ;
        RECT 800.710 5.690 801.010 6.990 ;
        RECT 807.630 5.870 808.810 7.050 ;
        RECT 820.015 6.990 832.290 7.290 ;
        RECT 820.015 6.975 820.345 6.990 ;
        RECT 800.270 4.510 801.450 5.690 ;
        RECT 831.990 5.250 832.290 6.990 ;
        RECT 859.590 6.610 859.890 8.350 ;
        RECT 866.030 7.970 866.330 8.350 ;
        RECT 974.575 8.335 974.905 8.665 ;
        RECT 1056.470 8.650 1056.770 11.750 ;
        RECT 1076.710 9.330 1077.010 11.750 ;
        RECT 1119.510 9.330 1120.690 9.770 ;
        RECT 1076.710 9.030 1080.690 9.330 ;
        RECT 1054.630 8.350 1056.770 8.650 ;
        RECT 1080.390 8.650 1080.690 9.030 ;
        RECT 1101.550 9.030 1120.690 9.330 ;
        RECT 1101.550 8.665 1101.850 9.030 ;
        RECT 1084.055 8.650 1084.385 8.665 ;
        RECT 1080.390 8.350 1084.385 8.650 ;
        RECT 866.030 7.670 878.290 7.970 ;
        RECT 851.310 6.310 859.890 6.610 ;
        RECT 851.310 5.250 851.610 6.310 ;
        RECT 831.990 4.950 851.610 5.250 ;
        RECT 877.990 5.250 878.290 7.670 ;
        RECT 952.495 7.655 952.825 7.985 ;
        RECT 992.055 7.970 992.385 7.985 ;
        RECT 992.055 7.670 1002.490 7.970 ;
        RECT 992.055 7.655 992.385 7.670 ;
        RECT 952.510 7.290 952.810 7.655 ;
        RECT 1002.190 7.305 1002.490 7.670 ;
        RECT 1054.630 7.305 1054.930 8.350 ;
        RECT 1084.055 8.335 1084.385 8.350 ;
        RECT 1101.535 8.335 1101.865 8.665 ;
        RECT 1119.510 8.590 1120.690 9.030 ;
        RECT 955.255 7.290 955.585 7.305 ;
        RECT 952.510 6.990 955.585 7.290 ;
        RECT 955.255 6.975 955.585 6.990 ;
        RECT 1002.175 6.975 1002.505 7.305 ;
        RECT 1054.615 6.975 1054.945 7.305 ;
        RECT 881.655 6.295 881.985 6.625 ;
        RECT 1073.935 6.610 1074.265 6.625 ;
        RECT 1069.350 6.310 1074.265 6.610 ;
        RECT 881.670 5.250 881.970 6.295 ;
        RECT 877.990 4.950 881.970 5.250 ;
        RECT 1053.710 5.630 1058.610 5.930 ;
        RECT 818.175 3.210 818.505 3.225 ;
        RECT 809.910 2.910 818.505 3.210 ;
        RECT 789.655 1.850 789.985 1.865 ;
        RECT 759.310 1.550 789.985 1.850 ;
        RECT 789.655 1.535 789.985 1.550 ;
        RECT 806.215 1.850 806.545 1.865 ;
        RECT 809.910 1.850 810.210 2.910 ;
        RECT 818.175 2.895 818.505 2.910 ;
        RECT 1020.575 3.210 1020.905 3.225 ;
        RECT 1023.335 3.210 1023.665 3.225 ;
        RECT 1020.575 2.910 1023.665 3.210 ;
        RECT 1020.575 2.895 1020.905 2.910 ;
        RECT 1023.335 2.895 1023.665 2.910 ;
        RECT 991.135 2.215 991.465 2.545 ;
        RECT 806.215 1.550 810.210 1.850 ;
        RECT 991.150 1.850 991.450 2.215 ;
        RECT 1053.710 1.850 1054.010 5.630 ;
        RECT 1058.310 2.530 1058.610 5.630 ;
        RECT 1069.350 2.530 1069.650 6.310 ;
        RECT 1073.935 6.295 1074.265 6.310 ;
        RECT 1129.150 5.930 1129.450 13.210 ;
        RECT 1139.270 9.330 1139.570 14.710 ;
        RECT 1301.190 12.050 1301.490 14.710 ;
        RECT 1132.830 9.090 1139.570 9.330 ;
        RECT 1132.390 9.030 1139.570 9.090 ;
        RECT 1147.550 11.750 1170.850 12.050 ;
        RECT 1301.190 11.750 1307.010 12.050 ;
        RECT 1132.390 7.910 1133.570 9.030 ;
        RECT 1137.430 7.670 1138.650 7.970 ;
        RECT 1137.430 6.625 1137.730 7.670 ;
        RECT 1138.350 6.625 1138.650 7.670 ;
        RECT 1147.550 7.290 1147.850 11.750 ;
        RECT 1170.550 8.650 1170.850 11.750 ;
        RECT 1171.455 8.650 1171.785 8.665 ;
        RECT 1170.550 8.350 1171.785 8.650 ;
        RECT 1171.455 8.335 1171.785 8.350 ;
        RECT 1189.855 8.335 1190.185 8.665 ;
        RECT 1189.870 7.970 1190.170 8.335 ;
        RECT 1193.535 7.970 1193.865 7.985 ;
        RECT 1268.975 7.970 1269.305 7.985 ;
        RECT 1189.870 7.670 1193.865 7.970 ;
        RECT 1193.535 7.655 1193.865 7.670 ;
        RECT 1267.150 7.670 1269.305 7.970 ;
        RECT 1267.150 7.305 1267.450 7.670 ;
        RECT 1268.975 7.655 1269.305 7.670 ;
        RECT 1303.030 7.670 1305.170 7.970 ;
        RECT 1303.030 7.305 1303.330 7.670 ;
        RECT 1304.870 7.305 1305.170 7.670 ;
        RECT 1145.710 6.990 1147.850 7.290 ;
        RECT 1145.710 6.625 1146.010 6.990 ;
        RECT 1267.135 6.975 1267.465 7.305 ;
        RECT 1303.015 6.975 1303.345 7.305 ;
        RECT 1304.855 6.975 1305.185 7.305 ;
        RECT 1137.415 6.295 1137.745 6.625 ;
        RECT 1138.335 6.295 1138.665 6.625 ;
        RECT 1145.695 6.295 1146.025 6.625 ;
        RECT 1306.710 6.610 1307.010 11.750 ;
        RECT 1625.030 11.750 1641.890 12.050 ;
        RECT 1428.135 8.335 1428.465 8.665 ;
        RECT 1625.030 8.650 1625.330 11.750 ;
        RECT 1624.110 8.350 1625.330 8.650 ;
        RECT 1641.590 8.650 1641.890 11.750 ;
        RECT 1641.590 8.350 1643.730 8.650 ;
        RECT 1399.630 6.990 1400.850 7.290 ;
        RECT 1314.055 6.610 1314.385 6.625 ;
        RECT 1306.710 6.310 1314.385 6.610 ;
        RECT 1314.055 6.295 1314.385 6.310 ;
        RECT 1324.175 6.295 1324.505 6.625 ;
        RECT 1133.735 5.930 1134.065 5.945 ;
        RECT 1129.150 5.630 1134.065 5.930 ;
        RECT 1133.735 5.615 1134.065 5.630 ;
        RECT 1324.190 3.890 1324.490 6.295 ;
        RECT 1344.415 5.615 1344.745 5.945 ;
        RECT 1397.775 5.615 1398.105 5.945 ;
        RECT 1324.190 3.590 1326.330 3.890 ;
        RECT 1058.310 2.230 1069.650 2.530 ;
        RECT 991.150 1.550 1054.010 1.850 ;
        RECT 1326.030 1.850 1326.330 3.590 ;
        RECT 1344.430 3.210 1344.730 5.615 ;
        RECT 1397.790 5.250 1398.090 5.615 ;
        RECT 1369.270 4.950 1398.090 5.250 ;
        RECT 1369.270 3.210 1369.570 4.950 ;
        RECT 1399.630 3.210 1399.930 6.990 ;
        RECT 1400.550 6.610 1400.850 6.990 ;
        RECT 1402.375 6.975 1402.705 7.305 ;
        RECT 1428.150 7.290 1428.450 8.335 ;
        RECT 1428.150 6.990 1448.690 7.290 ;
        RECT 1402.390 6.610 1402.690 6.975 ;
        RECT 1400.550 6.310 1402.690 6.610 ;
        RECT 1448.390 5.945 1448.690 6.990 ;
        RECT 1450.230 6.990 1454.210 7.290 ;
        RECT 1450.230 5.945 1450.530 6.990 ;
        RECT 1453.910 6.610 1454.210 6.990 ;
        RECT 1624.110 6.625 1624.410 8.350 ;
        RECT 1474.135 6.610 1474.465 6.625 ;
        RECT 1589.135 6.610 1589.465 6.625 ;
        RECT 1453.910 6.310 1455.130 6.610 ;
        RECT 1448.375 5.615 1448.705 5.945 ;
        RECT 1450.215 5.615 1450.545 5.945 ;
        RECT 1454.830 3.890 1455.130 6.310 ;
        RECT 1469.550 6.310 1474.465 6.610 ;
        RECT 1469.550 3.890 1469.850 6.310 ;
        RECT 1474.135 6.295 1474.465 6.310 ;
        RECT 1587.310 6.310 1589.465 6.610 ;
        RECT 1516.470 5.630 1518.610 5.930 ;
        RECT 1516.470 5.265 1516.770 5.630 ;
        RECT 1516.455 4.935 1516.785 5.265 ;
        RECT 1454.830 3.590 1469.850 3.890 ;
        RECT 1344.430 2.910 1369.570 3.210 ;
        RECT 1370.190 2.910 1399.930 3.210 ;
        RECT 1370.190 1.850 1370.490 2.910 ;
        RECT 1326.030 1.550 1370.490 1.850 ;
        RECT 1518.310 1.850 1518.610 5.630 ;
        RECT 1587.310 4.570 1587.610 6.310 ;
        RECT 1589.135 6.295 1589.465 6.310 ;
        RECT 1624.095 6.295 1624.425 6.625 ;
        RECT 1643.430 5.930 1643.730 8.350 ;
        RECT 1643.430 5.630 1645.570 5.930 ;
        RECT 1852.255 5.690 1852.585 5.945 ;
        RECT 1645.270 4.585 1645.570 5.630 ;
        RECT 1575.350 4.270 1587.610 4.570 ;
        RECT 1575.350 1.850 1575.650 4.270 ;
        RECT 1645.255 4.255 1645.585 4.585 ;
        RECT 1697.270 4.510 1698.450 5.690 ;
        RECT 1749.710 4.510 1750.890 5.690 ;
        RECT 1769.030 4.510 1770.210 5.690 ;
        RECT 1851.830 4.510 1853.010 5.690 ;
        RECT 1693.095 2.895 1693.425 3.225 ;
        RECT 1518.310 1.550 1575.650 1.850 ;
        RECT 1693.110 1.850 1693.410 2.895 ;
        RECT 1697.710 1.850 1698.010 4.510 ;
        RECT 1750.150 3.225 1750.450 4.510 ;
        RECT 1769.470 3.905 1769.770 4.510 ;
        RECT 1769.455 3.575 1769.785 3.905 ;
        RECT 1750.135 2.895 1750.465 3.225 ;
        RECT 1952.535 2.895 1952.865 3.225 ;
        RECT 1952.550 1.865 1952.850 2.895 ;
        RECT 2134.710 1.865 2135.010 14.710 ;
        RECT 2365.630 11.750 2367.080 12.050 ;
        RECT 2365.630 1.865 2365.930 11.750 ;
        RECT 2366.780 8.650 2367.080 11.750 ;
        RECT 2566.190 8.665 2566.490 14.710 ;
        RECT 2366.780 8.350 2367.770 8.650 ;
        RECT 2367.470 2.545 2367.770 8.350 ;
        RECT 2566.175 8.335 2566.505 8.665 ;
        RECT 2794.350 7.985 2794.650 49.150 ;
        RECT 2795.270 7.985 2795.570 55.510 ;
        RECT 2800.350 22.250 2801.530 22.690 ;
        RECT 2798.950 21.950 2801.530 22.250 ;
        RECT 2794.335 7.655 2794.665 7.985 ;
        RECT 2795.255 7.655 2795.585 7.985 ;
        RECT 2697.735 3.575 2698.065 3.905 ;
        RECT 2697.750 2.545 2698.050 3.575 ;
        RECT 2798.950 3.225 2799.250 21.950 ;
        RECT 2800.350 21.510 2801.530 21.950 ;
        RECT 2807.230 5.945 2807.530 130.310 ;
        RECT 2845.870 8.665 2846.170 181.750 ;
        RECT 2851.375 61.375 2851.705 61.705 ;
        RECT 2851.390 56.690 2851.690 61.375 ;
        RECT 2850.950 55.510 2852.130 56.690 ;
        RECT 2851.870 21.510 2853.050 22.690 ;
        RECT 2845.855 8.335 2846.185 8.665 ;
        RECT 2807.215 5.615 2807.545 5.945 ;
        RECT 2798.935 2.895 2799.265 3.225 ;
        RECT 2367.455 2.215 2367.785 2.545 ;
        RECT 2697.735 2.215 2698.065 2.545 ;
        RECT 1693.110 1.550 1698.010 1.850 ;
        RECT 806.215 1.535 806.545 1.550 ;
        RECT 1952.535 1.535 1952.865 1.865 ;
        RECT 2134.695 1.535 2135.025 1.865 ;
        RECT 2365.615 1.535 2365.945 1.865 ;
        RECT 427.190 0.190 437.610 0.490 ;
        RECT 393.135 0.175 393.465 0.190 ;
        RECT 415.215 0.175 415.545 0.190 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
        RECT 2954.200 -32.220 2957.200 3551.900 ;
      LAYER via4 ;
        RECT -36.670 3550.610 -35.490 3551.790 ;
        RECT -36.670 3549.010 -35.490 3550.190 ;
        RECT 2955.110 3550.610 2956.290 3551.790 ;
        RECT 2955.110 3549.010 2956.290 3550.190 ;
        RECT -36.670 3485.090 -35.490 3486.270 ;
        RECT -36.670 3483.490 -35.490 3484.670 ;
        RECT -36.670 3305.090 -35.490 3306.270 ;
        RECT -36.670 3303.490 -35.490 3304.670 ;
        RECT -36.670 3125.090 -35.490 3126.270 ;
        RECT -36.670 3123.490 -35.490 3124.670 ;
        RECT -36.670 2945.090 -35.490 2946.270 ;
        RECT -36.670 2943.490 -35.490 2944.670 ;
        RECT -36.670 2765.090 -35.490 2766.270 ;
        RECT -36.670 2763.490 -35.490 2764.670 ;
        RECT -36.670 2585.090 -35.490 2586.270 ;
        RECT -36.670 2583.490 -35.490 2584.670 ;
        RECT -36.670 2405.090 -35.490 2406.270 ;
        RECT -36.670 2403.490 -35.490 2404.670 ;
        RECT -36.670 2225.090 -35.490 2226.270 ;
        RECT -36.670 2223.490 -35.490 2224.670 ;
        RECT -36.670 2045.090 -35.490 2046.270 ;
        RECT -36.670 2043.490 -35.490 2044.670 ;
        RECT -36.670 1865.090 -35.490 1866.270 ;
        RECT -36.670 1863.490 -35.490 1864.670 ;
        RECT -36.670 1685.090 -35.490 1686.270 ;
        RECT -36.670 1683.490 -35.490 1684.670 ;
        RECT -36.670 1505.090 -35.490 1506.270 ;
        RECT -36.670 1503.490 -35.490 1504.670 ;
        RECT -36.670 1325.090 -35.490 1326.270 ;
        RECT -36.670 1323.490 -35.490 1324.670 ;
        RECT -36.670 1145.090 -35.490 1146.270 ;
        RECT -36.670 1143.490 -35.490 1144.670 ;
        RECT -36.670 965.090 -35.490 966.270 ;
        RECT -36.670 963.490 -35.490 964.670 ;
        RECT -36.670 785.090 -35.490 786.270 ;
        RECT -36.670 783.490 -35.490 784.670 ;
        RECT -36.670 605.090 -35.490 606.270 ;
        RECT -36.670 603.490 -35.490 604.670 ;
        RECT -36.670 425.090 -35.490 426.270 ;
        RECT -36.670 423.490 -35.490 424.670 ;
        RECT -36.670 245.090 -35.490 246.270 ;
        RECT -36.670 243.490 -35.490 244.670 ;
        RECT -36.670 65.090 -35.490 66.270 ;
        RECT -36.670 63.490 -35.490 64.670 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
        RECT 2955.110 3485.090 2956.290 3486.270 ;
        RECT 2955.110 3483.490 2956.290 3484.670 ;
        RECT 2955.110 3305.090 2956.290 3306.270 ;
        RECT 2955.110 3303.490 2956.290 3304.670 ;
        RECT 2955.110 3125.090 2956.290 3126.270 ;
        RECT 2955.110 3123.490 2956.290 3124.670 ;
        RECT 2955.110 2945.090 2956.290 2946.270 ;
        RECT 2955.110 2943.490 2956.290 2944.670 ;
        RECT 2955.110 2765.090 2956.290 2766.270 ;
        RECT 2955.110 2763.490 2956.290 2764.670 ;
        RECT 2955.110 2585.090 2956.290 2586.270 ;
        RECT 2955.110 2583.490 2956.290 2584.670 ;
        RECT 2955.110 2405.090 2956.290 2406.270 ;
        RECT 2955.110 2403.490 2956.290 2404.670 ;
        RECT 2955.110 2225.090 2956.290 2226.270 ;
        RECT 2955.110 2223.490 2956.290 2224.670 ;
        RECT 2955.110 2045.090 2956.290 2046.270 ;
        RECT 2955.110 2043.490 2956.290 2044.670 ;
        RECT 2955.110 1865.090 2956.290 1866.270 ;
        RECT 2955.110 1863.490 2956.290 1864.670 ;
        RECT 2955.110 1685.090 2956.290 1686.270 ;
        RECT 2955.110 1683.490 2956.290 1684.670 ;
        RECT 2955.110 1505.090 2956.290 1506.270 ;
        RECT 2955.110 1503.490 2956.290 1504.670 ;
        RECT 2955.110 1325.090 2956.290 1326.270 ;
        RECT 2955.110 1323.490 2956.290 1324.670 ;
        RECT 2955.110 1145.090 2956.290 1146.270 ;
        RECT 2955.110 1143.490 2956.290 1144.670 ;
        RECT 2955.110 965.090 2956.290 966.270 ;
        RECT 2955.110 963.490 2956.290 964.670 ;
        RECT 2955.110 785.090 2956.290 786.270 ;
        RECT 2955.110 783.490 2956.290 784.670 ;
        RECT 2955.110 605.090 2956.290 606.270 ;
        RECT 2955.110 603.490 2956.290 604.670 ;
        RECT 2955.110 425.090 2956.290 426.270 ;
        RECT 2955.110 423.490 2956.290 424.670 ;
        RECT 2955.110 245.090 2956.290 246.270 ;
        RECT 2955.110 243.490 2956.290 244.670 ;
        RECT 2955.110 65.090 2956.290 66.270 ;
        RECT 2955.110 63.490 2956.290 64.670 ;
        RECT -36.670 -30.510 -35.490 -29.330 ;
        RECT -36.670 -32.110 -35.490 -30.930 ;
        RECT 2955.110 -30.510 2956.290 -29.330 ;
        RECT 2955.110 -32.110 2956.290 -30.930 ;
      LAYER met5 ;
        RECT -37.580 3551.900 -34.580 3551.910 ;
        RECT 2954.200 3551.900 2957.200 3551.910 ;
        RECT -37.580 3548.900 2957.200 3551.900 ;
        RECT -37.580 3548.890 -34.580 3548.900 ;
        RECT 2954.200 3548.890 2957.200 3548.900 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -37.580 3486.380 -34.580 3486.390 ;
        RECT 2954.200 3486.380 2957.200 3486.390 ;
        RECT -42.180 3483.380 2961.800 3486.380 ;
        RECT -37.580 3483.370 -34.580 3483.380 ;
        RECT 2954.200 3483.370 2957.200 3483.380 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.580 3429.380 2934.200 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT 2793.700 3380.500 2799.900 3382.100 ;
        RECT -37.580 3306.380 -34.580 3306.390 ;
        RECT 2954.200 3306.380 2957.200 3306.390 ;
        RECT -42.180 3303.380 2961.800 3306.380 ;
        RECT -37.580 3303.370 -34.580 3303.380 ;
        RECT 2954.200 3303.370 2957.200 3303.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.580 3249.380 2934.200 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -37.580 3126.380 -34.580 3126.390 ;
        RECT 2954.200 3126.380 2957.200 3126.390 ;
        RECT -42.180 3123.380 2961.800 3126.380 ;
        RECT -37.580 3123.370 -34.580 3123.380 ;
        RECT 2954.200 3123.370 2957.200 3123.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.580 3069.380 2934.200 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -37.580 2946.380 -34.580 2946.390 ;
        RECT 2954.200 2946.380 2957.200 2946.390 ;
        RECT -42.180 2943.380 2961.800 2946.380 ;
        RECT -37.580 2943.370 -34.580 2943.380 ;
        RECT 2954.200 2943.370 2957.200 2943.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.580 2889.380 2934.200 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -37.580 2766.380 -34.580 2766.390 ;
        RECT 2954.200 2766.380 2957.200 2766.390 ;
        RECT -42.180 2763.380 2961.800 2766.380 ;
        RECT -37.580 2763.370 -34.580 2763.380 ;
        RECT 2954.200 2763.370 2957.200 2763.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.580 2709.380 2934.200 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -37.580 2586.380 -34.580 2586.390 ;
        RECT 2954.200 2586.380 2957.200 2586.390 ;
        RECT -42.180 2583.380 2961.800 2586.380 ;
        RECT -37.580 2583.370 -34.580 2583.380 ;
        RECT 2954.200 2583.370 2957.200 2583.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.580 2529.380 2934.200 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -37.580 2406.380 -34.580 2406.390 ;
        RECT 2954.200 2406.380 2957.200 2406.390 ;
        RECT -42.180 2403.380 2961.800 2406.380 ;
        RECT -37.580 2403.370 -34.580 2403.380 ;
        RECT 2954.200 2403.370 2957.200 2403.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.580 2349.380 2934.200 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -37.580 2226.380 -34.580 2226.390 ;
        RECT 2954.200 2226.380 2957.200 2226.390 ;
        RECT -42.180 2223.380 2961.800 2226.380 ;
        RECT -37.580 2223.370 -34.580 2223.380 ;
        RECT 2954.200 2223.370 2957.200 2223.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.580 2169.380 2934.200 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -37.580 2046.380 -34.580 2046.390 ;
        RECT 2954.200 2046.380 2957.200 2046.390 ;
        RECT -42.180 2043.380 2961.800 2046.380 ;
        RECT -37.580 2043.370 -34.580 2043.380 ;
        RECT 2954.200 2043.370 2957.200 2043.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.580 1989.380 2934.200 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -37.580 1866.380 -34.580 1866.390 ;
        RECT 2954.200 1866.380 2957.200 1866.390 ;
        RECT -42.180 1863.380 2961.800 1866.380 ;
        RECT -37.580 1863.370 -34.580 1863.380 ;
        RECT 2954.200 1863.370 2957.200 1863.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.580 1809.380 2934.200 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -37.580 1686.380 -34.580 1686.390 ;
        RECT 2954.200 1686.380 2957.200 1686.390 ;
        RECT -42.180 1683.380 2961.800 1686.380 ;
        RECT -37.580 1683.370 -34.580 1683.380 ;
        RECT 2954.200 1683.370 2957.200 1683.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.580 1629.380 2934.200 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -37.580 1506.380 -34.580 1506.390 ;
        RECT 2954.200 1506.380 2957.200 1506.390 ;
        RECT -42.180 1503.380 2961.800 1506.380 ;
        RECT -37.580 1503.370 -34.580 1503.380 ;
        RECT 2954.200 1503.370 2957.200 1503.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.580 1449.380 2934.200 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -37.580 1326.380 -34.580 1326.390 ;
        RECT 2954.200 1326.380 2957.200 1326.390 ;
        RECT -42.180 1323.380 2961.800 1326.380 ;
        RECT -37.580 1323.370 -34.580 1323.380 ;
        RECT 2954.200 1323.370 2957.200 1323.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.580 1269.380 2934.200 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -37.580 1146.380 -34.580 1146.390 ;
        RECT 2954.200 1146.380 2957.200 1146.390 ;
        RECT -42.180 1143.380 2961.800 1146.380 ;
        RECT -37.580 1143.370 -34.580 1143.380 ;
        RECT 2954.200 1143.370 2957.200 1143.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.580 1089.380 2934.200 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -37.580 966.380 -34.580 966.390 ;
        RECT 2954.200 966.380 2957.200 966.390 ;
        RECT -42.180 963.380 2961.800 966.380 ;
        RECT -37.580 963.370 -34.580 963.380 ;
        RECT 2954.200 963.370 2957.200 963.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.580 909.380 2934.200 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -37.580 786.380 -34.580 786.390 ;
        RECT 2954.200 786.380 2957.200 786.390 ;
        RECT -42.180 783.380 2961.800 786.380 ;
        RECT -37.580 783.370 -34.580 783.380 ;
        RECT 2954.200 783.370 2957.200 783.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.580 729.380 2934.200 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -37.580 606.380 -34.580 606.390 ;
        RECT 2954.200 606.380 2957.200 606.390 ;
        RECT -42.180 603.380 2961.800 606.380 ;
        RECT -37.580 603.370 -34.580 603.380 ;
        RECT 2954.200 603.370 2957.200 603.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.580 549.380 2934.200 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -37.580 426.380 -34.580 426.390 ;
        RECT 2954.200 426.380 2957.200 426.390 ;
        RECT -42.180 423.380 2961.800 426.380 ;
        RECT -37.580 423.370 -34.580 423.380 ;
        RECT 2954.200 423.370 2957.200 423.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.580 369.380 2934.200 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -37.580 246.380 -34.580 246.390 ;
        RECT 2954.200 246.380 2957.200 246.390 ;
        RECT -42.180 243.380 2961.800 246.380 ;
        RECT -37.580 243.370 -34.580 243.380 ;
        RECT 2954.200 243.370 2957.200 243.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.580 189.380 2934.200 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT 8.860 130.100 2808.180 131.700 ;
        RECT 996.940 96.100 1030.740 97.700 ;
        RECT 996.940 94.300 998.540 96.100 ;
        RECT 281.180 92.700 316.820 94.300 ;
        RECT 130.300 85.900 211.940 87.500 ;
        RECT 130.300 80.700 131.900 85.900 ;
        RECT 104.540 79.100 131.900 80.700 ;
        RECT 133.980 79.100 186.180 80.700 ;
        RECT 104.540 77.300 106.140 79.100 ;
        RECT 4.260 75.700 106.140 77.300 ;
        RECT 133.980 73.900 135.580 79.100 ;
        RECT 116.500 72.300 135.580 73.900 ;
        RECT 184.580 73.900 186.180 79.100 ;
        RECT 210.340 77.300 211.940 85.900 ;
        RECT 281.180 84.100 282.780 92.700 ;
        RECT 261.860 82.500 282.780 84.100 ;
        RECT 261.860 77.300 263.460 82.500 ;
        RECT 315.220 80.700 316.820 92.700 ;
        RECT 995.100 92.700 998.540 94.300 ;
        RECT 1001.540 92.700 1023.380 94.300 ;
        RECT 605.940 84.100 608.460 87.500 ;
        RECT 702.540 84.100 705.060 87.500 ;
        RECT 799.140 84.100 801.660 87.500 ;
        RECT 995.100 84.100 996.700 92.700 ;
        RECT 490.020 82.500 537.620 84.100 ;
        RECT 315.220 79.100 469.540 80.700 ;
        RECT 210.340 75.700 263.460 77.300 ;
        RECT 467.940 77.300 469.540 79.100 ;
        RECT 490.020 77.300 491.620 82.500 ;
        RECT 467.940 75.700 491.620 77.300 ;
        RECT 536.020 77.300 537.620 82.500 ;
        RECT 570.980 82.500 608.460 84.100 ;
        RECT 570.980 77.300 572.580 82.500 ;
        RECT 606.860 80.700 608.460 82.500 ;
        RECT 667.580 82.500 705.060 84.100 ;
        RECT 606.860 79.100 622.260 80.700 ;
        RECT 536.020 75.700 572.580 77.300 ;
        RECT 620.660 77.300 622.260 79.100 ;
        RECT 667.580 77.300 669.180 82.500 ;
        RECT 703.460 80.700 705.060 82.500 ;
        RECT 727.380 82.500 745.540 84.100 ;
        RECT 727.380 80.700 728.980 82.500 ;
        RECT 703.460 79.100 728.980 80.700 ;
        RECT 743.940 80.700 745.540 82.500 ;
        RECT 747.620 82.500 866.980 84.100 ;
        RECT 747.620 80.700 749.220 82.500 ;
        RECT 743.940 79.100 749.220 80.700 ;
        RECT 865.380 80.700 866.980 82.500 ;
        RECT 972.100 82.500 996.700 84.100 ;
        RECT 865.380 79.100 930.460 80.700 ;
        RECT 620.660 75.700 669.180 77.300 ;
        RECT 743.940 75.700 746.460 79.100 ;
        RECT 928.860 77.300 930.460 79.100 ;
        RECT 972.100 77.300 973.700 82.500 ;
        RECT 1001.540 80.700 1003.140 92.700 ;
        RECT 928.860 75.700 973.700 77.300 ;
        RECT 995.100 79.100 1003.140 80.700 ;
        RECT 995.100 73.900 996.700 79.100 ;
        RECT 184.580 72.300 190.780 73.900 ;
        RECT 116.500 70.500 118.100 72.300 ;
        RECT 8.860 68.900 25.180 70.500 ;
        RECT 103.620 69.800 118.100 70.500 ;
        RECT 99.940 68.900 118.100 69.800 ;
        RECT 189.180 70.500 190.780 72.300 ;
        RECT 244.380 72.300 263.460 73.900 ;
        RECT 244.380 70.500 245.980 72.300 ;
        RECT 189.180 68.900 245.980 70.500 ;
        RECT 261.860 70.500 263.460 72.300 ;
        RECT 324.420 72.300 367.420 73.900 ;
        RECT 324.420 70.500 326.020 72.300 ;
        RECT 261.860 68.900 326.020 70.500 ;
        RECT 365.820 70.500 367.420 72.300 ;
        RECT 459.660 72.300 996.700 73.900 ;
        RECT 1021.780 73.900 1023.380 92.700 ;
        RECT 1029.140 87.500 1030.740 96.100 ;
        RECT 2737.580 96.100 2756.660 97.700 ;
        RECT 1331.820 89.300 1380.340 90.900 ;
        RECT 1029.140 85.900 1033.500 87.500 ;
        RECT 1031.900 80.700 1033.500 85.900 ;
        RECT 1062.260 82.500 1131.940 84.100 ;
        RECT 1062.260 80.700 1063.860 82.500 ;
        RECT 1031.900 79.100 1063.860 80.700 ;
        RECT 1130.340 77.300 1131.940 82.500 ;
        RECT 1134.020 82.500 1180.700 84.100 ;
        RECT 1134.020 77.300 1135.620 82.500 ;
        RECT 1179.100 80.700 1180.700 82.500 ;
        RECT 1230.620 82.500 1274.540 84.100 ;
        RECT 1130.340 75.700 1135.620 77.300 ;
        RECT 1137.700 79.100 1174.260 80.700 ;
        RECT 1179.100 79.100 1228.540 80.700 ;
        RECT 1137.700 73.900 1139.300 79.100 ;
        RECT 1172.660 77.300 1174.260 79.100 ;
        RECT 1226.940 77.300 1228.540 79.100 ;
        RECT 1230.620 77.300 1232.220 82.500 ;
        RECT 1272.940 80.700 1274.540 82.500 ;
        RECT 1284.900 82.500 1315.020 84.100 ;
        RECT 1272.940 79.100 1275.460 80.700 ;
        RECT 1172.660 75.700 1177.020 77.300 ;
        RECT 1226.940 75.700 1232.220 77.300 ;
        RECT 1273.860 77.300 1275.460 79.100 ;
        RECT 1284.900 77.300 1286.500 82.500 ;
        RECT 1273.860 75.700 1286.500 77.300 ;
        RECT 1313.420 77.300 1315.020 82.500 ;
        RECT 1331.820 77.300 1333.420 89.300 ;
        RECT 1313.420 75.700 1333.420 77.300 ;
        RECT 1378.740 77.300 1380.340 89.300 ;
        RECT 2737.580 87.500 2739.180 96.100 ;
        RECT 2755.060 94.300 2756.660 96.100 ;
        RECT 2755.060 92.700 2799.900 94.300 ;
        RECT 2728.380 85.900 2739.180 87.500 ;
        RECT 1444.980 79.100 1466.820 80.700 ;
        RECT 1444.980 77.300 1446.580 79.100 ;
        RECT 1378.740 75.700 1446.580 77.300 ;
        RECT 1465.220 77.300 1466.820 79.100 ;
        RECT 1541.580 79.100 1563.420 80.700 ;
        RECT 1541.580 77.300 1543.180 79.100 ;
        RECT 1465.220 75.700 1543.180 77.300 ;
        RECT 1561.820 77.300 1563.420 79.100 ;
        RECT 1638.180 79.100 1660.020 80.700 ;
        RECT 1638.180 77.300 1639.780 79.100 ;
        RECT 1561.820 75.700 1639.780 77.300 ;
        RECT 1658.420 77.300 1660.020 79.100 ;
        RECT 1734.780 79.100 1756.620 80.700 ;
        RECT 1734.780 77.300 1736.380 79.100 ;
        RECT 1658.420 75.700 1736.380 77.300 ;
        RECT 1755.020 77.300 1756.620 79.100 ;
        RECT 1831.380 79.100 1853.220 80.700 ;
        RECT 1831.380 77.300 1832.980 79.100 ;
        RECT 1755.020 75.700 1832.980 77.300 ;
        RECT 1851.620 77.300 1853.220 79.100 ;
        RECT 1927.980 79.100 1949.820 80.700 ;
        RECT 1927.980 77.300 1929.580 79.100 ;
        RECT 1851.620 75.700 1929.580 77.300 ;
        RECT 1948.220 77.300 1949.820 79.100 ;
        RECT 2024.580 79.100 2046.420 80.700 ;
        RECT 2024.580 77.300 2026.180 79.100 ;
        RECT 1948.220 75.700 2026.180 77.300 ;
        RECT 2044.820 77.300 2046.420 79.100 ;
        RECT 2121.180 79.100 2143.020 80.700 ;
        RECT 2121.180 77.300 2122.780 79.100 ;
        RECT 2044.820 75.700 2122.780 77.300 ;
        RECT 2141.420 77.300 2143.020 79.100 ;
        RECT 2217.780 79.100 2239.620 80.700 ;
        RECT 2217.780 77.300 2219.380 79.100 ;
        RECT 2141.420 75.700 2219.380 77.300 ;
        RECT 2238.020 77.300 2239.620 79.100 ;
        RECT 2314.380 79.100 2336.220 80.700 ;
        RECT 2314.380 77.300 2315.980 79.100 ;
        RECT 2238.020 75.700 2315.980 77.300 ;
        RECT 2334.620 77.300 2336.220 79.100 ;
        RECT 2410.980 79.100 2432.820 80.700 ;
        RECT 2410.980 77.300 2412.580 79.100 ;
        RECT 2334.620 75.700 2412.580 77.300 ;
        RECT 2431.220 77.300 2432.820 79.100 ;
        RECT 2507.580 79.100 2529.420 80.700 ;
        RECT 2507.580 77.300 2509.180 79.100 ;
        RECT 2431.220 75.700 2509.180 77.300 ;
        RECT 2527.820 77.300 2529.420 79.100 ;
        RECT 2604.180 79.100 2626.020 80.700 ;
        RECT 2604.180 77.300 2605.780 79.100 ;
        RECT 2527.820 75.700 2605.780 77.300 ;
        RECT 2624.420 77.300 2626.020 79.100 ;
        RECT 2728.380 77.300 2729.980 85.900 ;
        RECT 2744.940 79.100 2795.300 80.700 ;
        RECT 2744.940 77.300 2746.540 79.100 ;
        RECT 2624.420 75.700 2729.980 77.300 ;
        RECT 2743.100 75.700 2746.540 77.300 ;
        RECT 1021.780 72.300 1139.300 73.900 ;
        RECT 459.660 70.500 461.260 72.300 ;
        RECT 365.820 68.900 461.260 70.500 ;
        RECT 1175.420 70.500 1177.020 75.700 ;
        RECT 1186.460 72.300 2691.340 73.900 ;
        RECT 1186.460 70.500 1188.060 72.300 ;
        RECT 1175.420 68.900 1188.060 70.500 ;
        RECT 2282.180 68.900 2284.700 72.300 ;
        RECT 2378.780 68.900 2381.300 72.300 ;
        RECT 2475.380 68.900 2477.900 72.300 ;
        RECT 2571.980 68.900 2574.500 72.300 ;
        RECT 2689.740 70.500 2691.340 72.300 ;
        RECT 2743.100 70.500 2744.700 75.700 ;
        RECT 2689.740 68.900 2744.700 70.500 ;
        RECT 99.940 68.200 105.220 68.900 ;
        RECT -37.580 66.380 -34.580 66.390 ;
        RECT 99.940 66.380 101.540 68.200 ;
        RECT 2954.200 66.380 2957.200 66.390 ;
        RECT -42.180 63.380 2961.800 66.380 ;
        RECT -37.580 63.370 -34.580 63.380 ;
        RECT 391.580 62.100 406.060 63.380 ;
        RECT 2954.200 63.370 2957.200 63.380 ;
        RECT 391.580 60.300 393.180 62.100 ;
        RECT 23.580 58.700 52.780 60.300 ;
        RECT 51.180 56.900 52.780 58.700 ;
        RECT 56.700 58.700 152.140 60.300 ;
        RECT 56.700 56.900 58.300 58.700 ;
        RECT 150.540 56.900 152.140 58.700 ;
        RECT 169.860 58.700 234.940 60.300 ;
        RECT 51.180 55.300 58.300 56.900 ;
        RECT 63.140 55.300 142.940 56.900 ;
        RECT 63.140 53.500 64.740 55.300 ;
        RECT 7.020 51.900 64.740 53.500 ;
        RECT 141.340 53.500 142.940 55.300 ;
        RECT 145.020 55.300 155.820 56.900 ;
        RECT 145.020 53.500 146.620 55.300 ;
        RECT 141.340 51.900 146.620 53.500 ;
        RECT 150.540 50.100 152.140 55.300 ;
        RECT 154.220 53.500 155.820 55.300 ;
        RECT 169.860 53.500 171.460 58.700 ;
        RECT 233.340 56.900 234.940 58.700 ;
        RECT 310.620 58.700 324.180 60.300 ;
        RECT 310.620 56.900 312.220 58.700 ;
        RECT 322.580 56.900 324.180 58.700 ;
        RECT 329.020 58.700 393.180 60.300 ;
        RECT 404.460 60.300 406.060 62.100 ;
        RECT 404.460 58.700 416.180 60.300 ;
        RECT 329.020 56.900 330.620 58.700 ;
        RECT 414.580 56.900 416.180 58.700 ;
        RECT 459.660 58.700 528.420 60.300 ;
        RECT 459.660 56.900 461.260 58.700 ;
        RECT 526.820 56.900 528.420 58.700 ;
        RECT 559.940 58.700 589.140 60.300 ;
        RECT 559.940 56.900 561.540 58.700 ;
        RECT 154.220 51.900 171.460 53.500 ;
        RECT 174.460 55.300 312.220 56.900 ;
        RECT 315.220 55.300 330.620 56.900 ;
        RECT 336.380 55.300 362.820 56.900 ;
        RECT 414.580 55.300 461.260 56.900 ;
        RECT 463.340 55.300 520.140 56.900 ;
        RECT 526.820 55.300 561.540 56.900 ;
        RECT 587.540 56.900 589.140 58.700 ;
        RECT 592.140 58.700 751.980 60.300 ;
        RECT 592.140 56.900 593.740 58.700 ;
        RECT 750.380 56.900 751.980 58.700 ;
        RECT 754.980 58.700 764.860 60.300 ;
        RECT 754.980 56.900 756.580 58.700 ;
        RECT 763.260 56.900 764.860 58.700 ;
        RECT 766.940 58.700 773.140 60.300 ;
        RECT 766.940 56.900 768.540 58.700 ;
        RECT 587.540 55.300 593.740 56.900 ;
        RECT 598.580 55.300 644.340 56.900 ;
        RECT 174.460 50.100 176.060 55.300 ;
        RECT 233.340 53.500 234.940 55.300 ;
        RECT 315.220 53.500 316.820 55.300 ;
        RECT 233.340 51.900 316.820 53.500 ;
        RECT 322.580 53.500 324.180 55.300 ;
        RECT 336.380 53.500 337.980 55.300 ;
        RECT 322.580 51.900 337.980 53.500 ;
        RECT 361.220 53.500 362.820 55.300 ;
        RECT 463.340 53.500 464.940 55.300 ;
        RECT 361.220 51.900 464.940 53.500 ;
        RECT 518.540 53.500 520.140 55.300 ;
        RECT 598.580 53.500 600.180 55.300 ;
        RECT 518.540 51.900 600.180 53.500 ;
        RECT 642.740 53.500 644.340 55.300 ;
        RECT 654.700 55.300 663.660 56.900 ;
        RECT 750.380 55.300 758.420 56.900 ;
        RECT 763.260 55.300 768.540 56.900 ;
        RECT 771.540 56.900 773.140 58.700 ;
        RECT 893.900 58.700 911.140 60.300 ;
        RECT 893.900 56.900 895.500 58.700 ;
        RECT 909.540 56.900 911.140 58.700 ;
        RECT 924.260 58.700 935.060 60.300 ;
        RECT 924.260 56.900 925.860 58.700 ;
        RECT 771.540 55.300 899.180 56.900 ;
        RECT 909.540 55.300 925.860 56.900 ;
        RECT 933.460 56.900 935.060 58.700 ;
        RECT 937.140 56.900 939.660 60.300 ;
        RECT 1009.820 58.700 1091.460 60.300 ;
        RECT 1009.820 56.900 1011.420 58.700 ;
        RECT 1089.860 56.900 1091.460 58.700 ;
        RECT 1127.580 58.700 1146.660 60.300 ;
        RECT 1127.580 56.900 1129.180 58.700 ;
        RECT 933.460 55.300 1011.420 56.900 ;
        RECT 1037.420 55.300 1084.100 56.900 ;
        RECT 1089.860 55.300 1129.180 56.900 ;
        RECT 1145.060 56.900 1146.660 58.700 ;
        RECT 1235.220 58.700 1248.780 60.300 ;
        RECT 1235.220 56.900 1236.820 58.700 ;
        RECT 1247.180 56.900 1248.780 58.700 ;
        RECT 1251.780 58.700 1310.420 60.300 ;
        RECT 1251.780 56.900 1253.380 58.700 ;
        RECT 1145.060 55.300 1236.820 56.900 ;
        RECT 1238.900 55.300 1245.100 56.900 ;
        RECT 1247.180 55.300 1253.380 56.900 ;
        RECT 1308.820 56.900 1310.420 58.700 ;
        RECT 1329.980 58.700 1576.300 60.300 ;
        RECT 1329.980 56.900 1331.580 58.700 ;
        RECT 1574.700 56.900 1576.300 58.700 ;
        RECT 1619.780 58.700 1671.060 60.300 ;
        RECT 1619.780 56.900 1621.380 58.700 ;
        RECT 1669.460 56.900 1671.060 58.700 ;
        RECT 1699.820 58.700 1724.420 60.300 ;
        RECT 1699.820 56.900 1701.420 58.700 ;
        RECT 1722.820 56.900 1724.420 58.700 ;
        RECT 1728.340 58.700 1869.780 60.300 ;
        RECT 1728.340 56.900 1729.940 58.700 ;
        RECT 1868.180 56.900 1869.780 58.700 ;
        RECT 1904.060 58.700 2794.380 60.300 ;
        RECT 1904.060 56.900 1905.660 58.700 ;
        RECT 1308.820 55.300 1331.580 56.900 ;
        RECT 1348.380 55.300 1443.820 56.900 ;
        RECT 1574.700 55.300 1621.380 56.900 ;
        RECT 1644.620 55.300 1658.180 56.900 ;
        RECT 1669.460 55.300 1701.420 56.900 ;
        RECT 1713.620 55.300 1719.820 56.900 ;
        RECT 1722.820 55.300 1729.940 56.900 ;
        RECT 1736.620 55.300 1866.100 56.900 ;
        RECT 1868.180 55.300 1905.660 56.900 ;
        RECT 1907.740 55.300 2161.420 56.900 ;
        RECT 654.700 53.500 656.300 55.300 ;
        RECT 642.740 51.900 656.300 53.500 ;
        RECT 662.060 53.500 663.660 55.300 ;
        RECT 752.220 53.500 753.820 55.300 ;
        RECT 662.060 51.900 753.820 53.500 ;
        RECT 756.820 53.500 758.420 55.300 ;
        RECT 893.900 53.500 895.500 55.300 ;
        RECT 756.820 51.900 895.500 53.500 ;
        RECT 897.580 53.500 899.180 55.300 ;
        RECT 1037.420 53.500 1039.020 55.300 ;
        RECT 897.580 51.900 1039.020 53.500 ;
        RECT 1082.500 53.500 1084.100 55.300 ;
        RECT 1238.900 53.500 1240.500 55.300 ;
        RECT 1082.500 51.900 1240.500 53.500 ;
        RECT 1243.500 53.500 1245.100 55.300 ;
        RECT 1348.380 53.500 1349.980 55.300 ;
        RECT 1243.500 51.900 1349.980 53.500 ;
        RECT 1442.220 53.500 1443.820 55.300 ;
        RECT 1644.620 53.500 1646.220 55.300 ;
        RECT 1442.220 51.900 1646.220 53.500 ;
        RECT 1656.580 53.500 1658.180 55.300 ;
        RECT 1713.620 53.500 1715.220 55.300 ;
        RECT 1656.580 51.900 1715.220 53.500 ;
        RECT 1718.220 53.500 1719.820 55.300 ;
        RECT 1736.620 53.500 1738.220 55.300 ;
        RECT 1718.220 51.900 1738.220 53.500 ;
        RECT 1864.500 53.500 1866.100 55.300 ;
        RECT 1907.740 53.500 1909.340 55.300 ;
        RECT 1864.500 51.900 1909.340 53.500 ;
        RECT 2159.820 53.500 2161.420 55.300 ;
        RECT 2217.780 55.300 2223.060 56.900 ;
        RECT 2217.780 53.500 2219.380 55.300 ;
        RECT 2159.820 51.900 2219.380 53.500 ;
        RECT 2221.460 53.500 2223.060 55.300 ;
        RECT 2268.380 55.300 2273.660 56.900 ;
        RECT 2268.380 53.500 2269.980 55.300 ;
        RECT 2221.460 51.900 2269.980 53.500 ;
        RECT 2272.060 53.500 2273.660 55.300 ;
        RECT 2314.380 55.300 2319.660 56.900 ;
        RECT 2314.380 53.500 2315.980 55.300 ;
        RECT 2272.060 51.900 2315.980 53.500 ;
        RECT 2318.060 53.500 2319.660 55.300 ;
        RECT 2364.980 55.300 2370.260 56.900 ;
        RECT 2364.980 53.500 2366.580 55.300 ;
        RECT 2318.060 51.900 2366.580 53.500 ;
        RECT 2368.660 53.500 2370.260 55.300 ;
        RECT 2410.980 55.300 2416.260 56.900 ;
        RECT 2410.980 53.500 2412.580 55.300 ;
        RECT 2368.660 51.900 2412.580 53.500 ;
        RECT 2414.660 53.500 2416.260 55.300 ;
        RECT 2461.580 55.300 2466.860 56.900 ;
        RECT 2461.580 53.500 2463.180 55.300 ;
        RECT 2414.660 51.900 2463.180 53.500 ;
        RECT 2465.260 53.500 2466.860 55.300 ;
        RECT 2507.580 55.300 2512.860 56.900 ;
        RECT 2507.580 53.500 2509.180 55.300 ;
        RECT 2465.260 51.900 2509.180 53.500 ;
        RECT 2511.260 53.500 2512.860 55.300 ;
        RECT 2558.180 55.300 2654.540 56.900 ;
        RECT 2558.180 53.500 2559.780 55.300 ;
        RECT 2511.260 51.900 2559.780 53.500 ;
        RECT 2652.940 53.500 2654.540 55.300 ;
        RECT 2701.700 55.300 2796.220 56.900 ;
        RECT 2798.300 55.300 2852.340 56.900 ;
        RECT 2701.700 53.500 2703.300 55.300 ;
        RECT 2652.940 51.900 2703.300 53.500 ;
        RECT 150.540 48.500 176.060 50.100 ;
        RECT 776.140 21.300 975.540 22.900 ;
        RECT 678.620 17.900 735.650 19.500 ;
        RECT 260.940 14.500 375.700 16.100 ;
        RECT 513.020 14.500 627.780 16.100 ;
        RECT 678.620 14.500 680.220 17.900 ;
        RECT 734.050 16.100 735.650 17.900 ;
        RECT 734.050 14.500 769.460 16.100 ;
        RECT 776.140 14.500 777.740 21.300 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 973.940 12.380 975.540 21.300 ;
        RECT 1128.500 13.000 1130.100 26.300 ;
        RECT 2288.620 21.300 2443.630 22.900 ;
        RECT 2288.620 19.500 2290.220 21.300 ;
        RECT 1138.620 17.900 1285.580 19.500 ;
        RECT 1138.620 14.500 1140.220 17.900 ;
        RECT 1283.980 16.100 1285.580 17.900 ;
        RECT 2134.060 17.900 2290.220 19.500 ;
        RECT 2442.030 19.500 2443.630 21.300 ;
        RECT 2445.940 21.300 2451.910 22.900 ;
        RECT 2445.940 19.500 2447.540 21.300 ;
        RECT 2442.030 17.900 2447.540 19.500 ;
        RECT 2450.310 19.500 2451.910 21.300 ;
        RECT 2454.220 21.300 2497.220 22.900 ;
        RECT 2800.140 21.300 2853.260 22.900 ;
        RECT 2450.310 17.900 2452.140 19.500 ;
        RECT 1283.980 14.500 1302.140 16.100 ;
        RECT 2134.060 14.500 2135.660 17.900 ;
        RECT 2450.540 16.100 2452.140 17.900 ;
        RECT 2454.220 16.100 2455.820 21.300 ;
        RECT 2495.620 19.500 2497.220 21.300 ;
        RECT 2495.620 17.900 2567.140 19.500 ;
        RECT 2450.540 14.500 2455.820 16.100 ;
        RECT 2565.540 14.500 2567.140 17.900 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.580 9.380 2934.200 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 769.930 8.380 796.140 9.380 ;
        RECT 1119.300 9.300 1120.900 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT 1119.300 7.700 1133.780 9.300 ;
        RECT 807.420 5.900 809.020 7.260 ;
        RECT 800.060 4.300 809.020 5.900 ;
        RECT 1697.060 4.300 1751.100 5.900 ;
        RECT 1768.820 4.300 1853.220 5.900 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
        RECT -37.580 -29.220 -34.580 -29.210 ;
        RECT 2954.200 -29.220 2957.200 -29.210 ;
        RECT -37.580 -32.220 2957.200 -29.220 ;
        RECT -37.580 -32.230 -34.580 -32.220 ;
        RECT 2954.200 -32.230 2957.200 -32.220 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2849.845 2755.105 2850.015 2760.375 ;
        RECT 2850.305 2643.585 2850.475 2655.655 ;
        RECT 2849.845 2592.245 2850.015 2613.155 ;
        RECT 2849.845 2515.065 2850.015 2525.775 ;
        RECT 2849.385 2342.685 2850.015 2342.855 ;
        RECT 2849.385 2307.155 2849.555 2342.685 ;
        RECT 2849.385 2306.985 2850.015 2307.155 ;
        RECT 2850.305 2183.905 2850.475 2208.215 ;
        RECT 2849.845 2011.185 2850.015 2090.235 ;
        RECT 2849.385 1788.145 2850.015 1788.315 ;
        RECT 2851.225 1788.145 2851.395 1883.515 ;
        RECT 2849.385 1724.395 2849.555 1788.145 ;
        RECT 2849.385 1724.225 2850.015 1724.395 ;
        RECT 2849.845 1656.225 2850.015 1711.135 ;
        RECT 2849.845 1605.565 2850.015 1655.375 ;
        RECT 2849.845 1589.585 2850.015 1603.695 ;
        RECT 2850.305 1482.825 2850.475 1500.675 ;
        RECT 2850.305 1418.395 2850.475 1448.995 ;
        RECT 2850.765 1448.825 2850.935 1459.875 ;
        RECT 2851.685 1459.705 2851.855 1482.995 ;
        RECT 2849.845 1418.225 2850.475 1418.395 ;
        RECT 2849.845 1371.135 2850.015 1418.225 ;
        RECT 2849.845 1370.965 2850.475 1371.135 ;
        RECT 2850.305 1369.775 2850.475 1370.965 ;
        RECT 2849.385 1369.605 2850.475 1369.775 ;
        RECT 2849.385 1228.505 2849.555 1369.605 ;
        RECT 2849.845 1205.555 2850.015 1228.675 ;
        RECT 2849.845 1205.385 2850.935 1205.555 ;
        RECT 2850.765 1149.285 2850.935 1205.385 ;
        RECT 2850.765 899.045 2850.935 969.595 ;
        RECT 2849.845 672.605 2850.015 741.795 ;
        RECT 2850.305 268.685 2850.475 386.495 ;
        RECT 9.805 47.005 9.975 93.755 ;
        RECT 26.825 3.315 26.995 3.655 ;
        RECT 25.445 3.145 26.995 3.315 ;
        RECT 65.925 0.085 66.095 3.655 ;
        RECT 72.365 0.085 72.535 1.955 ;
        RECT 193.345 1.105 193.515 1.955 ;
      LAYER mcon ;
        RECT 2849.845 2760.205 2850.015 2760.375 ;
        RECT 2850.305 2655.485 2850.475 2655.655 ;
        RECT 2849.845 2612.985 2850.015 2613.155 ;
        RECT 2849.845 2525.605 2850.015 2525.775 ;
        RECT 2849.845 2342.685 2850.015 2342.855 ;
        RECT 2849.845 2306.985 2850.015 2307.155 ;
        RECT 2850.305 2208.045 2850.475 2208.215 ;
        RECT 2849.845 2090.065 2850.015 2090.235 ;
        RECT 2851.225 1883.345 2851.395 1883.515 ;
        RECT 2849.845 1788.145 2850.015 1788.315 ;
        RECT 2849.845 1724.225 2850.015 1724.395 ;
        RECT 2849.845 1710.965 2850.015 1711.135 ;
        RECT 2849.845 1655.205 2850.015 1655.375 ;
        RECT 2849.845 1603.525 2850.015 1603.695 ;
        RECT 2850.305 1500.505 2850.475 1500.675 ;
        RECT 2851.685 1482.825 2851.855 1482.995 ;
        RECT 2850.765 1459.705 2850.935 1459.875 ;
        RECT 2850.305 1448.825 2850.475 1448.995 ;
        RECT 2849.845 1228.505 2850.015 1228.675 ;
        RECT 2850.765 969.425 2850.935 969.595 ;
        RECT 2849.845 741.625 2850.015 741.795 ;
        RECT 2850.305 386.325 2850.475 386.495 ;
        RECT 9.805 93.585 9.975 93.755 ;
        RECT 26.825 3.485 26.995 3.655 ;
        RECT 65.925 3.485 66.095 3.655 ;
        RECT 72.365 1.785 72.535 1.955 ;
        RECT 193.345 1.785 193.515 1.955 ;
      LAYER met1 ;
        RECT 2873.690 2873.920 2874.010 2873.980 ;
        RECT 2901.290 2873.920 2901.610 2873.980 ;
        RECT 2873.690 2873.780 2901.610 2873.920 ;
        RECT 2873.690 2873.720 2874.010 2873.780 ;
        RECT 2901.290 2873.720 2901.610 2873.780 ;
        RECT 2849.770 2815.440 2850.090 2815.500 ;
        RECT 2873.690 2815.440 2874.010 2815.500 ;
        RECT 2849.770 2815.300 2874.010 2815.440 ;
        RECT 2849.770 2815.240 2850.090 2815.300 ;
        RECT 2873.690 2815.240 2874.010 2815.300 ;
        RECT 2849.770 2760.360 2850.090 2760.420 ;
        RECT 2849.575 2760.220 2850.090 2760.360 ;
        RECT 2849.770 2760.160 2850.090 2760.220 ;
        RECT 2849.770 2755.260 2850.090 2755.320 ;
        RECT 2849.575 2755.120 2850.090 2755.260 ;
        RECT 2849.770 2755.060 2850.090 2755.120 ;
        RECT 2849.770 2655.640 2850.090 2655.700 ;
        RECT 2850.245 2655.640 2850.535 2655.685 ;
        RECT 2849.770 2655.500 2850.535 2655.640 ;
        RECT 2849.770 2655.440 2850.090 2655.500 ;
        RECT 2850.245 2655.455 2850.535 2655.500 ;
        RECT 2849.770 2643.740 2850.090 2643.800 ;
        RECT 2850.245 2643.740 2850.535 2643.785 ;
        RECT 2849.770 2643.600 2850.535 2643.740 ;
        RECT 2849.770 2643.540 2850.090 2643.600 ;
        RECT 2850.245 2643.555 2850.535 2643.600 ;
        RECT 2849.770 2613.140 2850.090 2613.200 ;
        RECT 2849.575 2613.000 2850.090 2613.140 ;
        RECT 2849.770 2612.940 2850.090 2613.000 ;
        RECT 2849.770 2592.400 2850.090 2592.460 ;
        RECT 2849.575 2592.260 2850.090 2592.400 ;
        RECT 2849.770 2592.200 2850.090 2592.260 ;
        RECT 2849.770 2525.760 2850.090 2525.820 ;
        RECT 2849.575 2525.620 2850.090 2525.760 ;
        RECT 2849.770 2525.560 2850.090 2525.620 ;
        RECT 2849.770 2515.220 2850.090 2515.280 ;
        RECT 2849.575 2515.080 2850.090 2515.220 ;
        RECT 2849.770 2515.020 2850.090 2515.080 ;
        RECT 2849.770 2434.980 2850.090 2435.040 ;
        RECT 2850.690 2434.980 2851.010 2435.040 ;
        RECT 2849.770 2434.840 2851.010 2434.980 ;
        RECT 2849.770 2434.780 2850.090 2434.840 ;
        RECT 2850.690 2434.780 2851.010 2434.840 ;
        RECT 2849.770 2342.840 2850.090 2342.900 ;
        RECT 2849.575 2342.700 2850.090 2342.840 ;
        RECT 2849.770 2342.640 2850.090 2342.700 ;
        RECT 2849.770 2307.140 2850.090 2307.200 ;
        RECT 2849.575 2307.000 2850.090 2307.140 ;
        RECT 2849.770 2306.940 2850.090 2307.000 ;
        RECT 2849.770 2246.760 2850.090 2247.020 ;
        RECT 2849.860 2246.000 2850.000 2246.760 ;
        RECT 2849.770 2245.740 2850.090 2246.000 ;
        RECT 2849.770 2208.200 2850.090 2208.260 ;
        RECT 2850.245 2208.200 2850.535 2208.245 ;
        RECT 2849.770 2208.060 2850.535 2208.200 ;
        RECT 2849.770 2208.000 2850.090 2208.060 ;
        RECT 2850.245 2208.015 2850.535 2208.060 ;
        RECT 2850.230 2184.060 2850.550 2184.120 ;
        RECT 2850.035 2183.920 2850.550 2184.060 ;
        RECT 2850.230 2183.860 2850.550 2183.920 ;
        RECT 2849.770 2091.580 2850.090 2091.640 ;
        RECT 2849.770 2091.440 2850.460 2091.580 ;
        RECT 2849.770 2091.380 2850.090 2091.440 ;
        RECT 2849.785 2090.220 2850.075 2090.265 ;
        RECT 2850.320 2090.220 2850.460 2091.440 ;
        RECT 2849.785 2090.080 2850.460 2090.220 ;
        RECT 2849.785 2090.035 2850.075 2090.080 ;
        RECT 2849.770 2011.340 2850.090 2011.400 ;
        RECT 2849.575 2011.200 2850.090 2011.340 ;
        RECT 2849.770 2011.140 2850.090 2011.200 ;
        RECT 2850.690 1883.500 2851.010 1883.560 ;
        RECT 2851.165 1883.500 2851.455 1883.545 ;
        RECT 2850.690 1883.360 2851.455 1883.500 ;
        RECT 2850.690 1883.300 2851.010 1883.360 ;
        RECT 2851.165 1883.315 2851.455 1883.360 ;
        RECT 2849.785 1788.300 2850.075 1788.345 ;
        RECT 2851.165 1788.300 2851.455 1788.345 ;
        RECT 2849.785 1788.160 2851.455 1788.300 ;
        RECT 2849.785 1788.115 2850.075 1788.160 ;
        RECT 2851.165 1788.115 2851.455 1788.160 ;
        RECT 2849.770 1724.380 2850.090 1724.440 ;
        RECT 2849.575 1724.240 2850.090 1724.380 ;
        RECT 2849.770 1724.180 2850.090 1724.240 ;
        RECT 2849.770 1711.120 2850.090 1711.180 ;
        RECT 2849.770 1710.980 2850.285 1711.120 ;
        RECT 2849.770 1710.920 2850.090 1710.980 ;
        RECT 2849.770 1656.380 2850.090 1656.440 ;
        RECT 2849.575 1656.240 2850.090 1656.380 ;
        RECT 2849.770 1656.180 2850.090 1656.240 ;
        RECT 2849.770 1655.360 2850.090 1655.420 ;
        RECT 2849.575 1655.220 2850.090 1655.360 ;
        RECT 2849.770 1655.160 2850.090 1655.220 ;
        RECT 2849.785 1605.720 2850.075 1605.765 ;
        RECT 2849.400 1605.580 2850.075 1605.720 ;
        RECT 2849.400 1603.680 2849.540 1605.580 ;
        RECT 2849.785 1605.535 2850.075 1605.580 ;
        RECT 2849.785 1603.680 2850.075 1603.725 ;
        RECT 2849.400 1603.540 2850.075 1603.680 ;
        RECT 2849.785 1603.495 2850.075 1603.540 ;
        RECT 2849.770 1589.740 2850.090 1589.800 ;
        RECT 2849.575 1589.600 2850.090 1589.740 ;
        RECT 2849.770 1589.540 2850.090 1589.600 ;
        RECT 2850.245 1500.660 2850.535 1500.705 ;
        RECT 2850.690 1500.660 2851.010 1500.720 ;
        RECT 2850.245 1500.520 2851.010 1500.660 ;
        RECT 2850.245 1500.475 2850.535 1500.520 ;
        RECT 2850.690 1500.460 2851.010 1500.520 ;
        RECT 2850.245 1482.980 2850.535 1483.025 ;
        RECT 2851.625 1482.980 2851.915 1483.025 ;
        RECT 2850.245 1482.840 2851.915 1482.980 ;
        RECT 2850.245 1482.795 2850.535 1482.840 ;
        RECT 2851.625 1482.795 2851.915 1482.840 ;
        RECT 2850.705 1459.860 2850.995 1459.905 ;
        RECT 2851.625 1459.860 2851.915 1459.905 ;
        RECT 2850.705 1459.720 2851.915 1459.860 ;
        RECT 2850.705 1459.675 2850.995 1459.720 ;
        RECT 2851.625 1459.675 2851.915 1459.720 ;
        RECT 2850.245 1448.980 2850.535 1449.025 ;
        RECT 2850.705 1448.980 2850.995 1449.025 ;
        RECT 2850.245 1448.840 2850.995 1448.980 ;
        RECT 2850.245 1448.795 2850.535 1448.840 ;
        RECT 2850.705 1448.795 2850.995 1448.840 ;
        RECT 2849.325 1228.660 2849.615 1228.705 ;
        RECT 2849.785 1228.660 2850.075 1228.705 ;
        RECT 2849.325 1228.520 2850.075 1228.660 ;
        RECT 2849.325 1228.475 2849.615 1228.520 ;
        RECT 2849.785 1228.475 2850.075 1228.520 ;
        RECT 2850.705 1149.440 2850.995 1149.485 ;
        RECT 2852.070 1149.440 2852.390 1149.500 ;
        RECT 2850.705 1149.300 2852.390 1149.440 ;
        RECT 2850.705 1149.255 2850.995 1149.300 ;
        RECT 2852.070 1149.240 2852.390 1149.300 ;
        RECT 2850.690 1042.000 2851.010 1042.060 ;
        RECT 2852.070 1042.000 2852.390 1042.060 ;
        RECT 2850.690 1041.860 2852.390 1042.000 ;
        RECT 2850.690 1041.800 2851.010 1041.860 ;
        RECT 2852.070 1041.800 2852.390 1041.860 ;
        RECT 2849.770 969.580 2850.090 969.640 ;
        RECT 2850.705 969.580 2850.995 969.625 ;
        RECT 2849.770 969.440 2850.995 969.580 ;
        RECT 2849.770 969.380 2850.090 969.440 ;
        RECT 2850.705 969.395 2850.995 969.440 ;
        RECT 2849.770 899.200 2850.090 899.260 ;
        RECT 2850.705 899.200 2850.995 899.245 ;
        RECT 2849.770 899.060 2850.995 899.200 ;
        RECT 2849.770 899.000 2850.090 899.060 ;
        RECT 2850.705 899.015 2850.995 899.060 ;
        RECT 2849.770 888.660 2850.090 888.720 ;
        RECT 2851.610 888.660 2851.930 888.720 ;
        RECT 2849.770 888.520 2851.930 888.660 ;
        RECT 2849.770 888.460 2850.090 888.520 ;
        RECT 2851.610 888.460 2851.930 888.520 ;
        RECT 2850.230 747.220 2850.550 747.280 ;
        RECT 2851.610 747.220 2851.930 747.280 ;
        RECT 2850.230 747.080 2851.930 747.220 ;
        RECT 2850.230 747.020 2850.550 747.080 ;
        RECT 2851.610 747.020 2851.930 747.080 ;
        RECT 2849.785 741.780 2850.075 741.825 ;
        RECT 2850.230 741.780 2850.550 741.840 ;
        RECT 2849.785 741.640 2850.550 741.780 ;
        RECT 2849.785 741.595 2850.075 741.640 ;
        RECT 2850.230 741.580 2850.550 741.640 ;
        RECT 2849.785 672.760 2850.075 672.805 ;
        RECT 2850.230 672.760 2850.550 672.820 ;
        RECT 2849.785 672.620 2850.550 672.760 ;
        RECT 2849.785 672.575 2850.075 672.620 ;
        RECT 2850.230 672.560 2850.550 672.620 ;
        RECT 2849.770 386.480 2850.090 386.540 ;
        RECT 2850.245 386.480 2850.535 386.525 ;
        RECT 2849.770 386.340 2850.535 386.480 ;
        RECT 2849.770 386.280 2850.090 386.340 ;
        RECT 2850.245 386.295 2850.535 386.340 ;
        RECT 2849.770 268.840 2850.090 268.900 ;
        RECT 2850.245 268.840 2850.535 268.885 ;
        RECT 2849.770 268.700 2850.535 268.840 ;
        RECT 2849.770 268.640 2850.090 268.700 ;
        RECT 2850.245 268.655 2850.535 268.700 ;
        RECT 2849.770 227.700 2850.090 227.760 ;
        RECT 2851.610 227.700 2851.930 227.760 ;
        RECT 2849.770 227.560 2851.930 227.700 ;
        RECT 2849.770 227.500 2850.090 227.560 ;
        RECT 2851.610 227.500 2851.930 227.560 ;
        RECT 6.970 93.740 7.290 93.800 ;
        RECT 9.745 93.740 10.035 93.785 ;
        RECT 6.970 93.600 10.035 93.740 ;
        RECT 6.970 93.540 7.290 93.600 ;
        RECT 9.745 93.555 10.035 93.600 ;
        RECT 6.510 47.160 6.830 47.220 ;
        RECT 9.745 47.160 10.035 47.205 ;
        RECT 6.510 47.020 10.035 47.160 ;
        RECT 6.510 46.960 6.830 47.020 ;
        RECT 9.745 46.975 10.035 47.020 ;
        RECT 26.765 3.640 27.055 3.685 ;
        RECT 65.865 3.640 66.155 3.685 ;
        RECT 26.765 3.500 66.155 3.640 ;
        RECT 26.765 3.455 27.055 3.500 ;
        RECT 65.865 3.455 66.155 3.500 ;
        RECT 6.510 3.300 6.830 3.360 ;
        RECT 25.385 3.300 25.675 3.345 ;
        RECT 6.510 3.160 25.675 3.300 ;
        RECT 6.510 3.100 6.830 3.160 ;
        RECT 25.385 3.115 25.675 3.160 ;
        RECT 72.305 1.940 72.595 1.985 ;
        RECT 193.285 1.940 193.575 1.985 ;
        RECT 72.305 1.800 193.575 1.940 ;
        RECT 72.305 1.755 72.595 1.800 ;
        RECT 193.285 1.755 193.575 1.800 ;
        RECT 193.285 1.260 193.575 1.305 ;
        RECT 265.950 1.260 266.270 1.320 ;
        RECT 193.285 1.120 266.270 1.260 ;
        RECT 193.285 1.075 193.575 1.120 ;
        RECT 265.950 1.060 266.270 1.120 ;
        RECT 65.865 0.240 66.155 0.285 ;
        RECT 72.305 0.240 72.595 0.285 ;
        RECT 65.865 0.100 72.595 0.240 ;
        RECT 65.865 0.055 66.155 0.100 ;
        RECT 72.305 0.055 72.595 0.100 ;
      LAYER via ;
        RECT 2873.720 2873.720 2873.980 2873.980 ;
        RECT 2901.320 2873.720 2901.580 2873.980 ;
        RECT 2849.800 2815.240 2850.060 2815.500 ;
        RECT 2873.720 2815.240 2873.980 2815.500 ;
        RECT 2849.800 2760.160 2850.060 2760.420 ;
        RECT 2849.800 2755.060 2850.060 2755.320 ;
        RECT 2849.800 2655.440 2850.060 2655.700 ;
        RECT 2849.800 2643.540 2850.060 2643.800 ;
        RECT 2849.800 2612.940 2850.060 2613.200 ;
        RECT 2849.800 2592.200 2850.060 2592.460 ;
        RECT 2849.800 2525.560 2850.060 2525.820 ;
        RECT 2849.800 2515.020 2850.060 2515.280 ;
        RECT 2849.800 2434.780 2850.060 2435.040 ;
        RECT 2850.720 2434.780 2850.980 2435.040 ;
        RECT 2849.800 2342.640 2850.060 2342.900 ;
        RECT 2849.800 2306.940 2850.060 2307.200 ;
        RECT 2849.800 2246.760 2850.060 2247.020 ;
        RECT 2849.800 2245.740 2850.060 2246.000 ;
        RECT 2849.800 2208.000 2850.060 2208.260 ;
        RECT 2850.260 2183.860 2850.520 2184.120 ;
        RECT 2849.800 2091.380 2850.060 2091.640 ;
        RECT 2849.800 2011.140 2850.060 2011.400 ;
        RECT 2850.720 1883.300 2850.980 1883.560 ;
        RECT 2849.800 1724.180 2850.060 1724.440 ;
        RECT 2849.800 1710.920 2850.060 1711.180 ;
        RECT 2849.800 1656.180 2850.060 1656.440 ;
        RECT 2849.800 1655.160 2850.060 1655.420 ;
        RECT 2849.800 1589.540 2850.060 1589.800 ;
        RECT 2850.720 1500.460 2850.980 1500.720 ;
        RECT 2852.100 1149.240 2852.360 1149.500 ;
        RECT 2850.720 1041.800 2850.980 1042.060 ;
        RECT 2852.100 1041.800 2852.360 1042.060 ;
        RECT 2849.800 969.380 2850.060 969.640 ;
        RECT 2849.800 899.000 2850.060 899.260 ;
        RECT 2849.800 888.460 2850.060 888.720 ;
        RECT 2851.640 888.460 2851.900 888.720 ;
        RECT 2850.260 747.020 2850.520 747.280 ;
        RECT 2851.640 747.020 2851.900 747.280 ;
        RECT 2850.260 741.580 2850.520 741.840 ;
        RECT 2850.260 672.560 2850.520 672.820 ;
        RECT 2849.800 386.280 2850.060 386.540 ;
        RECT 2849.800 268.640 2850.060 268.900 ;
        RECT 2849.800 227.500 2850.060 227.760 ;
        RECT 2851.640 227.500 2851.900 227.760 ;
        RECT 7.000 93.540 7.260 93.800 ;
        RECT 6.540 46.960 6.800 47.220 ;
        RECT 6.540 3.100 6.800 3.360 ;
        RECT 265.980 1.060 266.240 1.320 ;
      LAYER met2 ;
        RECT 2901.310 2903.755 2901.590 2904.125 ;
        RECT 2901.380 2874.010 2901.520 2903.755 ;
        RECT 2873.720 2873.690 2873.980 2874.010 ;
        RECT 2901.320 2873.690 2901.580 2874.010 ;
        RECT 2873.780 2815.530 2873.920 2873.690 ;
        RECT 2849.800 2815.210 2850.060 2815.530 ;
        RECT 2873.720 2815.210 2873.980 2815.530 ;
        RECT 2849.860 2814.930 2850.000 2815.210 ;
        RECT 2849.400 2814.790 2850.000 2814.930 ;
        RECT 2849.400 2760.530 2849.540 2814.790 ;
        RECT 2849.400 2760.450 2850.000 2760.530 ;
        RECT 2849.400 2760.390 2850.060 2760.450 ;
        RECT 2849.800 2760.130 2850.060 2760.390 ;
        RECT 2849.800 2755.090 2850.060 2755.350 ;
        RECT 2849.400 2755.030 2850.060 2755.090 ;
        RECT 2849.400 2754.950 2850.000 2755.030 ;
        RECT 2849.400 2666.690 2849.540 2754.950 ;
        RECT 2849.400 2666.550 2850.000 2666.690 ;
        RECT 2849.860 2655.730 2850.000 2666.550 ;
        RECT 2849.800 2655.410 2850.060 2655.730 ;
        RECT 2849.800 2643.570 2850.060 2643.830 ;
        RECT 2849.400 2643.510 2850.060 2643.570 ;
        RECT 2849.400 2643.430 2850.000 2643.510 ;
        RECT 2849.400 2635.410 2849.540 2643.430 ;
        RECT 2849.400 2635.270 2850.000 2635.410 ;
        RECT 2849.860 2613.230 2850.000 2635.270 ;
        RECT 2849.800 2612.910 2850.060 2613.230 ;
        RECT 2849.800 2592.170 2850.060 2592.490 ;
        RECT 2849.860 2587.130 2850.000 2592.170 ;
        RECT 2849.400 2586.990 2850.000 2587.130 ;
        RECT 2849.400 2538.850 2849.540 2586.990 ;
        RECT 2849.400 2538.710 2850.000 2538.850 ;
        RECT 2849.860 2525.850 2850.000 2538.710 ;
        RECT 2849.800 2525.530 2850.060 2525.850 ;
        RECT 2849.800 2515.050 2850.060 2515.310 ;
        RECT 2849.400 2514.990 2850.060 2515.050 ;
        RECT 2849.400 2514.910 2850.000 2514.990 ;
        RECT 2849.400 2456.570 2849.540 2514.910 ;
        RECT 2849.400 2456.430 2850.920 2456.570 ;
        RECT 2850.780 2435.070 2850.920 2456.430 ;
        RECT 2849.800 2434.810 2850.060 2435.070 ;
        RECT 2848.940 2434.750 2850.060 2434.810 ;
        RECT 2850.720 2434.750 2850.980 2435.070 ;
        RECT 2848.940 2434.670 2850.000 2434.750 ;
        RECT 2848.940 2343.010 2849.080 2434.670 ;
        RECT 2848.940 2342.930 2850.000 2343.010 ;
        RECT 2848.940 2342.870 2850.060 2342.930 ;
        RECT 2849.800 2342.610 2850.060 2342.870 ;
        RECT 2849.800 2306.910 2850.060 2307.230 ;
        RECT 2849.860 2247.050 2850.000 2306.910 ;
        RECT 2849.800 2246.730 2850.060 2247.050 ;
        RECT 2849.800 2245.710 2850.060 2246.030 ;
        RECT 2849.860 2239.650 2850.000 2245.710 ;
        RECT 2849.400 2239.510 2850.000 2239.650 ;
        RECT 2849.400 2208.370 2849.540 2239.510 ;
        RECT 2849.400 2208.290 2850.000 2208.370 ;
        RECT 2849.400 2208.230 2850.060 2208.290 ;
        RECT 2849.800 2207.970 2850.060 2208.230 ;
        RECT 2850.260 2183.830 2850.520 2184.150 ;
        RECT 2850.320 2143.770 2850.460 2183.830 ;
        RECT 2849.400 2143.630 2850.460 2143.770 ;
        RECT 2849.400 2142.410 2849.540 2143.630 ;
        RECT 2848.940 2142.270 2849.540 2142.410 ;
        RECT 2848.940 2092.090 2849.080 2142.270 ;
        RECT 2848.940 2091.950 2850.000 2092.090 ;
        RECT 2849.860 2091.670 2850.000 2091.950 ;
        RECT 2849.800 2091.350 2850.060 2091.670 ;
        RECT 2849.800 2011.170 2850.060 2011.430 ;
        RECT 2849.400 2011.110 2850.060 2011.170 ;
        RECT 2849.400 2011.030 2850.000 2011.110 ;
        RECT 2849.400 1983.290 2849.540 2011.030 ;
        RECT 2849.400 1983.150 2850.460 1983.290 ;
        RECT 2850.320 1982.440 2850.460 1983.150 ;
        RECT 2850.320 1982.300 2850.920 1982.440 ;
        RECT 2850.780 1883.590 2850.920 1982.300 ;
        RECT 2850.720 1883.270 2850.980 1883.590 ;
        RECT 2849.800 1724.150 2850.060 1724.470 ;
        RECT 2849.860 1711.210 2850.000 1724.150 ;
        RECT 2849.800 1710.890 2850.060 1711.210 ;
        RECT 2849.800 1656.210 2850.060 1656.470 ;
        RECT 2849.400 1656.150 2850.060 1656.210 ;
        RECT 2849.400 1656.070 2850.000 1656.150 ;
        RECT 2849.400 1655.530 2849.540 1656.070 ;
        RECT 2849.400 1655.450 2850.000 1655.530 ;
        RECT 2849.400 1655.390 2850.060 1655.450 ;
        RECT 2849.800 1655.130 2850.060 1655.390 ;
        RECT 2849.800 1589.570 2850.060 1589.830 ;
        RECT 2849.400 1589.510 2850.060 1589.570 ;
        RECT 2849.400 1589.430 2850.000 1589.510 ;
        RECT 2849.400 1578.860 2849.540 1589.430 ;
        RECT 2849.400 1578.720 2850.000 1578.860 ;
        RECT 2849.860 1578.690 2850.000 1578.720 ;
        RECT 2849.860 1578.550 2850.920 1578.690 ;
        RECT 2850.780 1500.750 2850.920 1578.550 ;
        RECT 2850.720 1500.430 2850.980 1500.750 ;
        RECT 2852.100 1149.210 2852.360 1149.530 ;
        RECT 2852.160 1042.090 2852.300 1149.210 ;
        RECT 2850.720 1041.770 2850.980 1042.090 ;
        RECT 2852.100 1041.770 2852.360 1042.090 ;
        RECT 2850.780 993.890 2850.920 1041.770 ;
        RECT 2849.400 993.750 2850.920 993.890 ;
        RECT 2849.400 983.010 2849.540 993.750 ;
        RECT 2849.400 982.870 2850.000 983.010 ;
        RECT 2849.860 969.670 2850.000 982.870 ;
        RECT 2849.800 969.350 2850.060 969.670 ;
        RECT 2849.800 898.970 2850.060 899.290 ;
        RECT 2849.860 888.750 2850.000 898.970 ;
        RECT 2849.800 888.430 2850.060 888.750 ;
        RECT 2851.640 888.430 2851.900 888.750 ;
        RECT 2851.700 747.310 2851.840 888.430 ;
        RECT 2850.260 746.990 2850.520 747.310 ;
        RECT 2851.640 746.990 2851.900 747.310 ;
        RECT 2850.320 741.870 2850.460 746.990 ;
        RECT 2850.260 741.550 2850.520 741.870 ;
        RECT 2850.260 672.530 2850.520 672.850 ;
        RECT 2850.320 521.290 2850.460 672.530 ;
        RECT 2849.400 521.150 2850.460 521.290 ;
        RECT 2849.400 386.480 2849.540 521.150 ;
        RECT 2849.800 386.480 2850.060 386.570 ;
        RECT 2849.400 386.340 2850.060 386.480 ;
        RECT 2849.800 386.250 2850.060 386.340 ;
        RECT 2849.400 268.930 2850.000 269.010 ;
        RECT 2849.400 268.870 2850.060 268.930 ;
        RECT 2849.400 227.700 2849.540 268.870 ;
        RECT 2849.800 268.610 2850.060 268.870 ;
        RECT 2849.800 227.700 2850.060 227.790 ;
        RECT 2849.400 227.560 2850.060 227.700 ;
        RECT 2849.800 227.470 2850.060 227.560 ;
        RECT 2851.640 227.470 2851.900 227.790 ;
        RECT 2851.700 174.605 2851.840 227.470 ;
        RECT 2851.630 174.235 2851.910 174.605 ;
        RECT 6.990 98.755 7.270 99.125 ;
        RECT 7.060 93.830 7.200 98.755 ;
        RECT 7.000 93.510 7.260 93.830 ;
        RECT 6.540 46.930 6.800 47.250 ;
        RECT 6.600 3.390 6.740 46.930 ;
        RECT 265.910 5.000 266.190 9.000 ;
        RECT 6.540 3.070 6.800 3.390 ;
        RECT 266.040 1.350 266.180 5.000 ;
        RECT 265.980 1.030 266.240 1.350 ;
      LAYER via2 ;
        RECT 2901.310 2903.800 2901.590 2904.080 ;
        RECT 2851.630 174.280 2851.910 174.560 ;
        RECT 6.990 98.800 7.270 99.080 ;
      LAYER met3 ;
        RECT 2901.285 2904.090 2901.615 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2901.285 2903.790 2924.800 2904.090 ;
        RECT 2901.285 2903.775 2901.615 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
        RECT 2851.605 174.580 2851.935 174.585 ;
        RECT 2851.350 174.570 2851.935 174.580 ;
        RECT 2851.350 174.270 2852.160 174.570 ;
        RECT 2851.350 174.260 2851.935 174.270 ;
        RECT 2851.605 174.255 2851.935 174.260 ;
        RECT 5.790 99.090 6.170 99.100 ;
        RECT 6.965 99.090 7.295 99.105 ;
        RECT 5.790 98.790 7.295 99.090 ;
        RECT 5.790 98.780 6.170 98.790 ;
        RECT 6.965 98.775 7.295 98.790 ;
      LAYER via3 ;
        RECT 2851.380 174.260 2851.700 174.580 ;
        RECT 5.820 98.780 6.140 99.100 ;
      LAYER met4 ;
        RECT 2851.375 174.255 2851.705 174.585 ;
        RECT 2851.390 162.090 2851.690 174.255 ;
        RECT 2810.470 160.910 2811.650 162.090 ;
        RECT 2850.950 160.910 2852.130 162.090 ;
        RECT 2810.910 128.090 2811.210 160.910 ;
        RECT 5.390 126.910 6.570 128.090 ;
        RECT 2810.470 126.910 2811.650 128.090 ;
        RECT 5.830 99.105 6.130 126.910 ;
        RECT 5.815 98.775 6.145 99.105 ;
      LAYER met5 ;
        RECT 2810.260 160.700 2852.340 162.300 ;
        RECT 5.180 126.700 2811.860 128.300 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 8.885 2998.545 9.055 3009.935 ;
        RECT 8.885 2815.625 9.055 2827.695 ;
        RECT 8.885 2612.305 9.055 2635.935 ;
        RECT 7.965 2508.945 8.135 2536.655 ;
        RECT 8.885 2238.985 9.055 2250.375 ;
        RECT 8.425 1894.905 8.595 1903.575 ;
        RECT 9.345 1790.525 9.515 1851.895 ;
        RECT 8.425 1648.745 8.595 1728.815 ;
        RECT 7.965 1558.305 8.135 1594.855 ;
        RECT 9.345 1481.125 9.515 1526.855 ;
        RECT 4.745 773.925 4.915 838.355 ;
        RECT 8.425 673.115 8.595 743.155 ;
        RECT 8.425 672.945 9.055 673.115 ;
        RECT 8.885 671.925 9.055 672.945 ;
        RECT 55.805 6.205 55.975 8.075 ;
      LAYER mcon ;
        RECT 8.885 3009.765 9.055 3009.935 ;
        RECT 8.885 2827.525 9.055 2827.695 ;
        RECT 8.885 2635.765 9.055 2635.935 ;
        RECT 7.965 2536.485 8.135 2536.655 ;
        RECT 8.885 2250.205 9.055 2250.375 ;
        RECT 8.425 1903.405 8.595 1903.575 ;
        RECT 9.345 1851.725 9.515 1851.895 ;
        RECT 8.425 1728.645 8.595 1728.815 ;
        RECT 7.965 1594.685 8.135 1594.855 ;
        RECT 9.345 1526.685 9.515 1526.855 ;
        RECT 4.745 838.185 4.915 838.355 ;
        RECT 8.425 742.985 8.595 743.155 ;
        RECT 55.805 7.905 55.975 8.075 ;
      LAYER met1 ;
        RECT 11.110 3395.480 11.430 3395.540 ;
        RECT 2846.090 3395.480 2846.410 3395.540 ;
        RECT 11.110 3395.340 2846.410 3395.480 ;
        RECT 11.110 3395.280 11.430 3395.340 ;
        RECT 2846.090 3395.280 2846.410 3395.340 ;
        RECT 2849.770 3271.040 2850.090 3271.100 ;
        RECT 2887.490 3271.040 2887.810 3271.100 ;
        RECT 2849.770 3270.900 2887.810 3271.040 ;
        RECT 2849.770 3270.840 2850.090 3270.900 ;
        RECT 2887.490 3270.840 2887.810 3270.900 ;
        RECT 9.730 3208.960 10.050 3209.220 ;
        RECT 9.820 3208.200 9.960 3208.960 ;
        RECT 9.730 3207.940 10.050 3208.200 ;
        RECT 2887.490 3139.460 2887.810 3139.520 ;
        RECT 2898.530 3139.460 2898.850 3139.520 ;
        RECT 2887.490 3139.320 2898.850 3139.460 ;
        RECT 2887.490 3139.260 2887.810 3139.320 ;
        RECT 2898.530 3139.260 2898.850 3139.320 ;
        RECT 8.825 3009.920 9.115 3009.965 ;
        RECT 9.730 3009.920 10.050 3009.980 ;
        RECT 8.825 3009.780 10.050 3009.920 ;
        RECT 8.825 3009.735 9.115 3009.780 ;
        RECT 9.730 3009.720 10.050 3009.780 ;
        RECT 8.825 2998.700 9.115 2998.745 ;
        RECT 9.730 2998.700 10.050 2998.760 ;
        RECT 8.825 2998.560 10.050 2998.700 ;
        RECT 8.825 2998.515 9.115 2998.560 ;
        RECT 9.730 2998.500 10.050 2998.560 ;
        RECT 8.825 2827.680 9.115 2827.725 ;
        RECT 9.730 2827.680 10.050 2827.740 ;
        RECT 8.825 2827.540 10.050 2827.680 ;
        RECT 8.825 2827.495 9.115 2827.540 ;
        RECT 9.730 2827.480 10.050 2827.540 ;
        RECT 8.825 2815.780 9.115 2815.825 ;
        RECT 9.730 2815.780 10.050 2815.840 ;
        RECT 8.825 2815.640 10.050 2815.780 ;
        RECT 8.825 2815.595 9.115 2815.640 ;
        RECT 9.730 2815.580 10.050 2815.640 ;
        RECT 8.825 2635.920 9.115 2635.965 ;
        RECT 9.730 2635.920 10.050 2635.980 ;
        RECT 8.825 2635.780 10.050 2635.920 ;
        RECT 8.825 2635.735 9.115 2635.780 ;
        RECT 9.730 2635.720 10.050 2635.780 ;
        RECT 8.825 2612.460 9.115 2612.505 ;
        RECT 9.730 2612.460 10.050 2612.520 ;
        RECT 8.825 2612.320 10.050 2612.460 ;
        RECT 8.825 2612.275 9.115 2612.320 ;
        RECT 9.730 2612.260 10.050 2612.320 ;
        RECT 7.905 2536.640 8.195 2536.685 ;
        RECT 9.730 2536.640 10.050 2536.700 ;
        RECT 7.905 2536.500 10.050 2536.640 ;
        RECT 7.905 2536.455 8.195 2536.500 ;
        RECT 9.730 2536.440 10.050 2536.500 ;
        RECT 7.905 2509.100 8.195 2509.145 ;
        RECT 9.730 2509.100 10.050 2509.160 ;
        RECT 7.905 2508.960 10.050 2509.100 ;
        RECT 7.905 2508.915 8.195 2508.960 ;
        RECT 9.730 2508.900 10.050 2508.960 ;
        RECT 8.350 2363.920 8.670 2363.980 ;
        RECT 9.730 2363.920 10.050 2363.980 ;
        RECT 8.350 2363.780 10.050 2363.920 ;
        RECT 8.350 2363.720 8.670 2363.780 ;
        RECT 9.730 2363.720 10.050 2363.780 ;
        RECT 8.825 2250.360 9.115 2250.405 ;
        RECT 9.730 2250.360 10.050 2250.420 ;
        RECT 8.825 2250.220 10.050 2250.360 ;
        RECT 8.825 2250.175 9.115 2250.220 ;
        RECT 9.730 2250.160 10.050 2250.220 ;
        RECT 8.825 2239.140 9.115 2239.185 ;
        RECT 9.730 2239.140 10.050 2239.200 ;
        RECT 8.825 2239.000 10.050 2239.140 ;
        RECT 8.825 2238.955 9.115 2239.000 ;
        RECT 9.730 2238.940 10.050 2239.000 ;
        RECT 8.810 1934.840 9.130 1934.900 ;
        RECT 9.730 1934.840 10.050 1934.900 ;
        RECT 8.810 1934.700 10.050 1934.840 ;
        RECT 8.810 1934.640 9.130 1934.700 ;
        RECT 9.730 1934.640 10.050 1934.700 ;
        RECT 8.365 1903.560 8.655 1903.605 ;
        RECT 8.810 1903.560 9.130 1903.620 ;
        RECT 8.365 1903.420 9.130 1903.560 ;
        RECT 8.365 1903.375 8.655 1903.420 ;
        RECT 8.810 1903.360 9.130 1903.420 ;
        RECT 8.365 1895.060 8.655 1895.105 ;
        RECT 9.730 1895.060 10.050 1895.120 ;
        RECT 8.365 1894.920 10.050 1895.060 ;
        RECT 8.365 1894.875 8.655 1894.920 ;
        RECT 9.730 1894.860 10.050 1894.920 ;
        RECT 9.285 1851.880 9.575 1851.925 ;
        RECT 9.730 1851.880 10.050 1851.940 ;
        RECT 9.285 1851.740 10.050 1851.880 ;
        RECT 9.285 1851.695 9.575 1851.740 ;
        RECT 9.730 1851.680 10.050 1851.740 ;
        RECT 9.270 1790.680 9.590 1790.740 ;
        RECT 9.075 1790.540 9.590 1790.680 ;
        RECT 9.270 1790.480 9.590 1790.540 ;
        RECT 8.365 1728.800 8.655 1728.845 ;
        RECT 9.730 1728.800 10.050 1728.860 ;
        RECT 8.365 1728.660 10.050 1728.800 ;
        RECT 8.365 1728.615 8.655 1728.660 ;
        RECT 9.730 1728.600 10.050 1728.660 ;
        RECT 8.365 1648.900 8.655 1648.945 ;
        RECT 9.730 1648.900 10.050 1648.960 ;
        RECT 8.365 1648.760 10.050 1648.900 ;
        RECT 8.365 1648.715 8.655 1648.760 ;
        RECT 9.730 1648.700 10.050 1648.760 ;
        RECT 7.905 1594.840 8.195 1594.885 ;
        RECT 9.730 1594.840 10.050 1594.900 ;
        RECT 7.905 1594.700 10.050 1594.840 ;
        RECT 7.905 1594.655 8.195 1594.700 ;
        RECT 9.730 1594.640 10.050 1594.700 ;
        RECT 7.905 1558.460 8.195 1558.505 ;
        RECT 9.730 1558.460 10.050 1558.520 ;
        RECT 7.905 1558.320 10.050 1558.460 ;
        RECT 7.905 1558.275 8.195 1558.320 ;
        RECT 9.730 1558.260 10.050 1558.320 ;
        RECT 9.285 1526.840 9.575 1526.885 ;
        RECT 9.730 1526.840 10.050 1526.900 ;
        RECT 9.285 1526.700 10.050 1526.840 ;
        RECT 9.285 1526.655 9.575 1526.700 ;
        RECT 9.730 1526.640 10.050 1526.700 ;
        RECT 6.510 1481.280 6.830 1481.340 ;
        RECT 9.285 1481.280 9.575 1481.325 ;
        RECT 6.510 1481.140 9.575 1481.280 ;
        RECT 6.510 1481.080 6.830 1481.140 ;
        RECT 9.285 1481.095 9.575 1481.140 ;
        RECT 6.510 1320.120 6.830 1320.180 ;
        RECT 9.730 1320.120 10.050 1320.180 ;
        RECT 6.510 1319.980 10.050 1320.120 ;
        RECT 6.510 1319.920 6.830 1319.980 ;
        RECT 9.730 1319.920 10.050 1319.980 ;
        RECT 2.370 1177.320 2.690 1177.380 ;
        RECT 8.810 1177.320 9.130 1177.380 ;
        RECT 2.370 1177.180 9.130 1177.320 ;
        RECT 2.370 1177.120 2.690 1177.180 ;
        RECT 8.810 1177.120 9.130 1177.180 ;
        RECT 1.910 838.340 2.230 838.400 ;
        RECT 4.685 838.340 4.975 838.385 ;
        RECT 1.910 838.200 4.975 838.340 ;
        RECT 1.910 838.140 2.230 838.200 ;
        RECT 4.685 838.155 4.975 838.200 ;
        RECT 4.685 774.080 4.975 774.125 ;
        RECT 6.970 774.080 7.290 774.140 ;
        RECT 4.685 773.940 7.290 774.080 ;
        RECT 4.685 773.895 4.975 773.940 ;
        RECT 6.970 773.880 7.290 773.940 ;
        RECT 6.970 743.140 7.290 743.200 ;
        RECT 8.365 743.140 8.655 743.185 ;
        RECT 6.970 743.000 8.655 743.140 ;
        RECT 6.970 742.940 7.290 743.000 ;
        RECT 8.365 742.955 8.655 743.000 ;
        RECT 4.670 672.080 4.990 672.140 ;
        RECT 8.825 672.080 9.115 672.125 ;
        RECT 4.670 671.940 9.115 672.080 ;
        RECT 4.670 671.880 4.990 671.940 ;
        RECT 8.825 671.895 9.115 671.940 ;
        RECT 3.750 606.120 4.070 606.180 ;
        RECT 4.670 606.120 4.990 606.180 ;
        RECT 3.750 605.980 4.990 606.120 ;
        RECT 3.750 605.920 4.070 605.980 ;
        RECT 4.670 605.920 4.990 605.980 ;
        RECT 52.050 8.060 52.370 8.120 ;
        RECT 55.745 8.060 56.035 8.105 ;
        RECT 52.050 7.920 56.035 8.060 ;
        RECT 52.050 7.860 52.370 7.920 ;
        RECT 55.745 7.875 56.035 7.920 ;
        RECT 282.970 7.720 283.290 7.780 ;
        RECT 244.880 7.580 283.290 7.720 ;
        RECT 244.880 7.440 245.020 7.580 ;
        RECT 282.970 7.520 283.290 7.580 ;
        RECT 244.790 7.180 245.110 7.440 ;
        RECT 55.745 6.360 56.035 6.405 ;
        RECT 139.450 6.360 139.770 6.420 ;
        RECT 55.745 6.220 139.770 6.360 ;
        RECT 55.745 6.175 56.035 6.220 ;
        RECT 139.450 6.160 139.770 6.220 ;
      LAYER via ;
        RECT 11.140 3395.280 11.400 3395.540 ;
        RECT 2846.120 3395.280 2846.380 3395.540 ;
        RECT 2849.800 3270.840 2850.060 3271.100 ;
        RECT 2887.520 3270.840 2887.780 3271.100 ;
        RECT 9.760 3208.960 10.020 3209.220 ;
        RECT 9.760 3207.940 10.020 3208.200 ;
        RECT 2887.520 3139.260 2887.780 3139.520 ;
        RECT 2898.560 3139.260 2898.820 3139.520 ;
        RECT 9.760 3009.720 10.020 3009.980 ;
        RECT 9.760 2998.500 10.020 2998.760 ;
        RECT 9.760 2827.480 10.020 2827.740 ;
        RECT 9.760 2815.580 10.020 2815.840 ;
        RECT 9.760 2635.720 10.020 2635.980 ;
        RECT 9.760 2612.260 10.020 2612.520 ;
        RECT 9.760 2536.440 10.020 2536.700 ;
        RECT 9.760 2508.900 10.020 2509.160 ;
        RECT 8.380 2363.720 8.640 2363.980 ;
        RECT 9.760 2363.720 10.020 2363.980 ;
        RECT 9.760 2250.160 10.020 2250.420 ;
        RECT 9.760 2238.940 10.020 2239.200 ;
        RECT 8.840 1934.640 9.100 1934.900 ;
        RECT 9.760 1934.640 10.020 1934.900 ;
        RECT 8.840 1903.360 9.100 1903.620 ;
        RECT 9.760 1894.860 10.020 1895.120 ;
        RECT 9.760 1851.680 10.020 1851.940 ;
        RECT 9.300 1790.480 9.560 1790.740 ;
        RECT 9.760 1728.600 10.020 1728.860 ;
        RECT 9.760 1648.700 10.020 1648.960 ;
        RECT 9.760 1594.640 10.020 1594.900 ;
        RECT 9.760 1558.260 10.020 1558.520 ;
        RECT 9.760 1526.640 10.020 1526.900 ;
        RECT 6.540 1481.080 6.800 1481.340 ;
        RECT 6.540 1319.920 6.800 1320.180 ;
        RECT 9.760 1319.920 10.020 1320.180 ;
        RECT 2.400 1177.120 2.660 1177.380 ;
        RECT 8.840 1177.120 9.100 1177.380 ;
        RECT 1.940 838.140 2.200 838.400 ;
        RECT 7.000 773.880 7.260 774.140 ;
        RECT 7.000 742.940 7.260 743.200 ;
        RECT 4.700 671.880 4.960 672.140 ;
        RECT 3.780 605.920 4.040 606.180 ;
        RECT 4.700 605.920 4.960 606.180 ;
        RECT 52.080 7.860 52.340 8.120 ;
        RECT 283.000 7.520 283.260 7.780 ;
        RECT 244.820 7.180 245.080 7.440 ;
        RECT 139.480 6.160 139.740 6.420 ;
      LAYER met2 ;
        RECT 11.140 3395.250 11.400 3395.570 ;
        RECT 2846.120 3395.250 2846.380 3395.570 ;
        RECT 11.200 3234.490 11.340 3395.250 ;
        RECT 2846.180 3295.690 2846.320 3395.250 ;
        RECT 2846.180 3295.550 2850.000 3295.690 ;
        RECT 2849.860 3271.130 2850.000 3295.550 ;
        RECT 2849.800 3270.810 2850.060 3271.130 ;
        RECT 2887.520 3270.810 2887.780 3271.130 ;
        RECT 10.280 3234.350 11.340 3234.490 ;
        RECT 10.280 3209.330 10.420 3234.350 ;
        RECT 9.820 3209.250 10.420 3209.330 ;
        RECT 9.760 3209.190 10.420 3209.250 ;
        RECT 9.760 3208.930 10.020 3209.190 ;
        RECT 9.760 3207.910 10.020 3208.230 ;
        RECT 9.820 3205.930 9.960 3207.910 ;
        RECT 9.820 3205.790 11.800 3205.930 ;
        RECT 11.660 3164.450 11.800 3205.790 ;
        RECT 11.660 3164.310 13.180 3164.450 ;
        RECT 13.040 3091.690 13.180 3164.310 ;
        RECT 2887.580 3139.550 2887.720 3270.810 ;
        RECT 2887.520 3139.230 2887.780 3139.550 ;
        RECT 2898.560 3139.230 2898.820 3139.550 ;
        RECT 2898.620 3138.725 2898.760 3139.230 ;
        RECT 2898.550 3138.355 2898.830 3138.725 ;
        RECT 12.120 3091.550 13.180 3091.690 ;
        RECT 12.120 3010.090 12.260 3091.550 ;
        RECT 9.820 3010.010 12.260 3010.090 ;
        RECT 9.760 3009.950 12.260 3010.010 ;
        RECT 9.760 3009.690 10.020 3009.950 ;
        RECT 9.760 2998.470 10.020 2998.790 ;
        RECT 9.820 2995.810 9.960 2998.470 ;
        RECT 9.820 2995.670 12.260 2995.810 ;
        RECT 12.120 2986.290 12.260 2995.670 ;
        RECT 11.200 2986.150 12.260 2986.290 ;
        RECT 11.200 2982.890 11.340 2986.150 ;
        RECT 11.200 2982.750 12.260 2982.890 ;
        RECT 12.120 2959.940 12.260 2982.750 ;
        RECT 12.120 2959.800 12.720 2959.940 ;
        RECT 12.580 2891.770 12.720 2959.800 ;
        RECT 9.360 2891.630 12.720 2891.770 ;
        RECT 9.360 2846.210 9.500 2891.630 ;
        RECT 9.360 2846.070 10.880 2846.210 ;
        RECT 10.740 2836.010 10.880 2846.070 ;
        RECT 10.740 2835.870 11.340 2836.010 ;
        RECT 11.200 2827.850 11.340 2835.870 ;
        RECT 9.820 2827.770 11.340 2827.850 ;
        RECT 9.760 2827.710 11.340 2827.770 ;
        RECT 9.760 2827.450 10.020 2827.710 ;
        RECT 9.760 2815.610 10.020 2815.870 ;
        RECT 9.760 2815.550 11.340 2815.610 ;
        RECT 9.820 2815.470 11.340 2815.550 ;
        RECT 11.200 2780.250 11.340 2815.470 ;
        RECT 11.200 2780.110 11.800 2780.250 ;
        RECT 11.660 2705.450 11.800 2780.110 ;
        RECT 11.200 2705.310 11.800 2705.450 ;
        RECT 11.200 2636.090 11.340 2705.310 ;
        RECT 9.820 2636.010 11.340 2636.090 ;
        RECT 9.760 2635.950 11.340 2636.010 ;
        RECT 9.760 2635.690 10.020 2635.950 ;
        RECT 9.760 2612.290 10.020 2612.550 ;
        RECT 9.760 2612.230 11.340 2612.290 ;
        RECT 9.820 2612.150 11.340 2612.230 ;
        RECT 11.200 2536.810 11.340 2612.150 ;
        RECT 9.820 2536.730 11.340 2536.810 ;
        RECT 9.760 2536.670 11.340 2536.730 ;
        RECT 9.760 2536.410 10.020 2536.670 ;
        RECT 9.760 2508.930 10.020 2509.190 ;
        RECT 9.760 2508.870 11.800 2508.930 ;
        RECT 9.820 2508.790 11.800 2508.870 ;
        RECT 11.660 2445.010 11.800 2508.790 ;
        RECT 10.740 2444.870 11.800 2445.010 ;
        RECT 10.740 2438.890 10.880 2444.870 ;
        RECT 10.740 2438.750 11.340 2438.890 ;
        RECT 8.380 2363.690 8.640 2364.010 ;
        RECT 9.760 2363.920 10.020 2364.010 ;
        RECT 11.200 2363.920 11.340 2438.750 ;
        RECT 9.760 2363.780 11.340 2363.920 ;
        RECT 9.760 2363.690 10.020 2363.780 ;
        RECT 8.440 2338.930 8.580 2363.690 ;
        RECT 8.440 2338.790 11.340 2338.930 ;
        RECT 11.200 2250.530 11.340 2338.790 ;
        RECT 9.820 2250.450 11.340 2250.530 ;
        RECT 9.760 2250.390 11.340 2250.450 ;
        RECT 9.760 2250.130 10.020 2250.390 ;
        RECT 9.760 2238.910 10.020 2239.230 ;
        RECT 9.820 2211.770 9.960 2238.910 ;
        RECT 9.820 2211.630 10.880 2211.770 ;
        RECT 10.740 2207.690 10.880 2211.630 ;
        RECT 10.740 2207.550 11.800 2207.690 ;
        RECT 11.660 2090.730 11.800 2207.550 ;
        RECT 11.200 2090.590 11.800 2090.730 ;
        RECT 11.200 1935.010 11.340 2090.590 ;
        RECT 9.820 1934.930 11.340 1935.010 ;
        RECT 8.840 1934.610 9.100 1934.930 ;
        RECT 9.760 1934.870 11.340 1934.930 ;
        RECT 9.760 1934.610 10.020 1934.870 ;
        RECT 8.900 1903.650 9.040 1934.610 ;
        RECT 8.840 1903.330 9.100 1903.650 ;
        RECT 9.760 1894.890 10.020 1895.150 ;
        RECT 9.760 1894.830 10.420 1894.890 ;
        RECT 9.820 1894.750 10.420 1894.830 ;
        RECT 10.280 1852.730 10.420 1894.750 ;
        RECT 9.820 1852.590 10.420 1852.730 ;
        RECT 9.820 1851.970 9.960 1852.590 ;
        RECT 9.760 1851.650 10.020 1851.970 ;
        RECT 9.300 1790.450 9.560 1790.770 ;
        RECT 9.360 1756.170 9.500 1790.450 ;
        RECT 9.360 1756.030 9.960 1756.170 ;
        RECT 9.820 1728.890 9.960 1756.030 ;
        RECT 9.760 1728.570 10.020 1728.890 ;
        RECT 9.760 1648.730 10.020 1648.990 ;
        RECT 9.760 1648.670 11.340 1648.730 ;
        RECT 9.820 1648.590 11.340 1648.670 ;
        RECT 11.200 1626.970 11.340 1648.590 ;
        RECT 10.280 1626.830 11.340 1626.970 ;
        RECT 9.760 1594.840 10.020 1594.930 ;
        RECT 10.280 1594.840 10.420 1626.830 ;
        RECT 9.760 1594.700 10.420 1594.840 ;
        RECT 9.760 1594.610 10.020 1594.700 ;
        RECT 9.760 1558.290 10.020 1558.550 ;
        RECT 9.760 1558.230 11.340 1558.290 ;
        RECT 9.820 1558.150 11.340 1558.230 ;
        RECT 11.200 1527.010 11.340 1558.150 ;
        RECT 9.820 1526.930 11.340 1527.010 ;
        RECT 9.760 1526.870 11.340 1526.930 ;
        RECT 9.760 1526.610 10.020 1526.870 ;
        RECT 6.540 1481.050 6.800 1481.370 ;
        RECT 6.600 1320.210 6.740 1481.050 ;
        RECT 6.540 1319.890 6.800 1320.210 ;
        RECT 9.760 1319.890 10.020 1320.210 ;
        RECT 9.820 1287.650 9.960 1319.890 ;
        RECT 9.820 1287.510 12.260 1287.650 ;
        RECT 12.120 1238.690 12.260 1287.510 ;
        RECT 10.740 1238.550 12.260 1238.690 ;
        RECT 10.740 1210.810 10.880 1238.550 ;
        RECT 9.360 1210.670 10.880 1210.810 ;
        RECT 9.360 1190.410 9.500 1210.670 ;
        RECT 8.900 1190.270 9.500 1190.410 ;
        RECT 8.900 1177.410 9.040 1190.270 ;
        RECT 2.400 1177.090 2.660 1177.410 ;
        RECT 8.840 1177.090 9.100 1177.410 ;
        RECT 2.460 872.850 2.600 1177.090 ;
        RECT 2.000 872.710 2.600 872.850 ;
        RECT 2.000 838.430 2.140 872.710 ;
        RECT 1.940 838.110 2.200 838.430 ;
        RECT 7.000 773.850 7.260 774.170 ;
        RECT 7.060 743.230 7.200 773.850 ;
        RECT 7.000 742.910 7.260 743.230 ;
        RECT 4.700 671.850 4.960 672.170 ;
        RECT 4.760 606.210 4.900 671.850 ;
        RECT 3.780 605.890 4.040 606.210 ;
        RECT 4.700 605.890 4.960 606.210 ;
        RECT 3.840 99.805 3.980 605.890 ;
        RECT 3.770 99.435 4.050 99.805 ;
        RECT 52.080 7.830 52.340 8.150 ;
        RECT 292.190 7.890 292.470 8.005 ;
        RECT 52.140 5.965 52.280 7.830 ;
        RECT 283.000 7.490 283.260 7.810 ;
        RECT 292.190 7.750 292.860 7.890 ;
        RECT 292.190 7.635 292.470 7.750 ;
        RECT 244.820 7.150 245.080 7.470 ;
        RECT 283.060 7.325 283.200 7.490 ;
        RECT 292.720 7.325 292.860 7.750 ;
        RECT 139.480 6.130 139.740 6.450 ;
        RECT 52.070 5.595 52.350 5.965 ;
        RECT 139.540 5.285 139.680 6.130 ;
        RECT 139.470 4.915 139.750 5.285 ;
        RECT 232.850 4.915 233.130 5.285 ;
        RECT 232.920 3.925 233.060 4.915 ;
        RECT 244.880 3.925 245.020 7.150 ;
        RECT 282.990 6.955 283.270 7.325 ;
        RECT 292.650 6.955 292.930 7.325 ;
        RECT 311.970 7.210 312.250 7.325 ;
        RECT 313.290 7.210 313.570 9.000 ;
        RECT 311.970 7.070 313.570 7.210 ;
        RECT 311.970 6.955 312.250 7.070 ;
        RECT 313.290 5.000 313.570 7.070 ;
        RECT 232.850 3.555 233.130 3.925 ;
        RECT 244.810 3.555 245.090 3.925 ;
      LAYER via2 ;
        RECT 2898.550 3138.400 2898.830 3138.680 ;
        RECT 3.770 99.480 4.050 99.760 ;
        RECT 292.190 7.680 292.470 7.960 ;
        RECT 52.070 5.640 52.350 5.920 ;
        RECT 139.470 4.960 139.750 5.240 ;
        RECT 232.850 4.960 233.130 5.240 ;
        RECT 282.990 7.000 283.270 7.280 ;
        RECT 292.650 7.000 292.930 7.280 ;
        RECT 311.970 7.000 312.250 7.280 ;
        RECT 232.850 3.600 233.130 3.880 ;
        RECT 244.810 3.600 245.090 3.880 ;
      LAYER met3 ;
        RECT 2898.525 3138.690 2898.855 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2898.525 3138.390 2924.800 3138.690 ;
        RECT 2898.525 3138.375 2898.855 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
        RECT 3.745 99.770 4.075 99.785 ;
        RECT 6.710 99.770 7.090 99.780 ;
        RECT 3.745 99.470 7.090 99.770 ;
        RECT 3.745 99.455 4.075 99.470 ;
        RECT 6.710 99.460 7.090 99.470 ;
        RECT 292.165 7.970 292.495 7.985 ;
        RECT 290.110 7.670 292.495 7.970 ;
        RECT 282.965 7.290 283.295 7.305 ;
        RECT 290.110 7.290 290.410 7.670 ;
        RECT 292.165 7.655 292.495 7.670 ;
        RECT 282.965 6.990 290.410 7.290 ;
        RECT 292.625 7.290 292.955 7.305 ;
        RECT 311.945 7.290 312.275 7.305 ;
        RECT 292.625 6.990 312.275 7.290 ;
        RECT 282.965 6.975 283.295 6.990 ;
        RECT 292.625 6.975 292.955 6.990 ;
        RECT 311.945 6.975 312.275 6.990 ;
        RECT 14.070 5.930 14.450 5.940 ;
        RECT 52.045 5.930 52.375 5.945 ;
        RECT 14.070 5.630 52.375 5.930 ;
        RECT 14.070 5.620 14.450 5.630 ;
        RECT 52.045 5.615 52.375 5.630 ;
        RECT 139.445 5.250 139.775 5.265 ;
        RECT 232.825 5.250 233.155 5.265 ;
        RECT 139.445 4.950 233.155 5.250 ;
        RECT 139.445 4.935 139.775 4.950 ;
        RECT 232.825 4.935 233.155 4.950 ;
        RECT 232.825 3.890 233.155 3.905 ;
        RECT 244.785 3.890 245.115 3.905 ;
        RECT 232.825 3.590 245.115 3.890 ;
        RECT 232.825 3.575 233.155 3.590 ;
        RECT 244.785 3.575 245.115 3.590 ;
      LAYER via3 ;
        RECT 6.740 99.460 7.060 99.780 ;
        RECT 14.100 5.620 14.420 5.940 ;
      LAYER met4 ;
        RECT 6.735 99.455 7.065 99.785 ;
        RECT 6.750 80.050 7.050 99.455 ;
        RECT 6.750 79.750 11.650 80.050 ;
        RECT 11.350 49.450 11.650 79.750 ;
        RECT 11.350 49.150 14.410 49.450 ;
        RECT 14.110 5.945 14.410 49.150 ;
        RECT 14.095 5.615 14.425 5.945 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 9.345 3167.185 9.515 3213.255 ;
        RECT 9.345 2832.965 9.515 2902.495 ;
        RECT 9.805 2738.445 9.975 2818.855 ;
        RECT 8.885 2487.525 9.055 2520.675 ;
        RECT 8.425 2324.665 8.595 2418.675 ;
        RECT 9.345 1903.405 9.515 1936.215 ;
        RECT 7.045 1790.185 7.215 1846.455 ;
        RECT 8.885 1679.855 9.055 1703.655 ;
        RECT 8.885 1679.685 9.515 1679.855 ;
        RECT 7.505 1563.405 7.675 1632.595 ;
        RECT 9.345 1632.425 9.515 1679.685 ;
        RECT 9.805 1549.125 9.975 1563.575 ;
        RECT 8.425 1507.305 8.595 1528.215 ;
        RECT 8.885 1416.865 9.055 1480.615 ;
        RECT 9.805 1250.605 9.975 1323.535 ;
        RECT 9.345 1113.415 9.515 1209.975 ;
        RECT 8.885 1113.245 9.515 1113.415 ;
        RECT 8.885 1106.445 9.055 1113.245 ;
        RECT 8.885 1028.755 9.055 1087.235 ;
        RECT 8.885 1028.585 9.515 1028.755 ;
        RECT 7.505 975.885 7.675 1003.595 ;
        RECT 9.345 1003.425 9.515 1028.585 ;
        RECT 8.885 895.305 9.055 976.055 ;
        RECT 8.425 865.045 8.595 884.935 ;
        RECT 7.965 817.105 8.135 840.055 ;
        RECT 9.805 734.825 9.975 817.275 ;
        RECT 7.505 689.605 7.675 706.775 ;
        RECT 6.125 541.705 6.295 672.435 ;
        RECT 6.125 458.745 6.295 468.095 ;
        RECT 6.585 403.665 6.755 419.135 ;
        RECT 7.045 314.925 7.215 346.715 ;
        RECT 7.045 275.825 7.215 283.815 ;
        RECT 303.745 7.225 304.835 7.395 ;
        RECT 246.245 1.445 246.415 2.975 ;
        RECT 303.745 0.765 303.915 7.225 ;
        RECT 310.645 6.545 310.815 7.395 ;
        RECT 316.625 6.545 316.795 8.415 ;
      LAYER mcon ;
        RECT 9.345 3213.085 9.515 3213.255 ;
        RECT 9.345 2902.325 9.515 2902.495 ;
        RECT 9.805 2818.685 9.975 2818.855 ;
        RECT 8.885 2520.505 9.055 2520.675 ;
        RECT 8.425 2418.505 8.595 2418.675 ;
        RECT 9.345 1936.045 9.515 1936.215 ;
        RECT 7.045 1846.285 7.215 1846.455 ;
        RECT 8.885 1703.485 9.055 1703.655 ;
        RECT 7.505 1632.425 7.675 1632.595 ;
        RECT 9.805 1563.405 9.975 1563.575 ;
        RECT 8.425 1528.045 8.595 1528.215 ;
        RECT 8.885 1480.445 9.055 1480.615 ;
        RECT 9.805 1323.365 9.975 1323.535 ;
        RECT 9.345 1209.805 9.515 1209.975 ;
        RECT 8.885 1087.065 9.055 1087.235 ;
        RECT 7.505 1003.425 7.675 1003.595 ;
        RECT 8.885 975.885 9.055 976.055 ;
        RECT 8.425 884.765 8.595 884.935 ;
        RECT 7.965 839.885 8.135 840.055 ;
        RECT 9.805 817.105 9.975 817.275 ;
        RECT 7.505 706.605 7.675 706.775 ;
        RECT 6.125 672.265 6.295 672.435 ;
        RECT 6.125 467.925 6.295 468.095 ;
        RECT 6.585 418.965 6.755 419.135 ;
        RECT 7.045 346.545 7.215 346.715 ;
        RECT 7.045 283.645 7.215 283.815 ;
        RECT 316.625 8.245 316.795 8.415 ;
        RECT 304.665 7.225 304.835 7.395 ;
        RECT 310.645 7.225 310.815 7.395 ;
        RECT 246.245 2.805 246.415 2.975 ;
      LAYER met1 ;
        RECT 9.270 3395.140 9.590 3395.200 ;
        RECT 2857.130 3395.140 2857.450 3395.200 ;
        RECT 9.270 3395.000 2857.450 3395.140 ;
        RECT 9.270 3394.940 9.590 3395.000 ;
        RECT 2857.130 3394.940 2857.450 3395.000 ;
        RECT 2857.130 3387.660 2857.450 3387.720 ;
        RECT 2890.710 3387.660 2891.030 3387.720 ;
        RECT 2857.130 3387.520 2891.030 3387.660 ;
        RECT 2857.130 3387.460 2857.450 3387.520 ;
        RECT 2890.710 3387.460 2891.030 3387.520 ;
        RECT 2890.710 3374.060 2891.030 3374.120 ;
        RECT 2900.830 3374.060 2901.150 3374.120 ;
        RECT 2890.710 3373.920 2901.150 3374.060 ;
        RECT 2890.710 3373.860 2891.030 3373.920 ;
        RECT 2900.830 3373.860 2901.150 3373.920 ;
        RECT 9.270 3243.160 9.590 3243.220 ;
        RECT 9.730 3243.160 10.050 3243.220 ;
        RECT 9.270 3243.020 10.050 3243.160 ;
        RECT 9.270 3242.960 9.590 3243.020 ;
        RECT 9.730 3242.960 10.050 3243.020 ;
        RECT 9.285 3213.240 9.575 3213.285 ;
        RECT 9.730 3213.240 10.050 3213.300 ;
        RECT 9.285 3213.100 10.050 3213.240 ;
        RECT 9.285 3213.055 9.575 3213.100 ;
        RECT 9.730 3213.040 10.050 3213.100 ;
        RECT 9.270 3167.340 9.590 3167.400 ;
        RECT 9.075 3167.200 9.590 3167.340 ;
        RECT 9.270 3167.140 9.590 3167.200 ;
        RECT 9.270 3091.520 9.590 3091.580 ;
        RECT 9.730 3091.520 10.050 3091.580 ;
        RECT 9.270 3091.380 10.050 3091.520 ;
        RECT 9.270 3091.320 9.590 3091.380 ;
        RECT 9.730 3091.320 10.050 3091.380 ;
        RECT 9.730 3043.580 10.050 3043.640 ;
        RECT 9.360 3043.440 10.050 3043.580 ;
        RECT 9.360 3042.960 9.500 3043.440 ;
        RECT 9.730 3043.380 10.050 3043.440 ;
        RECT 9.270 3042.700 9.590 3042.960 ;
        RECT 9.285 2902.480 9.575 2902.525 ;
        RECT 9.730 2902.480 10.050 2902.540 ;
        RECT 9.285 2902.340 10.050 2902.480 ;
        RECT 9.285 2902.295 9.575 2902.340 ;
        RECT 9.730 2902.280 10.050 2902.340 ;
        RECT 9.270 2833.120 9.590 2833.180 ;
        RECT 9.075 2832.980 9.590 2833.120 ;
        RECT 9.270 2832.920 9.590 2832.980 ;
        RECT 9.270 2818.840 9.590 2818.900 ;
        RECT 9.745 2818.840 10.035 2818.885 ;
        RECT 9.270 2818.700 10.035 2818.840 ;
        RECT 9.270 2818.640 9.590 2818.700 ;
        RECT 9.745 2818.655 10.035 2818.700 ;
        RECT 9.270 2738.600 9.590 2738.660 ;
        RECT 9.745 2738.600 10.035 2738.645 ;
        RECT 9.270 2738.460 10.035 2738.600 ;
        RECT 9.270 2738.400 9.590 2738.460 ;
        RECT 9.745 2738.415 10.035 2738.460 ;
        RECT 9.270 2670.060 9.590 2670.320 ;
        RECT 9.360 2669.300 9.500 2670.060 ;
        RECT 9.270 2669.040 9.590 2669.300 ;
        RECT 8.810 2520.660 9.130 2520.720 ;
        RECT 8.615 2520.520 9.130 2520.660 ;
        RECT 8.810 2520.460 9.130 2520.520 ;
        RECT 8.810 2487.680 9.130 2487.740 ;
        RECT 8.615 2487.540 9.130 2487.680 ;
        RECT 8.810 2487.480 9.130 2487.540 ;
        RECT 8.365 2418.660 8.655 2418.705 ;
        RECT 8.810 2418.660 9.130 2418.720 ;
        RECT 8.365 2418.520 9.130 2418.660 ;
        RECT 8.365 2418.475 8.655 2418.520 ;
        RECT 8.810 2418.460 9.130 2418.520 ;
        RECT 8.365 2324.820 8.655 2324.865 ;
        RECT 9.730 2324.820 10.050 2324.880 ;
        RECT 8.365 2324.680 10.050 2324.820 ;
        RECT 8.365 2324.635 8.655 2324.680 ;
        RECT 9.730 2324.620 10.050 2324.680 ;
        RECT 8.810 2254.440 9.130 2254.500 ;
        RECT 9.730 2254.440 10.050 2254.500 ;
        RECT 8.810 2254.300 10.050 2254.440 ;
        RECT 8.810 2254.240 9.130 2254.300 ;
        RECT 9.730 2254.240 10.050 2254.300 ;
        RECT 8.350 2161.280 8.670 2161.340 ;
        RECT 9.730 2161.280 10.050 2161.340 ;
        RECT 8.350 2161.140 10.050 2161.280 ;
        RECT 8.350 2161.080 8.670 2161.140 ;
        RECT 9.730 2161.080 10.050 2161.140 ;
        RECT 9.285 1936.200 9.575 1936.245 ;
        RECT 9.730 1936.200 10.050 1936.260 ;
        RECT 9.285 1936.060 10.050 1936.200 ;
        RECT 9.285 1936.015 9.575 1936.060 ;
        RECT 9.730 1936.000 10.050 1936.060 ;
        RECT 9.285 1903.560 9.575 1903.605 ;
        RECT 9.730 1903.560 10.050 1903.620 ;
        RECT 9.285 1903.420 10.050 1903.560 ;
        RECT 9.285 1903.375 9.575 1903.420 ;
        RECT 9.730 1903.360 10.050 1903.420 ;
        RECT 6.985 1846.440 7.275 1846.485 ;
        RECT 9.730 1846.440 10.050 1846.500 ;
        RECT 6.985 1846.300 10.050 1846.440 ;
        RECT 6.985 1846.255 7.275 1846.300 ;
        RECT 9.730 1846.240 10.050 1846.300 ;
        RECT 6.985 1790.340 7.275 1790.385 ;
        RECT 8.810 1790.340 9.130 1790.400 ;
        RECT 6.985 1790.200 9.130 1790.340 ;
        RECT 6.985 1790.155 7.275 1790.200 ;
        RECT 8.810 1790.140 9.130 1790.200 ;
        RECT 8.810 1765.520 9.130 1765.580 ;
        RECT 9.730 1765.520 10.050 1765.580 ;
        RECT 8.810 1765.380 10.050 1765.520 ;
        RECT 8.810 1765.320 9.130 1765.380 ;
        RECT 9.730 1765.320 10.050 1765.380 ;
        RECT 8.825 1703.640 9.115 1703.685 ;
        RECT 9.730 1703.640 10.050 1703.700 ;
        RECT 8.825 1703.500 10.050 1703.640 ;
        RECT 8.825 1703.455 9.115 1703.500 ;
        RECT 9.730 1703.440 10.050 1703.500 ;
        RECT 7.445 1632.580 7.735 1632.625 ;
        RECT 9.285 1632.580 9.575 1632.625 ;
        RECT 7.445 1632.440 9.575 1632.580 ;
        RECT 7.445 1632.395 7.735 1632.440 ;
        RECT 9.285 1632.395 9.575 1632.440 ;
        RECT 7.445 1563.560 7.735 1563.605 ;
        RECT 9.745 1563.560 10.035 1563.605 ;
        RECT 7.445 1563.420 10.035 1563.560 ;
        RECT 7.445 1563.375 7.735 1563.420 ;
        RECT 9.745 1563.375 10.035 1563.420 ;
        RECT 9.730 1549.280 10.050 1549.340 ;
        RECT 9.535 1549.140 10.050 1549.280 ;
        RECT 9.730 1549.080 10.050 1549.140 ;
        RECT 8.365 1528.200 8.655 1528.245 ;
        RECT 9.730 1528.200 10.050 1528.260 ;
        RECT 8.365 1528.060 10.050 1528.200 ;
        RECT 8.365 1528.015 8.655 1528.060 ;
        RECT 9.730 1528.000 10.050 1528.060 ;
        RECT 8.365 1507.460 8.655 1507.505 ;
        RECT 9.730 1507.460 10.050 1507.520 ;
        RECT 8.365 1507.320 10.050 1507.460 ;
        RECT 8.365 1507.275 8.655 1507.320 ;
        RECT 9.730 1507.260 10.050 1507.320 ;
        RECT 8.825 1480.600 9.115 1480.645 ;
        RECT 9.730 1480.600 10.050 1480.660 ;
        RECT 8.825 1480.460 10.050 1480.600 ;
        RECT 8.825 1480.415 9.115 1480.460 ;
        RECT 9.730 1480.400 10.050 1480.460 ;
        RECT 8.825 1417.020 9.115 1417.065 ;
        RECT 9.730 1417.020 10.050 1417.080 ;
        RECT 8.825 1416.880 10.050 1417.020 ;
        RECT 8.825 1416.835 9.115 1416.880 ;
        RECT 9.730 1416.820 10.050 1416.880 ;
        RECT 9.730 1323.520 10.050 1323.580 ;
        RECT 9.535 1323.380 10.050 1323.520 ;
        RECT 9.730 1323.320 10.050 1323.380 ;
        RECT 9.730 1250.760 10.050 1250.820 ;
        RECT 9.535 1250.620 10.050 1250.760 ;
        RECT 9.730 1250.560 10.050 1250.620 ;
        RECT 9.730 1211.120 10.050 1211.380 ;
        RECT 9.285 1209.960 9.575 1210.005 ;
        RECT 9.820 1209.960 9.960 1211.120 ;
        RECT 9.285 1209.820 9.960 1209.960 ;
        RECT 9.285 1209.775 9.575 1209.820 ;
        RECT 6.970 1106.600 7.290 1106.660 ;
        RECT 8.825 1106.600 9.115 1106.645 ;
        RECT 6.970 1106.460 9.115 1106.600 ;
        RECT 6.970 1106.400 7.290 1106.460 ;
        RECT 8.825 1106.415 9.115 1106.460 ;
        RECT 6.970 1087.220 7.290 1087.280 ;
        RECT 8.825 1087.220 9.115 1087.265 ;
        RECT 6.970 1087.080 9.115 1087.220 ;
        RECT 6.970 1087.020 7.290 1087.080 ;
        RECT 8.825 1087.035 9.115 1087.080 ;
        RECT 7.445 1003.580 7.735 1003.625 ;
        RECT 9.285 1003.580 9.575 1003.625 ;
        RECT 7.445 1003.440 9.575 1003.580 ;
        RECT 7.445 1003.395 7.735 1003.440 ;
        RECT 9.285 1003.395 9.575 1003.440 ;
        RECT 7.445 976.040 7.735 976.085 ;
        RECT 8.825 976.040 9.115 976.085 ;
        RECT 7.445 975.900 9.115 976.040 ;
        RECT 7.445 975.855 7.735 975.900 ;
        RECT 8.825 975.855 9.115 975.900 ;
        RECT 8.825 895.460 9.115 895.505 ;
        RECT 9.270 895.460 9.590 895.520 ;
        RECT 8.825 895.320 9.590 895.460 ;
        RECT 8.825 895.275 9.115 895.320 ;
        RECT 9.270 895.260 9.590 895.320 ;
        RECT 8.365 884.920 8.655 884.965 ;
        RECT 9.270 884.920 9.590 884.980 ;
        RECT 8.365 884.780 9.590 884.920 ;
        RECT 8.365 884.735 8.655 884.780 ;
        RECT 9.270 884.720 9.590 884.780 ;
        RECT 8.365 865.200 8.655 865.245 ;
        RECT 9.270 865.200 9.590 865.260 ;
        RECT 8.365 865.060 9.590 865.200 ;
        RECT 8.365 865.015 8.655 865.060 ;
        RECT 9.270 865.000 9.590 865.060 ;
        RECT 7.905 840.040 8.195 840.085 ;
        RECT 9.730 840.040 10.050 840.100 ;
        RECT 7.905 839.900 10.050 840.040 ;
        RECT 7.905 839.855 8.195 839.900 ;
        RECT 9.730 839.840 10.050 839.900 ;
        RECT 7.905 817.260 8.195 817.305 ;
        RECT 9.745 817.260 10.035 817.305 ;
        RECT 7.905 817.120 10.035 817.260 ;
        RECT 7.905 817.075 8.195 817.120 ;
        RECT 9.745 817.075 10.035 817.120 ;
        RECT 9.730 734.980 10.050 735.040 ;
        RECT 9.535 734.840 10.050 734.980 ;
        RECT 9.730 734.780 10.050 734.840 ;
        RECT 9.730 729.000 10.050 729.260 ;
        RECT 9.820 728.240 9.960 729.000 ;
        RECT 9.730 727.980 10.050 728.240 ;
        RECT 7.445 706.760 7.735 706.805 ;
        RECT 9.730 706.760 10.050 706.820 ;
        RECT 7.445 706.620 10.050 706.760 ;
        RECT 7.445 706.575 7.735 706.620 ;
        RECT 9.730 706.560 10.050 706.620 ;
        RECT 7.445 689.760 7.735 689.805 ;
        RECT 9.730 689.760 10.050 689.820 ;
        RECT 7.445 689.620 10.050 689.760 ;
        RECT 7.445 689.575 7.735 689.620 ;
        RECT 9.730 689.560 10.050 689.620 ;
        RECT 6.065 672.420 6.355 672.465 ;
        RECT 9.730 672.420 10.050 672.480 ;
        RECT 6.065 672.280 10.050 672.420 ;
        RECT 6.065 672.235 6.355 672.280 ;
        RECT 9.730 672.220 10.050 672.280 ;
        RECT 6.065 541.860 6.355 541.905 ;
        RECT 9.730 541.860 10.050 541.920 ;
        RECT 6.065 541.720 10.050 541.860 ;
        RECT 6.065 541.675 6.355 541.720 ;
        RECT 9.730 541.660 10.050 541.720 ;
        RECT 6.065 468.080 6.355 468.125 ;
        RECT 9.730 468.080 10.050 468.140 ;
        RECT 6.065 467.940 10.050 468.080 ;
        RECT 6.065 467.895 6.355 467.940 ;
        RECT 9.730 467.880 10.050 467.940 ;
        RECT 6.065 458.900 6.355 458.945 ;
        RECT 9.730 458.900 10.050 458.960 ;
        RECT 6.065 458.760 10.050 458.900 ;
        RECT 6.065 458.715 6.355 458.760 ;
        RECT 9.730 458.700 10.050 458.760 ;
        RECT 6.525 419.120 6.815 419.165 ;
        RECT 9.730 419.120 10.050 419.180 ;
        RECT 6.525 418.980 10.050 419.120 ;
        RECT 6.525 418.935 6.815 418.980 ;
        RECT 9.730 418.920 10.050 418.980 ;
        RECT 6.525 403.820 6.815 403.865 ;
        RECT 9.730 403.820 10.050 403.880 ;
        RECT 6.525 403.680 10.050 403.820 ;
        RECT 6.525 403.635 6.815 403.680 ;
        RECT 9.730 403.620 10.050 403.680 ;
        RECT 6.510 360.980 6.830 361.040 ;
        RECT 9.730 360.980 10.050 361.040 ;
        RECT 6.510 360.840 10.050 360.980 ;
        RECT 6.510 360.780 6.830 360.840 ;
        RECT 9.730 360.780 10.050 360.840 ;
        RECT 6.510 346.700 6.830 346.760 ;
        RECT 6.985 346.700 7.275 346.745 ;
        RECT 6.510 346.560 7.275 346.700 ;
        RECT 6.510 346.500 6.830 346.560 ;
        RECT 6.985 346.515 7.275 346.560 ;
        RECT 6.985 315.080 7.275 315.125 ;
        RECT 9.730 315.080 10.050 315.140 ;
        RECT 6.985 314.940 10.050 315.080 ;
        RECT 6.985 314.895 7.275 314.940 ;
        RECT 9.730 314.880 10.050 314.940 ;
        RECT 6.985 283.800 7.275 283.845 ;
        RECT 9.730 283.800 10.050 283.860 ;
        RECT 6.985 283.660 10.050 283.800 ;
        RECT 6.985 283.615 7.275 283.660 ;
        RECT 9.730 283.600 10.050 283.660 ;
        RECT 6.985 275.980 7.275 276.025 ;
        RECT 9.730 275.980 10.050 276.040 ;
        RECT 6.985 275.840 10.050 275.980 ;
        RECT 6.985 275.795 7.275 275.840 ;
        RECT 9.730 275.780 10.050 275.840 ;
        RECT 1.910 176.360 2.230 176.420 ;
        RECT 9.730 176.360 10.050 176.420 ;
        RECT 1.910 176.220 10.050 176.360 ;
        RECT 1.910 176.160 2.230 176.220 ;
        RECT 9.730 176.160 10.050 176.220 ;
        RECT 316.565 8.400 316.855 8.445 ;
        RECT 358.870 8.400 359.190 8.460 ;
        RECT 316.565 8.260 359.190 8.400 ;
        RECT 316.565 8.215 316.855 8.260 ;
        RECT 358.870 8.200 359.190 8.260 ;
        RECT 304.605 7.380 304.895 7.425 ;
        RECT 310.585 7.380 310.875 7.425 ;
        RECT 304.605 7.240 310.875 7.380 ;
        RECT 304.605 7.195 304.895 7.240 ;
        RECT 310.585 7.195 310.875 7.240 ;
        RECT 310.585 6.700 310.875 6.745 ;
        RECT 316.565 6.700 316.855 6.745 ;
        RECT 310.585 6.560 316.855 6.700 ;
        RECT 310.585 6.515 310.875 6.560 ;
        RECT 316.565 6.515 316.855 6.560 ;
        RECT 36.870 3.300 37.190 3.360 ;
        RECT 36.870 3.160 133.240 3.300 ;
        RECT 36.870 3.100 37.190 3.160 ;
        RECT 133.100 2.960 133.240 3.160 ;
        RECT 246.185 2.960 246.475 3.005 ;
        RECT 133.100 2.820 246.475 2.960 ;
        RECT 246.185 2.775 246.475 2.820 ;
        RECT 246.185 1.600 246.475 1.645 ;
        RECT 294.930 1.600 295.250 1.660 ;
        RECT 246.185 1.460 295.250 1.600 ;
        RECT 246.185 1.415 246.475 1.460 ;
        RECT 294.930 1.400 295.250 1.460 ;
        RECT 294.930 0.920 295.250 0.980 ;
        RECT 303.685 0.920 303.975 0.965 ;
        RECT 294.930 0.780 303.975 0.920 ;
        RECT 294.930 0.720 295.250 0.780 ;
        RECT 303.685 0.735 303.975 0.780 ;
      LAYER via ;
        RECT 9.300 3394.940 9.560 3395.200 ;
        RECT 2857.160 3394.940 2857.420 3395.200 ;
        RECT 2857.160 3387.460 2857.420 3387.720 ;
        RECT 2890.740 3387.460 2891.000 3387.720 ;
        RECT 2890.740 3373.860 2891.000 3374.120 ;
        RECT 2900.860 3373.860 2901.120 3374.120 ;
        RECT 9.300 3242.960 9.560 3243.220 ;
        RECT 9.760 3242.960 10.020 3243.220 ;
        RECT 9.760 3213.040 10.020 3213.300 ;
        RECT 9.300 3167.140 9.560 3167.400 ;
        RECT 9.300 3091.320 9.560 3091.580 ;
        RECT 9.760 3091.320 10.020 3091.580 ;
        RECT 9.760 3043.380 10.020 3043.640 ;
        RECT 9.300 3042.700 9.560 3042.960 ;
        RECT 9.760 2902.280 10.020 2902.540 ;
        RECT 9.300 2832.920 9.560 2833.180 ;
        RECT 9.300 2818.640 9.560 2818.900 ;
        RECT 9.300 2738.400 9.560 2738.660 ;
        RECT 9.300 2670.060 9.560 2670.320 ;
        RECT 9.300 2669.040 9.560 2669.300 ;
        RECT 8.840 2520.460 9.100 2520.720 ;
        RECT 8.840 2487.480 9.100 2487.740 ;
        RECT 8.840 2418.460 9.100 2418.720 ;
        RECT 9.760 2324.620 10.020 2324.880 ;
        RECT 8.840 2254.240 9.100 2254.500 ;
        RECT 9.760 2254.240 10.020 2254.500 ;
        RECT 8.380 2161.080 8.640 2161.340 ;
        RECT 9.760 2161.080 10.020 2161.340 ;
        RECT 9.760 1936.000 10.020 1936.260 ;
        RECT 9.760 1903.360 10.020 1903.620 ;
        RECT 9.760 1846.240 10.020 1846.500 ;
        RECT 8.840 1790.140 9.100 1790.400 ;
        RECT 8.840 1765.320 9.100 1765.580 ;
        RECT 9.760 1765.320 10.020 1765.580 ;
        RECT 9.760 1703.440 10.020 1703.700 ;
        RECT 9.760 1549.080 10.020 1549.340 ;
        RECT 9.760 1528.000 10.020 1528.260 ;
        RECT 9.760 1507.260 10.020 1507.520 ;
        RECT 9.760 1480.400 10.020 1480.660 ;
        RECT 9.760 1416.820 10.020 1417.080 ;
        RECT 9.760 1323.320 10.020 1323.580 ;
        RECT 9.760 1250.560 10.020 1250.820 ;
        RECT 9.760 1211.120 10.020 1211.380 ;
        RECT 7.000 1106.400 7.260 1106.660 ;
        RECT 7.000 1087.020 7.260 1087.280 ;
        RECT 9.300 895.260 9.560 895.520 ;
        RECT 9.300 884.720 9.560 884.980 ;
        RECT 9.300 865.000 9.560 865.260 ;
        RECT 9.760 839.840 10.020 840.100 ;
        RECT 9.760 734.780 10.020 735.040 ;
        RECT 9.760 729.000 10.020 729.260 ;
        RECT 9.760 727.980 10.020 728.240 ;
        RECT 9.760 706.560 10.020 706.820 ;
        RECT 9.760 689.560 10.020 689.820 ;
        RECT 9.760 672.220 10.020 672.480 ;
        RECT 9.760 541.660 10.020 541.920 ;
        RECT 9.760 467.880 10.020 468.140 ;
        RECT 9.760 458.700 10.020 458.960 ;
        RECT 9.760 418.920 10.020 419.180 ;
        RECT 9.760 403.620 10.020 403.880 ;
        RECT 6.540 360.780 6.800 361.040 ;
        RECT 9.760 360.780 10.020 361.040 ;
        RECT 6.540 346.500 6.800 346.760 ;
        RECT 9.760 314.880 10.020 315.140 ;
        RECT 9.760 283.600 10.020 283.860 ;
        RECT 9.760 275.780 10.020 276.040 ;
        RECT 1.940 176.160 2.200 176.420 ;
        RECT 9.760 176.160 10.020 176.420 ;
        RECT 358.900 8.200 359.160 8.460 ;
        RECT 36.900 3.100 37.160 3.360 ;
        RECT 294.960 1.400 295.220 1.660 ;
        RECT 294.960 0.720 295.220 0.980 ;
      LAYER met2 ;
        RECT 9.300 3394.910 9.560 3395.230 ;
        RECT 2857.160 3394.910 2857.420 3395.230 ;
        RECT 9.360 3362.330 9.500 3394.910 ;
        RECT 2857.220 3387.750 2857.360 3394.910 ;
        RECT 2857.160 3387.430 2857.420 3387.750 ;
        RECT 2890.740 3387.430 2891.000 3387.750 ;
        RECT 2890.800 3374.150 2890.940 3387.430 ;
        RECT 2890.740 3373.830 2891.000 3374.150 ;
        RECT 2900.860 3373.830 2901.120 3374.150 ;
        RECT 2900.920 3373.325 2901.060 3373.830 ;
        RECT 2900.850 3372.955 2901.130 3373.325 ;
        RECT 9.360 3362.190 10.420 3362.330 ;
        RECT 10.280 3290.930 10.420 3362.190 ;
        RECT 9.820 3290.790 10.420 3290.930 ;
        RECT 9.820 3243.250 9.960 3290.790 ;
        RECT 9.300 3242.930 9.560 3243.250 ;
        RECT 9.760 3242.930 10.020 3243.250 ;
        RECT 9.360 3239.930 9.500 3242.930 ;
        RECT 9.360 3239.790 9.960 3239.930 ;
        RECT 9.820 3213.330 9.960 3239.790 ;
        RECT 9.760 3213.010 10.020 3213.330 ;
        RECT 9.300 3167.110 9.560 3167.430 ;
        RECT 9.360 3091.610 9.500 3167.110 ;
        RECT 9.300 3091.290 9.560 3091.610 ;
        RECT 9.760 3091.290 10.020 3091.610 ;
        RECT 9.820 3043.670 9.960 3091.290 ;
        RECT 9.760 3043.350 10.020 3043.670 ;
        RECT 9.300 3042.670 9.560 3042.990 ;
        RECT 9.360 2981.530 9.500 3042.670 ;
        RECT 9.360 2981.390 9.960 2981.530 ;
        RECT 9.820 2902.570 9.960 2981.390 ;
        RECT 9.760 2902.250 10.020 2902.570 ;
        RECT 9.300 2832.890 9.560 2833.210 ;
        RECT 9.360 2818.930 9.500 2832.890 ;
        RECT 9.300 2818.610 9.560 2818.930 ;
        RECT 9.300 2738.370 9.560 2738.690 ;
        RECT 9.360 2670.350 9.500 2738.370 ;
        RECT 9.300 2670.030 9.560 2670.350 ;
        RECT 9.300 2669.010 9.560 2669.330 ;
        RECT 9.360 2549.050 9.500 2669.010 ;
        RECT 8.900 2548.910 9.500 2549.050 ;
        RECT 8.900 2520.750 9.040 2548.910 ;
        RECT 8.840 2520.430 9.100 2520.750 ;
        RECT 8.840 2487.450 9.100 2487.770 ;
        RECT 8.900 2418.750 9.040 2487.450 ;
        RECT 8.840 2418.430 9.100 2418.750 ;
        RECT 9.760 2324.820 10.020 2324.910 ;
        RECT 9.760 2324.680 10.420 2324.820 ;
        RECT 9.760 2324.590 10.020 2324.680 ;
        RECT 10.280 2254.610 10.420 2324.680 ;
        RECT 9.820 2254.530 10.420 2254.610 ;
        RECT 8.840 2254.210 9.100 2254.530 ;
        RECT 9.760 2254.470 10.420 2254.530 ;
        RECT 9.760 2254.210 10.020 2254.470 ;
        RECT 8.900 2211.090 9.040 2254.210 ;
        RECT 8.900 2210.950 9.500 2211.090 ;
        RECT 9.360 2206.330 9.500 2210.950 ;
        RECT 9.360 2206.190 10.420 2206.330 ;
        RECT 10.280 2161.450 10.420 2206.190 ;
        RECT 9.820 2161.370 10.420 2161.450 ;
        RECT 8.380 2161.050 8.640 2161.370 ;
        RECT 9.760 2161.310 10.420 2161.370 ;
        RECT 9.760 2161.050 10.020 2161.310 ;
        RECT 8.440 2127.450 8.580 2161.050 ;
        RECT 8.440 2127.310 9.040 2127.450 ;
        RECT 8.900 2074.410 9.040 2127.310 ;
        RECT 8.900 2074.270 10.420 2074.410 ;
        RECT 10.280 2012.530 10.420 2074.270 ;
        RECT 8.900 2012.390 10.420 2012.530 ;
        RECT 8.900 1992.810 9.040 2012.390 ;
        RECT 8.900 1992.670 10.420 1992.810 ;
        RECT 10.280 1936.370 10.420 1992.670 ;
        RECT 9.820 1936.290 10.420 1936.370 ;
        RECT 9.760 1936.230 10.420 1936.290 ;
        RECT 9.760 1935.970 10.020 1936.230 ;
        RECT 9.760 1903.560 10.020 1903.650 ;
        RECT 9.760 1903.420 11.800 1903.560 ;
        RECT 9.760 1903.330 10.020 1903.420 ;
        RECT 11.660 1896.250 11.800 1903.420 ;
        RECT 11.660 1896.110 12.260 1896.250 ;
        RECT 12.120 1876.530 12.260 1896.110 ;
        RECT 11.660 1876.390 12.260 1876.530 ;
        RECT 11.660 1851.880 11.800 1876.390 ;
        RECT 11.660 1851.740 12.260 1851.880 ;
        RECT 12.120 1850.010 12.260 1851.740 ;
        RECT 9.820 1849.870 12.260 1850.010 ;
        RECT 9.820 1846.530 9.960 1849.870 ;
        RECT 9.760 1846.210 10.020 1846.530 ;
        RECT 8.840 1790.110 9.100 1790.430 ;
        RECT 8.900 1765.610 9.040 1790.110 ;
        RECT 8.840 1765.290 9.100 1765.610 ;
        RECT 9.760 1765.520 10.020 1765.610 ;
        RECT 9.760 1765.380 10.420 1765.520 ;
        RECT 9.760 1765.290 10.020 1765.380 ;
        RECT 10.280 1765.010 10.420 1765.380 ;
        RECT 10.280 1764.870 10.880 1765.010 ;
        RECT 10.740 1703.810 10.880 1764.870 ;
        RECT 9.820 1703.730 10.880 1703.810 ;
        RECT 9.760 1703.670 10.880 1703.730 ;
        RECT 9.760 1703.410 10.020 1703.670 ;
        RECT 9.760 1549.050 10.020 1549.370 ;
        RECT 9.820 1548.770 9.960 1549.050 ;
        RECT 9.820 1548.630 10.420 1548.770 ;
        RECT 9.760 1528.200 10.020 1528.290 ;
        RECT 10.280 1528.200 10.420 1548.630 ;
        RECT 9.760 1528.060 10.420 1528.200 ;
        RECT 9.760 1527.970 10.020 1528.060 ;
        RECT 9.760 1507.230 10.020 1507.550 ;
        RECT 9.820 1480.690 9.960 1507.230 ;
        RECT 9.760 1480.370 10.020 1480.690 ;
        RECT 9.760 1416.850 10.020 1417.110 ;
        RECT 9.760 1416.790 10.420 1416.850 ;
        RECT 9.820 1416.710 10.420 1416.790 ;
        RECT 10.280 1351.570 10.420 1416.710 ;
        RECT 10.280 1351.430 11.800 1351.570 ;
        RECT 11.660 1323.690 11.800 1351.430 ;
        RECT 9.820 1323.610 11.800 1323.690 ;
        RECT 9.760 1323.550 11.800 1323.610 ;
        RECT 9.760 1323.290 10.020 1323.550 ;
        RECT 9.760 1250.530 10.020 1250.850 ;
        RECT 9.820 1245.490 9.960 1250.530 ;
        RECT 9.820 1245.350 10.420 1245.490 ;
        RECT 10.280 1211.490 10.420 1245.350 ;
        RECT 9.820 1211.410 10.420 1211.490 ;
        RECT 9.760 1211.350 10.420 1211.410 ;
        RECT 9.760 1211.090 10.020 1211.350 ;
        RECT 7.000 1106.370 7.260 1106.690 ;
        RECT 7.060 1087.310 7.200 1106.370 ;
        RECT 7.000 1086.990 7.260 1087.310 ;
        RECT 9.300 895.230 9.560 895.550 ;
        RECT 9.360 885.010 9.500 895.230 ;
        RECT 9.300 884.690 9.560 885.010 ;
        RECT 9.300 864.970 9.560 865.290 ;
        RECT 9.360 844.970 9.500 864.970 ;
        RECT 9.360 844.830 10.420 844.970 ;
        RECT 9.760 840.040 10.020 840.130 ;
        RECT 10.280 840.040 10.420 844.830 ;
        RECT 9.760 839.900 10.420 840.040 ;
        RECT 9.760 839.810 10.020 839.900 ;
        RECT 9.760 734.750 10.020 735.070 ;
        RECT 9.820 729.290 9.960 734.750 ;
        RECT 9.760 728.970 10.020 729.290 ;
        RECT 9.760 727.950 10.020 728.270 ;
        RECT 9.820 706.850 9.960 727.950 ;
        RECT 9.760 706.530 10.020 706.850 ;
        RECT 9.760 689.530 10.020 689.850 ;
        RECT 9.820 672.510 9.960 689.530 ;
        RECT 9.760 672.190 10.020 672.510 ;
        RECT 9.760 541.860 10.020 541.950 ;
        RECT 9.760 541.720 13.640 541.860 ;
        RECT 9.760 541.630 10.020 541.720 ;
        RECT 9.760 468.080 10.020 468.170 ;
        RECT 13.500 468.080 13.640 541.720 ;
        RECT 9.760 467.940 13.640 468.080 ;
        RECT 9.760 467.850 10.020 467.940 ;
        RECT 9.760 458.900 10.020 458.990 ;
        RECT 9.760 458.760 13.640 458.900 ;
        RECT 9.760 458.670 10.020 458.760 ;
        RECT 9.760 419.120 10.020 419.210 ;
        RECT 13.500 419.120 13.640 458.760 ;
        RECT 9.760 418.980 13.640 419.120 ;
        RECT 9.760 418.890 10.020 418.980 ;
        RECT 9.760 403.590 10.020 403.910 ;
        RECT 9.820 361.070 9.960 403.590 ;
        RECT 6.540 360.750 6.800 361.070 ;
        RECT 9.760 360.750 10.020 361.070 ;
        RECT 6.600 346.790 6.740 360.750 ;
        RECT 6.540 346.470 6.800 346.790 ;
        RECT 9.760 315.080 10.020 315.170 ;
        RECT 9.760 314.940 12.260 315.080 ;
        RECT 9.760 314.850 10.020 314.940 ;
        RECT 9.760 283.800 10.020 283.890 ;
        RECT 9.760 283.660 10.420 283.800 ;
        RECT 9.760 283.570 10.020 283.660 ;
        RECT 10.280 283.290 10.420 283.660 ;
        RECT 12.120 283.290 12.260 314.940 ;
        RECT 10.280 283.150 12.260 283.290 ;
        RECT 9.760 275.810 10.020 276.070 ;
        RECT 9.760 275.750 12.260 275.810 ;
        RECT 9.820 275.670 12.260 275.750 ;
        RECT 12.120 217.330 12.260 275.670 ;
        RECT 12.120 217.190 12.720 217.330 ;
        RECT 12.580 216.650 12.720 217.190 ;
        RECT 12.580 216.510 13.640 216.650 ;
        RECT 13.500 176.530 13.640 216.510 ;
        RECT 9.820 176.450 13.640 176.530 ;
        RECT 1.940 176.130 2.200 176.450 ;
        RECT 9.760 176.390 13.640 176.450 ;
        RECT 9.760 176.130 10.020 176.390 ;
        RECT 2.000 2.565 2.140 176.130 ;
        RECT 360.670 8.570 360.950 9.000 ;
        RECT 358.960 8.490 360.950 8.570 ;
        RECT 358.900 8.430 360.950 8.490 ;
        RECT 358.900 8.170 359.160 8.430 ;
        RECT 360.670 5.000 360.950 8.430 ;
        RECT 36.900 3.070 37.160 3.390 ;
        RECT 36.960 2.565 37.100 3.070 ;
        RECT 1.930 2.195 2.210 2.565 ;
        RECT 36.890 2.195 37.170 2.565 ;
        RECT 294.960 1.370 295.220 1.690 ;
        RECT 295.020 1.010 295.160 1.370 ;
        RECT 294.960 0.690 295.220 1.010 ;
      LAYER via2 ;
        RECT 2900.850 3373.000 2901.130 3373.280 ;
        RECT 1.930 2.240 2.210 2.520 ;
        RECT 36.890 2.240 37.170 2.520 ;
      LAYER met3 ;
        RECT 2900.825 3373.290 2901.155 3373.305 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2900.825 3372.990 2924.800 3373.290 ;
        RECT 2900.825 3372.975 2901.155 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
        RECT 1.905 2.530 2.235 2.545 ;
        RECT 36.865 2.530 37.195 2.545 ;
        RECT 1.905 2.230 37.195 2.530 ;
        RECT 1.905 2.215 2.235 2.230 ;
        RECT 36.865 2.215 37.195 2.230 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 54.810 3501.560 55.130 3501.620 ;
        RECT 2798.250 3501.560 2798.570 3501.620 ;
        RECT 54.810 3501.420 2798.570 3501.560 ;
        RECT 54.810 3501.360 55.130 3501.420 ;
        RECT 2798.250 3501.360 2798.570 3501.420 ;
      LAYER via ;
        RECT 54.840 3501.360 55.100 3501.620 ;
        RECT 2798.280 3501.360 2798.540 3501.620 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3501.650 2798.480 3517.600 ;
        RECT 54.840 3501.330 55.100 3501.650 ;
        RECT 2798.280 3501.330 2798.540 3501.650 ;
        RECT 53.850 3404.490 54.130 3405.000 ;
        RECT 54.900 3404.490 55.040 3501.330 ;
        RECT 53.850 3404.350 55.040 3404.490 ;
        RECT 53.850 3401.000 54.130 3404.350 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 158.310 3501.900 158.630 3501.960 ;
        RECT 2473.950 3501.900 2474.270 3501.960 ;
        RECT 158.310 3501.760 2474.270 3501.900 ;
        RECT 158.310 3501.700 158.630 3501.760 ;
        RECT 2473.950 3501.700 2474.270 3501.760 ;
        RECT 151.870 3422.340 152.190 3422.400 ;
        RECT 158.310 3422.340 158.630 3422.400 ;
        RECT 151.870 3422.200 158.630 3422.340 ;
        RECT 151.870 3422.140 152.190 3422.200 ;
        RECT 158.310 3422.140 158.630 3422.200 ;
      LAYER via ;
        RECT 158.340 3501.700 158.600 3501.960 ;
        RECT 2473.980 3501.700 2474.240 3501.960 ;
        RECT 151.900 3422.140 152.160 3422.400 ;
        RECT 158.340 3422.140 158.600 3422.400 ;
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3501.990 2474.180 3517.600 ;
        RECT 158.340 3501.670 158.600 3501.990 ;
        RECT 2473.980 3501.670 2474.240 3501.990 ;
        RECT 158.400 3422.430 158.540 3501.670 ;
        RECT 151.900 3422.110 152.160 3422.430 ;
        RECT 158.340 3422.110 158.600 3422.430 ;
        RECT 151.960 3405.000 152.100 3422.110 ;
        RECT 151.830 3401.000 152.110 3405.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 254.910 3502.240 255.230 3502.300 ;
        RECT 2149.190 3502.240 2149.510 3502.300 ;
        RECT 254.910 3502.100 2149.510 3502.240 ;
        RECT 254.910 3502.040 255.230 3502.100 ;
        RECT 2149.190 3502.040 2149.510 3502.100 ;
        RECT 250.310 3422.340 250.630 3422.400 ;
        RECT 254.910 3422.340 255.230 3422.400 ;
        RECT 250.310 3422.200 255.230 3422.340 ;
        RECT 250.310 3422.140 250.630 3422.200 ;
        RECT 254.910 3422.140 255.230 3422.200 ;
      LAYER via ;
        RECT 254.940 3502.040 255.200 3502.300 ;
        RECT 2149.220 3502.040 2149.480 3502.300 ;
        RECT 250.340 3422.140 250.600 3422.400 ;
        RECT 254.940 3422.140 255.200 3422.400 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3502.330 2149.420 3517.600 ;
        RECT 254.940 3502.010 255.200 3502.330 ;
        RECT 2149.220 3502.010 2149.480 3502.330 ;
        RECT 255.000 3422.430 255.140 3502.010 ;
        RECT 250.340 3422.110 250.600 3422.430 ;
        RECT 254.940 3422.110 255.200 3422.430 ;
        RECT 250.400 3405.000 250.540 3422.110 ;
        RECT 250.270 3401.000 250.550 3405.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 351.510 3502.580 351.830 3502.640 ;
        RECT 1824.890 3502.580 1825.210 3502.640 ;
        RECT 351.510 3502.440 1825.210 3502.580 ;
        RECT 351.510 3502.380 351.830 3502.440 ;
        RECT 1824.890 3502.380 1825.210 3502.440 ;
      LAYER via ;
        RECT 351.540 3502.380 351.800 3502.640 ;
        RECT 1824.920 3502.380 1825.180 3502.640 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3502.670 1825.120 3517.600 ;
        RECT 351.540 3502.350 351.800 3502.670 ;
        RECT 1824.920 3502.350 1825.180 3502.670 ;
        RECT 348.250 3403.810 348.530 3405.000 ;
        RECT 351.600 3403.810 351.740 3502.350 ;
        RECT 348.250 3403.670 351.740 3403.810 ;
        RECT 348.250 3401.000 348.530 3403.670 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 448.110 3502.920 448.430 3502.980 ;
        RECT 1500.590 3502.920 1500.910 3502.980 ;
        RECT 448.110 3502.780 1500.910 3502.920 ;
        RECT 448.110 3502.720 448.430 3502.780 ;
        RECT 1500.590 3502.720 1500.910 3502.780 ;
      LAYER via ;
        RECT 448.140 3502.720 448.400 3502.980 ;
        RECT 1500.620 3502.720 1500.880 3502.980 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3503.010 1500.820 3517.600 ;
        RECT 448.140 3502.690 448.400 3503.010 ;
        RECT 1500.620 3502.690 1500.880 3503.010 ;
        RECT 446.690 3404.490 446.970 3405.000 ;
        RECT 448.200 3404.490 448.340 3502.690 ;
        RECT 446.690 3404.350 448.340 3404.490 ;
        RECT 446.690 3401.000 446.970 3404.350 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2873.690 317.800 2874.010 317.860 ;
        RECT 2900.830 317.800 2901.150 317.860 ;
        RECT 2873.690 317.660 2901.150 317.800 ;
        RECT 2873.690 317.600 2874.010 317.660 ;
        RECT 2900.830 317.600 2901.150 317.660 ;
      LAYER via ;
        RECT 2873.720 317.600 2873.980 317.860 ;
        RECT 2900.860 317.600 2901.120 317.860 ;
      LAYER met2 ;
        RECT 2900.850 322.475 2901.130 322.845 ;
        RECT 2900.920 317.890 2901.060 322.475 ;
        RECT 2873.720 317.570 2873.980 317.890 ;
        RECT 2900.860 317.570 2901.120 317.890 ;
        RECT 2873.780 209.285 2873.920 317.570 ;
        RECT 2873.710 208.915 2873.990 209.285 ;
      LAYER via2 ;
        RECT 2900.850 322.520 2901.130 322.800 ;
        RECT 2873.710 208.960 2873.990 209.240 ;
      LAYER met3 ;
        RECT 2900.825 322.810 2901.155 322.825 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2900.825 322.510 2924.800 322.810 ;
        RECT 2900.825 322.495 2901.155 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
        RECT 2851.000 209.250 2855.000 209.640 ;
        RECT 2873.685 209.250 2874.015 209.265 ;
        RECT 2851.000 209.040 2874.015 209.250 ;
        RECT 2854.300 208.950 2874.015 209.040 ;
        RECT 2873.685 208.935 2874.015 208.950 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 551.610 3503.260 551.930 3503.320 ;
        RECT 1175.830 3503.260 1176.150 3503.320 ;
        RECT 551.610 3503.120 1176.150 3503.260 ;
        RECT 551.610 3503.060 551.930 3503.120 ;
        RECT 1175.830 3503.060 1176.150 3503.120 ;
        RECT 545.170 3420.300 545.490 3420.360 ;
        RECT 551.610 3420.300 551.930 3420.360 ;
        RECT 545.170 3420.160 551.930 3420.300 ;
        RECT 545.170 3420.100 545.490 3420.160 ;
        RECT 551.610 3420.100 551.930 3420.160 ;
      LAYER via ;
        RECT 551.640 3503.060 551.900 3503.320 ;
        RECT 1175.860 3503.060 1176.120 3503.320 ;
        RECT 545.200 3420.100 545.460 3420.360 ;
        RECT 551.640 3420.100 551.900 3420.360 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3503.350 1176.060 3517.600 ;
        RECT 551.640 3503.030 551.900 3503.350 ;
        RECT 1175.860 3503.030 1176.120 3503.350 ;
        RECT 551.700 3420.390 551.840 3503.030 ;
        RECT 545.200 3420.070 545.460 3420.390 ;
        RECT 551.640 3420.070 551.900 3420.390 ;
        RECT 545.260 3405.000 545.400 3420.070 ;
        RECT 545.130 3401.000 545.410 3405.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 648.210 3503.600 648.530 3503.660 ;
        RECT 851.530 3503.600 851.850 3503.660 ;
        RECT 648.210 3503.460 851.850 3503.600 ;
        RECT 648.210 3503.400 648.530 3503.460 ;
        RECT 851.530 3503.400 851.850 3503.460 ;
        RECT 643.150 3422.340 643.470 3422.400 ;
        RECT 648.210 3422.340 648.530 3422.400 ;
        RECT 643.150 3422.200 648.530 3422.340 ;
        RECT 643.150 3422.140 643.470 3422.200 ;
        RECT 648.210 3422.140 648.530 3422.200 ;
      LAYER via ;
        RECT 648.240 3503.400 648.500 3503.660 ;
        RECT 851.560 3503.400 851.820 3503.660 ;
        RECT 643.180 3422.140 643.440 3422.400 ;
        RECT 648.240 3422.140 648.500 3422.400 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3503.690 851.760 3517.600 ;
        RECT 648.240 3503.370 648.500 3503.690 ;
        RECT 851.560 3503.370 851.820 3503.690 ;
        RECT 648.300 3422.430 648.440 3503.370 ;
        RECT 643.180 3422.110 643.440 3422.430 ;
        RECT 648.240 3422.110 648.500 3422.430 ;
        RECT 643.240 3405.000 643.380 3422.110 ;
        RECT 643.110 3401.000 643.390 3405.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 527.230 3503.260 527.550 3503.320 ;
        RECT 530.910 3503.260 531.230 3503.320 ;
        RECT 527.230 3503.120 531.230 3503.260 ;
        RECT 527.230 3503.060 527.550 3503.120 ;
        RECT 530.910 3503.060 531.230 3503.120 ;
        RECT 530.910 3419.280 531.230 3419.340 ;
        RECT 741.590 3419.280 741.910 3419.340 ;
        RECT 530.910 3419.140 741.910 3419.280 ;
        RECT 530.910 3419.080 531.230 3419.140 ;
        RECT 741.590 3419.080 741.910 3419.140 ;
      LAYER via ;
        RECT 527.260 3503.060 527.520 3503.320 ;
        RECT 530.940 3503.060 531.200 3503.320 ;
        RECT 530.940 3419.080 531.200 3419.340 ;
        RECT 741.620 3419.080 741.880 3419.340 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3503.350 527.460 3517.600 ;
        RECT 527.260 3503.030 527.520 3503.350 ;
        RECT 530.940 3503.030 531.200 3503.350 ;
        RECT 531.000 3419.370 531.140 3503.030 ;
        RECT 530.940 3419.050 531.200 3419.370 ;
        RECT 741.620 3419.050 741.880 3419.370 ;
        RECT 741.680 3405.000 741.820 3419.050 ;
        RECT 741.550 3401.000 741.830 3405.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 202.470 3502.580 202.790 3502.640 ;
        RECT 206.610 3502.580 206.930 3502.640 ;
        RECT 202.470 3502.440 206.930 3502.580 ;
        RECT 202.470 3502.380 202.790 3502.440 ;
        RECT 206.610 3502.380 206.930 3502.440 ;
        RECT 206.610 3418.940 206.930 3419.000 ;
        RECT 840.030 3418.940 840.350 3419.000 ;
        RECT 206.610 3418.800 840.350 3418.940 ;
        RECT 206.610 3418.740 206.930 3418.800 ;
        RECT 840.030 3418.740 840.350 3418.800 ;
      LAYER via ;
        RECT 202.500 3502.380 202.760 3502.640 ;
        RECT 206.640 3502.380 206.900 3502.640 ;
        RECT 206.640 3418.740 206.900 3419.000 ;
        RECT 840.060 3418.740 840.320 3419.000 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3502.670 202.700 3517.600 ;
        RECT 202.500 3502.350 202.760 3502.670 ;
        RECT 206.640 3502.350 206.900 3502.670 ;
        RECT 206.700 3419.030 206.840 3502.350 ;
        RECT 206.640 3418.710 206.900 3419.030 ;
        RECT 840.060 3418.710 840.320 3419.030 ;
        RECT 840.120 3405.000 840.260 3418.710 ;
        RECT 839.990 3401.000 840.270 3405.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1.065 829.345 1.235 873.035 ;
        RECT 1.985 734.825 2.155 769.335 ;
        RECT 6.585 7.565 6.755 59.415 ;
        RECT 25.445 8.925 27.455 9.095 ;
        RECT 25.445 7.565 25.615 8.925 ;
        RECT 27.285 8.245 27.455 8.925 ;
      LAYER mcon ;
        RECT 1.065 872.865 1.235 873.035 ;
        RECT 1.985 769.165 2.155 769.335 ;
        RECT 6.585 59.245 6.755 59.415 ;
      LAYER met1 ;
        RECT 0.990 3387.660 1.310 3387.720 ;
        RECT 6.970 3387.660 7.290 3387.720 ;
        RECT 0.990 3387.520 7.290 3387.660 ;
        RECT 0.990 3387.460 1.310 3387.520 ;
        RECT 6.970 3387.460 7.290 3387.520 ;
        RECT 0.990 873.020 1.310 873.080 ;
        RECT 0.795 872.880 1.310 873.020 ;
        RECT 0.990 872.820 1.310 872.880 ;
        RECT 1.005 829.500 1.295 829.545 ;
        RECT 1.910 829.500 2.230 829.560 ;
        RECT 1.005 829.360 2.230 829.500 ;
        RECT 1.005 829.315 1.295 829.360 ;
        RECT 1.910 829.300 2.230 829.360 ;
        RECT 1.910 769.320 2.230 769.380 ;
        RECT 1.715 769.180 2.230 769.320 ;
        RECT 1.910 769.120 2.230 769.180 ;
        RECT 1.910 734.980 2.230 735.040 ;
        RECT 1.715 734.840 2.230 734.980 ;
        RECT 1.910 734.780 2.230 734.840 ;
        RECT 1.910 631.620 2.230 631.680 ;
        RECT 4.210 631.620 4.530 631.680 ;
        RECT 1.910 631.480 4.530 631.620 ;
        RECT 1.910 631.420 2.230 631.480 ;
        RECT 4.210 631.420 4.530 631.480 ;
        RECT 4.210 59.400 4.530 59.460 ;
        RECT 6.525 59.400 6.815 59.445 ;
        RECT 4.210 59.260 6.815 59.400 ;
        RECT 4.210 59.200 4.530 59.260 ;
        RECT 6.525 59.215 6.815 59.260 ;
        RECT 27.210 8.400 27.530 8.460 ;
        RECT 27.015 8.260 27.530 8.400 ;
        RECT 27.210 8.200 27.530 8.260 ;
        RECT 6.525 7.720 6.815 7.765 ;
        RECT 25.385 7.720 25.675 7.765 ;
        RECT 6.525 7.580 25.675 7.720 ;
        RECT 6.525 7.535 6.815 7.580 ;
        RECT 25.385 7.535 25.675 7.580 ;
      LAYER via ;
        RECT 1.020 3387.460 1.280 3387.720 ;
        RECT 7.000 3387.460 7.260 3387.720 ;
        RECT 1.020 872.820 1.280 873.080 ;
        RECT 1.940 829.300 2.200 829.560 ;
        RECT 1.940 769.120 2.200 769.380 ;
        RECT 1.940 734.780 2.200 735.040 ;
        RECT 1.940 631.420 2.200 631.680 ;
        RECT 4.240 631.420 4.500 631.680 ;
        RECT 4.240 59.200 4.500 59.460 ;
        RECT 27.240 8.200 27.500 8.460 ;
      LAYER met2 ;
        RECT 6.990 3411.035 7.270 3411.405 ;
        RECT 7.060 3387.750 7.200 3411.035 ;
        RECT 1.020 3387.430 1.280 3387.750 ;
        RECT 7.000 3387.430 7.260 3387.750 ;
        RECT 1.080 873.110 1.220 3387.430 ;
        RECT 1.020 872.790 1.280 873.110 ;
        RECT 1.940 829.270 2.200 829.590 ;
        RECT 2.000 769.410 2.140 829.270 ;
        RECT 1.940 769.090 2.200 769.410 ;
        RECT 1.940 734.750 2.200 735.070 ;
        RECT 2.000 631.710 2.140 734.750 ;
        RECT 1.940 631.390 2.200 631.710 ;
        RECT 4.240 631.390 4.500 631.710 ;
        RECT 4.300 59.490 4.440 631.390 ;
        RECT 4.240 59.170 4.500 59.490 ;
        RECT 28.550 8.570 28.830 9.000 ;
        RECT 27.300 8.490 28.830 8.570 ;
        RECT 27.240 8.430 28.830 8.490 ;
        RECT 27.240 8.170 27.500 8.430 ;
        RECT 28.550 5.000 28.830 8.430 ;
      LAYER via2 ;
        RECT 6.990 3411.080 7.270 3411.360 ;
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 6.965 3411.370 7.295 3411.385 ;
        RECT -4.800 3411.070 7.295 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 6.965 3411.055 7.295 3411.070 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 7.965 1416.185 8.135 1435.055 ;
        RECT 8.425 1350.905 8.595 1369.775 ;
        RECT 7.505 797.385 7.675 817.955 ;
        RECT 9.345 817.785 9.515 880.515 ;
        RECT 8.425 743.495 8.595 797.555 ;
        RECT 7.965 743.325 8.595 743.495 ;
        RECT 7.965 729.725 8.135 743.325 ;
        RECT 8.425 5.525 8.595 51.255 ;
      LAYER mcon ;
        RECT 7.965 1434.885 8.135 1435.055 ;
        RECT 8.425 1369.605 8.595 1369.775 ;
        RECT 9.345 880.345 9.515 880.515 ;
        RECT 7.505 817.785 7.675 817.955 ;
        RECT 8.425 797.385 8.595 797.555 ;
        RECT 8.425 51.085 8.595 51.255 ;
      LAYER met1 ;
        RECT 0.070 1435.040 0.390 1435.100 ;
        RECT 7.905 1435.040 8.195 1435.085 ;
        RECT 0.070 1434.900 8.195 1435.040 ;
        RECT 0.070 1434.840 0.390 1434.900 ;
        RECT 7.905 1434.855 8.195 1434.900 ;
        RECT 7.905 1416.340 8.195 1416.385 ;
        RECT 9.730 1416.340 10.050 1416.400 ;
        RECT 7.905 1416.200 10.050 1416.340 ;
        RECT 7.905 1416.155 8.195 1416.200 ;
        RECT 9.730 1416.140 10.050 1416.200 ;
        RECT 8.365 1369.760 8.655 1369.805 ;
        RECT 9.730 1369.760 10.050 1369.820 ;
        RECT 8.365 1369.620 10.050 1369.760 ;
        RECT 8.365 1369.575 8.655 1369.620 ;
        RECT 9.730 1369.560 10.050 1369.620 ;
        RECT 8.365 1351.060 8.655 1351.105 ;
        RECT 9.730 1351.060 10.050 1351.120 ;
        RECT 8.365 1350.920 10.050 1351.060 ;
        RECT 8.365 1350.875 8.655 1350.920 ;
        RECT 9.730 1350.860 10.050 1350.920 ;
        RECT 1.450 1331.680 1.770 1331.740 ;
        RECT 9.730 1331.680 10.050 1331.740 ;
        RECT 1.450 1331.540 10.050 1331.680 ;
        RECT 1.450 1331.480 1.770 1331.540 ;
        RECT 9.730 1331.480 10.050 1331.540 ;
        RECT 1.910 880.500 2.230 880.560 ;
        RECT 9.285 880.500 9.575 880.545 ;
        RECT 1.910 880.360 9.575 880.500 ;
        RECT 1.910 880.300 2.230 880.360 ;
        RECT 9.285 880.315 9.575 880.360 ;
        RECT 7.445 817.940 7.735 817.985 ;
        RECT 9.285 817.940 9.575 817.985 ;
        RECT 7.445 817.800 9.575 817.940 ;
        RECT 7.445 817.755 7.735 817.800 ;
        RECT 9.285 817.755 9.575 817.800 ;
        RECT 7.445 797.540 7.735 797.585 ;
        RECT 8.365 797.540 8.655 797.585 ;
        RECT 7.445 797.400 8.655 797.540 ;
        RECT 7.445 797.355 7.735 797.400 ;
        RECT 8.365 797.355 8.655 797.400 ;
        RECT 6.050 729.880 6.370 729.940 ;
        RECT 7.905 729.880 8.195 729.925 ;
        RECT 6.050 729.740 8.195 729.880 ;
        RECT 6.050 729.680 6.370 729.740 ;
        RECT 7.905 729.695 8.195 729.740 ;
        RECT 4.670 605.440 4.990 605.500 ;
        RECT 6.050 605.440 6.370 605.500 ;
        RECT 4.670 605.300 6.370 605.440 ;
        RECT 4.670 605.240 4.990 605.300 ;
        RECT 6.050 605.240 6.370 605.300 ;
        RECT 4.670 51.240 4.990 51.300 ;
        RECT 8.365 51.240 8.655 51.285 ;
        RECT 4.670 51.100 8.655 51.240 ;
        RECT 4.670 51.040 4.990 51.100 ;
        RECT 8.365 51.055 8.655 51.100 ;
        RECT 8.365 5.680 8.655 5.725 ;
        RECT 24.910 5.680 25.230 5.740 ;
        RECT 8.365 5.540 25.230 5.680 ;
        RECT 8.365 5.495 8.655 5.540 ;
        RECT 24.910 5.480 25.230 5.540 ;
        RECT 66.310 3.640 66.630 3.700 ;
        RECT 75.970 3.640 76.290 3.700 ;
        RECT 66.310 3.500 76.290 3.640 ;
        RECT 66.310 3.440 66.630 3.500 ;
        RECT 75.970 3.440 76.290 3.500 ;
      LAYER via ;
        RECT 0.100 1434.840 0.360 1435.100 ;
        RECT 9.760 1416.140 10.020 1416.400 ;
        RECT 9.760 1369.560 10.020 1369.820 ;
        RECT 9.760 1350.860 10.020 1351.120 ;
        RECT 1.480 1331.480 1.740 1331.740 ;
        RECT 9.760 1331.480 10.020 1331.740 ;
        RECT 1.940 880.300 2.200 880.560 ;
        RECT 6.080 729.680 6.340 729.940 ;
        RECT 4.700 605.240 4.960 605.500 ;
        RECT 6.080 605.240 6.340 605.500 ;
        RECT 4.700 51.040 4.960 51.300 ;
        RECT 24.940 5.480 25.200 5.740 ;
        RECT 66.340 3.440 66.600 3.700 ;
        RECT 76.000 3.440 76.260 3.700 ;
      LAYER met2 ;
        RECT 0.090 3122.715 0.370 3123.085 ;
        RECT 0.160 1435.130 0.300 3122.715 ;
        RECT 0.100 1434.810 0.360 1435.130 ;
        RECT 9.760 1416.110 10.020 1416.430 ;
        RECT 9.820 1369.850 9.960 1416.110 ;
        RECT 9.760 1369.530 10.020 1369.850 ;
        RECT 9.760 1350.890 10.020 1351.150 ;
        RECT 9.760 1350.830 11.340 1350.890 ;
        RECT 9.820 1350.750 11.340 1350.830 ;
        RECT 1.480 1331.450 1.740 1331.770 ;
        RECT 9.760 1331.680 10.020 1331.770 ;
        RECT 11.200 1331.680 11.340 1350.750 ;
        RECT 9.760 1331.540 11.340 1331.680 ;
        RECT 9.760 1331.450 10.020 1331.540 ;
        RECT 1.540 1106.090 1.680 1331.450 ;
        RECT 1.540 1105.950 2.140 1106.090 ;
        RECT 2.000 880.590 2.140 1105.950 ;
        RECT 1.940 880.270 2.200 880.590 ;
        RECT 6.080 729.650 6.340 729.970 ;
        RECT 6.140 605.530 6.280 729.650 ;
        RECT 4.700 605.210 4.960 605.530 ;
        RECT 6.080 605.210 6.340 605.530 ;
        RECT 4.760 51.330 4.900 605.210 ;
        RECT 4.700 51.010 4.960 51.330 ;
        RECT 25.000 5.770 28.360 5.850 ;
        RECT 24.940 5.710 28.360 5.770 ;
        RECT 24.940 5.450 25.200 5.710 ;
        RECT 28.220 4.490 28.360 5.710 ;
        RECT 75.930 5.000 76.210 9.000 ;
        RECT 27.760 4.350 28.360 4.490 ;
        RECT 27.760 3.130 27.900 4.350 ;
        RECT 76.060 3.730 76.200 5.000 ;
        RECT 66.340 3.410 66.600 3.730 ;
        RECT 76.000 3.410 76.260 3.730 ;
        RECT 66.400 3.245 66.540 3.410 ;
        RECT 28.150 3.130 28.430 3.245 ;
        RECT 27.760 2.990 28.430 3.130 ;
        RECT 28.150 2.875 28.430 2.990 ;
        RECT 66.330 2.875 66.610 3.245 ;
      LAYER via2 ;
        RECT 0.090 3122.760 0.370 3123.040 ;
        RECT 28.150 2.920 28.430 3.200 ;
        RECT 66.330 2.920 66.610 3.200 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT -4.800 3124.110 3.370 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 0.065 3123.050 0.395 3123.065 ;
        RECT 3.070 3123.050 3.370 3124.110 ;
        RECT 0.065 3122.750 3.370 3123.050 ;
        RECT 0.065 3122.735 0.395 3122.750 ;
        RECT 28.125 3.210 28.455 3.225 ;
        RECT 66.305 3.210 66.635 3.225 ;
        RECT 28.125 2.910 66.635 3.210 ;
        RECT 28.125 2.895 28.455 2.910 ;
        RECT 66.305 2.895 66.635 2.910 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1035.145 3395.665 1035.315 3401.615 ;
        RECT 1082.985 3398.725 1083.155 3401.955 ;
        RECT 2718.745 3398.725 2718.915 3401.955 ;
        RECT 2807.985 3399.405 2808.155 3401.615 ;
        RECT 8.425 3002.625 8.595 3005.515 ;
        RECT 9.805 2999.225 9.975 3010.615 ;
        RECT 8.425 2816.985 8.595 2822.255 ;
        RECT 8.425 2630.665 8.595 2632.535 ;
        RECT 7.505 2510.985 7.675 2535.975 ;
        RECT 8.885 2524.245 9.055 2530.535 ;
        RECT 7.045 2239.665 7.215 2249.695 ;
        RECT 7.965 2242.385 8.135 2243.915 ;
        RECT 7.045 1667.105 7.215 1671.015 ;
        RECT 8.885 1659.965 9.055 1670.335 ;
        RECT 6.125 1520.565 6.295 1560.855 ;
        RECT 6.585 1558.985 6.755 1575.815 ;
        RECT 7.045 1560.685 7.215 1561.535 ;
        RECT 5.665 1472.285 5.835 1490.475 ;
        RECT 6.125 1465.485 6.295 1516.995 ;
        RECT 6.585 1490.305 6.755 1522.775 ;
        RECT 7.045 1519.885 7.215 1560.175 ;
        RECT 7.505 1542.155 7.675 1562.215 ;
        RECT 7.505 1541.985 8.135 1542.155 ;
        RECT 6.585 1460.725 6.755 1480.275 ;
        RECT 7.965 1480.105 8.135 1541.985 ;
        RECT 6.585 1422.985 6.755 1435.735 ;
        RECT 7.045 1423.665 7.215 1467.015 ;
        RECT 7.505 1435.565 7.675 1472.455 ;
        RECT 7.965 1435.395 8.135 1460.895 ;
        RECT 7.505 1435.225 8.135 1435.395 ;
        RECT 7.505 1421.625 7.675 1435.225 ;
        RECT 7.045 1417.205 7.215 1419.755 ;
        RECT 9.345 1332.715 9.515 1417.375 ;
        RECT 8.885 1332.545 9.515 1332.715 ;
        RECT 8.885 1320.645 9.055 1332.545 ;
        RECT 3.365 969.765 3.535 1009.375 ;
        RECT 5.205 1004.615 5.375 1024.675 ;
        RECT 4.745 1004.445 5.375 1004.615 ;
        RECT 4.745 997.135 4.915 1004.445 ;
        RECT 4.285 996.965 4.915 997.135 ;
        RECT 4.285 980.985 4.455 996.965 ;
        RECT 5.665 989.485 5.835 1038.955 ;
        RECT 7.965 1038.785 8.135 1099.815 ;
        RECT 8.885 1088.425 9.055 1091.655 ;
        RECT 5.665 973.505 5.835 988.975 ;
        RECT 6.585 978.945 6.755 989.655 ;
        RECT 9.805 981.665 9.975 988.295 ;
        RECT 7.505 942.565 7.675 948.175 ;
        RECT 7.505 883.745 7.675 942.055 ;
        RECT 6.585 797.045 6.755 836.315 ;
        RECT 7.045 827.305 7.215 832.235 ;
        RECT 4.745 714.085 4.915 734.995 ;
        RECT 6.125 734.825 6.295 768.995 ;
        RECT 8.885 731.765 9.055 797.215 ;
        RECT 1.525 651.185 1.695 694.875 ;
        RECT 2.445 647.105 2.615 652.035 ;
        RECT 2.905 546.465 3.075 653.055 ;
        RECT 3.365 631.125 3.535 660.535 ;
        RECT 3.825 651.865 3.995 706.095 ;
        RECT 8.885 694.705 9.055 699.975 ;
        RECT 3.825 587.265 3.995 651.355 ;
        RECT 4.745 641.665 4.915 672.775 ;
        RECT 9.345 666.485 9.515 714.935 ;
        RECT 7.965 645.745 8.135 654.415 ;
        RECT 4.745 586.925 4.915 631.295 ;
        RECT 5.205 597.805 5.375 632.655 ;
        RECT 7.965 632.485 8.135 644.555 ;
        RECT 5.205 576.045 5.375 587.435 ;
        RECT 3.365 545.785 3.535 547.315 ;
        RECT 3.825 543.745 3.995 548.675 ;
        RECT 4.745 544.425 4.915 575.535 ;
        RECT 5.205 540.345 5.375 555.135 ;
        RECT 7.505 542.385 7.675 576.215 ;
        RECT 7.965 543.065 8.135 631.975 ;
        RECT 8.885 512.805 9.055 597.975 ;
        RECT 6.585 467.585 6.755 491.555 ;
        RECT 4.745 430.525 4.915 460.275 ;
        RECT 6.585 457.385 6.755 467.075 ;
        RECT 4.745 410.465 4.915 423.895 ;
        RECT 5.205 417.945 5.375 438.175 ;
        RECT 7.505 438.005 7.675 467.755 ;
        RECT 3.825 323.085 3.995 333.795 ;
        RECT 4.285 289.425 4.455 333.115 ;
        RECT 4.745 315.605 4.915 336.175 ;
        RECT 5.205 314.245 5.375 337.535 ;
        RECT 7.965 331.415 8.135 359.975 ;
        RECT 7.505 331.245 8.135 331.415 ;
        RECT 5.665 311.185 5.835 327.335 ;
        RECT 6.125 279.225 6.295 285.515 ;
        RECT 7.505 262.905 7.675 331.245 ;
        RECT 5.205 185.045 5.375 251.855 ;
        RECT 6.125 136.595 6.295 177.735 ;
        RECT 5.665 136.425 6.295 136.595 ;
        RECT 3.365 50.405 3.535 82.875 ;
        RECT 4.745 37.485 4.915 100.215 ;
        RECT 5.205 72.845 5.375 89.675 ;
        RECT 5.665 75.905 5.835 136.425 ;
        RECT 6.125 76.585 6.295 136.255 ;
        RECT 7.045 110.925 7.215 141.695 ;
        RECT 7.505 135.405 7.675 147.475 ;
        RECT 9.805 94.265 9.975 148.835 ;
        RECT 5.665 72.675 5.835 74.035 ;
        RECT 5.205 72.505 5.835 72.675 ;
        RECT 5.205 66.725 5.375 72.505 ;
        RECT 5.665 6.545 5.835 72.335 ;
        RECT 6.125 16.405 6.295 67.575 ;
        RECT 6.585 61.625 6.755 82.195 ;
        RECT 8.885 0.085 9.055 61.115 ;
        RECT 283.965 8.245 284.135 9.095 ;
        RECT 26.365 3.485 26.535 5.355 ;
        RECT 36.485 3.145 36.655 7.055 ;
        RECT 52.125 5.525 52.295 6.375 ;
        RECT 52.585 5.525 52.755 7.055 ;
        RECT 55.345 6.035 55.515 6.375 ;
        RECT 56.265 6.035 56.435 8.075 ;
        RECT 141.365 6.205 141.535 7.735 ;
        RECT 55.345 5.865 56.435 6.035 ;
        RECT 212.205 4.165 212.375 8.075 ;
        RECT 327.205 7.055 327.375 9.095 ;
        RECT 507.985 8.245 511.375 8.415 ;
        RECT 334.105 7.905 335.655 8.075 ;
        RECT 334.105 7.735 334.275 7.905 ;
        RECT 333.645 7.565 334.275 7.735 ;
        RECT 328.125 7.055 328.295 7.395 ;
        RECT 333.645 7.225 333.815 7.565 ;
        RECT 327.205 6.885 328.295 7.055 ;
        RECT 335.485 6.545 335.655 7.905 ;
        RECT 507.985 7.225 508.155 8.245 ;
        RECT 511.205 8.075 511.375 8.245 ;
        RECT 511.205 7.905 518.735 8.075 ;
        RECT 462.905 6.885 465.375 7.055 ;
        RECT 364.005 5.695 364.175 6.715 ;
        RECT 364.005 5.525 365.555 5.695 ;
        RECT 365.385 5.185 365.555 5.525 ;
        RECT 417.825 5.355 417.995 6.715 ;
        RECT 417.365 5.185 417.995 5.355 ;
        RECT 422.885 6.205 428.575 6.375 ;
        RECT 417.365 4.845 417.535 5.185 ;
        RECT 23.605 2.805 26.075 2.975 ;
        RECT 23.605 2.125 23.775 2.805 ;
        RECT 30.045 1.105 30.215 2.635 ;
        RECT 422.885 0.765 423.055 6.205 ;
        RECT 428.405 0.595 428.575 6.205 ;
        RECT 518.565 5.525 518.735 7.905 ;
        RECT 448.185 0.595 448.355 1.955 ;
        RECT 27.285 0.425 28.375 0.595 ;
        RECT 428.405 0.425 448.355 0.595 ;
      LAYER mcon ;
        RECT 1082.985 3401.785 1083.155 3401.955 ;
        RECT 1035.145 3401.445 1035.315 3401.615 ;
        RECT 2718.745 3401.785 2718.915 3401.955 ;
        RECT 2807.985 3401.445 2808.155 3401.615 ;
        RECT 9.805 3010.445 9.975 3010.615 ;
        RECT 8.425 3005.345 8.595 3005.515 ;
        RECT 8.425 2822.085 8.595 2822.255 ;
        RECT 8.425 2632.365 8.595 2632.535 ;
        RECT 7.505 2535.805 7.675 2535.975 ;
        RECT 8.885 2530.365 9.055 2530.535 ;
        RECT 7.045 2249.525 7.215 2249.695 ;
        RECT 7.965 2243.745 8.135 2243.915 ;
        RECT 7.045 1670.845 7.215 1671.015 ;
        RECT 8.885 1670.165 9.055 1670.335 ;
        RECT 6.585 1575.645 6.755 1575.815 ;
        RECT 6.125 1560.685 6.295 1560.855 ;
        RECT 7.505 1562.045 7.675 1562.215 ;
        RECT 7.045 1561.365 7.215 1561.535 ;
        RECT 7.045 1560.005 7.215 1560.175 ;
        RECT 6.585 1522.605 6.755 1522.775 ;
        RECT 6.125 1516.825 6.295 1516.995 ;
        RECT 5.665 1490.305 5.835 1490.475 ;
        RECT 6.585 1480.105 6.755 1480.275 ;
        RECT 7.505 1472.285 7.675 1472.455 ;
        RECT 7.045 1466.845 7.215 1467.015 ;
        RECT 6.585 1435.565 6.755 1435.735 ;
        RECT 7.965 1460.725 8.135 1460.895 ;
        RECT 7.045 1419.585 7.215 1419.755 ;
        RECT 9.345 1417.205 9.515 1417.375 ;
        RECT 7.965 1099.645 8.135 1099.815 ;
        RECT 8.885 1091.485 9.055 1091.655 ;
        RECT 5.665 1038.785 5.835 1038.955 ;
        RECT 5.205 1024.505 5.375 1024.675 ;
        RECT 3.365 1009.205 3.535 1009.375 ;
        RECT 6.585 989.485 6.755 989.655 ;
        RECT 5.665 988.805 5.835 988.975 ;
        RECT 9.805 988.125 9.975 988.295 ;
        RECT 7.505 948.005 7.675 948.175 ;
        RECT 7.505 941.885 7.675 942.055 ;
        RECT 6.585 836.145 6.755 836.315 ;
        RECT 7.045 832.065 7.215 832.235 ;
        RECT 8.885 797.045 9.055 797.215 ;
        RECT 6.125 768.825 6.295 768.995 ;
        RECT 4.745 734.825 4.915 734.995 ;
        RECT 9.345 714.765 9.515 714.935 ;
        RECT 3.825 705.925 3.995 706.095 ;
        RECT 1.525 694.705 1.695 694.875 ;
        RECT 3.365 660.365 3.535 660.535 ;
        RECT 2.905 652.885 3.075 653.055 ;
        RECT 2.445 651.865 2.615 652.035 ;
        RECT 8.885 699.805 9.055 699.975 ;
        RECT 4.745 672.605 4.915 672.775 ;
        RECT 3.825 651.185 3.995 651.355 ;
        RECT 7.965 654.245 8.135 654.415 ;
        RECT 7.965 644.385 8.135 644.555 ;
        RECT 5.205 632.485 5.375 632.655 ;
        RECT 4.745 631.125 4.915 631.295 ;
        RECT 7.965 631.805 8.135 631.975 ;
        RECT 5.205 587.265 5.375 587.435 ;
        RECT 7.505 576.045 7.675 576.215 ;
        RECT 4.745 575.365 4.915 575.535 ;
        RECT 3.825 548.505 3.995 548.675 ;
        RECT 3.365 547.145 3.535 547.315 ;
        RECT 5.205 554.965 5.375 555.135 ;
        RECT 8.885 597.805 9.055 597.975 ;
        RECT 6.585 491.385 6.755 491.555 ;
        RECT 7.505 467.585 7.675 467.755 ;
        RECT 6.585 466.905 6.755 467.075 ;
        RECT 4.745 460.105 4.915 460.275 ;
        RECT 5.205 438.005 5.375 438.175 ;
        RECT 4.745 423.725 4.915 423.895 ;
        RECT 7.965 359.805 8.135 359.975 ;
        RECT 5.205 337.365 5.375 337.535 ;
        RECT 4.745 336.005 4.915 336.175 ;
        RECT 3.825 333.625 3.995 333.795 ;
        RECT 4.285 332.945 4.455 333.115 ;
        RECT 5.665 327.165 5.835 327.335 ;
        RECT 6.125 285.345 6.295 285.515 ;
        RECT 5.205 251.685 5.375 251.855 ;
        RECT 6.125 177.565 6.295 177.735 ;
        RECT 9.805 148.665 9.975 148.835 ;
        RECT 7.505 147.305 7.675 147.475 ;
        RECT 7.045 141.525 7.215 141.695 ;
        RECT 4.745 100.045 4.915 100.215 ;
        RECT 3.365 82.705 3.535 82.875 ;
        RECT 5.205 89.505 5.375 89.675 ;
        RECT 6.125 136.085 6.295 136.255 ;
        RECT 6.585 82.025 6.755 82.195 ;
        RECT 5.665 73.865 5.835 74.035 ;
        RECT 5.665 72.165 5.835 72.335 ;
        RECT 6.125 67.405 6.295 67.575 ;
        RECT 8.885 60.945 9.055 61.115 ;
        RECT 283.965 8.925 284.135 9.095 ;
        RECT 327.205 8.925 327.375 9.095 ;
        RECT 56.265 7.905 56.435 8.075 ;
        RECT 36.485 6.885 36.655 7.055 ;
        RECT 26.365 5.185 26.535 5.355 ;
        RECT 52.585 6.885 52.755 7.055 ;
        RECT 52.125 6.205 52.295 6.375 ;
        RECT 55.345 6.205 55.515 6.375 ;
        RECT 212.205 7.905 212.375 8.075 ;
        RECT 141.365 7.565 141.535 7.735 ;
        RECT 328.125 7.225 328.295 7.395 ;
        RECT 465.205 6.885 465.375 7.055 ;
        RECT 364.005 6.545 364.175 6.715 ;
        RECT 417.825 6.545 417.995 6.715 ;
        RECT 25.905 2.805 26.075 2.975 ;
        RECT 30.045 2.465 30.215 2.635 ;
        RECT 448.185 1.785 448.355 1.955 ;
        RECT 28.205 0.425 28.375 0.595 ;
      LAYER met1 ;
        RECT 1082.925 3401.940 1083.215 3401.985 ;
        RECT 1133.510 3401.940 1133.830 3402.000 ;
        RECT 1329.470 3401.940 1329.790 3402.000 ;
        RECT 1082.925 3401.800 1133.830 3401.940 ;
        RECT 1082.925 3401.755 1083.215 3401.800 ;
        RECT 1133.510 3401.740 1133.830 3401.800 ;
        RECT 1269.760 3401.800 1329.790 3401.940 ;
        RECT 1035.070 3401.600 1035.390 3401.660 ;
        RECT 1034.875 3401.460 1035.390 3401.600 ;
        RECT 1035.070 3401.400 1035.390 3401.460 ;
        RECT 17.090 3398.880 17.410 3398.940 ;
        RECT 1082.925 3398.880 1083.215 3398.925 ;
        RECT 17.090 3398.740 1083.215 3398.880 ;
        RECT 17.090 3398.680 17.410 3398.740 ;
        RECT 1082.925 3398.695 1083.215 3398.740 ;
        RECT 12.490 3398.200 12.810 3398.260 ;
        RECT 1269.760 3398.200 1269.900 3401.800 ;
        RECT 1329.470 3401.740 1329.790 3401.800 ;
        RECT 2709.010 3401.940 2709.330 3402.000 ;
        RECT 2718.685 3401.940 2718.975 3401.985 ;
        RECT 2709.010 3401.800 2718.975 3401.940 ;
        RECT 2709.010 3401.740 2709.330 3401.800 ;
        RECT 2718.685 3401.755 2718.975 3401.800 ;
        RECT 2807.910 3401.600 2808.230 3401.660 ;
        RECT 2807.715 3401.460 2808.230 3401.600 ;
        RECT 2807.910 3401.400 2808.230 3401.460 ;
        RECT 2807.925 3399.560 2808.215 3399.605 ;
        RECT 2734.860 3399.420 2808.215 3399.560 ;
        RECT 2718.685 3398.880 2718.975 3398.925 ;
        RECT 2734.860 3398.880 2735.000 3399.420 ;
        RECT 2807.925 3399.375 2808.215 3399.420 ;
        RECT 2718.685 3398.740 2735.000 3398.880 ;
        RECT 2718.685 3398.695 2718.975 3398.740 ;
        RECT 12.490 3398.060 1269.900 3398.200 ;
        RECT 12.490 3398.000 12.810 3398.060 ;
        RECT 18.470 3395.820 18.790 3395.880 ;
        RECT 1035.085 3395.820 1035.375 3395.865 ;
        RECT 18.470 3395.680 1035.375 3395.820 ;
        RECT 18.470 3395.620 18.790 3395.680 ;
        RECT 1035.085 3395.635 1035.375 3395.680 ;
        RECT 9.730 3010.600 10.050 3010.660 ;
        RECT 9.535 3010.460 10.050 3010.600 ;
        RECT 9.730 3010.400 10.050 3010.460 ;
        RECT 8.365 3005.500 8.655 3005.545 ;
        RECT 9.730 3005.500 10.050 3005.560 ;
        RECT 8.365 3005.360 10.050 3005.500 ;
        RECT 8.365 3005.315 8.655 3005.360 ;
        RECT 9.730 3005.300 10.050 3005.360 ;
        RECT 7.890 3004.820 8.210 3004.880 ;
        RECT 9.730 3004.820 10.050 3004.880 ;
        RECT 7.890 3004.680 10.050 3004.820 ;
        RECT 7.890 3004.620 8.210 3004.680 ;
        RECT 9.730 3004.620 10.050 3004.680 ;
        RECT 8.365 3002.780 8.655 3002.825 ;
        RECT 9.730 3002.780 10.050 3002.840 ;
        RECT 8.365 3002.640 10.050 3002.780 ;
        RECT 8.365 3002.595 8.655 3002.640 ;
        RECT 9.730 3002.580 10.050 3002.640 ;
        RECT 9.730 2999.380 10.050 2999.440 ;
        RECT 9.535 2999.240 10.050 2999.380 ;
        RECT 9.730 2999.180 10.050 2999.240 ;
        RECT 7.890 2886.500 8.210 2886.560 ;
        RECT 9.730 2886.500 10.050 2886.560 ;
        RECT 7.890 2886.360 10.050 2886.500 ;
        RECT 7.890 2886.300 8.210 2886.360 ;
        RECT 9.730 2886.300 10.050 2886.360 ;
        RECT 9.730 2846.520 10.050 2846.780 ;
        RECT 8.810 2845.700 9.130 2845.760 ;
        RECT 9.820 2845.700 9.960 2846.520 ;
        RECT 8.810 2845.560 9.960 2845.700 ;
        RECT 8.810 2845.500 9.130 2845.560 ;
        RECT 8.365 2822.240 8.655 2822.285 ;
        RECT 9.730 2822.240 10.050 2822.300 ;
        RECT 8.365 2822.100 10.050 2822.240 ;
        RECT 8.365 2822.055 8.655 2822.100 ;
        RECT 9.730 2822.040 10.050 2822.100 ;
        RECT 6.510 2820.540 6.830 2820.600 ;
        RECT 9.730 2820.540 10.050 2820.600 ;
        RECT 6.510 2820.400 10.050 2820.540 ;
        RECT 6.510 2820.340 6.830 2820.400 ;
        RECT 9.730 2820.340 10.050 2820.400 ;
        RECT 8.365 2817.140 8.655 2817.185 ;
        RECT 9.730 2817.140 10.050 2817.200 ;
        RECT 8.365 2817.000 10.050 2817.140 ;
        RECT 8.365 2816.955 8.655 2817.000 ;
        RECT 9.730 2816.940 10.050 2817.000 ;
        RECT 8.365 2632.520 8.655 2632.565 ;
        RECT 9.730 2632.520 10.050 2632.580 ;
        RECT 8.365 2632.380 10.050 2632.520 ;
        RECT 8.365 2632.335 8.655 2632.380 ;
        RECT 9.730 2632.320 10.050 2632.380 ;
        RECT 7.890 2631.840 8.210 2631.900 ;
        RECT 9.730 2631.840 10.050 2631.900 ;
        RECT 7.890 2631.700 10.050 2631.840 ;
        RECT 7.890 2631.640 8.210 2631.700 ;
        RECT 9.730 2631.640 10.050 2631.700 ;
        RECT 8.365 2630.820 8.655 2630.865 ;
        RECT 9.730 2630.820 10.050 2630.880 ;
        RECT 8.365 2630.680 10.050 2630.820 ;
        RECT 8.365 2630.635 8.655 2630.680 ;
        RECT 9.730 2630.620 10.050 2630.680 ;
        RECT 7.445 2535.960 7.735 2536.005 ;
        RECT 9.730 2535.960 10.050 2536.020 ;
        RECT 7.445 2535.820 10.050 2535.960 ;
        RECT 7.445 2535.775 7.735 2535.820 ;
        RECT 9.730 2535.760 10.050 2535.820 ;
        RECT 8.825 2530.520 9.115 2530.565 ;
        RECT 9.730 2530.520 10.050 2530.580 ;
        RECT 8.825 2530.380 10.050 2530.520 ;
        RECT 8.825 2530.335 9.115 2530.380 ;
        RECT 9.730 2530.320 10.050 2530.380 ;
        RECT 7.890 2526.100 8.210 2526.160 ;
        RECT 9.730 2526.100 10.050 2526.160 ;
        RECT 7.890 2525.960 10.050 2526.100 ;
        RECT 7.890 2525.900 8.210 2525.960 ;
        RECT 9.730 2525.900 10.050 2525.960 ;
        RECT 8.825 2524.400 9.115 2524.445 ;
        RECT 8.825 2524.260 9.960 2524.400 ;
        RECT 8.825 2524.215 9.115 2524.260 ;
        RECT 9.820 2524.120 9.960 2524.260 ;
        RECT 9.730 2523.860 10.050 2524.120 ;
        RECT 7.445 2511.140 7.735 2511.185 ;
        RECT 9.730 2511.140 10.050 2511.200 ;
        RECT 7.445 2511.000 10.050 2511.140 ;
        RECT 7.445 2510.955 7.735 2511.000 ;
        RECT 9.730 2510.940 10.050 2511.000 ;
        RECT 5.130 2348.960 5.450 2349.020 ;
        RECT 9.730 2348.960 10.050 2349.020 ;
        RECT 5.130 2348.820 10.050 2348.960 ;
        RECT 5.130 2348.760 5.450 2348.820 ;
        RECT 9.730 2348.760 10.050 2348.820 ;
        RECT 9.730 2341.280 10.050 2341.540 ;
        RECT 9.820 2340.520 9.960 2341.280 ;
        RECT 9.730 2340.260 10.050 2340.520 ;
        RECT 6.985 2249.680 7.275 2249.725 ;
        RECT 9.730 2249.680 10.050 2249.740 ;
        RECT 6.985 2249.540 10.050 2249.680 ;
        RECT 6.985 2249.495 7.275 2249.540 ;
        RECT 9.730 2249.480 10.050 2249.540 ;
        RECT 7.905 2243.900 8.195 2243.945 ;
        RECT 9.730 2243.900 10.050 2243.960 ;
        RECT 7.905 2243.760 10.050 2243.900 ;
        RECT 7.905 2243.715 8.195 2243.760 ;
        RECT 9.730 2243.700 10.050 2243.760 ;
        RECT 6.970 2243.220 7.290 2243.280 ;
        RECT 9.730 2243.220 10.050 2243.280 ;
        RECT 6.970 2243.080 10.050 2243.220 ;
        RECT 6.970 2243.020 7.290 2243.080 ;
        RECT 9.730 2243.020 10.050 2243.080 ;
        RECT 7.905 2242.540 8.195 2242.585 ;
        RECT 9.730 2242.540 10.050 2242.600 ;
        RECT 7.905 2242.400 10.050 2242.540 ;
        RECT 7.905 2242.355 8.195 2242.400 ;
        RECT 9.730 2242.340 10.050 2242.400 ;
        RECT 6.985 2239.820 7.275 2239.865 ;
        RECT 9.730 2239.820 10.050 2239.880 ;
        RECT 6.985 2239.680 10.050 2239.820 ;
        RECT 6.985 2239.635 7.275 2239.680 ;
        RECT 9.730 2239.620 10.050 2239.680 ;
        RECT 6.985 1671.000 7.275 1671.045 ;
        RECT 9.730 1671.000 10.050 1671.060 ;
        RECT 6.985 1670.860 10.050 1671.000 ;
        RECT 6.985 1670.815 7.275 1670.860 ;
        RECT 9.730 1670.800 10.050 1670.860 ;
        RECT 8.825 1670.320 9.115 1670.365 ;
        RECT 9.730 1670.320 10.050 1670.380 ;
        RECT 8.825 1670.180 10.050 1670.320 ;
        RECT 8.825 1670.135 9.115 1670.180 ;
        RECT 9.730 1670.120 10.050 1670.180 ;
        RECT 6.510 1668.620 6.830 1668.680 ;
        RECT 9.730 1668.620 10.050 1668.680 ;
        RECT 6.510 1668.480 10.050 1668.620 ;
        RECT 6.510 1668.420 6.830 1668.480 ;
        RECT 9.730 1668.420 10.050 1668.480 ;
        RECT 6.985 1667.260 7.275 1667.305 ;
        RECT 9.730 1667.260 10.050 1667.320 ;
        RECT 6.985 1667.120 10.050 1667.260 ;
        RECT 6.985 1667.075 7.275 1667.120 ;
        RECT 9.730 1667.060 10.050 1667.120 ;
        RECT 8.825 1660.120 9.115 1660.165 ;
        RECT 8.825 1659.980 9.960 1660.120 ;
        RECT 8.825 1659.935 9.115 1659.980 ;
        RECT 9.820 1659.160 9.960 1659.980 ;
        RECT 9.730 1658.900 10.050 1659.160 ;
        RECT 6.525 1575.800 6.815 1575.845 ;
        RECT 9.730 1575.800 10.050 1575.860 ;
        RECT 6.525 1575.660 10.050 1575.800 ;
        RECT 6.525 1575.615 6.815 1575.660 ;
        RECT 9.730 1575.600 10.050 1575.660 ;
        RECT 7.445 1562.200 7.735 1562.245 ;
        RECT 9.730 1562.200 10.050 1562.260 ;
        RECT 7.445 1562.060 10.050 1562.200 ;
        RECT 7.445 1562.015 7.735 1562.060 ;
        RECT 9.730 1562.000 10.050 1562.060 ;
        RECT 6.985 1561.520 7.275 1561.565 ;
        RECT 9.730 1561.520 10.050 1561.580 ;
        RECT 6.985 1561.380 10.050 1561.520 ;
        RECT 6.985 1561.335 7.275 1561.380 ;
        RECT 9.730 1561.320 10.050 1561.380 ;
        RECT 6.065 1560.840 6.355 1560.885 ;
        RECT 6.985 1560.840 7.275 1560.885 ;
        RECT 6.065 1560.700 7.275 1560.840 ;
        RECT 6.065 1560.655 6.355 1560.700 ;
        RECT 6.985 1560.655 7.275 1560.700 ;
        RECT 9.730 1560.640 10.050 1560.900 ;
        RECT 9.820 1560.500 9.960 1560.640 ;
        RECT 7.060 1560.360 9.960 1560.500 ;
        RECT 7.060 1560.205 7.200 1560.360 ;
        RECT 6.985 1559.975 7.275 1560.205 ;
        RECT 6.525 1559.140 6.815 1559.185 ;
        RECT 9.730 1559.140 10.050 1559.200 ;
        RECT 6.525 1559.000 10.050 1559.140 ;
        RECT 6.525 1558.955 6.815 1559.000 ;
        RECT 9.730 1558.940 10.050 1559.000 ;
        RECT 6.525 1522.760 6.815 1522.805 ;
        RECT 9.730 1522.760 10.050 1522.820 ;
        RECT 6.525 1522.620 10.050 1522.760 ;
        RECT 6.525 1522.575 6.815 1522.620 ;
        RECT 9.730 1522.560 10.050 1522.620 ;
        RECT 6.065 1520.720 6.355 1520.765 ;
        RECT 9.730 1520.720 10.050 1520.780 ;
        RECT 6.065 1520.580 10.050 1520.720 ;
        RECT 6.065 1520.535 6.355 1520.580 ;
        RECT 9.730 1520.520 10.050 1520.580 ;
        RECT 6.985 1520.040 7.275 1520.085 ;
        RECT 9.730 1520.040 10.050 1520.100 ;
        RECT 6.985 1519.900 10.050 1520.040 ;
        RECT 6.985 1519.855 7.275 1519.900 ;
        RECT 9.730 1519.840 10.050 1519.900 ;
        RECT 6.065 1516.980 6.355 1517.025 ;
        RECT 9.730 1516.980 10.050 1517.040 ;
        RECT 6.065 1516.840 10.050 1516.980 ;
        RECT 6.065 1516.795 6.355 1516.840 ;
        RECT 9.730 1516.780 10.050 1516.840 ;
        RECT 5.605 1490.460 5.895 1490.505 ;
        RECT 6.525 1490.460 6.815 1490.505 ;
        RECT 5.605 1490.320 6.815 1490.460 ;
        RECT 5.605 1490.275 5.895 1490.320 ;
        RECT 6.525 1490.275 6.815 1490.320 ;
        RECT 6.525 1480.260 6.815 1480.305 ;
        RECT 7.905 1480.260 8.195 1480.305 ;
        RECT 6.525 1480.120 8.195 1480.260 ;
        RECT 6.525 1480.075 6.815 1480.120 ;
        RECT 7.905 1480.075 8.195 1480.120 ;
        RECT 5.605 1472.440 5.895 1472.485 ;
        RECT 7.445 1472.440 7.735 1472.485 ;
        RECT 5.605 1472.300 7.735 1472.440 ;
        RECT 5.605 1472.255 5.895 1472.300 ;
        RECT 7.445 1472.255 7.735 1472.300 ;
        RECT 6.985 1467.000 7.275 1467.045 ;
        RECT 9.730 1467.000 10.050 1467.060 ;
        RECT 6.985 1466.860 10.050 1467.000 ;
        RECT 6.985 1466.815 7.275 1466.860 ;
        RECT 9.730 1466.800 10.050 1466.860 ;
        RECT 6.065 1465.640 6.355 1465.685 ;
        RECT 9.730 1465.640 10.050 1465.700 ;
        RECT 6.065 1465.500 10.050 1465.640 ;
        RECT 6.065 1465.455 6.355 1465.500 ;
        RECT 9.730 1465.440 10.050 1465.500 ;
        RECT 6.525 1460.880 6.815 1460.925 ;
        RECT 7.905 1460.880 8.195 1460.925 ;
        RECT 6.525 1460.740 8.195 1460.880 ;
        RECT 6.525 1460.695 6.815 1460.740 ;
        RECT 7.905 1460.695 8.195 1460.740 ;
        RECT 6.525 1435.720 6.815 1435.765 ;
        RECT 7.445 1435.720 7.735 1435.765 ;
        RECT 6.525 1435.580 7.735 1435.720 ;
        RECT 6.525 1435.535 6.815 1435.580 ;
        RECT 7.445 1435.535 7.735 1435.580 ;
        RECT 6.985 1423.820 7.275 1423.865 ;
        RECT 9.730 1423.820 10.050 1423.880 ;
        RECT 6.985 1423.680 10.050 1423.820 ;
        RECT 6.985 1423.635 7.275 1423.680 ;
        RECT 9.730 1423.620 10.050 1423.680 ;
        RECT 6.525 1423.140 6.815 1423.185 ;
        RECT 9.730 1423.140 10.050 1423.200 ;
        RECT 6.525 1423.000 10.050 1423.140 ;
        RECT 6.525 1422.955 6.815 1423.000 ;
        RECT 9.730 1422.940 10.050 1423.000 ;
        RECT 7.445 1421.780 7.735 1421.825 ;
        RECT 9.730 1421.780 10.050 1421.840 ;
        RECT 7.445 1421.640 10.050 1421.780 ;
        RECT 7.445 1421.595 7.735 1421.640 ;
        RECT 9.730 1421.580 10.050 1421.640 ;
        RECT 6.970 1419.740 7.290 1419.800 ;
        RECT 6.775 1419.600 7.290 1419.740 ;
        RECT 6.970 1419.540 7.290 1419.600 ;
        RECT 6.985 1417.360 7.275 1417.405 ;
        RECT 9.285 1417.360 9.575 1417.405 ;
        RECT 6.985 1417.220 9.575 1417.360 ;
        RECT 6.985 1417.175 7.275 1417.220 ;
        RECT 9.285 1417.175 9.575 1417.220 ;
        RECT 8.825 1320.800 9.115 1320.845 ;
        RECT 9.730 1320.800 10.050 1320.860 ;
        RECT 8.825 1320.660 10.050 1320.800 ;
        RECT 8.825 1320.615 9.115 1320.660 ;
        RECT 9.730 1320.600 10.050 1320.660 ;
        RECT 7.905 1099.800 8.195 1099.845 ;
        RECT 9.730 1099.800 10.050 1099.860 ;
        RECT 7.905 1099.660 10.050 1099.800 ;
        RECT 7.905 1099.615 8.195 1099.660 ;
        RECT 9.730 1099.600 10.050 1099.660 ;
        RECT 8.825 1091.640 9.115 1091.685 ;
        RECT 9.730 1091.640 10.050 1091.700 ;
        RECT 8.825 1091.500 10.050 1091.640 ;
        RECT 8.825 1091.455 9.115 1091.500 ;
        RECT 9.730 1091.440 10.050 1091.500 ;
        RECT 8.825 1088.580 9.115 1088.625 ;
        RECT 9.730 1088.580 10.050 1088.640 ;
        RECT 8.825 1088.440 10.050 1088.580 ;
        RECT 8.825 1088.395 9.115 1088.440 ;
        RECT 9.730 1088.380 10.050 1088.440 ;
        RECT 6.970 1071.580 7.290 1071.640 ;
        RECT 9.730 1071.580 10.050 1071.640 ;
        RECT 6.970 1071.440 10.050 1071.580 ;
        RECT 6.970 1071.380 7.290 1071.440 ;
        RECT 9.730 1071.380 10.050 1071.440 ;
        RECT 5.605 1038.940 5.895 1038.985 ;
        RECT 7.905 1038.940 8.195 1038.985 ;
        RECT 5.605 1038.800 8.195 1038.940 ;
        RECT 5.605 1038.755 5.895 1038.800 ;
        RECT 7.905 1038.755 8.195 1038.800 ;
        RECT 5.145 1024.660 5.435 1024.705 ;
        RECT 6.970 1024.660 7.290 1024.720 ;
        RECT 5.145 1024.520 7.290 1024.660 ;
        RECT 5.145 1024.475 5.435 1024.520 ;
        RECT 6.970 1024.460 7.290 1024.520 ;
        RECT 3.305 1009.360 3.595 1009.405 ;
        RECT 9.730 1009.360 10.050 1009.420 ;
        RECT 3.305 1009.220 10.050 1009.360 ;
        RECT 3.305 1009.175 3.595 1009.220 ;
        RECT 9.730 1009.160 10.050 1009.220 ;
        RECT 6.970 991.340 7.290 991.400 ;
        RECT 6.970 991.200 9.960 991.340 ;
        RECT 6.970 991.140 7.290 991.200 ;
        RECT 9.820 991.060 9.960 991.200 ;
        RECT 9.730 990.800 10.050 991.060 ;
        RECT 5.605 989.640 5.895 989.685 ;
        RECT 6.525 989.640 6.815 989.685 ;
        RECT 5.605 989.500 6.815 989.640 ;
        RECT 5.605 989.455 5.895 989.500 ;
        RECT 6.525 989.455 6.815 989.500 ;
        RECT 5.605 988.960 5.895 989.005 ;
        RECT 9.730 988.960 10.050 989.020 ;
        RECT 5.605 988.820 10.050 988.960 ;
        RECT 5.605 988.775 5.895 988.820 ;
        RECT 9.730 988.760 10.050 988.820 ;
        RECT 9.730 988.280 10.050 988.340 ;
        RECT 9.535 988.140 10.050 988.280 ;
        RECT 9.730 988.080 10.050 988.140 ;
        RECT 9.730 981.820 10.050 981.880 ;
        RECT 9.535 981.680 10.050 981.820 ;
        RECT 9.730 981.620 10.050 981.680 ;
        RECT 4.225 981.140 4.515 981.185 ;
        RECT 9.730 981.140 10.050 981.200 ;
        RECT 4.225 981.000 10.050 981.140 ;
        RECT 4.225 980.955 4.515 981.000 ;
        RECT 9.730 980.940 10.050 981.000 ;
        RECT 6.525 979.100 6.815 979.145 ;
        RECT 9.730 979.100 10.050 979.160 ;
        RECT 6.525 978.960 10.050 979.100 ;
        RECT 6.525 978.915 6.815 978.960 ;
        RECT 9.730 978.900 10.050 978.960 ;
        RECT 5.605 973.660 5.895 973.705 ;
        RECT 9.730 973.660 10.050 973.720 ;
        RECT 5.605 973.520 10.050 973.660 ;
        RECT 5.605 973.475 5.895 973.520 ;
        RECT 9.730 973.460 10.050 973.520 ;
        RECT 3.290 969.920 3.610 969.980 ;
        RECT 3.095 969.780 3.610 969.920 ;
        RECT 3.290 969.720 3.610 969.780 ;
        RECT 7.445 948.160 7.735 948.205 ;
        RECT 9.730 948.160 10.050 948.220 ;
        RECT 7.445 948.020 10.050 948.160 ;
        RECT 7.445 947.975 7.735 948.020 ;
        RECT 9.730 947.960 10.050 948.020 ;
        RECT 9.730 943.400 10.050 943.460 ;
        RECT 7.060 943.260 10.050 943.400 ;
        RECT 7.060 942.040 7.200 943.260 ;
        RECT 9.730 943.200 10.050 943.260 ;
        RECT 7.445 942.720 7.735 942.765 ;
        RECT 9.730 942.720 10.050 942.780 ;
        RECT 7.445 942.580 10.050 942.720 ;
        RECT 7.445 942.535 7.735 942.580 ;
        RECT 9.730 942.520 10.050 942.580 ;
        RECT 7.445 942.040 7.735 942.085 ;
        RECT 7.060 941.900 7.735 942.040 ;
        RECT 7.445 941.855 7.735 941.900 ;
        RECT 7.445 883.900 7.735 883.945 ;
        RECT 9.730 883.900 10.050 883.960 ;
        RECT 7.445 883.760 10.050 883.900 ;
        RECT 7.445 883.715 7.735 883.760 ;
        RECT 9.730 883.700 10.050 883.760 ;
        RECT 7.430 865.880 7.750 865.940 ;
        RECT 9.270 865.880 9.590 865.940 ;
        RECT 7.430 865.740 9.590 865.880 ;
        RECT 7.430 865.680 7.750 865.740 ;
        RECT 9.270 865.680 9.590 865.740 ;
        RECT 5.130 836.300 5.450 836.360 ;
        RECT 6.525 836.300 6.815 836.345 ;
        RECT 5.130 836.160 6.815 836.300 ;
        RECT 5.130 836.100 5.450 836.160 ;
        RECT 6.525 836.115 6.815 836.160 ;
        RECT 6.985 832.220 7.275 832.265 ;
        RECT 9.730 832.220 10.050 832.280 ;
        RECT 6.985 832.080 10.050 832.220 ;
        RECT 6.985 832.035 7.275 832.080 ;
        RECT 9.730 832.020 10.050 832.080 ;
        RECT 9.730 831.540 10.050 831.600 ;
        RECT 6.600 831.400 10.050 831.540 ;
        RECT 6.600 829.500 6.740 831.400 ;
        RECT 9.730 831.340 10.050 831.400 ;
        RECT 6.970 830.180 7.290 830.240 ;
        RECT 9.730 830.180 10.050 830.240 ;
        RECT 6.970 830.040 10.050 830.180 ;
        RECT 6.970 829.980 7.290 830.040 ;
        RECT 9.730 829.980 10.050 830.040 ;
        RECT 9.730 829.500 10.050 829.560 ;
        RECT 6.600 829.360 10.050 829.500 ;
        RECT 9.730 829.300 10.050 829.360 ;
        RECT 6.985 827.460 7.275 827.505 ;
        RECT 9.730 827.460 10.050 827.520 ;
        RECT 6.985 827.320 10.050 827.460 ;
        RECT 6.985 827.275 7.275 827.320 ;
        RECT 9.730 827.260 10.050 827.320 ;
        RECT 7.430 799.920 7.750 799.980 ;
        RECT 9.730 799.920 10.050 799.980 ;
        RECT 7.430 799.780 10.050 799.920 ;
        RECT 7.430 799.720 7.750 799.780 ;
        RECT 9.730 799.720 10.050 799.780 ;
        RECT 7.430 798.560 7.750 798.620 ;
        RECT 9.730 798.560 10.050 798.620 ;
        RECT 7.430 798.420 10.050 798.560 ;
        RECT 7.430 798.360 7.750 798.420 ;
        RECT 9.730 798.360 10.050 798.420 ;
        RECT 6.525 797.200 6.815 797.245 ;
        RECT 8.825 797.200 9.115 797.245 ;
        RECT 6.525 797.060 9.115 797.200 ;
        RECT 6.525 797.015 6.815 797.060 ;
        RECT 8.825 797.015 9.115 797.060 ;
        RECT 6.065 768.980 6.355 769.025 ;
        RECT 9.270 768.980 9.590 769.040 ;
        RECT 6.065 768.840 9.590 768.980 ;
        RECT 6.065 768.795 6.355 768.840 ;
        RECT 9.270 768.780 9.590 768.840 ;
        RECT 7.890 735.660 8.210 735.720 ;
        RECT 9.730 735.660 10.050 735.720 ;
        RECT 7.890 735.520 10.050 735.660 ;
        RECT 7.890 735.460 8.210 735.520 ;
        RECT 9.730 735.460 10.050 735.520 ;
        RECT 4.685 734.980 4.975 735.025 ;
        RECT 6.065 734.980 6.355 735.025 ;
        RECT 4.685 734.840 6.355 734.980 ;
        RECT 4.685 734.795 4.975 734.840 ;
        RECT 6.065 734.795 6.355 734.840 ;
        RECT 7.890 731.920 8.210 731.980 ;
        RECT 8.825 731.920 9.115 731.965 ;
        RECT 7.890 731.780 9.115 731.920 ;
        RECT 7.890 731.720 8.210 731.780 ;
        RECT 8.825 731.735 9.115 731.780 ;
        RECT 7.890 714.920 8.210 714.980 ;
        RECT 9.285 714.920 9.575 714.965 ;
        RECT 7.890 714.780 9.575 714.920 ;
        RECT 7.890 714.720 8.210 714.780 ;
        RECT 9.285 714.735 9.575 714.780 ;
        RECT 4.685 714.240 4.975 714.285 ;
        RECT 5.130 714.240 5.450 714.300 ;
        RECT 4.685 714.100 5.450 714.240 ;
        RECT 4.685 714.055 4.975 714.100 ;
        RECT 5.130 714.040 5.450 714.100 ;
        RECT 2.830 708.800 3.150 708.860 ;
        RECT 4.210 708.800 4.530 708.860 ;
        RECT 2.830 708.660 4.530 708.800 ;
        RECT 2.830 708.600 3.150 708.660 ;
        RECT 4.210 708.600 4.530 708.660 ;
        RECT 3.765 706.080 4.055 706.125 ;
        RECT 9.730 706.080 10.050 706.140 ;
        RECT 3.765 705.940 10.050 706.080 ;
        RECT 3.765 705.895 4.055 705.940 ;
        RECT 9.730 705.880 10.050 705.940 ;
        RECT 8.825 699.960 9.115 700.005 ;
        RECT 9.730 699.960 10.050 700.020 ;
        RECT 8.825 699.820 10.050 699.960 ;
        RECT 8.825 699.775 9.115 699.820 ;
        RECT 9.730 699.760 10.050 699.820 ;
        RECT 1.465 694.860 1.755 694.905 ;
        RECT 8.825 694.860 9.115 694.905 ;
        RECT 1.465 694.720 9.115 694.860 ;
        RECT 1.465 694.675 1.755 694.720 ;
        RECT 8.825 694.675 9.115 694.720 ;
        RECT 7.430 693.160 7.750 693.220 ;
        RECT 9.730 693.160 10.050 693.220 ;
        RECT 7.430 693.020 10.050 693.160 ;
        RECT 7.430 692.960 7.750 693.020 ;
        RECT 9.730 692.960 10.050 693.020 ;
        RECT 4.685 672.760 4.975 672.805 ;
        RECT 5.130 672.760 5.450 672.820 ;
        RECT 4.685 672.620 5.450 672.760 ;
        RECT 4.685 672.575 4.975 672.620 ;
        RECT 5.130 672.560 5.450 672.620 ;
        RECT 5.130 666.640 5.450 666.700 ;
        RECT 9.285 666.640 9.575 666.685 ;
        RECT 5.130 666.500 9.575 666.640 ;
        RECT 5.130 666.440 5.450 666.500 ;
        RECT 9.285 666.455 9.575 666.500 ;
        RECT 3.305 660.520 3.595 660.565 ;
        RECT 9.730 660.520 10.050 660.580 ;
        RECT 3.305 660.380 10.050 660.520 ;
        RECT 3.305 660.335 3.595 660.380 ;
        RECT 9.730 660.320 10.050 660.380 ;
        RECT 7.905 654.400 8.195 654.445 ;
        RECT 9.730 654.400 10.050 654.460 ;
        RECT 7.905 654.260 10.050 654.400 ;
        RECT 7.905 654.215 8.195 654.260 ;
        RECT 9.730 654.200 10.050 654.260 ;
        RECT 2.845 653.040 3.135 653.085 ;
        RECT 9.730 653.040 10.050 653.100 ;
        RECT 2.845 652.900 10.050 653.040 ;
        RECT 2.845 652.855 3.135 652.900 ;
        RECT 9.730 652.840 10.050 652.900 ;
        RECT 2.385 652.020 2.675 652.065 ;
        RECT 3.765 652.020 4.055 652.065 ;
        RECT 2.385 651.880 4.055 652.020 ;
        RECT 2.385 651.835 2.675 651.880 ;
        RECT 3.765 651.835 4.055 651.880 ;
        RECT 1.465 651.340 1.755 651.385 ;
        RECT 3.765 651.340 4.055 651.385 ;
        RECT 1.465 651.200 4.055 651.340 ;
        RECT 1.465 651.155 1.755 651.200 ;
        RECT 3.765 651.155 4.055 651.200 ;
        RECT 2.385 647.260 2.675 647.305 ;
        RECT 9.730 647.260 10.050 647.320 ;
        RECT 2.385 647.120 10.050 647.260 ;
        RECT 2.385 647.075 2.675 647.120 ;
        RECT 9.730 647.060 10.050 647.120 ;
        RECT 7.905 645.900 8.195 645.945 ;
        RECT 9.730 645.900 10.050 645.960 ;
        RECT 7.905 645.760 10.050 645.900 ;
        RECT 7.905 645.715 8.195 645.760 ;
        RECT 9.730 645.700 10.050 645.760 ;
        RECT 4.210 644.540 4.530 644.600 ;
        RECT 7.905 644.540 8.195 644.585 ;
        RECT 4.210 644.400 8.195 644.540 ;
        RECT 4.210 644.340 4.530 644.400 ;
        RECT 7.905 644.355 8.195 644.400 ;
        RECT 4.685 641.820 4.975 641.865 ;
        RECT 9.270 641.820 9.590 641.880 ;
        RECT 4.685 641.680 9.590 641.820 ;
        RECT 4.685 641.635 4.975 641.680 ;
        RECT 9.270 641.620 9.590 641.680 ;
        RECT 5.145 632.640 5.435 632.685 ;
        RECT 7.905 632.640 8.195 632.685 ;
        RECT 5.145 632.500 8.195 632.640 ;
        RECT 5.145 632.455 5.435 632.500 ;
        RECT 7.905 632.455 8.195 632.500 ;
        RECT 7.905 631.960 8.195 632.005 ;
        RECT 9.270 631.960 9.590 632.020 ;
        RECT 7.905 631.820 9.590 631.960 ;
        RECT 7.905 631.775 8.195 631.820 ;
        RECT 9.270 631.760 9.590 631.820 ;
        RECT 3.305 631.280 3.595 631.325 ;
        RECT 4.685 631.280 4.975 631.325 ;
        RECT 3.305 631.140 4.975 631.280 ;
        RECT 3.305 631.095 3.595 631.140 ;
        RECT 4.685 631.095 4.975 631.140 ;
        RECT 5.145 597.960 5.435 598.005 ;
        RECT 8.825 597.960 9.115 598.005 ;
        RECT 5.145 597.820 9.115 597.960 ;
        RECT 5.145 597.775 5.435 597.820 ;
        RECT 8.825 597.775 9.115 597.820 ;
        RECT 6.050 587.760 6.370 587.820 ;
        RECT 9.730 587.760 10.050 587.820 ;
        RECT 6.050 587.620 10.050 587.760 ;
        RECT 6.050 587.560 6.370 587.620 ;
        RECT 9.730 587.560 10.050 587.620 ;
        RECT 3.765 587.420 4.055 587.465 ;
        RECT 5.145 587.420 5.435 587.465 ;
        RECT 3.765 587.280 5.435 587.420 ;
        RECT 3.765 587.235 4.055 587.280 ;
        RECT 5.145 587.235 5.435 587.280 ;
        RECT 4.685 587.080 4.975 587.125 ;
        RECT 9.730 587.080 10.050 587.140 ;
        RECT 4.685 586.940 10.050 587.080 ;
        RECT 4.685 586.895 4.975 586.940 ;
        RECT 9.730 586.880 10.050 586.940 ;
        RECT 5.145 576.200 5.435 576.245 ;
        RECT 7.445 576.200 7.735 576.245 ;
        RECT 5.145 576.060 7.735 576.200 ;
        RECT 5.145 576.015 5.435 576.060 ;
        RECT 7.445 576.015 7.735 576.060 ;
        RECT 4.685 575.520 4.975 575.565 ;
        RECT 6.050 575.520 6.370 575.580 ;
        RECT 4.685 575.380 6.370 575.520 ;
        RECT 4.685 575.335 4.975 575.380 ;
        RECT 6.050 575.320 6.370 575.380 ;
        RECT 5.145 555.120 5.435 555.165 ;
        RECT 9.730 555.120 10.050 555.180 ;
        RECT 5.145 554.980 10.050 555.120 ;
        RECT 5.145 554.935 5.435 554.980 ;
        RECT 9.730 554.920 10.050 554.980 ;
        RECT 6.050 550.360 6.370 550.420 ;
        RECT 9.730 550.360 10.050 550.420 ;
        RECT 6.050 550.220 10.050 550.360 ;
        RECT 6.050 550.160 6.370 550.220 ;
        RECT 9.730 550.160 10.050 550.220 ;
        RECT 3.765 548.660 4.055 548.705 ;
        RECT 9.730 548.660 10.050 548.720 ;
        RECT 3.765 548.520 10.050 548.660 ;
        RECT 3.765 548.475 4.055 548.520 ;
        RECT 9.730 548.460 10.050 548.520 ;
        RECT 3.305 547.300 3.595 547.345 ;
        RECT 9.730 547.300 10.050 547.360 ;
        RECT 3.305 547.160 10.050 547.300 ;
        RECT 3.305 547.115 3.595 547.160 ;
        RECT 9.730 547.100 10.050 547.160 ;
        RECT 2.845 546.620 3.135 546.665 ;
        RECT 9.730 546.620 10.050 546.680 ;
        RECT 2.845 546.480 10.050 546.620 ;
        RECT 2.845 546.435 3.135 546.480 ;
        RECT 9.730 546.420 10.050 546.480 ;
        RECT 3.305 545.940 3.595 545.985 ;
        RECT 9.730 545.940 10.050 546.000 ;
        RECT 3.305 545.800 10.050 545.940 ;
        RECT 3.305 545.755 3.595 545.800 ;
        RECT 9.730 545.740 10.050 545.800 ;
        RECT 4.685 544.580 4.975 544.625 ;
        RECT 9.730 544.580 10.050 544.640 ;
        RECT 4.685 544.440 10.050 544.580 ;
        RECT 4.685 544.395 4.975 544.440 ;
        RECT 9.730 544.380 10.050 544.440 ;
        RECT 3.765 543.900 4.055 543.945 ;
        RECT 9.730 543.900 10.050 543.960 ;
        RECT 3.765 543.760 10.050 543.900 ;
        RECT 3.765 543.715 4.055 543.760 ;
        RECT 9.730 543.700 10.050 543.760 ;
        RECT 7.905 543.220 8.195 543.265 ;
        RECT 9.730 543.220 10.050 543.280 ;
        RECT 7.905 543.080 10.050 543.220 ;
        RECT 7.905 543.035 8.195 543.080 ;
        RECT 9.730 543.020 10.050 543.080 ;
        RECT 7.445 542.540 7.735 542.585 ;
        RECT 9.730 542.540 10.050 542.600 ;
        RECT 7.445 542.400 10.050 542.540 ;
        RECT 7.445 542.355 7.735 542.400 ;
        RECT 9.730 542.340 10.050 542.400 ;
        RECT 5.145 540.500 5.435 540.545 ;
        RECT 6.050 540.500 6.370 540.560 ;
        RECT 5.145 540.360 6.370 540.500 ;
        RECT 5.145 540.315 5.435 540.360 ;
        RECT 6.050 540.300 6.370 540.360 ;
        RECT 6.050 512.960 6.370 513.020 ;
        RECT 8.825 512.960 9.115 513.005 ;
        RECT 6.050 512.820 9.115 512.960 ;
        RECT 6.050 512.760 6.370 512.820 ;
        RECT 8.825 512.775 9.115 512.820 ;
        RECT 6.510 491.540 6.830 491.600 ;
        RECT 6.315 491.400 6.830 491.540 ;
        RECT 6.510 491.340 6.830 491.400 ;
        RECT 6.525 467.740 6.815 467.785 ;
        RECT 7.445 467.740 7.735 467.785 ;
        RECT 6.525 467.600 7.735 467.740 ;
        RECT 6.525 467.555 6.815 467.600 ;
        RECT 7.445 467.555 7.735 467.600 ;
        RECT 9.270 467.400 9.590 467.460 ;
        RECT 6.140 467.260 9.590 467.400 ;
        RECT 6.140 466.720 6.280 467.260 ;
        RECT 9.270 467.200 9.590 467.260 ;
        RECT 6.525 467.060 6.815 467.105 ;
        RECT 9.730 467.060 10.050 467.120 ;
        RECT 6.525 466.920 10.050 467.060 ;
        RECT 6.525 466.875 6.815 466.920 ;
        RECT 9.730 466.860 10.050 466.920 ;
        RECT 6.140 466.580 9.960 466.720 ;
        RECT 9.820 466.440 9.960 466.580 ;
        RECT 9.730 466.180 10.050 466.440 ;
        RECT 9.730 460.940 10.050 461.000 ;
        RECT 4.300 460.800 10.050 460.940 ;
        RECT 4.300 459.580 4.440 460.800 ;
        RECT 9.730 460.740 10.050 460.800 ;
        RECT 4.685 460.260 4.975 460.305 ;
        RECT 9.730 460.260 10.050 460.320 ;
        RECT 4.685 460.120 10.050 460.260 ;
        RECT 4.685 460.075 4.975 460.120 ;
        RECT 9.730 460.060 10.050 460.120 ;
        RECT 9.730 459.580 10.050 459.640 ;
        RECT 4.300 459.440 10.050 459.580 ;
        RECT 9.730 459.380 10.050 459.440 ;
        RECT 6.525 457.540 6.815 457.585 ;
        RECT 9.730 457.540 10.050 457.600 ;
        RECT 6.525 457.400 10.050 457.540 ;
        RECT 6.525 457.355 6.815 457.400 ;
        RECT 9.730 457.340 10.050 457.400 ;
        RECT 5.145 438.160 5.435 438.205 ;
        RECT 7.445 438.160 7.735 438.205 ;
        RECT 5.145 438.020 7.735 438.160 ;
        RECT 5.145 437.975 5.435 438.020 ;
        RECT 7.445 437.975 7.735 438.020 ;
        RECT 4.685 430.680 4.975 430.725 ;
        RECT 9.270 430.680 9.590 430.740 ;
        RECT 4.685 430.540 9.590 430.680 ;
        RECT 4.685 430.495 4.975 430.540 ;
        RECT 9.270 430.480 9.590 430.540 ;
        RECT 4.685 423.880 4.975 423.925 ;
        RECT 9.730 423.880 10.050 423.940 ;
        RECT 4.685 423.740 10.050 423.880 ;
        RECT 4.685 423.695 4.975 423.740 ;
        RECT 9.730 423.680 10.050 423.740 ;
        RECT 5.145 418.100 5.435 418.145 ;
        RECT 9.730 418.100 10.050 418.160 ;
        RECT 5.145 417.960 10.050 418.100 ;
        RECT 5.145 417.915 5.435 417.960 ;
        RECT 9.730 417.900 10.050 417.960 ;
        RECT 4.685 410.620 4.975 410.665 ;
        RECT 9.730 410.620 10.050 410.680 ;
        RECT 4.685 410.480 10.050 410.620 ;
        RECT 4.685 410.435 4.975 410.480 ;
        RECT 9.730 410.420 10.050 410.480 ;
        RECT 7.905 359.960 8.195 360.005 ;
        RECT 9.730 359.960 10.050 360.020 ;
        RECT 7.905 359.820 10.050 359.960 ;
        RECT 7.905 359.775 8.195 359.820 ;
        RECT 9.730 359.760 10.050 359.820 ;
        RECT 6.050 355.200 6.370 355.260 ;
        RECT 9.730 355.200 10.050 355.260 ;
        RECT 6.050 355.060 10.050 355.200 ;
        RECT 6.050 355.000 6.370 355.060 ;
        RECT 9.730 355.000 10.050 355.060 ;
        RECT 5.145 337.520 5.435 337.565 ;
        RECT 9.730 337.520 10.050 337.580 ;
        RECT 5.145 337.380 10.050 337.520 ;
        RECT 5.145 337.335 5.435 337.380 ;
        RECT 9.730 337.320 10.050 337.380 ;
        RECT 6.510 336.840 6.830 336.900 ;
        RECT 9.730 336.840 10.050 336.900 ;
        RECT 6.510 336.700 10.050 336.840 ;
        RECT 6.510 336.640 6.830 336.700 ;
        RECT 9.730 336.640 10.050 336.700 ;
        RECT 4.685 336.160 4.975 336.205 ;
        RECT 9.730 336.160 10.050 336.220 ;
        RECT 4.685 336.020 10.050 336.160 ;
        RECT 4.685 335.975 4.975 336.020 ;
        RECT 9.730 335.960 10.050 336.020 ;
        RECT 3.765 333.780 4.055 333.825 ;
        RECT 9.730 333.780 10.050 333.840 ;
        RECT 3.765 333.640 10.050 333.780 ;
        RECT 3.765 333.595 4.055 333.640 ;
        RECT 9.730 333.580 10.050 333.640 ;
        RECT 4.225 333.100 4.515 333.145 ;
        RECT 9.730 333.100 10.050 333.160 ;
        RECT 4.225 332.960 10.050 333.100 ;
        RECT 4.225 332.915 4.515 332.960 ;
        RECT 9.730 332.900 10.050 332.960 ;
        RECT 5.605 327.320 5.895 327.365 ;
        RECT 6.050 327.320 6.370 327.380 ;
        RECT 10.190 327.320 10.510 327.380 ;
        RECT 5.605 327.180 6.370 327.320 ;
        RECT 5.605 327.135 5.895 327.180 ;
        RECT 6.050 327.120 6.370 327.180 ;
        RECT 9.820 327.180 10.510 327.320 ;
        RECT 9.820 326.980 9.960 327.180 ;
        RECT 10.190 327.120 10.510 327.180 ;
        RECT 6.600 326.840 9.960 326.980 ;
        RECT 6.600 326.360 6.740 326.840 ;
        RECT 6.510 326.100 6.830 326.360 ;
        RECT 3.765 323.240 4.055 323.285 ;
        RECT 9.730 323.240 10.050 323.300 ;
        RECT 3.765 323.100 10.050 323.240 ;
        RECT 3.765 323.055 4.055 323.100 ;
        RECT 9.730 323.040 10.050 323.100 ;
        RECT 6.050 316.780 6.370 316.840 ;
        RECT 9.730 316.780 10.050 316.840 ;
        RECT 6.050 316.640 10.050 316.780 ;
        RECT 6.050 316.580 6.370 316.640 ;
        RECT 9.730 316.580 10.050 316.640 ;
        RECT 4.685 315.760 4.975 315.805 ;
        RECT 9.730 315.760 10.050 315.820 ;
        RECT 4.685 315.620 10.050 315.760 ;
        RECT 4.685 315.575 4.975 315.620 ;
        RECT 9.730 315.560 10.050 315.620 ;
        RECT 5.145 314.400 5.435 314.445 ;
        RECT 9.730 314.400 10.050 314.460 ;
        RECT 5.145 314.260 10.050 314.400 ;
        RECT 5.145 314.215 5.435 314.260 ;
        RECT 9.730 314.200 10.050 314.260 ;
        RECT 5.605 311.340 5.895 311.385 ;
        RECT 9.730 311.340 10.050 311.400 ;
        RECT 5.605 311.200 10.050 311.340 ;
        RECT 5.605 311.155 5.895 311.200 ;
        RECT 9.730 311.140 10.050 311.200 ;
        RECT 4.225 289.580 4.515 289.625 ;
        RECT 6.510 289.580 6.830 289.640 ;
        RECT 4.225 289.440 6.830 289.580 ;
        RECT 4.225 289.395 4.515 289.440 ;
        RECT 6.510 289.380 6.830 289.440 ;
        RECT 6.065 285.500 6.355 285.545 ;
        RECT 9.730 285.500 10.050 285.560 ;
        RECT 6.065 285.360 10.050 285.500 ;
        RECT 6.065 285.315 6.355 285.360 ;
        RECT 9.730 285.300 10.050 285.360 ;
        RECT 9.730 284.480 10.050 284.540 ;
        RECT 6.600 284.340 10.050 284.480 ;
        RECT 6.600 283.120 6.740 284.340 ;
        RECT 9.730 284.280 10.050 284.340 ;
        RECT 9.730 283.120 10.050 283.180 ;
        RECT 6.600 282.980 10.050 283.120 ;
        RECT 9.730 282.920 10.050 282.980 ;
        RECT 6.065 279.380 6.355 279.425 ;
        RECT 9.730 279.380 10.050 279.440 ;
        RECT 6.065 279.240 10.050 279.380 ;
        RECT 6.065 279.195 6.355 279.240 ;
        RECT 9.730 279.180 10.050 279.240 ;
        RECT 7.445 263.060 7.735 263.105 ;
        RECT 9.730 263.060 10.050 263.120 ;
        RECT 7.445 262.920 10.050 263.060 ;
        RECT 7.445 262.875 7.735 262.920 ;
        RECT 9.730 262.860 10.050 262.920 ;
        RECT 5.130 251.840 5.450 251.900 ;
        RECT 4.935 251.700 5.450 251.840 ;
        RECT 5.130 251.640 5.450 251.700 ;
        RECT 5.130 185.200 5.450 185.260 ;
        RECT 4.935 185.060 5.450 185.200 ;
        RECT 5.130 185.000 5.450 185.060 ;
        RECT 6.065 177.720 6.355 177.765 ;
        RECT 9.730 177.720 10.050 177.780 ;
        RECT 6.065 177.580 10.050 177.720 ;
        RECT 6.065 177.535 6.355 177.580 ;
        RECT 9.730 177.520 10.050 177.580 ;
        RECT 9.270 148.820 9.590 148.880 ;
        RECT 9.745 148.820 10.035 148.865 ;
        RECT 9.270 148.680 10.035 148.820 ;
        RECT 9.270 148.620 9.590 148.680 ;
        RECT 9.745 148.635 10.035 148.680 ;
        RECT 7.430 147.460 7.750 147.520 ;
        RECT 7.235 147.320 7.750 147.460 ;
        RECT 7.430 147.260 7.750 147.320 ;
        RECT 6.985 141.680 7.275 141.725 ;
        RECT 9.730 141.680 10.050 141.740 ;
        RECT 6.985 141.540 10.050 141.680 ;
        RECT 6.985 141.495 7.275 141.540 ;
        RECT 9.730 141.480 10.050 141.540 ;
        RECT 7.430 139.980 7.750 140.040 ;
        RECT 9.730 139.980 10.050 140.040 ;
        RECT 7.430 139.840 10.050 139.980 ;
        RECT 7.430 139.780 7.750 139.840 ;
        RECT 9.730 139.780 10.050 139.840 ;
        RECT 6.065 136.240 6.355 136.285 ;
        RECT 9.730 136.240 10.050 136.300 ;
        RECT 6.065 136.100 10.050 136.240 ;
        RECT 6.065 136.055 6.355 136.100 ;
        RECT 9.730 136.040 10.050 136.100 ;
        RECT 7.445 135.560 7.735 135.605 ;
        RECT 9.730 135.560 10.050 135.620 ;
        RECT 7.445 135.420 10.050 135.560 ;
        RECT 7.445 135.375 7.735 135.420 ;
        RECT 9.730 135.360 10.050 135.420 ;
        RECT 6.050 134.880 6.370 134.940 ;
        RECT 9.730 134.880 10.050 134.940 ;
        RECT 6.050 134.740 10.050 134.880 ;
        RECT 6.050 134.680 6.370 134.740 ;
        RECT 9.730 134.680 10.050 134.740 ;
        RECT 7.430 134.200 7.750 134.260 ;
        RECT 9.730 134.200 10.050 134.260 ;
        RECT 7.430 134.060 10.050 134.200 ;
        RECT 7.430 134.000 7.750 134.060 ;
        RECT 9.730 134.000 10.050 134.060 ;
        RECT 6.985 111.080 7.275 111.125 ;
        RECT 9.730 111.080 10.050 111.140 ;
        RECT 6.985 110.940 10.050 111.080 ;
        RECT 6.985 110.895 7.275 110.940 ;
        RECT 9.730 110.880 10.050 110.940 ;
        RECT 4.685 100.200 4.975 100.245 ;
        RECT 5.130 100.200 5.450 100.260 ;
        RECT 4.685 100.060 5.450 100.200 ;
        RECT 4.685 100.015 4.975 100.060 ;
        RECT 5.130 100.000 5.450 100.060 ;
        RECT 6.510 94.420 6.830 94.480 ;
        RECT 9.745 94.420 10.035 94.465 ;
        RECT 6.510 94.280 10.035 94.420 ;
        RECT 6.510 94.220 6.830 94.280 ;
        RECT 9.745 94.235 10.035 94.280 ;
        RECT 5.145 89.660 5.435 89.705 ;
        RECT 9.270 89.660 9.590 89.720 ;
        RECT 5.145 89.520 9.590 89.660 ;
        RECT 5.145 89.475 5.435 89.520 ;
        RECT 9.270 89.460 9.590 89.520 ;
        RECT 3.305 82.860 3.595 82.905 ;
        RECT 9.270 82.860 9.590 82.920 ;
        RECT 3.305 82.720 9.590 82.860 ;
        RECT 3.305 82.675 3.595 82.720 ;
        RECT 9.270 82.660 9.590 82.720 ;
        RECT 6.525 82.180 6.815 82.225 ;
        RECT 9.270 82.180 9.590 82.240 ;
        RECT 6.525 82.040 9.590 82.180 ;
        RECT 6.525 81.995 6.815 82.040 ;
        RECT 9.270 81.980 9.590 82.040 ;
        RECT 5.590 78.100 5.910 78.160 ;
        RECT 9.730 78.100 10.050 78.160 ;
        RECT 5.590 77.960 10.050 78.100 ;
        RECT 5.590 77.900 5.910 77.960 ;
        RECT 9.730 77.900 10.050 77.960 ;
        RECT 6.065 76.740 6.355 76.785 ;
        RECT 9.730 76.740 10.050 76.800 ;
        RECT 6.065 76.600 10.050 76.740 ;
        RECT 6.065 76.555 6.355 76.600 ;
        RECT 9.730 76.540 10.050 76.600 ;
        RECT 5.605 76.060 5.895 76.105 ;
        RECT 5.605 75.920 9.960 76.060 ;
        RECT 5.605 75.875 5.895 75.920 ;
        RECT 9.820 75.780 9.960 75.920 ;
        RECT 9.730 75.520 10.050 75.780 ;
        RECT 5.590 74.020 5.910 74.080 ;
        RECT 5.395 73.880 5.910 74.020 ;
        RECT 5.590 73.820 5.910 73.880 ;
        RECT 5.145 73.000 5.435 73.045 ;
        RECT 5.145 72.860 5.820 73.000 ;
        RECT 5.145 72.815 5.435 72.860 ;
        RECT 5.680 72.365 5.820 72.860 ;
        RECT 5.605 72.135 5.895 72.365 ;
        RECT 6.065 67.560 6.355 67.605 ;
        RECT 9.730 67.560 10.050 67.620 ;
        RECT 6.065 67.420 10.050 67.560 ;
        RECT 6.065 67.375 6.355 67.420 ;
        RECT 9.730 67.360 10.050 67.420 ;
        RECT 5.145 66.880 5.435 66.925 ;
        RECT 9.730 66.880 10.050 66.940 ;
        RECT 5.145 66.740 10.050 66.880 ;
        RECT 5.145 66.695 5.435 66.740 ;
        RECT 9.730 66.680 10.050 66.740 ;
        RECT 5.590 61.780 5.910 61.840 ;
        RECT 6.525 61.780 6.815 61.825 ;
        RECT 5.590 61.640 6.815 61.780 ;
        RECT 5.590 61.580 5.910 61.640 ;
        RECT 6.525 61.595 6.815 61.640 ;
        RECT 6.510 61.100 6.830 61.160 ;
        RECT 8.825 61.100 9.115 61.145 ;
        RECT 6.510 60.960 9.115 61.100 ;
        RECT 6.510 60.900 6.830 60.960 ;
        RECT 8.825 60.915 9.115 60.960 ;
        RECT 3.305 50.560 3.595 50.605 ;
        RECT 5.130 50.560 5.450 50.620 ;
        RECT 3.305 50.420 5.450 50.560 ;
        RECT 3.305 50.375 3.595 50.420 ;
        RECT 5.130 50.360 5.450 50.420 ;
        RECT 4.210 37.640 4.530 37.700 ;
        RECT 4.685 37.640 4.975 37.685 ;
        RECT 4.210 37.500 4.975 37.640 ;
        RECT 4.210 37.440 4.530 37.500 ;
        RECT 4.685 37.455 4.975 37.500 ;
        RECT 6.050 16.560 6.370 16.620 ;
        RECT 5.855 16.420 6.370 16.560 ;
        RECT 6.050 16.360 6.370 16.420 ;
        RECT 283.905 9.080 284.195 9.125 ;
        RECT 327.145 9.080 327.435 9.125 ;
        RECT 283.905 8.940 327.435 9.080 ;
        RECT 283.905 8.895 284.195 8.940 ;
        RECT 327.145 8.895 327.435 8.940 ;
        RECT 18.930 8.740 19.250 8.800 ;
        RECT 38.250 8.740 38.570 8.800 ;
        RECT 18.930 8.600 38.570 8.740 ;
        RECT 18.930 8.540 19.250 8.600 ;
        RECT 38.250 8.540 38.570 8.600 ;
        RECT 283.890 8.400 284.210 8.460 ;
        RECT 283.890 8.260 284.405 8.400 ;
        RECT 283.890 8.200 284.210 8.260 ;
        RECT 56.205 8.060 56.495 8.105 ;
        RECT 212.145 8.060 212.435 8.105 ;
        RECT 56.205 7.920 212.435 8.060 ;
        RECT 56.205 7.875 56.495 7.920 ;
        RECT 212.145 7.875 212.435 7.920 ;
        RECT 90.230 7.720 90.550 7.780 ;
        RECT 141.305 7.720 141.595 7.765 ;
        RECT 90.230 7.580 141.595 7.720 ;
        RECT 90.230 7.520 90.550 7.580 ;
        RECT 141.305 7.535 141.595 7.580 ;
        RECT 328.065 7.380 328.355 7.425 ;
        RECT 333.585 7.380 333.875 7.425 ;
        RECT 328.065 7.240 333.875 7.380 ;
        RECT 328.065 7.195 328.355 7.240 ;
        RECT 333.585 7.195 333.875 7.240 ;
        RECT 507.925 7.195 508.215 7.425 ;
        RECT 29.510 7.040 29.830 7.100 ;
        RECT 32.270 7.040 32.590 7.100 ;
        RECT 29.510 6.900 32.590 7.040 ;
        RECT 29.510 6.840 29.830 6.900 ;
        RECT 32.270 6.840 32.590 6.900 ;
        RECT 36.425 7.040 36.715 7.085 ;
        RECT 52.525 7.040 52.815 7.085 ;
        RECT 462.845 7.040 463.135 7.085 ;
        RECT 36.425 6.900 52.815 7.040 ;
        RECT 36.425 6.855 36.715 6.900 ;
        RECT 52.525 6.855 52.815 6.900 ;
        RECT 461.540 6.900 463.135 7.040 ;
        RECT 5.605 6.700 5.895 6.745 ;
        RECT 24.910 6.700 25.230 6.760 ;
        RECT 5.605 6.560 25.230 6.700 ;
        RECT 5.605 6.515 5.895 6.560 ;
        RECT 24.910 6.500 25.230 6.560 ;
        RECT 26.750 6.700 27.070 6.760 ;
        RECT 72.750 6.700 73.070 6.760 ;
        RECT 90.230 6.700 90.550 6.760 ;
        RECT 26.750 6.560 51.820 6.700 ;
        RECT 26.750 6.500 27.070 6.560 ;
        RECT 51.680 6.020 51.820 6.560 ;
        RECT 72.750 6.560 90.550 6.700 ;
        RECT 72.750 6.500 73.070 6.560 ;
        RECT 90.230 6.500 90.550 6.560 ;
        RECT 335.425 6.700 335.715 6.745 ;
        RECT 363.945 6.700 364.235 6.745 ;
        RECT 335.425 6.560 364.235 6.700 ;
        RECT 335.425 6.515 335.715 6.560 ;
        RECT 363.945 6.515 364.235 6.560 ;
        RECT 417.765 6.700 418.055 6.745 ;
        RECT 461.540 6.700 461.680 6.900 ;
        RECT 462.845 6.855 463.135 6.900 ;
        RECT 465.145 7.040 465.435 7.085 ;
        RECT 508.000 7.040 508.140 7.195 ;
        RECT 465.145 6.900 508.140 7.040 ;
        RECT 465.145 6.855 465.435 6.900 ;
        RECT 417.765 6.560 431.320 6.700 ;
        RECT 417.765 6.515 418.055 6.560 ;
        RECT 52.065 6.360 52.355 6.405 ;
        RECT 55.285 6.360 55.575 6.405 ;
        RECT 52.065 6.220 55.575 6.360 ;
        RECT 52.065 6.175 52.355 6.220 ;
        RECT 55.285 6.175 55.575 6.220 ;
        RECT 141.305 6.360 141.595 6.405 ;
        RECT 431.180 6.360 431.320 6.560 ;
        RECT 438.540 6.560 461.680 6.700 ;
        RECT 438.540 6.360 438.680 6.560 ;
        RECT 141.305 6.220 196.720 6.360 ;
        RECT 431.180 6.220 438.680 6.360 ;
        RECT 141.305 6.175 141.595 6.220 ;
        RECT 121.510 6.020 121.830 6.080 ;
        RECT 51.680 5.880 121.830 6.020 ;
        RECT 121.510 5.820 121.830 5.880 ;
        RECT 52.065 5.680 52.355 5.725 ;
        RECT 26.840 5.540 52.355 5.680 ;
        RECT 26.305 5.340 26.595 5.385 ;
        RECT 26.840 5.340 26.980 5.540 ;
        RECT 52.065 5.495 52.355 5.540 ;
        RECT 52.525 5.680 52.815 5.725 ;
        RECT 169.350 5.680 169.670 5.740 ;
        RECT 52.525 5.540 169.670 5.680 ;
        RECT 196.580 5.680 196.720 6.220 ;
        RECT 394.290 5.680 394.610 5.740 ;
        RECT 196.580 5.540 394.610 5.680 ;
        RECT 52.525 5.495 52.815 5.540 ;
        RECT 169.350 5.480 169.670 5.540 ;
        RECT 394.290 5.480 394.610 5.540 ;
        RECT 518.505 5.680 518.795 5.725 ;
        RECT 519.870 5.680 520.190 5.740 ;
        RECT 518.505 5.540 520.190 5.680 ;
        RECT 518.505 5.495 518.795 5.540 ;
        RECT 519.870 5.480 520.190 5.540 ;
        RECT 26.305 5.200 26.980 5.340 ;
        RECT 365.325 5.340 365.615 5.385 ;
        RECT 365.325 5.200 414.760 5.340 ;
        RECT 26.305 5.155 26.595 5.200 ;
        RECT 365.325 5.155 365.615 5.200 ;
        RECT 414.620 5.000 414.760 5.200 ;
        RECT 417.305 5.000 417.595 5.045 ;
        RECT 414.620 4.860 417.595 5.000 ;
        RECT 417.305 4.815 417.595 4.860 ;
        RECT 16.630 4.660 16.950 4.720 ;
        RECT 283.890 4.660 284.210 4.720 ;
        RECT 16.630 4.520 284.210 4.660 ;
        RECT 16.630 4.460 16.950 4.520 ;
        RECT 283.890 4.460 284.210 4.520 ;
        RECT 212.145 4.320 212.435 4.365 ;
        RECT 233.290 4.320 233.610 4.380 ;
        RECT 212.145 4.180 233.610 4.320 ;
        RECT 212.145 4.135 212.435 4.180 ;
        RECT 233.290 4.120 233.610 4.180 ;
        RECT 4.210 3.640 4.530 3.700 ;
        RECT 26.305 3.640 26.595 3.685 ;
        RECT 4.210 3.500 26.595 3.640 ;
        RECT 4.210 3.440 4.530 3.500 ;
        RECT 26.305 3.455 26.595 3.500 ;
        RECT 36.425 3.300 36.715 3.345 ;
        RECT 26.380 3.160 36.715 3.300 ;
        RECT 25.845 2.960 26.135 3.005 ;
        RECT 26.380 2.960 26.520 3.160 ;
        RECT 36.425 3.115 36.715 3.160 ;
        RECT 25.845 2.820 26.520 2.960 ;
        RECT 52.510 2.960 52.830 3.020 ;
        RECT 67.230 2.960 67.550 3.020 ;
        RECT 52.510 2.820 67.550 2.960 ;
        RECT 25.845 2.775 26.135 2.820 ;
        RECT 52.510 2.760 52.830 2.820 ;
        RECT 67.230 2.760 67.550 2.820 ;
        RECT 18.010 2.620 18.330 2.680 ;
        RECT 29.985 2.620 30.275 2.665 ;
        RECT 18.010 2.480 24.220 2.620 ;
        RECT 18.010 2.420 18.330 2.480 ;
        RECT 5.130 2.280 5.450 2.340 ;
        RECT 23.545 2.280 23.835 2.325 ;
        RECT 5.130 2.140 23.835 2.280 ;
        RECT 24.080 2.280 24.220 2.480 ;
        RECT 25.920 2.480 30.275 2.620 ;
        RECT 25.920 2.280 26.060 2.480 ;
        RECT 29.985 2.435 30.275 2.480 ;
        RECT 24.080 2.140 26.060 2.280 ;
        RECT 5.130 2.080 5.450 2.140 ;
        RECT 23.545 2.095 23.835 2.140 ;
        RECT 448.125 1.940 448.415 1.985 ;
        RECT 453.630 1.940 453.950 2.000 ;
        RECT 448.125 1.800 453.950 1.940 ;
        RECT 448.125 1.755 448.415 1.800 ;
        RECT 453.630 1.740 453.950 1.800 ;
        RECT 134.390 1.600 134.710 1.660 ;
        RECT 175.790 1.600 176.110 1.660 ;
        RECT 134.390 1.460 176.110 1.600 ;
        RECT 134.390 1.400 134.710 1.460 ;
        RECT 175.790 1.400 176.110 1.460 ;
        RECT 29.985 1.260 30.275 1.305 ;
        RECT 52.050 1.260 52.370 1.320 ;
        RECT 29.985 1.120 52.370 1.260 ;
        RECT 29.985 1.075 30.275 1.120 ;
        RECT 52.050 1.060 52.370 1.120 ;
        RECT 249.390 0.920 249.710 0.980 ;
        RECT 293.090 0.920 293.410 0.980 ;
        RECT 249.390 0.780 293.410 0.920 ;
        RECT 249.390 0.720 249.710 0.780 ;
        RECT 293.090 0.720 293.410 0.780 ;
        RECT 422.350 0.920 422.670 0.980 ;
        RECT 422.825 0.920 423.115 0.965 ;
        RECT 422.350 0.780 423.115 0.920 ;
        RECT 422.350 0.720 422.670 0.780 ;
        RECT 422.825 0.735 423.115 0.780 ;
        RECT 27.225 0.580 27.515 0.625 ;
        RECT 26.380 0.440 27.515 0.580 ;
        RECT 8.825 0.240 9.115 0.285 ;
        RECT 26.380 0.240 26.520 0.440 ;
        RECT 27.225 0.395 27.515 0.440 ;
        RECT 28.145 0.580 28.435 0.625 ;
        RECT 28.145 0.440 29.740 0.580 ;
        RECT 28.145 0.395 28.435 0.440 ;
        RECT 8.825 0.100 26.520 0.240 ;
        RECT 29.600 0.240 29.740 0.440 ;
        RECT 65.390 0.240 65.710 0.300 ;
        RECT 29.600 0.100 65.710 0.240 ;
        RECT 8.825 0.055 9.115 0.100 ;
        RECT 65.390 0.040 65.710 0.100 ;
      LAYER via ;
        RECT 1133.540 3401.740 1133.800 3402.000 ;
        RECT 1035.100 3401.400 1035.360 3401.660 ;
        RECT 17.120 3398.680 17.380 3398.940 ;
        RECT 12.520 3398.000 12.780 3398.260 ;
        RECT 1329.500 3401.740 1329.760 3402.000 ;
        RECT 2709.040 3401.740 2709.300 3402.000 ;
        RECT 2807.940 3401.400 2808.200 3401.660 ;
        RECT 18.500 3395.620 18.760 3395.880 ;
        RECT 9.760 3010.400 10.020 3010.660 ;
        RECT 9.760 3005.300 10.020 3005.560 ;
        RECT 7.920 3004.620 8.180 3004.880 ;
        RECT 9.760 3004.620 10.020 3004.880 ;
        RECT 9.760 3002.580 10.020 3002.840 ;
        RECT 9.760 2999.180 10.020 2999.440 ;
        RECT 7.920 2886.300 8.180 2886.560 ;
        RECT 9.760 2886.300 10.020 2886.560 ;
        RECT 9.760 2846.520 10.020 2846.780 ;
        RECT 8.840 2845.500 9.100 2845.760 ;
        RECT 9.760 2822.040 10.020 2822.300 ;
        RECT 6.540 2820.340 6.800 2820.600 ;
        RECT 9.760 2820.340 10.020 2820.600 ;
        RECT 9.760 2816.940 10.020 2817.200 ;
        RECT 9.760 2632.320 10.020 2632.580 ;
        RECT 7.920 2631.640 8.180 2631.900 ;
        RECT 9.760 2631.640 10.020 2631.900 ;
        RECT 9.760 2630.620 10.020 2630.880 ;
        RECT 9.760 2535.760 10.020 2536.020 ;
        RECT 9.760 2530.320 10.020 2530.580 ;
        RECT 7.920 2525.900 8.180 2526.160 ;
        RECT 9.760 2525.900 10.020 2526.160 ;
        RECT 9.760 2523.860 10.020 2524.120 ;
        RECT 9.760 2510.940 10.020 2511.200 ;
        RECT 5.160 2348.760 5.420 2349.020 ;
        RECT 9.760 2348.760 10.020 2349.020 ;
        RECT 9.760 2341.280 10.020 2341.540 ;
        RECT 9.760 2340.260 10.020 2340.520 ;
        RECT 9.760 2249.480 10.020 2249.740 ;
        RECT 9.760 2243.700 10.020 2243.960 ;
        RECT 7.000 2243.020 7.260 2243.280 ;
        RECT 9.760 2243.020 10.020 2243.280 ;
        RECT 9.760 2242.340 10.020 2242.600 ;
        RECT 9.760 2239.620 10.020 2239.880 ;
        RECT 9.760 1670.800 10.020 1671.060 ;
        RECT 9.760 1670.120 10.020 1670.380 ;
        RECT 6.540 1668.420 6.800 1668.680 ;
        RECT 9.760 1668.420 10.020 1668.680 ;
        RECT 9.760 1667.060 10.020 1667.320 ;
        RECT 9.760 1658.900 10.020 1659.160 ;
        RECT 9.760 1575.600 10.020 1575.860 ;
        RECT 9.760 1562.000 10.020 1562.260 ;
        RECT 9.760 1561.320 10.020 1561.580 ;
        RECT 9.760 1560.640 10.020 1560.900 ;
        RECT 9.760 1558.940 10.020 1559.200 ;
        RECT 9.760 1522.560 10.020 1522.820 ;
        RECT 9.760 1520.520 10.020 1520.780 ;
        RECT 9.760 1519.840 10.020 1520.100 ;
        RECT 9.760 1516.780 10.020 1517.040 ;
        RECT 9.760 1466.800 10.020 1467.060 ;
        RECT 9.760 1465.440 10.020 1465.700 ;
        RECT 9.760 1423.620 10.020 1423.880 ;
        RECT 9.760 1422.940 10.020 1423.200 ;
        RECT 9.760 1421.580 10.020 1421.840 ;
        RECT 7.000 1419.540 7.260 1419.800 ;
        RECT 9.760 1320.600 10.020 1320.860 ;
        RECT 9.760 1099.600 10.020 1099.860 ;
        RECT 9.760 1091.440 10.020 1091.700 ;
        RECT 9.760 1088.380 10.020 1088.640 ;
        RECT 7.000 1071.380 7.260 1071.640 ;
        RECT 9.760 1071.380 10.020 1071.640 ;
        RECT 7.000 1024.460 7.260 1024.720 ;
        RECT 9.760 1009.160 10.020 1009.420 ;
        RECT 7.000 991.140 7.260 991.400 ;
        RECT 9.760 990.800 10.020 991.060 ;
        RECT 9.760 988.760 10.020 989.020 ;
        RECT 9.760 988.080 10.020 988.340 ;
        RECT 9.760 981.620 10.020 981.880 ;
        RECT 9.760 980.940 10.020 981.200 ;
        RECT 9.760 978.900 10.020 979.160 ;
        RECT 9.760 973.460 10.020 973.720 ;
        RECT 3.320 969.720 3.580 969.980 ;
        RECT 9.760 947.960 10.020 948.220 ;
        RECT 9.760 943.200 10.020 943.460 ;
        RECT 9.760 942.520 10.020 942.780 ;
        RECT 9.760 883.700 10.020 883.960 ;
        RECT 7.460 865.680 7.720 865.940 ;
        RECT 9.300 865.680 9.560 865.940 ;
        RECT 5.160 836.100 5.420 836.360 ;
        RECT 9.760 832.020 10.020 832.280 ;
        RECT 9.760 831.340 10.020 831.600 ;
        RECT 7.000 829.980 7.260 830.240 ;
        RECT 9.760 829.980 10.020 830.240 ;
        RECT 9.760 829.300 10.020 829.560 ;
        RECT 9.760 827.260 10.020 827.520 ;
        RECT 7.460 799.720 7.720 799.980 ;
        RECT 9.760 799.720 10.020 799.980 ;
        RECT 7.460 798.360 7.720 798.620 ;
        RECT 9.760 798.360 10.020 798.620 ;
        RECT 9.300 768.780 9.560 769.040 ;
        RECT 7.920 735.460 8.180 735.720 ;
        RECT 9.760 735.460 10.020 735.720 ;
        RECT 7.920 731.720 8.180 731.980 ;
        RECT 7.920 714.720 8.180 714.980 ;
        RECT 5.160 714.040 5.420 714.300 ;
        RECT 2.860 708.600 3.120 708.860 ;
        RECT 4.240 708.600 4.500 708.860 ;
        RECT 9.760 705.880 10.020 706.140 ;
        RECT 9.760 699.760 10.020 700.020 ;
        RECT 7.460 692.960 7.720 693.220 ;
        RECT 9.760 692.960 10.020 693.220 ;
        RECT 5.160 672.560 5.420 672.820 ;
        RECT 5.160 666.440 5.420 666.700 ;
        RECT 9.760 660.320 10.020 660.580 ;
        RECT 9.760 654.200 10.020 654.460 ;
        RECT 9.760 652.840 10.020 653.100 ;
        RECT 9.760 647.060 10.020 647.320 ;
        RECT 9.760 645.700 10.020 645.960 ;
        RECT 4.240 644.340 4.500 644.600 ;
        RECT 9.300 641.620 9.560 641.880 ;
        RECT 9.300 631.760 9.560 632.020 ;
        RECT 6.080 587.560 6.340 587.820 ;
        RECT 9.760 587.560 10.020 587.820 ;
        RECT 9.760 586.880 10.020 587.140 ;
        RECT 6.080 575.320 6.340 575.580 ;
        RECT 9.760 554.920 10.020 555.180 ;
        RECT 6.080 550.160 6.340 550.420 ;
        RECT 9.760 550.160 10.020 550.420 ;
        RECT 9.760 548.460 10.020 548.720 ;
        RECT 9.760 547.100 10.020 547.360 ;
        RECT 9.760 546.420 10.020 546.680 ;
        RECT 9.760 545.740 10.020 546.000 ;
        RECT 9.760 544.380 10.020 544.640 ;
        RECT 9.760 543.700 10.020 543.960 ;
        RECT 9.760 543.020 10.020 543.280 ;
        RECT 9.760 542.340 10.020 542.600 ;
        RECT 6.080 540.300 6.340 540.560 ;
        RECT 6.080 512.760 6.340 513.020 ;
        RECT 6.540 491.340 6.800 491.600 ;
        RECT 9.300 467.200 9.560 467.460 ;
        RECT 9.760 466.860 10.020 467.120 ;
        RECT 9.760 466.180 10.020 466.440 ;
        RECT 9.760 460.740 10.020 461.000 ;
        RECT 9.760 460.060 10.020 460.320 ;
        RECT 9.760 459.380 10.020 459.640 ;
        RECT 9.760 457.340 10.020 457.600 ;
        RECT 9.300 430.480 9.560 430.740 ;
        RECT 9.760 423.680 10.020 423.940 ;
        RECT 9.760 417.900 10.020 418.160 ;
        RECT 9.760 410.420 10.020 410.680 ;
        RECT 9.760 359.760 10.020 360.020 ;
        RECT 6.080 355.000 6.340 355.260 ;
        RECT 9.760 355.000 10.020 355.260 ;
        RECT 9.760 337.320 10.020 337.580 ;
        RECT 6.540 336.640 6.800 336.900 ;
        RECT 9.760 336.640 10.020 336.900 ;
        RECT 9.760 335.960 10.020 336.220 ;
        RECT 9.760 333.580 10.020 333.840 ;
        RECT 9.760 332.900 10.020 333.160 ;
        RECT 6.080 327.120 6.340 327.380 ;
        RECT 10.220 327.120 10.480 327.380 ;
        RECT 6.540 326.100 6.800 326.360 ;
        RECT 9.760 323.040 10.020 323.300 ;
        RECT 6.080 316.580 6.340 316.840 ;
        RECT 9.760 316.580 10.020 316.840 ;
        RECT 9.760 315.560 10.020 315.820 ;
        RECT 9.760 314.200 10.020 314.460 ;
        RECT 9.760 311.140 10.020 311.400 ;
        RECT 6.540 289.380 6.800 289.640 ;
        RECT 9.760 285.300 10.020 285.560 ;
        RECT 9.760 284.280 10.020 284.540 ;
        RECT 9.760 282.920 10.020 283.180 ;
        RECT 9.760 279.180 10.020 279.440 ;
        RECT 9.760 262.860 10.020 263.120 ;
        RECT 5.160 251.640 5.420 251.900 ;
        RECT 5.160 185.000 5.420 185.260 ;
        RECT 9.760 177.520 10.020 177.780 ;
        RECT 9.300 148.620 9.560 148.880 ;
        RECT 7.460 147.260 7.720 147.520 ;
        RECT 9.760 141.480 10.020 141.740 ;
        RECT 7.460 139.780 7.720 140.040 ;
        RECT 9.760 139.780 10.020 140.040 ;
        RECT 9.760 136.040 10.020 136.300 ;
        RECT 9.760 135.360 10.020 135.620 ;
        RECT 6.080 134.680 6.340 134.940 ;
        RECT 9.760 134.680 10.020 134.940 ;
        RECT 7.460 134.000 7.720 134.260 ;
        RECT 9.760 134.000 10.020 134.260 ;
        RECT 9.760 110.880 10.020 111.140 ;
        RECT 5.160 100.000 5.420 100.260 ;
        RECT 6.540 94.220 6.800 94.480 ;
        RECT 9.300 89.460 9.560 89.720 ;
        RECT 9.300 82.660 9.560 82.920 ;
        RECT 9.300 81.980 9.560 82.240 ;
        RECT 5.620 77.900 5.880 78.160 ;
        RECT 9.760 77.900 10.020 78.160 ;
        RECT 9.760 76.540 10.020 76.800 ;
        RECT 9.760 75.520 10.020 75.780 ;
        RECT 5.620 73.820 5.880 74.080 ;
        RECT 9.760 67.360 10.020 67.620 ;
        RECT 9.760 66.680 10.020 66.940 ;
        RECT 5.620 61.580 5.880 61.840 ;
        RECT 6.540 60.900 6.800 61.160 ;
        RECT 5.160 50.360 5.420 50.620 ;
        RECT 4.240 37.440 4.500 37.700 ;
        RECT 6.080 16.360 6.340 16.620 ;
        RECT 18.960 8.540 19.220 8.800 ;
        RECT 38.280 8.540 38.540 8.800 ;
        RECT 283.920 8.200 284.180 8.460 ;
        RECT 90.260 7.520 90.520 7.780 ;
        RECT 29.540 6.840 29.800 7.100 ;
        RECT 32.300 6.840 32.560 7.100 ;
        RECT 24.940 6.500 25.200 6.760 ;
        RECT 26.780 6.500 27.040 6.760 ;
        RECT 72.780 6.500 73.040 6.760 ;
        RECT 90.260 6.500 90.520 6.760 ;
        RECT 121.540 5.820 121.800 6.080 ;
        RECT 169.380 5.480 169.640 5.740 ;
        RECT 394.320 5.480 394.580 5.740 ;
        RECT 519.900 5.480 520.160 5.740 ;
        RECT 16.660 4.460 16.920 4.720 ;
        RECT 283.920 4.460 284.180 4.720 ;
        RECT 233.320 4.120 233.580 4.380 ;
        RECT 4.240 3.440 4.500 3.700 ;
        RECT 52.540 2.760 52.800 3.020 ;
        RECT 67.260 2.760 67.520 3.020 ;
        RECT 18.040 2.420 18.300 2.680 ;
        RECT 5.160 2.080 5.420 2.340 ;
        RECT 453.660 1.740 453.920 2.000 ;
        RECT 134.420 1.400 134.680 1.660 ;
        RECT 175.820 1.400 176.080 1.660 ;
        RECT 52.080 1.060 52.340 1.320 ;
        RECT 249.420 0.720 249.680 0.980 ;
        RECT 293.120 0.720 293.380 0.980 ;
        RECT 422.380 0.720 422.640 0.980 ;
        RECT 65.420 0.040 65.680 0.300 ;
      LAYER met2 ;
        RECT 1036.410 3401.770 1036.690 3405.000 ;
        RECT 1035.160 3401.690 1036.690 3401.770 ;
        RECT 1133.540 3401.770 1133.800 3402.030 ;
        RECT 1134.850 3401.770 1135.130 3405.000 ;
        RECT 1133.540 3401.710 1135.130 3401.770 ;
        RECT 1329.500 3401.770 1329.760 3402.030 ;
        RECT 1331.270 3401.770 1331.550 3405.000 ;
        RECT 1329.500 3401.710 1331.550 3401.770 ;
        RECT 1035.100 3401.630 1036.690 3401.690 ;
        RECT 1133.600 3401.630 1135.130 3401.710 ;
        RECT 1329.560 3401.630 1331.550 3401.710 ;
        RECT 1035.100 3401.370 1035.360 3401.630 ;
        RECT 1036.410 3401.000 1036.690 3401.630 ;
        RECT 1134.850 3401.000 1135.130 3401.630 ;
        RECT 1331.270 3401.000 1331.550 3401.630 ;
        RECT 2707.130 3401.770 2707.410 3405.000 ;
        RECT 2709.040 3401.770 2709.300 3402.030 ;
        RECT 2707.130 3401.710 2709.300 3401.770 ;
        RECT 2805.570 3401.770 2805.850 3405.000 ;
        RECT 2807.930 3402.195 2808.210 3402.565 ;
        RECT 2806.090 3401.770 2806.370 3401.885 ;
        RECT 2707.130 3401.630 2709.240 3401.710 ;
        RECT 2805.570 3401.630 2806.370 3401.770 ;
        RECT 2808.000 3401.690 2808.140 3402.195 ;
        RECT 2707.130 3401.000 2707.410 3401.630 ;
        RECT 2805.570 3401.000 2805.850 3401.630 ;
        RECT 2806.090 3401.515 2806.370 3401.630 ;
        RECT 2807.940 3401.370 2808.200 3401.690 ;
        RECT 17.120 3398.650 17.380 3398.970 ;
        RECT 12.520 3397.970 12.780 3398.290 ;
        RECT 12.580 3385.450 12.720 3397.970 ;
        RECT 11.660 3385.310 12.720 3385.450 ;
        RECT 11.660 3263.730 11.800 3385.310 ;
        RECT 17.180 3275.970 17.320 3398.650 ;
        RECT 18.500 3395.590 18.760 3395.910 ;
        RECT 18.560 3381.370 18.700 3395.590 ;
        RECT 18.560 3381.230 19.160 3381.370 ;
        RECT 19.020 3333.090 19.160 3381.230 ;
        RECT 18.100 3332.950 19.160 3333.090 ;
        RECT 18.100 3298.410 18.240 3332.950 ;
        RECT 18.100 3298.270 19.160 3298.410 ;
        RECT 16.720 3275.830 17.320 3275.970 ;
        RECT 16.720 3267.130 16.860 3275.830 ;
        RECT 16.720 3266.990 17.780 3267.130 ;
        RECT 11.660 3263.590 12.720 3263.730 ;
        RECT 12.580 3208.650 12.720 3263.590 ;
        RECT 17.640 3243.330 17.780 3266.990 ;
        RECT 19.020 3243.330 19.160 3298.270 ;
        RECT 17.640 3243.190 18.240 3243.330 ;
        RECT 9.360 3208.510 12.720 3208.650 ;
        RECT 9.360 3205.250 9.500 3208.510 ;
        RECT 9.360 3205.110 10.880 3205.250 ;
        RECT 10.740 3163.090 10.880 3205.110 ;
        RECT 18.100 3195.730 18.240 3243.190 ;
        RECT 17.180 3195.590 18.240 3195.730 ;
        RECT 18.560 3243.190 19.160 3243.330 ;
        RECT 17.180 3195.050 17.320 3195.590 ;
        RECT 16.720 3194.910 17.320 3195.050 ;
        RECT 16.720 3177.370 16.860 3194.910 ;
        RECT 15.340 3177.230 16.860 3177.370 ;
        RECT 10.740 3162.950 11.800 3163.090 ;
        RECT 11.660 3010.770 11.800 3162.950 ;
        RECT 15.340 3114.130 15.480 3177.230 ;
        RECT 18.560 3173.290 18.700 3243.190 ;
        RECT 18.100 3173.150 18.700 3173.290 ;
        RECT 18.100 3118.890 18.240 3173.150 ;
        RECT 17.640 3118.750 18.240 3118.890 ;
        RECT 15.340 3113.990 16.860 3114.130 ;
        RECT 9.820 3010.690 11.800 3010.770 ;
        RECT 9.760 3010.630 11.800 3010.690 ;
        RECT 9.760 3010.370 10.020 3010.630 ;
        RECT 16.720 3009.410 16.860 3113.990 ;
        RECT 17.640 3067.890 17.780 3118.750 ;
        RECT 17.640 3067.750 18.700 3067.890 ;
        RECT 18.560 3063.810 18.700 3067.750 ;
        RECT 18.560 3063.670 19.160 3063.810 ;
        RECT 19.020 3012.130 19.160 3063.670 ;
        RECT 9.820 3009.270 16.860 3009.410 ;
        RECT 18.100 3011.990 19.160 3012.130 ;
        RECT 9.820 3005.590 9.960 3009.270 ;
        RECT 7.910 3005.075 8.190 3005.445 ;
        RECT 9.760 3005.270 10.020 3005.590 ;
        RECT 7.980 3004.910 8.120 3005.075 ;
        RECT 7.920 3004.590 8.180 3004.910 ;
        RECT 9.760 3004.820 10.020 3004.910 ;
        RECT 9.760 3004.680 10.880 3004.820 ;
        RECT 9.760 3004.590 10.020 3004.680 ;
        RECT 10.740 3003.970 10.880 3004.680 ;
        RECT 10.740 3003.830 12.720 3003.970 ;
        RECT 12.580 3003.290 12.720 3003.830 ;
        RECT 14.880 3003.830 16.860 3003.970 ;
        RECT 14.880 3003.290 15.020 3003.830 ;
        RECT 12.580 3003.150 15.020 3003.290 ;
        RECT 9.760 3002.610 10.020 3002.870 ;
        RECT 9.760 3002.550 11.800 3002.610 ;
        RECT 9.820 3002.470 11.800 3002.550 ;
        RECT 11.660 2999.890 11.800 3002.470 ;
        RECT 11.660 2999.750 13.640 2999.890 ;
        RECT 9.760 2999.380 10.020 2999.470 ;
        RECT 9.760 2999.240 13.180 2999.380 ;
        RECT 9.760 2999.150 10.020 2999.240 ;
        RECT 13.040 2994.450 13.180 2999.240 ;
        RECT 12.580 2994.310 13.180 2994.450 ;
        RECT 12.580 2967.250 12.720 2994.310 ;
        RECT 13.500 2990.370 13.640 2999.750 ;
        RECT 13.500 2990.230 14.100 2990.370 ;
        RECT 12.580 2967.110 13.640 2967.250 ;
        RECT 7.910 2891.515 8.190 2891.885 ;
        RECT 7.980 2886.590 8.120 2891.515 ;
        RECT 7.920 2886.270 8.180 2886.590 ;
        RECT 9.760 2886.500 10.020 2886.590 ;
        RECT 9.760 2886.360 13.180 2886.500 ;
        RECT 9.760 2886.270 10.020 2886.360 ;
        RECT 9.820 2846.810 11.340 2846.890 ;
        RECT 9.760 2846.750 11.340 2846.810 ;
        RECT 9.760 2846.490 10.020 2846.750 ;
        RECT 11.200 2846.210 11.340 2846.750 ;
        RECT 13.040 2846.210 13.180 2886.360 ;
        RECT 11.200 2846.070 13.180 2846.210 ;
        RECT 8.840 2845.470 9.100 2845.790 ;
        RECT 6.530 2836.435 6.810 2836.805 ;
        RECT 6.600 2820.630 6.740 2836.435 ;
        RECT 6.540 2820.310 6.800 2820.630 ;
        RECT 8.900 2817.650 9.040 2845.470 ;
        RECT 13.500 2827.170 13.640 2967.110 ;
        RECT 13.960 2898.570 14.100 2990.230 ;
        RECT 16.720 2974.050 16.860 3003.830 ;
        RECT 16.260 2973.910 16.860 2974.050 ;
        RECT 16.260 2964.530 16.400 2973.910 ;
        RECT 16.260 2964.390 17.320 2964.530 ;
        RECT 13.960 2898.430 14.560 2898.570 ;
        RECT 14.420 2897.890 14.560 2898.430 ;
        RECT 14.420 2897.750 15.940 2897.890 ;
        RECT 15.800 2883.610 15.940 2897.750 ;
        RECT 15.340 2883.470 15.940 2883.610 ;
        RECT 15.340 2882.930 15.480 2883.470 ;
        RECT 14.880 2882.790 15.480 2882.930 ;
        RECT 14.880 2861.850 15.020 2882.790 ;
        RECT 17.180 2861.850 17.320 2964.390 ;
        RECT 18.100 2959.940 18.240 3011.990 ;
        RECT 18.100 2959.800 18.700 2959.940 ;
        RECT 18.560 2959.090 18.700 2959.800 ;
        RECT 18.560 2958.950 19.160 2959.090 ;
        RECT 14.420 2861.710 15.020 2861.850 ;
        RECT 16.260 2861.710 17.320 2861.850 ;
        RECT 14.420 2852.330 14.560 2861.710 ;
        RECT 16.260 2853.690 16.400 2861.710 ;
        RECT 15.340 2853.550 16.400 2853.690 ;
        RECT 14.420 2852.190 15.020 2852.330 ;
        RECT 14.880 2850.290 15.020 2852.190 ;
        RECT 15.340 2850.970 15.480 2853.550 ;
        RECT 15.340 2850.830 15.940 2850.970 ;
        RECT 15.800 2850.290 15.940 2850.830 ;
        RECT 14.880 2850.150 18.700 2850.290 ;
        RECT 15.800 2829.890 15.940 2850.150 ;
        RECT 15.800 2829.750 16.860 2829.890 ;
        RECT 9.820 2827.030 13.640 2827.170 ;
        RECT 9.820 2822.330 9.960 2827.030 ;
        RECT 9.760 2822.010 10.020 2822.330 ;
        RECT 9.760 2820.370 10.020 2820.630 ;
        RECT 9.760 2820.310 13.640 2820.370 ;
        RECT 9.820 2820.230 13.640 2820.310 ;
        RECT 8.900 2817.510 12.720 2817.650 ;
        RECT 9.760 2816.910 10.020 2817.230 ;
        RECT 9.820 2816.290 9.960 2816.910 ;
        RECT 9.820 2816.150 12.260 2816.290 ;
        RECT 12.120 2683.690 12.260 2816.150 ;
        RECT 12.580 2753.730 12.720 2817.510 ;
        RECT 13.500 2774.130 13.640 2820.230 ;
        RECT 13.500 2773.990 15.480 2774.130 ;
        RECT 12.580 2753.590 15.020 2753.730 ;
        RECT 14.880 2752.370 15.020 2753.590 ;
        RECT 15.340 2753.050 15.480 2773.990 ;
        RECT 15.340 2752.910 16.400 2753.050 ;
        RECT 11.660 2683.550 12.260 2683.690 ;
        RECT 13.960 2752.230 15.020 2752.370 ;
        RECT 7.910 2665.075 8.190 2665.445 ;
        RECT 7.980 2631.930 8.120 2665.075 ;
        RECT 11.660 2632.690 11.800 2683.550 ;
        RECT 9.820 2632.610 11.800 2632.690 ;
        RECT 9.760 2632.550 11.800 2632.610 ;
        RECT 9.760 2632.290 10.020 2632.550 ;
        RECT 9.820 2631.930 13.640 2632.010 ;
        RECT 7.920 2631.610 8.180 2631.930 ;
        RECT 9.760 2631.870 13.640 2631.930 ;
        RECT 9.760 2631.610 10.020 2631.870 ;
        RECT 9.760 2630.650 10.020 2630.910 ;
        RECT 9.760 2630.590 12.720 2630.650 ;
        RECT 9.820 2630.510 12.720 2630.590 ;
        RECT 12.580 2574.210 12.720 2630.510 ;
        RECT 13.500 2581.010 13.640 2631.870 ;
        RECT 11.660 2574.070 12.720 2574.210 ;
        RECT 13.040 2580.870 13.640 2581.010 ;
        RECT 7.910 2549.475 8.190 2549.845 ;
        RECT 7.980 2526.190 8.120 2549.475 ;
        RECT 11.660 2536.130 11.800 2574.070 ;
        RECT 9.820 2536.050 11.800 2536.130 ;
        RECT 9.760 2535.990 11.800 2536.050 ;
        RECT 9.760 2535.730 10.020 2535.990 ;
        RECT 13.040 2532.730 13.180 2580.870 ;
        RECT 9.820 2532.590 13.180 2532.730 ;
        RECT 9.820 2530.610 9.960 2532.590 ;
        RECT 9.760 2530.290 10.020 2530.610 ;
        RECT 13.960 2527.290 14.100 2752.230 ;
        RECT 16.260 2728.570 16.400 2752.910 ;
        RECT 15.340 2728.430 16.400 2728.570 ;
        RECT 15.340 2553.810 15.480 2728.430 ;
        RECT 15.340 2553.670 16.400 2553.810 ;
        RECT 9.360 2527.150 14.100 2527.290 ;
        RECT 7.920 2525.870 8.180 2526.190 ;
        RECT 9.360 2524.570 9.500 2527.150 ;
        RECT 9.760 2525.930 10.020 2526.190 ;
        RECT 9.760 2525.870 15.020 2525.930 ;
        RECT 9.820 2525.790 15.020 2525.870 ;
        RECT 9.360 2524.430 14.100 2524.570 ;
        RECT 9.760 2524.060 10.020 2524.150 ;
        RECT 9.760 2523.920 10.420 2524.060 ;
        RECT 9.760 2523.830 10.020 2523.920 ;
        RECT 9.760 2510.910 10.020 2511.230 ;
        RECT 9.820 2509.610 9.960 2510.910 ;
        RECT 10.280 2510.290 10.420 2523.920 ;
        RECT 10.280 2510.150 13.640 2510.290 ;
        RECT 9.820 2509.470 12.720 2509.610 ;
        RECT 12.580 2444.330 12.720 2509.470 ;
        RECT 13.500 2445.010 13.640 2510.150 ;
        RECT 13.960 2446.370 14.100 2524.430 ;
        RECT 14.880 2476.970 15.020 2525.790 ;
        RECT 14.880 2476.830 15.480 2476.970 ;
        RECT 13.960 2446.230 15.020 2446.370 ;
        RECT 14.880 2445.010 15.020 2446.230 ;
        RECT 15.340 2445.690 15.480 2476.830 ;
        RECT 16.260 2446.370 16.400 2553.670 ;
        RECT 15.800 2446.230 16.400 2446.370 ;
        RECT 15.800 2445.690 15.940 2446.230 ;
        RECT 15.340 2445.550 16.400 2445.690 ;
        RECT 13.500 2444.870 15.020 2445.010 ;
        RECT 14.880 2444.330 15.020 2444.870 ;
        RECT 11.660 2444.190 15.020 2444.330 ;
        RECT 11.660 2362.050 11.800 2444.190 ;
        RECT 12.580 2438.890 12.720 2444.190 ;
        RECT 14.880 2442.970 15.020 2444.190 ;
        RECT 14.420 2442.830 15.020 2442.970 ;
        RECT 12.580 2438.750 13.180 2438.890 ;
        RECT 13.040 2390.610 13.180 2438.750 ;
        RECT 14.420 2414.410 14.560 2442.830 ;
        RECT 15.800 2439.570 15.940 2445.550 ;
        RECT 14.880 2439.430 15.940 2439.570 ;
        RECT 14.880 2435.490 15.020 2439.430 ;
        RECT 14.880 2435.350 15.480 2435.490 ;
        RECT 15.340 2415.090 15.480 2435.350 ;
        RECT 15.340 2414.950 15.940 2415.090 ;
        RECT 13.500 2414.270 14.560 2414.410 ;
        RECT 13.500 2391.290 13.640 2414.270 ;
        RECT 15.800 2412.370 15.940 2414.950 ;
        RECT 15.340 2412.230 15.940 2412.370 ;
        RECT 13.500 2391.150 15.020 2391.290 ;
        RECT 13.040 2390.470 13.640 2390.610 ;
        RECT 9.360 2361.910 11.800 2362.050 ;
        RECT 5.160 2348.730 5.420 2349.050 ;
        RECT 3.320 969.690 3.580 970.010 ;
        RECT 3.380 730.730 3.520 969.690 ;
        RECT 5.220 836.390 5.360 2348.730 ;
        RECT 9.360 2340.970 9.500 2361.910 ;
        RECT 13.500 2361.370 13.640 2390.470 ;
        RECT 14.880 2366.810 15.020 2391.150 ;
        RECT 9.820 2361.230 13.640 2361.370 ;
        RECT 13.960 2366.670 15.020 2366.810 ;
        RECT 9.820 2349.050 9.960 2361.230 ;
        RECT 13.960 2360.690 14.100 2366.670 ;
        RECT 12.120 2360.550 14.100 2360.690 ;
        RECT 12.120 2349.810 12.260 2360.550 ;
        RECT 10.280 2349.670 12.260 2349.810 ;
        RECT 9.760 2348.730 10.020 2349.050 ;
        RECT 10.280 2341.650 10.420 2349.670 ;
        RECT 9.820 2341.570 10.420 2341.650 ;
        RECT 9.760 2341.510 10.420 2341.570 ;
        RECT 10.740 2341.510 14.100 2341.650 ;
        RECT 9.760 2341.250 10.020 2341.510 ;
        RECT 10.740 2340.970 10.880 2341.510 ;
        RECT 9.360 2340.830 10.880 2340.970 ;
        RECT 9.760 2340.290 10.020 2340.550 ;
        RECT 9.760 2340.230 12.260 2340.290 ;
        RECT 9.820 2340.150 12.260 2340.230 ;
        RECT 12.120 2335.530 12.260 2340.150 ;
        RECT 11.660 2335.390 12.260 2335.530 ;
        RECT 6.990 2261.835 7.270 2262.205 ;
        RECT 7.060 2243.310 7.200 2261.835 ;
        RECT 11.660 2249.850 11.800 2335.390 ;
        RECT 13.960 2300.170 14.100 2341.510 ;
        RECT 15.340 2315.130 15.480 2412.230 ;
        RECT 16.260 2370.890 16.400 2445.550 ;
        RECT 12.580 2300.030 14.100 2300.170 ;
        RECT 14.880 2314.990 15.480 2315.130 ;
        RECT 15.800 2370.750 16.400 2370.890 ;
        RECT 12.580 2270.250 12.720 2300.030 ;
        RECT 9.820 2249.770 11.800 2249.850 ;
        RECT 9.760 2249.710 11.800 2249.770 ;
        RECT 12.120 2270.110 12.720 2270.250 ;
        RECT 9.760 2249.450 10.020 2249.710 ;
        RECT 12.120 2249.170 12.260 2270.110 ;
        RECT 14.880 2256.650 15.020 2314.990 ;
        RECT 15.800 2276.370 15.940 2370.750 ;
        RECT 16.720 2370.380 16.860 2829.750 ;
        RECT 18.560 2774.130 18.700 2850.150 ;
        RECT 18.100 2773.990 18.700 2774.130 ;
        RECT 18.100 2729.250 18.240 2773.990 ;
        RECT 19.020 2746.250 19.160 2958.950 ;
        RECT 17.180 2729.110 18.240 2729.250 ;
        RECT 18.560 2746.110 19.160 2746.250 ;
        RECT 17.180 2683.690 17.320 2729.110 ;
        RECT 17.180 2683.550 18.240 2683.690 ;
        RECT 18.100 2632.520 18.240 2683.550 ;
        RECT 18.560 2670.090 18.700 2746.110 ;
        RECT 18.560 2669.950 19.160 2670.090 ;
        RECT 17.180 2632.380 18.240 2632.520 ;
        RECT 17.180 2608.210 17.320 2632.380 ;
        RECT 17.180 2608.070 18.240 2608.210 ;
        RECT 18.100 2560.610 18.240 2608.070 ;
        RECT 17.180 2560.470 18.240 2560.610 ;
        RECT 17.180 2487.850 17.320 2560.470 ;
        RECT 17.180 2487.710 18.700 2487.850 ;
        RECT 18.560 2435.490 18.700 2487.710 ;
        RECT 18.100 2435.350 18.700 2435.490 ;
        RECT 18.100 2415.090 18.240 2435.350 ;
        RECT 17.640 2414.950 18.240 2415.090 ;
        RECT 17.640 2394.690 17.780 2414.950 ;
        RECT 17.180 2394.550 17.780 2394.690 ;
        RECT 17.180 2374.290 17.320 2394.550 ;
        RECT 17.180 2374.150 18.700 2374.290 ;
        RECT 16.720 2370.240 17.320 2370.380 ;
        RECT 17.180 2369.530 17.320 2370.240 ;
        RECT 16.720 2369.390 17.320 2369.530 ;
        RECT 15.800 2276.230 16.400 2276.370 ;
        RECT 14.880 2256.510 15.940 2256.650 ;
        RECT 15.800 2255.970 15.940 2256.510 ;
        RECT 16.260 2255.970 16.400 2276.230 ;
        RECT 14.880 2255.830 16.400 2255.970 ;
        RECT 14.880 2253.760 15.020 2255.830 ;
        RECT 9.820 2249.030 12.260 2249.170 ;
        RECT 13.500 2253.620 15.020 2253.760 ;
        RECT 9.820 2243.990 9.960 2249.030 ;
        RECT 9.760 2243.670 10.020 2243.990 ;
        RECT 7.000 2242.990 7.260 2243.310 ;
        RECT 9.760 2243.220 10.020 2243.310 ;
        RECT 9.760 2243.080 11.800 2243.220 ;
        RECT 9.760 2242.990 10.020 2243.080 ;
        RECT 9.760 2242.540 10.020 2242.630 ;
        RECT 9.760 2242.400 10.880 2242.540 ;
        RECT 9.760 2242.310 10.020 2242.400 ;
        RECT 9.760 2239.820 10.020 2239.910 ;
        RECT 9.760 2239.680 10.420 2239.820 ;
        RECT 9.760 2239.590 10.020 2239.680 ;
        RECT 10.280 2223.330 10.420 2239.680 ;
        RECT 10.740 2224.010 10.880 2242.400 ;
        RECT 11.660 2224.690 11.800 2243.080 ;
        RECT 11.660 2224.550 13.180 2224.690 ;
        RECT 10.740 2223.870 12.720 2224.010 ;
        RECT 10.280 2223.190 12.260 2223.330 ;
        RECT 12.120 2045.850 12.260 2223.190 ;
        RECT 12.580 2207.690 12.720 2223.870 ;
        RECT 13.040 2208.370 13.180 2224.550 ;
        RECT 13.500 2219.930 13.640 2253.620 ;
        RECT 15.800 2253.250 15.940 2255.830 ;
        RECT 15.340 2253.110 15.940 2253.250 ;
        RECT 13.500 2219.790 14.560 2219.930 ;
        RECT 13.040 2208.230 13.640 2208.370 ;
        RECT 12.580 2207.550 13.180 2207.690 ;
        RECT 13.040 2097.530 13.180 2207.550 ;
        RECT 13.500 2196.810 13.640 2208.230 ;
        RECT 13.500 2196.670 14.100 2196.810 ;
        RECT 13.960 2122.010 14.100 2196.670 ;
        RECT 14.420 2123.370 14.560 2219.790 ;
        RECT 15.340 2196.130 15.480 2253.110 ;
        RECT 16.720 2240.330 16.860 2369.390 ;
        RECT 18.560 2317.850 18.700 2374.150 ;
        RECT 17.180 2317.710 18.700 2317.850 ;
        RECT 17.180 2297.450 17.320 2317.710 ;
        RECT 17.180 2297.310 18.700 2297.450 ;
        RECT 18.560 2270.250 18.700 2297.310 ;
        RECT 17.180 2270.110 18.700 2270.250 ;
        RECT 17.180 2241.690 17.320 2270.110 ;
        RECT 19.020 2269.570 19.160 2669.950 ;
        RECT 18.100 2269.430 19.160 2269.570 ;
        RECT 18.100 2249.170 18.240 2269.430 ;
        RECT 18.100 2249.030 19.160 2249.170 ;
        RECT 17.180 2241.550 18.700 2241.690 ;
        RECT 16.720 2240.190 17.780 2240.330 ;
        RECT 17.640 2238.290 17.780 2240.190 ;
        RECT 17.180 2238.150 17.780 2238.290 ;
        RECT 17.180 2197.490 17.320 2238.150 ;
        RECT 18.560 2224.690 18.700 2241.550 ;
        RECT 17.640 2224.550 18.700 2224.690 ;
        RECT 17.640 2198.170 17.780 2224.550 ;
        RECT 17.640 2198.030 18.700 2198.170 ;
        RECT 17.180 2197.350 17.780 2197.490 ;
        RECT 15.340 2195.990 17.320 2196.130 ;
        RECT 14.420 2123.230 15.480 2123.370 ;
        RECT 13.960 2121.870 14.560 2122.010 ;
        RECT 11.660 2045.710 12.260 2045.850 ;
        RECT 12.580 2097.390 13.180 2097.530 ;
        RECT 11.660 1990.090 11.800 2045.710 ;
        RECT 12.580 1997.570 12.720 2097.390 ;
        RECT 14.420 2083.250 14.560 2121.870 ;
        RECT 15.340 2113.170 15.480 2123.230 ;
        RECT 17.180 2113.170 17.320 2195.990 ;
        RECT 14.880 2113.030 17.320 2113.170 ;
        RECT 14.880 2083.250 15.020 2113.030 ;
        RECT 15.340 2083.930 15.480 2113.030 ;
        RECT 17.640 2111.810 17.780 2197.350 ;
        RECT 17.180 2111.670 17.780 2111.810 ;
        RECT 17.180 2110.450 17.320 2111.670 ;
        RECT 18.560 2110.450 18.700 2198.030 ;
        RECT 16.720 2110.310 17.320 2110.450 ;
        RECT 17.640 2110.310 18.700 2110.450 ;
        RECT 15.340 2083.790 16.400 2083.930 ;
        RECT 14.420 2083.110 15.480 2083.250 ;
        RECT 14.880 2081.890 15.020 2083.110 ;
        RECT 13.040 2081.750 15.020 2081.890 ;
        RECT 13.040 1998.250 13.180 2081.750 ;
        RECT 15.340 2067.610 15.480 2083.110 ;
        RECT 16.260 2076.450 16.400 2083.790 ;
        RECT 15.800 2076.310 16.400 2076.450 ;
        RECT 15.800 2068.290 15.940 2076.310 ;
        RECT 16.720 2069.650 16.860 2110.310 ;
        RECT 17.640 2109.770 17.780 2110.310 ;
        RECT 17.180 2109.630 17.780 2109.770 ;
        RECT 17.180 2071.010 17.320 2109.630 ;
        RECT 17.180 2070.870 18.700 2071.010 ;
        RECT 16.720 2069.510 17.780 2069.650 ;
        RECT 15.800 2068.150 17.320 2068.290 ;
        RECT 14.880 2067.470 15.480 2067.610 ;
        RECT 13.040 1998.110 13.640 1998.250 ;
        RECT 13.500 1997.570 13.640 1998.110 ;
        RECT 12.580 1997.430 13.180 1997.570 ;
        RECT 13.500 1997.430 14.560 1997.570 ;
        RECT 13.040 1996.890 13.180 1997.430 ;
        RECT 13.040 1996.750 13.640 1996.890 ;
        RECT 11.660 1989.950 12.260 1990.090 ;
        RECT 12.120 1934.330 12.260 1989.950 ;
        RECT 13.500 1973.770 13.640 1996.750 ;
        RECT 10.280 1934.190 12.260 1934.330 ;
        RECT 12.580 1973.630 13.640 1973.770 ;
        RECT 10.280 1911.890 10.420 1934.190 ;
        RECT 12.580 1932.970 12.720 1973.630 ;
        RECT 14.420 1973.090 14.560 1997.430 ;
        RECT 10.740 1932.830 12.720 1932.970 ;
        RECT 13.040 1972.950 14.560 1973.090 ;
        RECT 14.880 1973.090 15.020 2067.470 ;
        RECT 17.180 2022.050 17.320 2068.150 ;
        RECT 15.340 2021.910 17.320 2022.050 ;
        RECT 15.340 1973.770 15.480 2021.910 ;
        RECT 17.640 2013.890 17.780 2069.510 ;
        RECT 16.720 2013.750 17.780 2013.890 ;
        RECT 16.720 2001.650 16.860 2013.750 ;
        RECT 16.720 2001.510 17.780 2001.650 ;
        RECT 17.640 1999.610 17.780 2001.510 ;
        RECT 16.720 1999.470 17.780 1999.610 ;
        RECT 16.720 1979.890 16.860 1999.470 ;
        RECT 16.720 1979.750 17.780 1979.890 ;
        RECT 15.340 1973.630 16.860 1973.770 ;
        RECT 14.880 1972.950 15.940 1973.090 ;
        RECT 10.740 1912.570 10.880 1932.830 ;
        RECT 13.040 1932.290 13.180 1972.950 ;
        RECT 15.800 1971.730 15.940 1972.950 ;
        RECT 15.340 1971.590 15.940 1971.730 ;
        RECT 15.340 1970.370 15.480 1971.590 ;
        RECT 14.880 1970.230 15.480 1970.370 ;
        RECT 14.880 1956.090 15.020 1970.230 ;
        RECT 16.720 1969.860 16.860 1973.630 ;
        RECT 15.800 1969.720 16.860 1969.860 ;
        RECT 14.880 1955.950 15.480 1956.090 ;
        RECT 11.660 1932.150 13.180 1932.290 ;
        RECT 11.660 1913.250 11.800 1932.150 ;
        RECT 15.340 1931.610 15.480 1955.950 ;
        RECT 14.420 1931.470 15.480 1931.610 ;
        RECT 15.800 1931.610 15.940 1969.720 ;
        RECT 17.640 1934.840 17.780 1979.750 ;
        RECT 17.640 1934.700 18.240 1934.840 ;
        RECT 15.800 1931.470 16.400 1931.610 ;
        RECT 14.420 1930.930 14.560 1931.470 ;
        RECT 13.500 1930.790 14.560 1930.930 ;
        RECT 13.500 1914.610 13.640 1930.790 ;
        RECT 16.260 1928.890 16.400 1931.470 ;
        RECT 15.340 1928.750 16.400 1928.890 ;
        RECT 15.340 1927.530 15.480 1928.750 ;
        RECT 15.340 1927.390 16.400 1927.530 ;
        RECT 16.260 1925.490 16.400 1927.390 ;
        RECT 16.260 1925.350 17.320 1925.490 ;
        RECT 13.500 1914.470 15.020 1914.610 ;
        RECT 11.660 1913.110 14.560 1913.250 ;
        RECT 10.740 1912.430 14.100 1912.570 ;
        RECT 10.280 1911.750 13.180 1911.890 ;
        RECT 13.040 1841.170 13.180 1911.750 ;
        RECT 13.960 1852.560 14.100 1912.430 ;
        RECT 11.200 1841.030 13.180 1841.170 ;
        RECT 13.500 1852.420 14.100 1852.560 ;
        RECT 11.200 1735.090 11.340 1841.030 ;
        RECT 13.500 1824.850 13.640 1852.420 ;
        RECT 12.580 1824.710 13.640 1824.850 ;
        RECT 12.580 1822.130 12.720 1824.710 ;
        RECT 14.420 1824.170 14.560 1913.110 ;
        RECT 13.960 1824.030 14.560 1824.170 ;
        RECT 13.960 1822.130 14.100 1824.030 ;
        RECT 12.580 1821.990 14.560 1822.130 ;
        RECT 13.960 1819.410 14.100 1821.990 ;
        RECT 11.660 1819.270 14.100 1819.410 ;
        RECT 11.660 1815.330 11.800 1819.270 ;
        RECT 14.420 1816.690 14.560 1821.990 ;
        RECT 14.880 1817.370 15.020 1914.470 ;
        RECT 17.180 1913.250 17.320 1925.350 ;
        RECT 16.720 1913.110 17.320 1913.250 ;
        RECT 16.720 1890.130 16.860 1913.110 ;
        RECT 15.340 1889.990 16.860 1890.130 ;
        RECT 15.340 1824.850 15.480 1889.990 ;
        RECT 18.100 1881.290 18.240 1934.700 ;
        RECT 16.260 1881.150 18.240 1881.290 ;
        RECT 16.260 1878.570 16.400 1881.150 ;
        RECT 16.260 1878.430 16.860 1878.570 ;
        RECT 16.720 1827.570 16.860 1878.430 ;
        RECT 16.720 1827.430 17.780 1827.570 ;
        RECT 15.340 1824.710 17.320 1824.850 ;
        RECT 14.880 1817.230 15.480 1817.370 ;
        RECT 13.960 1816.550 14.560 1816.690 ;
        RECT 11.660 1815.190 12.260 1815.330 ;
        RECT 11.200 1734.950 11.800 1735.090 ;
        RECT 11.660 1703.130 11.800 1734.950 ;
        RECT 12.120 1730.330 12.260 1815.190 ;
        RECT 13.960 1733.050 14.100 1816.550 ;
        RECT 15.340 1761.610 15.480 1817.230 ;
        RECT 17.180 1816.690 17.320 1824.710 ;
        RECT 14.420 1761.470 15.480 1761.610 ;
        RECT 16.260 1816.550 17.320 1816.690 ;
        RECT 14.420 1750.050 14.560 1761.470 ;
        RECT 16.260 1760.930 16.400 1816.550 ;
        RECT 17.640 1806.490 17.780 1827.430 ;
        RECT 15.340 1760.790 16.400 1760.930 ;
        RECT 16.720 1806.350 17.780 1806.490 ;
        RECT 14.420 1749.910 15.020 1750.050 ;
        RECT 12.580 1732.910 14.100 1733.050 ;
        RECT 12.580 1730.330 12.720 1732.910 ;
        RECT 12.120 1730.190 13.640 1730.330 ;
        RECT 12.580 1724.890 12.720 1730.190 ;
        RECT 13.500 1727.610 13.640 1730.190 ;
        RECT 13.500 1727.470 14.560 1727.610 ;
        RECT 12.580 1724.750 13.640 1724.890 ;
        RECT 10.740 1702.990 11.800 1703.130 ;
        RECT 6.530 1687.235 6.810 1687.605 ;
        RECT 6.600 1668.710 6.740 1687.235 ;
        RECT 10.740 1682.730 10.880 1702.990 ;
        RECT 13.500 1698.370 13.640 1724.750 ;
        RECT 9.820 1682.590 10.880 1682.730 ;
        RECT 11.200 1698.230 13.640 1698.370 ;
        RECT 9.820 1671.090 9.960 1682.590 ;
        RECT 11.200 1682.050 11.340 1698.230 ;
        RECT 10.280 1681.910 11.340 1682.050 ;
        RECT 9.760 1670.770 10.020 1671.090 ;
        RECT 9.760 1670.320 10.020 1670.410 ;
        RECT 10.280 1670.320 10.420 1681.910 ;
        RECT 14.420 1670.320 14.560 1727.470 ;
        RECT 14.880 1724.890 15.020 1749.910 ;
        RECT 15.340 1726.930 15.480 1760.790 ;
        RECT 16.720 1731.010 16.860 1806.350 ;
        RECT 18.560 1772.490 18.700 2070.870 ;
        RECT 17.640 1772.350 18.700 1772.490 ;
        RECT 17.640 1737.130 17.780 1772.350 ;
        RECT 17.640 1736.990 18.700 1737.130 ;
        RECT 16.720 1730.870 18.240 1731.010 ;
        RECT 15.340 1726.790 17.320 1726.930 ;
        RECT 17.180 1726.250 17.320 1726.790 ;
        RECT 18.100 1726.250 18.240 1730.870 ;
        RECT 16.720 1726.110 18.240 1726.250 ;
        RECT 14.880 1724.750 15.480 1724.890 ;
        RECT 9.760 1670.180 10.420 1670.320 ;
        RECT 10.740 1670.180 14.560 1670.320 ;
        RECT 15.340 1670.320 15.480 1724.750 ;
        RECT 16.720 1722.850 16.860 1726.110 ;
        RECT 17.180 1725.570 17.320 1726.110 ;
        RECT 17.180 1725.430 18.240 1725.570 ;
        RECT 16.260 1722.710 16.860 1722.850 ;
        RECT 16.260 1721.490 16.400 1722.710 ;
        RECT 16.260 1721.350 16.860 1721.490 ;
        RECT 15.730 1698.370 16.010 1698.485 ;
        RECT 16.720 1698.370 16.860 1721.350 ;
        RECT 15.730 1698.230 16.860 1698.370 ;
        RECT 15.730 1698.115 16.010 1698.230 ;
        RECT 18.100 1670.320 18.240 1725.430 ;
        RECT 15.340 1670.180 15.940 1670.320 ;
        RECT 9.760 1670.090 10.020 1670.180 ;
        RECT 10.740 1669.130 10.880 1670.180 ;
        RECT 9.360 1668.990 10.880 1669.130 ;
        RECT 6.540 1668.390 6.800 1668.710 ;
        RECT 9.360 1667.770 9.500 1668.990 ;
        RECT 9.760 1668.450 10.020 1668.710 ;
        RECT 9.760 1668.390 14.560 1668.450 ;
        RECT 9.820 1668.310 14.560 1668.390 ;
        RECT 14.420 1668.280 14.560 1668.310 ;
        RECT 14.420 1668.140 15.020 1668.280 ;
        RECT 9.360 1667.630 14.560 1667.770 ;
        RECT 9.760 1667.030 10.020 1667.350 ;
        RECT 9.820 1660.290 9.960 1667.030 ;
        RECT 9.820 1660.150 14.100 1660.290 ;
        RECT 9.760 1658.930 10.020 1659.190 ;
        RECT 9.760 1658.870 13.180 1658.930 ;
        RECT 9.820 1658.790 13.180 1658.870 ;
        RECT 13.040 1624.930 13.180 1658.790 ;
        RECT 10.740 1624.790 13.180 1624.930 ;
        RECT 10.740 1594.330 10.880 1624.790 ;
        RECT 13.960 1624.250 14.100 1660.150 ;
        RECT 12.580 1624.110 14.100 1624.250 ;
        RECT 12.580 1605.210 12.720 1624.110 ;
        RECT 14.420 1623.570 14.560 1667.630 ;
        RECT 13.040 1623.430 14.560 1623.570 ;
        RECT 13.040 1605.890 13.180 1623.430 ;
        RECT 13.040 1605.750 14.100 1605.890 ;
        RECT 12.580 1605.070 13.180 1605.210 ;
        RECT 9.820 1594.190 10.880 1594.330 ;
        RECT 9.820 1575.890 9.960 1594.190 ;
        RECT 13.040 1589.570 13.180 1605.070 ;
        RECT 13.960 1590.250 14.100 1605.750 ;
        RECT 14.880 1592.290 15.020 1668.140 ;
        RECT 15.800 1637.170 15.940 1670.180 ;
        RECT 17.640 1670.180 18.240 1670.320 ;
        RECT 15.800 1637.030 16.400 1637.170 ;
        RECT 16.260 1635.810 16.400 1637.030 ;
        RECT 15.340 1635.670 16.400 1635.810 ;
        RECT 15.340 1605.890 15.480 1635.670 ;
        RECT 17.640 1610.650 17.780 1670.180 ;
        RECT 17.180 1610.510 17.780 1610.650 ;
        RECT 15.340 1605.750 16.400 1605.890 ;
        RECT 15.730 1604.955 16.010 1605.325 ;
        RECT 14.880 1592.150 15.480 1592.290 ;
        RECT 15.340 1590.250 15.480 1592.150 ;
        RECT 13.960 1590.110 14.560 1590.250 ;
        RECT 10.280 1589.430 13.180 1589.570 ;
        RECT 9.760 1575.570 10.020 1575.890 ;
        RECT 9.760 1562.200 10.020 1562.290 ;
        RECT 10.280 1562.200 10.420 1589.430 ;
        RECT 14.420 1588.890 14.560 1590.110 ;
        RECT 13.040 1588.750 14.560 1588.890 ;
        RECT 14.880 1590.110 15.480 1590.250 ;
        RECT 13.040 1588.210 13.180 1588.750 ;
        RECT 9.760 1562.060 10.420 1562.200 ;
        RECT 12.120 1588.070 13.180 1588.210 ;
        RECT 9.760 1561.970 10.020 1562.060 ;
        RECT 12.120 1561.690 12.260 1588.070 ;
        RECT 14.880 1586.170 15.020 1590.110 ;
        RECT 13.960 1586.030 15.020 1586.170 ;
        RECT 13.960 1570.530 14.100 1586.030 ;
        RECT 9.820 1561.610 12.260 1561.690 ;
        RECT 9.760 1561.550 12.260 1561.610 ;
        RECT 13.040 1570.390 14.100 1570.530 ;
        RECT 9.760 1561.290 10.020 1561.550 ;
        RECT 13.040 1561.010 13.180 1570.390 ;
        RECT 15.800 1569.170 15.940 1604.955 ;
        RECT 9.820 1560.930 13.180 1561.010 ;
        RECT 9.760 1560.870 13.180 1560.930 ;
        RECT 14.880 1569.030 15.940 1569.170 ;
        RECT 9.760 1560.610 10.020 1560.870 ;
        RECT 14.880 1560.330 15.020 1569.030 ;
        RECT 13.040 1560.190 15.020 1560.330 ;
        RECT 9.760 1558.970 10.020 1559.230 ;
        RECT 9.760 1558.910 11.800 1558.970 ;
        RECT 9.820 1558.830 11.800 1558.910 ;
        RECT 11.660 1522.930 11.800 1558.830 ;
        RECT 13.040 1552.170 13.180 1560.190 ;
        RECT 16.260 1552.850 16.400 1605.750 ;
        RECT 17.180 1602.490 17.320 1610.510 ;
        RECT 16.720 1602.350 17.320 1602.490 ;
        RECT 16.720 1573.930 16.860 1602.350 ;
        RECT 18.560 1601.810 18.700 1736.990 ;
        RECT 17.180 1601.670 18.700 1601.810 ;
        RECT 17.180 1600.450 17.320 1601.670 ;
        RECT 17.180 1600.310 18.700 1600.450 ;
        RECT 18.560 1575.290 18.700 1600.310 ;
        RECT 17.180 1575.150 18.700 1575.290 ;
        RECT 17.180 1573.930 17.320 1575.150 ;
        RECT 16.720 1573.790 17.780 1573.930 ;
        RECT 16.260 1552.710 16.860 1552.850 ;
        RECT 16.720 1552.170 16.860 1552.710 ;
        RECT 13.040 1552.030 14.100 1552.170 ;
        RECT 9.820 1522.850 11.800 1522.930 ;
        RECT 9.760 1522.790 11.800 1522.850 ;
        RECT 9.760 1522.530 10.020 1522.790 ;
        RECT 9.820 1521.430 11.800 1521.570 ;
        RECT 9.820 1520.810 9.960 1521.430 ;
        RECT 9.760 1520.490 10.020 1520.810 ;
        RECT 9.760 1519.810 10.020 1520.130 ;
        RECT 9.820 1519.530 9.960 1519.810 ;
        RECT 9.820 1519.390 11.340 1519.530 ;
        RECT 9.760 1516.810 10.020 1517.070 ;
        RECT 11.200 1516.810 11.340 1519.390 ;
        RECT 9.760 1516.750 11.340 1516.810 ;
        RECT 9.820 1516.670 11.340 1516.750 ;
        RECT 11.660 1478.730 11.800 1521.430 ;
        RECT 9.820 1478.590 11.800 1478.730 ;
        RECT 6.990 1471.675 7.270 1472.045 ;
        RECT 7.060 1419.830 7.200 1471.675 ;
        RECT 9.820 1467.090 9.960 1478.590 ;
        RECT 13.960 1477.370 14.100 1552.030 ;
        RECT 14.880 1552.030 16.860 1552.170 ;
        RECT 14.880 1525.650 15.020 1552.030 ;
        RECT 17.180 1529.050 17.320 1573.790 ;
        RECT 16.260 1528.910 17.320 1529.050 ;
        RECT 14.880 1525.510 15.940 1525.650 ;
        RECT 15.800 1493.690 15.940 1525.510 ;
        RECT 16.260 1509.160 16.400 1528.910 ;
        RECT 16.660 1509.160 16.920 1509.250 ;
        RECT 16.260 1509.020 16.920 1509.160 ;
        RECT 16.660 1508.930 16.920 1509.020 ;
        RECT 17.640 1508.650 17.780 1573.790 ;
        RECT 19.020 1513.410 19.160 2249.030 ;
        RECT 11.200 1477.230 14.100 1477.370 ;
        RECT 14.880 1493.550 15.940 1493.690 ;
        RECT 16.720 1508.510 17.780 1508.650 ;
        RECT 18.100 1513.270 19.160 1513.410 ;
        RECT 9.760 1466.770 10.020 1467.090 ;
        RECT 9.760 1465.410 10.020 1465.730 ;
        RECT 9.820 1424.330 9.960 1465.410 ;
        RECT 11.200 1440.650 11.340 1477.230 ;
        RECT 14.880 1441.330 15.020 1493.550 ;
        RECT 16.720 1490.290 16.860 1508.510 ;
        RECT 16.720 1490.150 17.320 1490.290 ;
        RECT 17.180 1483.490 17.320 1490.150 ;
        RECT 15.800 1483.350 17.320 1483.490 ;
        RECT 15.800 1480.600 15.940 1483.350 ;
        RECT 18.100 1482.810 18.240 1513.270 ;
        RECT 18.500 1509.160 18.760 1509.250 ;
        RECT 18.500 1509.020 19.160 1509.160 ;
        RECT 18.500 1508.930 18.760 1509.020 ;
        RECT 16.720 1482.670 18.240 1482.810 ;
        RECT 16.720 1480.600 16.860 1482.670 ;
        RECT 15.340 1480.460 16.860 1480.600 ;
        RECT 15.340 1476.010 15.480 1480.460 ;
        RECT 15.800 1480.090 15.940 1480.460 ;
        RECT 15.800 1479.950 17.320 1480.090 ;
        RECT 17.180 1479.920 17.320 1479.950 ;
        RECT 17.180 1479.780 18.240 1479.920 ;
        RECT 15.340 1475.870 15.940 1476.010 ;
        RECT 14.880 1441.190 15.480 1441.330 ;
        RECT 11.200 1440.510 15.020 1440.650 ;
        RECT 9.820 1424.190 14.560 1424.330 ;
        RECT 9.760 1423.820 10.020 1423.910 ;
        RECT 9.760 1423.680 14.100 1423.820 ;
        RECT 9.760 1423.590 10.020 1423.680 ;
        RECT 9.760 1423.140 10.020 1423.230 ;
        RECT 9.760 1423.000 12.720 1423.140 ;
        RECT 9.760 1422.910 10.020 1423.000 ;
        RECT 9.760 1421.610 10.020 1421.870 ;
        RECT 9.760 1421.550 12.260 1421.610 ;
        RECT 9.820 1421.470 12.260 1421.550 ;
        RECT 7.000 1419.510 7.260 1419.830 ;
        RECT 12.120 1383.530 12.260 1421.470 ;
        RECT 12.580 1384.210 12.720 1423.000 ;
        RECT 12.580 1384.070 13.640 1384.210 ;
        RECT 11.200 1383.390 12.260 1383.530 ;
        RECT 11.200 1374.690 11.340 1383.390 ;
        RECT 13.500 1382.850 13.640 1384.070 ;
        RECT 13.040 1382.710 13.640 1382.850 ;
        RECT 13.040 1382.170 13.180 1382.710 ;
        RECT 12.580 1382.030 13.180 1382.170 ;
        RECT 12.580 1378.770 12.720 1382.030 ;
        RECT 13.960 1380.810 14.100 1423.680 ;
        RECT 14.420 1408.010 14.560 1424.190 ;
        RECT 14.880 1408.690 15.020 1440.510 ;
        RECT 15.340 1412.770 15.480 1441.190 ;
        RECT 15.800 1417.020 15.940 1475.870 ;
        RECT 18.100 1417.020 18.240 1479.780 ;
        RECT 19.020 1417.020 19.160 1509.020 ;
        RECT 15.800 1416.880 17.320 1417.020 ;
        RECT 17.180 1414.810 17.320 1416.880 ;
        RECT 17.640 1416.880 19.160 1417.020 ;
        RECT 17.640 1414.810 17.780 1416.880 ;
        RECT 18.100 1415.490 18.240 1416.880 ;
        RECT 18.100 1415.350 18.700 1415.490 ;
        RECT 18.560 1414.810 18.700 1415.350 ;
        RECT 17.180 1414.670 19.160 1414.810 ;
        RECT 15.340 1412.630 17.320 1412.770 ;
        RECT 17.180 1410.730 17.320 1412.630 ;
        RECT 17.640 1411.410 17.780 1414.670 ;
        RECT 17.640 1411.270 18.240 1411.410 ;
        RECT 16.720 1410.590 17.320 1410.730 ;
        RECT 16.720 1410.050 16.860 1410.590 ;
        RECT 16.260 1409.910 16.860 1410.050 ;
        RECT 14.880 1408.550 15.940 1408.690 ;
        RECT 14.420 1407.870 15.480 1408.010 ;
        RECT 15.340 1407.330 15.480 1407.870 ;
        RECT 14.420 1407.190 15.480 1407.330 ;
        RECT 14.420 1381.490 14.560 1407.190 ;
        RECT 15.800 1389.650 15.940 1408.550 ;
        RECT 16.260 1389.650 16.400 1409.910 ;
        RECT 14.880 1389.510 16.400 1389.650 ;
        RECT 14.880 1383.530 15.020 1389.510 ;
        RECT 15.800 1387.610 15.940 1389.510 ;
        RECT 15.800 1387.470 17.320 1387.610 ;
        RECT 14.880 1383.390 16.400 1383.530 ;
        RECT 14.420 1381.350 15.020 1381.490 ;
        RECT 13.040 1380.670 14.100 1380.810 ;
        RECT 13.040 1378.770 13.180 1380.670 ;
        RECT 12.580 1378.630 14.560 1378.770 ;
        RECT 13.040 1376.730 13.180 1378.630 ;
        RECT 13.040 1376.590 14.100 1376.730 ;
        RECT 11.200 1374.550 13.640 1374.690 ;
        RECT 9.820 1320.890 10.880 1320.970 ;
        RECT 9.760 1320.830 10.880 1320.890 ;
        RECT 9.760 1320.570 10.020 1320.830 ;
        RECT 10.740 1307.370 10.880 1320.830 ;
        RECT 13.500 1319.610 13.640 1374.550 ;
        RECT 12.120 1319.470 13.640 1319.610 ;
        RECT 12.120 1310.770 12.260 1319.470 ;
        RECT 13.960 1318.250 14.100 1376.590 ;
        RECT 14.420 1335.930 14.560 1378.630 ;
        RECT 14.880 1345.450 15.020 1381.350 ;
        RECT 16.260 1346.130 16.400 1383.390 ;
        RECT 17.180 1382.170 17.320 1387.470 ;
        RECT 15.800 1345.990 16.400 1346.130 ;
        RECT 16.720 1382.030 17.320 1382.170 ;
        RECT 15.800 1345.450 15.940 1345.990 ;
        RECT 14.880 1345.310 16.400 1345.450 ;
        RECT 15.800 1343.410 15.940 1345.310 ;
        RECT 15.340 1343.270 15.940 1343.410 ;
        RECT 15.340 1341.370 15.480 1343.270 ;
        RECT 14.880 1341.230 15.480 1341.370 ;
        RECT 14.880 1340.010 15.020 1341.230 ;
        RECT 14.880 1339.870 15.480 1340.010 ;
        RECT 15.340 1335.930 15.480 1339.870 ;
        RECT 14.420 1335.790 15.940 1335.930 ;
        RECT 13.040 1318.110 14.100 1318.250 ;
        RECT 13.040 1310.770 13.180 1318.110 ;
        RECT 15.340 1316.890 15.480 1335.790 ;
        RECT 13.960 1316.750 15.480 1316.890 ;
        RECT 13.960 1311.450 14.100 1316.750 ;
        RECT 15.800 1312.810 15.940 1335.790 ;
        RECT 15.340 1312.670 15.940 1312.810 ;
        RECT 13.960 1311.310 15.020 1311.450 ;
        RECT 14.880 1310.770 15.020 1311.310 ;
        RECT 15.340 1310.770 15.480 1312.670 ;
        RECT 12.120 1310.630 12.720 1310.770 ;
        RECT 13.040 1310.630 14.100 1310.770 ;
        RECT 14.880 1310.630 15.940 1310.770 ;
        RECT 12.580 1310.090 12.720 1310.630 ;
        RECT 12.580 1309.950 13.180 1310.090 ;
        RECT 10.280 1307.230 10.880 1307.370 ;
        RECT 10.280 1291.050 10.420 1307.230 ;
        RECT 13.040 1291.050 13.180 1309.950 ;
        RECT 10.280 1290.910 13.640 1291.050 ;
        RECT 13.040 1214.890 13.180 1290.910 ;
        RECT 11.660 1214.750 13.180 1214.890 ;
        RECT 9.760 1099.800 10.020 1099.890 ;
        RECT 11.660 1099.800 11.800 1214.750 ;
        RECT 13.500 1171.370 13.640 1290.910 ;
        RECT 12.120 1171.230 13.640 1171.370 ;
        RECT 12.120 1168.650 12.260 1171.230 ;
        RECT 13.960 1170.010 14.100 1310.630 ;
        RECT 15.340 1284.930 15.480 1310.630 ;
        RECT 14.420 1284.790 15.480 1284.930 ;
        RECT 14.420 1170.010 14.560 1284.790 ;
        RECT 15.800 1284.250 15.940 1310.630 ;
        RECT 13.500 1169.870 14.560 1170.010 ;
        RECT 14.880 1284.110 15.940 1284.250 ;
        RECT 13.500 1169.330 13.640 1169.870 ;
        RECT 13.040 1169.190 13.640 1169.330 ;
        RECT 13.960 1169.330 14.100 1169.870 ;
        RECT 13.960 1169.190 14.560 1169.330 ;
        RECT 13.040 1168.650 13.180 1169.190 ;
        RECT 12.120 1168.510 14.100 1168.650 ;
        RECT 13.040 1161.170 13.180 1168.510 ;
        RECT 9.760 1099.660 11.800 1099.800 ;
        RECT 12.580 1161.030 13.180 1161.170 ;
        RECT 9.760 1099.570 10.020 1099.660 ;
        RECT 12.580 1091.810 12.720 1161.030 ;
        RECT 9.820 1091.730 12.720 1091.810 ;
        RECT 9.760 1091.670 12.720 1091.730 ;
        RECT 9.760 1091.410 10.020 1091.670 ;
        RECT 9.760 1088.410 10.020 1088.670 ;
        RECT 9.760 1088.350 11.800 1088.410 ;
        RECT 9.820 1088.270 11.800 1088.350 ;
        RECT 11.660 1087.220 11.800 1088.270 ;
        RECT 11.660 1087.080 12.260 1087.220 ;
        RECT 12.120 1082.970 12.260 1087.080 ;
        RECT 13.960 1087.050 14.100 1168.510 ;
        RECT 9.820 1082.830 12.260 1082.970 ;
        RECT 13.040 1086.910 14.100 1087.050 ;
        RECT 9.820 1071.670 9.960 1082.830 ;
        RECT 7.000 1071.350 7.260 1071.670 ;
        RECT 9.760 1071.350 10.020 1071.670 ;
        RECT 7.060 1024.750 7.200 1071.350 ;
        RECT 13.040 1039.450 13.180 1086.910 ;
        RECT 10.740 1039.310 13.180 1039.450 ;
        RECT 7.000 1024.430 7.260 1024.750 ;
        RECT 10.740 1018.370 10.880 1039.310 ;
        RECT 14.420 1019.730 14.560 1169.190 ;
        RECT 14.880 1163.210 15.020 1284.110 ;
        RECT 16.260 1283.570 16.400 1345.310 ;
        RECT 15.340 1283.430 16.400 1283.570 ;
        RECT 15.340 1276.090 15.480 1283.430 ;
        RECT 16.720 1280.000 16.860 1382.030 ;
        RECT 18.100 1371.970 18.240 1411.270 ;
        RECT 15.800 1279.860 16.860 1280.000 ;
        RECT 17.180 1371.830 18.240 1371.970 ;
        RECT 15.800 1276.770 15.940 1279.860 ;
        RECT 15.800 1276.630 16.860 1276.770 ;
        RECT 16.720 1276.090 16.860 1276.630 ;
        RECT 17.180 1276.090 17.320 1371.830 ;
        RECT 18.560 1371.290 18.700 1414.670 ;
        RECT 17.640 1371.150 18.700 1371.290 ;
        RECT 17.640 1316.890 17.780 1371.150 ;
        RECT 17.640 1316.750 18.240 1316.890 ;
        RECT 18.100 1314.850 18.240 1316.750 ;
        RECT 18.100 1314.710 18.700 1314.850 ;
        RECT 18.560 1313.490 18.700 1314.710 ;
        RECT 19.020 1313.490 19.160 1414.670 ;
        RECT 17.640 1313.350 19.160 1313.490 ;
        RECT 17.640 1286.290 17.780 1313.350 ;
        RECT 18.560 1286.970 18.700 1313.350 ;
        RECT 18.560 1286.830 19.160 1286.970 ;
        RECT 17.640 1286.150 18.700 1286.290 ;
        RECT 15.340 1275.950 18.240 1276.090 ;
        RECT 16.720 1257.050 16.860 1275.950 ;
        RECT 15.340 1256.910 16.860 1257.050 ;
        RECT 15.340 1163.890 15.480 1256.910 ;
        RECT 17.180 1229.170 17.320 1275.950 ;
        RECT 15.800 1229.030 17.320 1229.170 ;
        RECT 15.800 1199.250 15.940 1229.030 ;
        RECT 18.100 1206.730 18.240 1275.950 ;
        RECT 16.720 1206.590 18.240 1206.730 ;
        RECT 16.720 1200.610 16.860 1206.590 ;
        RECT 18.560 1204.690 18.700 1286.150 ;
        RECT 18.100 1204.550 18.700 1204.690 ;
        RECT 18.100 1203.330 18.240 1204.550 ;
        RECT 19.020 1204.010 19.160 1286.830 ;
        RECT 18.560 1203.870 19.160 1204.010 ;
        RECT 18.560 1203.330 18.700 1203.870 ;
        RECT 18.100 1203.190 19.160 1203.330 ;
        RECT 16.720 1200.470 18.240 1200.610 ;
        RECT 15.800 1199.110 17.780 1199.250 ;
        RECT 17.640 1198.570 17.780 1199.110 ;
        RECT 18.100 1198.570 18.240 1200.470 ;
        RECT 16.260 1198.430 18.240 1198.570 ;
        RECT 16.260 1170.690 16.400 1198.430 ;
        RECT 17.640 1197.210 17.780 1198.430 ;
        RECT 18.560 1197.210 18.700 1203.190 ;
        RECT 17.180 1197.070 18.700 1197.210 ;
        RECT 17.180 1172.050 17.320 1197.070 ;
        RECT 15.800 1170.550 16.400 1170.690 ;
        RECT 16.720 1171.910 17.320 1172.050 ;
        RECT 15.800 1168.650 15.940 1170.550 ;
        RECT 16.720 1170.010 16.860 1171.910 ;
        RECT 17.640 1170.010 17.780 1197.070 ;
        RECT 16.260 1169.870 17.780 1170.010 ;
        RECT 16.260 1168.650 16.400 1169.870 ;
        RECT 16.720 1169.330 16.860 1169.870 ;
        RECT 16.720 1169.190 17.780 1169.330 ;
        RECT 15.800 1168.510 17.320 1168.650 ;
        RECT 16.260 1163.890 16.400 1168.510 ;
        RECT 15.340 1163.750 16.860 1163.890 ;
        RECT 14.880 1163.070 15.940 1163.210 ;
        RECT 15.800 1129.890 15.940 1163.070 ;
        RECT 9.820 1018.230 10.880 1018.370 ;
        RECT 11.200 1019.590 14.560 1019.730 ;
        RECT 14.880 1129.750 15.940 1129.890 ;
        RECT 9.820 1009.450 9.960 1018.230 ;
        RECT 9.760 1009.130 10.020 1009.450 ;
        RECT 7.000 991.285 7.260 991.430 ;
        RECT 6.990 990.915 7.270 991.285 ;
        RECT 11.200 991.170 11.340 1019.590 ;
        RECT 14.880 1017.690 15.020 1129.750 ;
        RECT 16.260 1128.530 16.400 1163.750 ;
        RECT 15.800 1128.390 16.400 1128.530 ;
        RECT 15.800 1127.170 15.940 1128.390 ;
        RECT 16.720 1127.850 16.860 1163.750 ;
        RECT 17.180 1131.930 17.320 1168.510 ;
        RECT 17.640 1131.930 17.780 1169.190 ;
        RECT 19.020 1158.450 19.160 1203.190 ;
        RECT 18.100 1158.310 19.160 1158.450 ;
        RECT 18.100 1132.610 18.240 1158.310 ;
        RECT 18.100 1132.470 19.160 1132.610 ;
        RECT 17.180 1131.790 18.700 1131.930 ;
        RECT 17.640 1131.250 17.780 1131.790 ;
        RECT 17.640 1131.110 18.240 1131.250 ;
        RECT 9.820 991.090 11.340 991.170 ;
        RECT 9.760 991.030 11.340 991.090 ;
        RECT 11.660 1017.550 15.020 1017.690 ;
        RECT 15.340 1127.030 15.940 1127.170 ;
        RECT 16.260 1127.710 16.860 1127.850 ;
        RECT 9.760 990.770 10.020 991.030 ;
        RECT 11.660 989.130 11.800 1017.550 ;
        RECT 15.340 1015.650 15.480 1127.030 ;
        RECT 16.260 1126.490 16.400 1127.710 ;
        RECT 15.800 1126.350 16.400 1126.490 ;
        RECT 15.800 1093.850 15.940 1126.350 ;
        RECT 18.100 1099.290 18.240 1131.110 ;
        RECT 17.180 1099.150 18.240 1099.290 ;
        RECT 17.180 1097.930 17.320 1099.150 ;
        RECT 16.260 1097.790 17.320 1097.930 ;
        RECT 16.260 1095.210 16.400 1097.790 ;
        RECT 16.260 1095.070 16.860 1095.210 ;
        RECT 16.720 1093.850 16.860 1095.070 ;
        RECT 17.180 1095.070 18.240 1095.210 ;
        RECT 17.180 1093.850 17.320 1095.070 ;
        RECT 15.800 1093.710 17.320 1093.850 ;
        RECT 16.720 1091.130 16.860 1093.710 ;
        RECT 16.260 1090.990 16.860 1091.130 ;
        RECT 16.260 1054.410 16.400 1090.990 ;
        RECT 16.260 1054.270 17.320 1054.410 ;
        RECT 17.180 1015.650 17.320 1054.270 ;
        RECT 9.820 989.050 11.800 989.130 ;
        RECT 9.760 988.990 11.800 989.050 ;
        RECT 14.880 1015.510 15.480 1015.650 ;
        RECT 16.260 1015.510 17.320 1015.650 ;
        RECT 9.760 988.730 10.020 988.990 ;
        RECT 14.880 988.450 15.020 1015.510 ;
        RECT 16.260 1014.970 16.400 1015.510 ;
        RECT 18.100 1014.970 18.240 1095.070 ;
        RECT 9.820 988.370 15.020 988.450 ;
        RECT 9.760 988.310 15.020 988.370 ;
        RECT 15.340 1014.830 16.400 1014.970 ;
        RECT 17.180 1014.830 18.240 1014.970 ;
        RECT 9.760 988.050 10.020 988.310 ;
        RECT 9.760 981.650 10.020 981.910 ;
        RECT 9.760 981.590 14.560 981.650 ;
        RECT 9.820 981.510 14.560 981.590 ;
        RECT 9.760 981.140 10.020 981.230 ;
        RECT 9.760 981.000 14.100 981.140 ;
        RECT 9.760 980.910 10.020 981.000 ;
        RECT 9.760 978.930 10.020 979.190 ;
        RECT 9.760 978.870 10.880 978.930 ;
        RECT 9.820 978.790 10.880 978.870 ;
        RECT 10.740 976.210 10.880 978.790 ;
        RECT 10.740 976.070 12.720 976.210 ;
        RECT 9.760 973.660 10.020 973.750 ;
        RECT 9.760 973.520 10.880 973.660 ;
        RECT 9.760 973.430 10.020 973.520 ;
        RECT 9.760 948.160 10.020 948.250 ;
        RECT 10.740 948.160 10.880 973.520 ;
        RECT 9.760 948.020 10.880 948.160 ;
        RECT 9.760 947.930 10.020 948.020 ;
        RECT 12.580 946.120 12.720 976.070 ;
        RECT 12.120 945.980 12.720 946.120 ;
        RECT 9.760 943.400 10.020 943.490 ;
        RECT 12.120 943.400 12.260 945.980 ;
        RECT 9.760 943.260 12.260 943.400 ;
        RECT 9.760 943.170 10.020 943.260 ;
        RECT 9.760 942.720 10.020 942.810 ;
        RECT 9.760 942.580 10.420 942.720 ;
        RECT 9.760 942.490 10.020 942.580 ;
        RECT 10.280 884.410 10.420 942.580 ;
        RECT 13.960 929.970 14.100 981.000 ;
        RECT 13.500 929.830 14.100 929.970 ;
        RECT 13.500 889.850 13.640 929.830 ;
        RECT 14.420 927.930 14.560 981.510 ;
        RECT 15.340 966.690 15.480 1014.830 ;
        RECT 17.180 966.690 17.320 1014.830 ;
        RECT 18.560 978.250 18.700 1131.790 ;
        RECT 14.880 966.550 17.320 966.690 ;
        RECT 18.100 978.110 18.700 978.250 ;
        RECT 14.880 960.570 15.020 966.550 ;
        RECT 15.340 961.250 15.480 966.550 ;
        RECT 15.340 961.110 17.780 961.250 ;
        RECT 14.880 960.430 15.940 960.570 ;
        RECT 14.420 927.790 15.480 927.930 ;
        RECT 14.350 926.315 14.630 926.685 ;
        RECT 13.500 889.710 14.100 889.850 ;
        RECT 9.360 884.270 10.420 884.410 ;
        RECT 9.360 865.970 9.500 884.270 ;
        RECT 9.760 883.730 10.020 883.990 ;
        RECT 9.760 883.670 12.260 883.730 ;
        RECT 9.820 883.590 12.260 883.670 ;
        RECT 12.120 883.050 12.260 883.590 ;
        RECT 12.120 882.910 12.720 883.050 ;
        RECT 7.460 865.650 7.720 865.970 ;
        RECT 9.300 865.650 9.560 865.970 ;
        RECT 7.520 865.485 7.660 865.650 ;
        RECT 7.450 865.115 7.730 865.485 ;
        RECT 6.990 837.915 7.270 838.285 ;
        RECT 5.160 836.070 5.420 836.390 ;
        RECT 7.060 830.270 7.200 837.915 ;
        RECT 12.580 835.450 12.720 882.910 ;
        RECT 9.360 835.310 12.720 835.450 ;
        RECT 7.000 829.950 7.260 830.270 ;
        RECT 7.460 799.690 7.720 800.010 ;
        RECT 7.520 798.650 7.660 799.690 ;
        RECT 7.460 798.330 7.720 798.650 ;
        RECT 9.360 769.070 9.500 835.310 ;
        RECT 13.960 833.410 14.100 889.710 ;
        RECT 9.820 833.270 14.100 833.410 ;
        RECT 9.820 832.310 9.960 833.270 ;
        RECT 9.760 831.990 10.020 832.310 ;
        RECT 9.760 831.370 10.020 831.630 ;
        RECT 9.760 831.310 11.800 831.370 ;
        RECT 9.820 831.230 11.800 831.310 ;
        RECT 9.760 830.010 10.020 830.270 ;
        RECT 11.660 830.010 11.800 831.230 ;
        RECT 14.420 830.010 14.560 926.315 ;
        RECT 15.340 925.890 15.480 927.790 ;
        RECT 14.880 925.750 15.480 925.890 ;
        RECT 14.880 863.330 15.020 925.750 ;
        RECT 15.800 921.130 15.940 960.430 ;
        RECT 17.640 956.490 17.780 961.110 ;
        RECT 16.720 956.350 17.780 956.490 ;
        RECT 16.720 955.810 16.860 956.350 ;
        RECT 15.340 920.990 15.940 921.130 ;
        RECT 16.260 955.670 16.860 955.810 ;
        RECT 15.340 864.010 15.480 920.990 ;
        RECT 16.260 915.010 16.400 955.670 ;
        RECT 18.100 945.610 18.240 978.110 ;
        RECT 19.020 976.890 19.160 1132.470 ;
        RECT 15.800 914.870 16.400 915.010 ;
        RECT 17.640 945.470 18.240 945.610 ;
        RECT 18.560 976.750 19.160 976.890 ;
        RECT 15.800 900.730 15.940 914.870 ;
        RECT 17.640 901.410 17.780 945.470 ;
        RECT 18.560 924.530 18.700 976.750 ;
        RECT 18.560 924.390 19.160 924.530 ;
        RECT 17.640 901.270 18.700 901.410 ;
        RECT 15.800 900.590 16.400 900.730 ;
        RECT 16.260 900.050 16.400 900.590 ;
        RECT 16.260 899.910 17.320 900.050 ;
        RECT 17.180 898.010 17.320 899.910 ;
        RECT 17.180 897.870 17.780 898.010 ;
        RECT 15.800 896.510 17.320 896.650 ;
        RECT 15.800 865.370 15.940 896.510 ;
        RECT 17.180 894.610 17.320 896.510 ;
        RECT 17.640 895.290 17.780 897.870 ;
        RECT 17.640 895.150 18.240 895.290 ;
        RECT 18.100 894.610 18.240 895.150 ;
        RECT 18.560 894.610 18.700 901.270 ;
        RECT 17.180 894.470 18.700 894.610 ;
        RECT 18.100 893.930 18.240 894.470 ;
        RECT 16.260 893.790 18.240 893.930 ;
        RECT 16.260 871.490 16.400 893.790 ;
        RECT 19.020 885.090 19.160 924.390 ;
        RECT 18.100 884.950 19.160 885.090 ;
        RECT 18.100 871.490 18.240 884.950 ;
        RECT 16.260 871.350 19.160 871.490 ;
        RECT 18.100 865.370 18.240 871.350 ;
        RECT 15.800 865.230 18.700 865.370 ;
        RECT 15.340 863.870 16.860 864.010 ;
        RECT 16.720 863.330 16.860 863.870 ;
        RECT 14.880 863.190 17.780 863.330 ;
        RECT 16.720 861.970 16.860 863.190 ;
        RECT 9.760 829.950 10.880 830.010 ;
        RECT 9.820 829.870 10.880 829.950 ;
        RECT 11.660 829.870 14.560 830.010 ;
        RECT 14.880 861.830 16.860 861.970 ;
        RECT 9.760 829.270 10.020 829.590 ;
        RECT 9.820 827.970 9.960 829.270 ;
        RECT 10.740 828.650 10.880 829.870 ;
        RECT 10.740 828.510 14.100 828.650 ;
        RECT 9.820 827.830 13.640 827.970 ;
        RECT 9.760 827.230 10.020 827.550 ;
        RECT 9.820 800.010 9.960 827.230 ;
        RECT 13.500 801.450 13.640 827.830 ;
        RECT 12.120 801.310 13.640 801.450 ;
        RECT 9.760 799.690 10.020 800.010 ;
        RECT 9.760 798.330 10.020 798.650 ;
        RECT 9.820 797.370 9.960 798.330 ;
        RECT 9.820 797.230 10.880 797.370 ;
        RECT 9.300 768.750 9.560 769.070 ;
        RECT 10.740 755.210 10.880 797.230 ;
        RECT 12.120 766.090 12.260 801.310 ;
        RECT 13.960 800.600 14.100 828.510 ;
        RECT 9.820 755.070 10.880 755.210 ;
        RECT 11.660 765.950 12.260 766.090 ;
        RECT 13.040 800.460 14.100 800.600 ;
        RECT 9.820 735.750 9.960 755.070 ;
        RECT 11.660 741.610 11.800 765.950 ;
        RECT 11.200 741.470 11.800 741.610 ;
        RECT 7.920 735.430 8.180 735.750 ;
        RECT 9.760 735.430 10.020 735.750 ;
        RECT 7.980 734.925 8.120 735.430 ;
        RECT 7.910 734.555 8.190 734.925 ;
        RECT 7.920 731.690 8.180 732.010 ;
        RECT 2.920 730.590 3.520 730.730 ;
        RECT 2.920 708.890 3.060 730.590 ;
        RECT 7.980 715.010 8.120 731.690 ;
        RECT 7.920 714.690 8.180 715.010 ;
        RECT 5.160 714.010 5.420 714.330 ;
        RECT 2.860 708.570 3.120 708.890 ;
        RECT 4.240 708.570 4.500 708.890 ;
        RECT 4.300 644.630 4.440 708.570 ;
        RECT 5.220 672.850 5.360 714.010 ;
        RECT 11.200 706.250 11.340 741.470 ;
        RECT 13.040 733.450 13.180 800.460 ;
        RECT 14.880 800.090 15.020 861.830 ;
        RECT 13.500 799.950 15.020 800.090 ;
        RECT 15.340 861.150 16.860 861.290 ;
        RECT 13.500 740.250 13.640 799.950 ;
        RECT 15.340 793.970 15.480 861.150 ;
        RECT 16.720 859.250 16.860 861.150 ;
        RECT 17.640 859.250 17.780 863.190 ;
        RECT 18.100 859.250 18.240 865.230 ;
        RECT 16.720 859.110 18.240 859.250 ;
        RECT 17.640 858.570 17.780 859.110 ;
        RECT 17.640 858.430 18.240 858.570 ;
        RECT 15.340 793.830 16.400 793.970 ;
        RECT 16.260 755.890 16.400 793.830 ;
        RECT 15.340 755.750 16.400 755.890 ;
        RECT 13.500 740.110 14.560 740.250 ;
        RECT 13.040 733.310 13.640 733.450 ;
        RECT 9.820 706.170 11.340 706.250 ;
        RECT 9.760 706.110 11.340 706.170 ;
        RECT 9.760 705.850 10.020 706.110 ;
        RECT 9.760 699.960 10.020 700.050 ;
        RECT 13.500 699.960 13.640 733.310 ;
        RECT 13.900 718.090 14.160 718.410 ;
        RECT 9.760 699.820 13.640 699.960 ;
        RECT 9.760 699.730 10.020 699.820 ;
        RECT 13.960 699.280 14.100 718.090 ;
        RECT 12.580 699.140 14.100 699.280 ;
        RECT 7.450 693.075 7.730 693.445 ;
        RECT 9.760 693.160 10.020 693.250 ;
        RECT 7.460 692.930 7.720 693.075 ;
        RECT 9.760 693.020 11.340 693.160 ;
        RECT 9.760 692.930 10.020 693.020 ;
        RECT 5.160 672.530 5.420 672.850 ;
        RECT 5.160 666.410 5.420 666.730 ;
        RECT 4.240 644.310 4.500 644.630 ;
        RECT 5.220 251.930 5.360 666.410 ;
        RECT 11.200 660.690 11.340 693.020 ;
        RECT 9.820 660.610 11.340 660.690 ;
        RECT 9.760 660.550 11.340 660.610 ;
        RECT 9.760 660.290 10.020 660.550 ;
        RECT 12.580 657.970 12.720 699.140 ;
        RECT 9.360 657.830 12.720 657.970 ;
        RECT 9.360 646.410 9.500 657.830 ;
        RECT 9.760 654.400 10.020 654.490 ;
        RECT 14.420 654.400 14.560 740.110 ;
        RECT 15.340 711.010 15.480 755.750 ;
        RECT 18.100 753.850 18.240 858.430 ;
        RECT 17.180 753.710 18.240 753.850 ;
        RECT 17.180 753.170 17.320 753.710 ;
        RECT 18.560 753.170 18.700 865.230 ;
        RECT 15.800 753.030 17.320 753.170 ;
        RECT 17.640 753.030 18.700 753.170 ;
        RECT 15.800 718.410 15.940 753.030 ;
        RECT 17.640 751.810 17.780 753.030 ;
        RECT 19.020 751.810 19.160 871.350 ;
        RECT 16.260 751.670 19.160 751.810 ;
        RECT 15.740 718.090 16.000 718.410 ;
        RECT 16.260 717.670 16.400 751.670 ;
        RECT 17.640 751.130 17.780 751.670 ;
        RECT 17.640 750.990 18.240 751.130 ;
        RECT 18.100 717.810 18.240 750.990 ;
        RECT 17.640 717.670 18.240 717.810 ;
        RECT 16.260 717.530 16.860 717.670 ;
        RECT 16.720 711.010 16.860 717.530 ;
        RECT 9.760 654.260 14.560 654.400 ;
        RECT 14.880 710.870 16.860 711.010 ;
        RECT 9.760 654.170 10.020 654.260 ;
        RECT 14.880 653.890 15.020 710.870 ;
        RECT 15.340 694.690 15.480 710.870 ;
        RECT 17.640 698.770 17.780 717.670 ;
        RECT 16.720 698.630 17.780 698.770 ;
        RECT 16.720 696.050 16.860 698.630 ;
        RECT 16.720 695.910 17.320 696.050 ;
        RECT 17.180 694.690 17.320 695.910 ;
        RECT 15.340 694.550 19.160 694.690 ;
        RECT 17.180 694.180 17.320 694.550 ;
        RECT 17.180 694.040 17.780 694.180 ;
        RECT 17.640 692.650 17.780 694.040 ;
        RECT 17.640 692.510 18.240 692.650 ;
        RECT 9.820 653.750 15.020 653.890 ;
        RECT 9.820 653.130 9.960 653.750 ;
        RECT 9.760 652.810 10.020 653.130 ;
        RECT 9.760 647.090 10.020 647.350 ;
        RECT 9.760 647.030 14.560 647.090 ;
        RECT 9.820 646.950 14.560 647.030 ;
        RECT 9.360 646.270 10.880 646.410 ;
        RECT 9.760 645.900 10.020 645.990 ;
        RECT 10.740 645.900 10.880 646.270 ;
        RECT 14.420 645.900 14.560 646.950 ;
        RECT 9.760 645.760 10.420 645.900 ;
        RECT 10.740 645.760 14.100 645.900 ;
        RECT 14.420 645.760 15.480 645.900 ;
        RECT 9.760 645.670 10.020 645.760 ;
        RECT 9.300 641.590 9.560 641.910 ;
        RECT 9.360 632.050 9.500 641.590 ;
        RECT 10.280 640.290 10.420 645.760 ;
        RECT 10.280 640.150 11.800 640.290 ;
        RECT 9.300 631.730 9.560 632.050 ;
        RECT 11.660 601.530 11.800 640.150 ;
        RECT 13.960 624.480 14.100 645.760 ;
        RECT 13.960 624.340 14.560 624.480 ;
        RECT 11.660 601.390 14.100 601.530 ;
        RECT 6.080 587.530 6.340 587.850 ;
        RECT 9.760 587.760 10.020 587.850 ;
        RECT 13.960 587.760 14.100 601.390 ;
        RECT 9.760 587.620 14.100 587.760 ;
        RECT 9.760 587.530 10.020 587.620 ;
        RECT 6.140 575.610 6.280 587.530 ;
        RECT 9.760 586.850 10.020 587.170 ;
        RECT 6.080 575.290 6.340 575.610 ;
        RECT 9.820 555.210 9.960 586.850 ;
        RECT 9.760 554.890 10.020 555.210 ;
        RECT 14.420 551.890 14.560 624.340 ;
        RECT 15.340 623.290 15.480 645.760 ;
        RECT 18.100 624.820 18.240 692.510 ;
        RECT 17.640 624.680 18.240 624.820 ;
        RECT 15.340 623.150 17.320 623.290 ;
        RECT 17.180 589.120 17.320 623.150 ;
        RECT 11.200 551.750 14.560 551.890 ;
        RECT 16.260 588.980 17.320 589.120 ;
        RECT 11.200 551.210 11.340 551.750 ;
        RECT 16.260 551.210 16.400 588.980 ;
        RECT 17.640 584.530 17.780 624.680 ;
        RECT 19.020 620.570 19.160 694.550 ;
        RECT 10.280 551.070 11.340 551.210 ;
        RECT 11.660 551.070 16.400 551.210 ;
        RECT 16.720 584.390 17.780 584.530 ;
        RECT 18.100 620.430 19.160 620.570 ;
        RECT 10.280 550.530 10.420 551.070 ;
        RECT 9.820 550.450 10.420 550.530 ;
        RECT 6.080 550.130 6.340 550.450 ;
        RECT 9.760 550.390 10.420 550.450 ;
        RECT 9.760 550.130 10.020 550.390 ;
        RECT 6.140 541.125 6.280 550.130 ;
        RECT 9.760 548.660 10.020 548.750 ;
        RECT 11.660 548.660 11.800 551.070 ;
        RECT 16.720 549.850 16.860 584.390 ;
        RECT 18.100 572.970 18.240 620.430 ;
        RECT 18.100 572.830 18.700 572.970 ;
        RECT 15.340 549.710 16.860 549.850 ;
        RECT 9.760 548.520 11.800 548.660 ;
        RECT 12.120 548.860 13.640 549.000 ;
        RECT 9.760 548.430 10.020 548.520 ;
        RECT 12.120 547.810 12.260 548.860 ;
        RECT 9.820 547.670 12.260 547.810 ;
        RECT 13.500 547.810 13.640 548.860 ;
        RECT 15.340 547.810 15.480 549.710 ;
        RECT 18.560 549.000 18.700 572.830 ;
        RECT 18.560 548.860 19.160 549.000 ;
        RECT 13.500 547.670 15.480 547.810 ;
        RECT 9.820 547.390 9.960 547.670 ;
        RECT 9.760 547.070 10.020 547.390 ;
        RECT 12.580 546.990 18.700 547.130 ;
        RECT 9.760 546.620 10.020 546.710 ;
        RECT 12.580 546.620 12.720 546.990 ;
        RECT 9.760 546.480 12.720 546.620 ;
        RECT 9.760 546.390 10.020 546.480 ;
        RECT 13.500 546.310 16.860 546.450 ;
        RECT 9.760 545.770 10.020 546.030 ;
        RECT 13.500 545.770 13.640 546.310 ;
        RECT 9.760 545.710 13.640 545.770 ;
        RECT 9.820 545.630 13.640 545.710 ;
        RECT 9.760 544.410 10.020 544.670 ;
        RECT 16.720 544.410 16.860 546.310 ;
        RECT 9.760 544.350 16.400 544.410 ;
        RECT 9.820 544.270 16.400 544.350 ;
        RECT 16.720 544.270 17.320 544.410 ;
        RECT 9.760 543.730 10.020 543.990 ;
        RECT 16.260 543.730 16.400 544.270 ;
        RECT 9.760 543.670 15.480 543.730 ;
        RECT 9.820 543.590 15.480 543.670 ;
        RECT 16.260 543.590 16.860 543.730 ;
        RECT 9.760 543.050 10.020 543.310 ;
        RECT 9.760 542.990 14.560 543.050 ;
        RECT 9.820 542.910 14.560 542.990 ;
        RECT 9.760 542.370 10.020 542.630 ;
        RECT 9.760 542.310 14.100 542.370 ;
        RECT 9.820 542.230 14.100 542.310 ;
        RECT 6.070 540.755 6.350 541.125 ;
        RECT 6.080 540.270 6.340 540.590 ;
        RECT 6.140 535.685 6.280 540.270 ;
        RECT 6.070 535.315 6.350 535.685 ;
        RECT 6.080 512.730 6.340 513.050 ;
        RECT 6.140 404.445 6.280 512.730 ;
        RECT 6.530 497.915 6.810 498.285 ;
        RECT 6.600 491.630 6.740 497.915 ;
        RECT 6.540 491.310 6.800 491.630 ;
        RECT 13.960 467.570 14.100 542.230 ;
        RECT 9.360 467.490 14.100 467.570 ;
        RECT 9.300 467.430 14.100 467.490 ;
        RECT 9.300 467.170 9.560 467.430 ;
        RECT 9.760 467.060 10.020 467.150 ;
        RECT 14.420 467.060 14.560 542.910 ;
        RECT 15.340 528.090 15.480 543.590 ;
        RECT 15.340 527.950 16.400 528.090 ;
        RECT 16.260 503.610 16.400 527.950 ;
        RECT 9.760 466.920 14.560 467.060 ;
        RECT 15.340 503.470 16.400 503.610 ;
        RECT 9.760 466.830 10.020 466.920 ;
        RECT 9.760 466.380 10.020 466.470 ;
        RECT 9.760 466.240 14.100 466.380 ;
        RECT 9.760 466.150 10.020 466.240 ;
        RECT 9.760 460.940 10.020 461.030 ;
        RECT 13.960 460.940 14.100 466.240 ;
        RECT 9.760 460.800 14.100 460.940 ;
        RECT 9.760 460.710 10.020 460.800 ;
        RECT 9.760 460.090 10.020 460.350 ;
        RECT 15.340 460.090 15.480 503.470 ;
        RECT 9.760 460.030 15.480 460.090 ;
        RECT 9.820 459.950 15.480 460.030 ;
        RECT 9.760 459.410 10.020 459.670 ;
        RECT 9.760 459.350 14.100 459.410 ;
        RECT 9.820 459.270 14.100 459.350 ;
        RECT 9.760 457.540 10.020 457.630 ;
        RECT 9.760 457.400 11.800 457.540 ;
        RECT 9.760 457.310 10.020 457.400 ;
        RECT 9.300 430.450 9.560 430.770 ;
        RECT 9.360 418.610 9.500 430.450 ;
        RECT 11.660 424.730 11.800 457.400 ;
        RECT 9.820 424.590 11.800 424.730 ;
        RECT 9.820 423.970 9.960 424.590 ;
        RECT 9.760 423.650 10.020 423.970 ;
        RECT 13.960 419.970 14.100 459.270 ;
        RECT 16.720 448.530 16.860 543.590 ;
        RECT 14.880 448.390 16.860 448.530 ;
        RECT 14.880 420.650 15.020 448.390 ;
        RECT 17.180 441.050 17.320 544.270 ;
        RECT 17.570 480.235 17.850 480.605 ;
        RECT 15.340 440.910 17.320 441.050 ;
        RECT 15.340 421.330 15.480 440.910 ;
        RECT 17.640 439.010 17.780 480.235 ;
        RECT 18.560 474.370 18.700 546.990 ;
        RECT 19.020 474.370 19.160 548.860 ;
        RECT 17.180 438.870 17.780 439.010 ;
        RECT 18.100 474.230 19.160 474.370 ;
        RECT 15.340 421.190 16.400 421.330 ;
        RECT 14.880 420.510 15.940 420.650 ;
        RECT 13.960 419.830 15.020 419.970 ;
        RECT 9.360 418.470 14.560 418.610 ;
        RECT 9.760 417.930 10.020 418.190 ;
        RECT 9.760 417.870 14.100 417.930 ;
        RECT 9.820 417.790 14.100 417.870 ;
        RECT 13.960 413.170 14.100 417.790 ;
        RECT 11.660 413.030 14.100 413.170 ;
        RECT 9.760 410.450 10.020 410.710 ;
        RECT 9.760 410.390 10.420 410.450 ;
        RECT 9.820 410.310 10.420 410.390 ;
        RECT 6.070 404.075 6.350 404.445 ;
        RECT 10.280 360.130 10.420 410.310 ;
        RECT 9.820 360.050 10.420 360.130 ;
        RECT 9.760 359.990 10.420 360.050 ;
        RECT 9.760 359.730 10.020 359.990 ;
        RECT 11.660 355.370 11.800 413.030 ;
        RECT 14.420 412.490 14.560 418.470 ;
        RECT 9.820 355.290 11.800 355.370 ;
        RECT 6.080 354.970 6.340 355.290 ;
        RECT 9.760 355.230 11.800 355.290 ;
        RECT 12.580 412.350 14.560 412.490 ;
        RECT 9.760 354.970 10.020 355.230 ;
        RECT 6.140 327.410 6.280 354.970 ;
        RECT 12.580 338.370 12.720 412.350 ;
        RECT 14.880 394.130 15.020 419.830 ;
        RECT 15.800 419.290 15.940 420.510 ;
        RECT 16.260 419.970 16.400 421.190 ;
        RECT 16.260 419.830 16.860 419.970 ;
        RECT 15.800 419.150 16.400 419.290 ;
        RECT 13.040 393.990 15.020 394.130 ;
        RECT 13.040 380.530 13.180 393.990 ;
        RECT 16.260 387.330 16.400 419.150 ;
        RECT 16.720 415.210 16.860 419.830 ;
        RECT 17.180 417.930 17.320 438.870 ;
        RECT 18.100 424.730 18.240 474.230 ;
        RECT 18.560 451.930 18.700 474.230 ;
        RECT 18.560 451.790 19.160 451.930 ;
        RECT 17.640 424.590 18.240 424.730 ;
        RECT 17.640 417.930 17.780 424.590 ;
        RECT 17.180 417.790 18.240 417.930 ;
        RECT 16.720 415.070 17.320 415.210 ;
        RECT 14.880 387.190 16.400 387.330 ;
        RECT 13.040 380.390 14.560 380.530 ;
        RECT 14.420 377.810 14.560 380.390 ;
        RECT 14.880 377.810 15.020 387.190 ;
        RECT 17.180 385.290 17.320 415.070 ;
        RECT 13.500 377.670 15.020 377.810 ;
        RECT 15.340 385.150 17.320 385.290 ;
        RECT 13.500 359.960 13.640 377.670 ;
        RECT 10.280 338.230 12.720 338.370 ;
        RECT 13.040 359.820 13.640 359.960 ;
        RECT 10.280 337.690 10.420 338.230 ;
        RECT 9.820 337.610 10.420 337.690 ;
        RECT 9.760 337.550 10.420 337.610 ;
        RECT 9.760 337.290 10.020 337.550 ;
        RECT 13.040 337.010 13.180 359.820 ;
        RECT 14.420 359.450 14.560 377.670 ;
        RECT 9.820 336.930 13.180 337.010 ;
        RECT 6.540 336.610 6.800 336.930 ;
        RECT 9.760 336.870 13.180 336.930 ;
        RECT 13.500 359.310 14.560 359.450 ;
        RECT 9.760 336.610 10.020 336.870 ;
        RECT 6.080 327.090 6.340 327.410 ;
        RECT 6.600 326.810 6.740 336.610 ;
        RECT 13.500 336.330 13.640 359.310 ;
        RECT 9.820 336.250 13.640 336.330 ;
        RECT 9.760 336.190 13.640 336.250 ;
        RECT 9.760 335.930 10.020 336.190 ;
        RECT 9.760 333.780 10.020 333.870 ;
        RECT 9.760 333.640 13.640 333.780 ;
        RECT 9.760 333.550 10.020 333.640 ;
        RECT 9.760 332.930 10.020 333.190 ;
        RECT 9.760 332.870 13.180 332.930 ;
        RECT 9.820 332.790 13.180 332.870 ;
        RECT 13.040 331.570 13.180 332.790 ;
        RECT 13.500 332.250 13.640 333.640 ;
        RECT 15.340 333.610 15.480 385.150 ;
        RECT 17.640 365.570 17.780 417.790 ;
        RECT 17.180 365.430 17.780 365.570 ;
        RECT 17.180 345.170 17.320 365.430 ;
        RECT 14.880 333.470 15.480 333.610 ;
        RECT 16.720 345.030 17.320 345.170 ;
        RECT 14.880 332.250 15.020 333.470 ;
        RECT 13.500 332.110 15.020 332.250 ;
        RECT 16.720 331.570 16.860 345.030 ;
        RECT 13.040 331.430 16.860 331.570 ;
        RECT 10.220 327.090 10.480 327.410 ;
        RECT 6.140 326.670 6.740 326.810 ;
        RECT 6.140 316.870 6.280 326.670 ;
        RECT 6.540 326.070 6.800 326.390 ;
        RECT 6.080 316.550 6.340 316.870 ;
        RECT 6.600 290.205 6.740 326.070 ;
        RECT 10.280 324.770 10.420 327.090 ;
        RECT 18.100 324.770 18.240 417.790 ;
        RECT 19.020 377.130 19.160 451.790 ;
        RECT 18.560 376.990 19.160 377.130 ;
        RECT 18.560 374.410 18.700 376.990 ;
        RECT 18.560 374.270 19.160 374.410 ;
        RECT 10.280 324.630 18.240 324.770 ;
        RECT 19.020 324.090 19.160 374.270 ;
        RECT 18.100 323.950 19.160 324.090 ;
        RECT 9.760 323.240 10.020 323.330 ;
        RECT 9.760 323.100 15.020 323.240 ;
        RECT 9.760 323.010 10.020 323.100 ;
        RECT 9.760 316.610 10.020 316.870 ;
        RECT 9.760 316.550 14.100 316.610 ;
        RECT 9.820 316.470 14.100 316.550 ;
        RECT 9.760 315.760 10.020 315.850 ;
        RECT 9.760 315.620 13.640 315.760 ;
        RECT 9.760 315.530 10.020 315.620 ;
        RECT 9.760 314.170 10.020 314.490 ;
        RECT 9.820 313.890 9.960 314.170 ;
        RECT 9.820 313.750 11.340 313.890 ;
        RECT 9.760 311.340 10.020 311.430 ;
        RECT 9.760 311.200 10.880 311.340 ;
        RECT 9.760 311.110 10.020 311.200 ;
        RECT 6.530 289.835 6.810 290.205 ;
        RECT 6.540 289.350 6.800 289.670 ;
        RECT 5.160 251.610 5.420 251.930 ;
        RECT 6.600 229.685 6.740 289.350 ;
        RECT 9.760 285.500 10.020 285.590 ;
        RECT 10.740 285.500 10.880 311.200 ;
        RECT 9.760 285.360 10.880 285.500 ;
        RECT 9.760 285.270 10.020 285.360 ;
        RECT 9.760 284.480 10.020 284.570 ;
        RECT 11.200 284.480 11.340 313.750 ;
        RECT 9.760 284.340 11.340 284.480 ;
        RECT 9.760 284.250 10.020 284.340 ;
        RECT 9.760 282.890 10.020 283.210 ;
        RECT 9.820 279.890 9.960 282.890 ;
        RECT 9.820 279.750 13.180 279.890 ;
        RECT 9.760 279.380 10.020 279.470 ;
        RECT 9.760 279.240 12.720 279.380 ;
        RECT 9.760 279.150 10.020 279.240 ;
        RECT 9.760 262.830 10.020 263.150 ;
        RECT 6.530 229.315 6.810 229.685 ;
        RECT 9.820 215.970 9.960 262.830 ;
        RECT 12.580 218.010 12.720 279.240 ;
        RECT 13.040 218.690 13.180 279.750 ;
        RECT 13.500 222.770 13.640 315.620 ;
        RECT 13.960 315.080 14.100 316.470 ;
        RECT 14.880 315.760 15.020 323.100 ;
        RECT 14.880 315.620 17.780 315.760 ;
        RECT 13.960 314.940 15.940 315.080 ;
        RECT 15.800 255.410 15.940 314.940 ;
        RECT 17.640 255.410 17.780 315.620 ;
        RECT 18.100 282.610 18.240 323.950 ;
        RECT 18.100 282.470 18.700 282.610 ;
        RECT 13.960 255.270 15.940 255.410 ;
        RECT 16.720 255.270 17.780 255.410 ;
        RECT 13.960 224.130 14.100 255.270 ;
        RECT 16.720 254.050 16.860 255.270 ;
        RECT 18.560 254.730 18.700 282.470 ;
        RECT 18.560 254.590 19.160 254.730 ;
        RECT 16.720 253.910 17.780 254.050 ;
        RECT 13.960 223.990 16.400 224.130 ;
        RECT 13.500 222.630 15.480 222.770 ;
        RECT 13.040 218.550 14.100 218.690 ;
        RECT 13.960 218.010 14.100 218.550 ;
        RECT 12.580 217.870 13.180 218.010 ;
        RECT 13.960 217.870 14.560 218.010 ;
        RECT 13.040 217.330 13.180 217.870 ;
        RECT 13.040 217.190 14.100 217.330 ;
        RECT 9.820 215.830 10.880 215.970 ;
        RECT 10.740 215.290 10.880 215.830 ;
        RECT 10.740 215.150 12.720 215.290 ;
        RECT 5.160 184.970 5.420 185.290 ;
        RECT 5.220 100.290 5.360 184.970 ;
        RECT 12.580 177.890 12.720 215.150 ;
        RECT 9.820 177.810 12.720 177.890 ;
        RECT 9.760 177.750 12.720 177.810 ;
        RECT 9.760 177.490 10.020 177.750 ;
        RECT 13.960 173.130 14.100 217.190 ;
        RECT 9.360 172.990 14.100 173.130 ;
        RECT 7.450 151.115 7.730 151.485 ;
        RECT 7.520 147.550 7.660 151.115 ;
        RECT 9.360 148.910 9.500 172.990 ;
        RECT 14.420 149.330 14.560 217.870 ;
        RECT 15.340 202.370 15.480 222.630 ;
        RECT 16.260 203.050 16.400 223.990 ;
        RECT 17.640 213.930 17.780 253.910 ;
        RECT 17.640 213.790 18.240 213.930 ;
        RECT 18.100 203.730 18.240 213.790 ;
        RECT 19.020 203.730 19.160 254.590 ;
        RECT 17.180 203.590 19.160 203.730 ;
        RECT 17.180 203.050 17.320 203.590 ;
        RECT 18.100 203.050 18.240 203.590 ;
        RECT 16.260 202.910 18.700 203.050 ;
        RECT 15.340 202.230 16.860 202.370 ;
        RECT 16.720 178.400 16.860 202.230 ;
        RECT 10.280 149.190 14.560 149.330 ;
        RECT 15.340 178.260 16.860 178.400 ;
        RECT 9.300 148.590 9.560 148.910 ;
        RECT 7.460 147.230 7.720 147.550 ;
        RECT 10.280 141.850 10.420 149.190 ;
        RECT 9.820 141.770 10.420 141.850 ;
        RECT 9.760 141.710 10.420 141.770 ;
        RECT 9.760 141.450 10.020 141.710 ;
        RECT 15.340 140.490 15.480 178.260 ;
        RECT 17.180 177.720 17.320 202.910 ;
        RECT 18.100 200.330 18.240 202.910 ;
        RECT 17.640 200.190 18.240 200.330 ;
        RECT 17.640 186.050 17.780 200.190 ;
        RECT 17.640 185.910 18.240 186.050 ;
        RECT 9.820 140.350 15.480 140.490 ;
        RECT 16.260 177.580 17.320 177.720 ;
        RECT 9.820 140.070 9.960 140.350 ;
        RECT 7.460 139.750 7.720 140.070 ;
        RECT 9.760 139.750 10.020 140.070 ;
        RECT 6.070 134.795 6.350 135.165 ;
        RECT 6.080 134.650 6.340 134.795 ;
        RECT 7.520 134.290 7.660 139.750 ;
        RECT 16.260 139.130 16.400 177.580 ;
        RECT 18.100 177.040 18.240 185.910 ;
        RECT 9.360 138.990 16.400 139.130 ;
        RECT 17.180 176.900 18.240 177.040 ;
        RECT 7.460 133.970 7.720 134.290 ;
        RECT 9.360 118.730 9.500 138.990 ;
        RECT 17.180 138.450 17.320 176.900 ;
        RECT 18.560 169.050 18.700 202.910 ;
        RECT 18.950 201.435 19.230 201.805 ;
        RECT 16.720 138.310 17.320 138.450 ;
        RECT 18.100 168.910 18.700 169.050 ;
        RECT 16.720 136.410 16.860 138.310 ;
        RECT 9.820 136.330 16.860 136.410 ;
        RECT 9.760 136.270 16.860 136.330 ;
        RECT 9.760 136.010 10.020 136.270 ;
        RECT 9.760 135.560 10.020 135.650 ;
        RECT 9.760 135.420 15.480 135.560 ;
        RECT 9.760 135.330 10.020 135.420 ;
        RECT 9.760 134.880 10.020 134.970 ;
        RECT 9.760 134.740 14.100 134.880 ;
        RECT 9.760 134.650 10.020 134.740 ;
        RECT 13.960 134.370 14.100 134.740 ;
        RECT 9.760 133.970 10.020 134.290 ;
        RECT 13.960 134.230 14.560 134.370 ;
        RECT 9.820 133.690 9.960 133.970 ;
        RECT 9.820 133.550 14.100 133.690 ;
        RECT 9.360 118.590 12.720 118.730 ;
        RECT 9.760 111.080 10.020 111.170 ;
        RECT 9.760 110.940 11.340 111.080 ;
        RECT 9.760 110.850 10.020 110.940 ;
        RECT 5.160 99.970 5.420 100.290 ;
        RECT 6.540 94.190 6.800 94.510 ;
        RECT 5.620 77.870 5.880 78.190 ;
        RECT 5.680 74.110 5.820 77.870 ;
        RECT 5.620 73.790 5.880 74.110 ;
        RECT 5.620 61.550 5.880 61.870 ;
        RECT 5.680 61.045 5.820 61.550 ;
        RECT 6.600 61.190 6.740 94.190 ;
        RECT 11.200 90.170 11.340 110.940 ;
        RECT 9.360 90.030 11.340 90.170 ;
        RECT 9.360 89.750 9.500 90.030 ;
        RECT 9.300 89.430 9.560 89.750 ;
        RECT 9.300 82.690 9.560 82.950 ;
        RECT 12.580 82.690 12.720 118.590 ;
        RECT 13.960 107.850 14.100 133.550 ;
        RECT 13.500 107.710 14.100 107.850 ;
        RECT 13.500 88.130 13.640 107.710 ;
        RECT 13.500 87.990 14.100 88.130 ;
        RECT 9.300 82.630 12.720 82.690 ;
        RECT 9.360 82.550 12.720 82.630 ;
        RECT 9.300 82.010 9.560 82.270 ;
        RECT 9.300 81.950 10.420 82.010 ;
        RECT 9.360 81.870 10.420 81.950 ;
        RECT 10.280 81.330 10.420 81.870 ;
        RECT 13.960 81.330 14.100 87.990 ;
        RECT 10.280 81.190 14.100 81.330 ;
        RECT 14.420 80.480 14.560 134.230 ;
        RECT 15.340 83.370 15.480 135.420 ;
        RECT 18.100 83.370 18.240 168.910 ;
        RECT 13.040 80.340 14.560 80.480 ;
        RECT 14.880 83.230 18.240 83.370 ;
        RECT 13.040 79.800 13.180 80.340 ;
        RECT 14.880 79.800 15.020 83.230 ;
        RECT 15.340 82.860 15.480 83.230 ;
        RECT 15.340 82.720 18.700 82.860 ;
        RECT 10.280 79.660 15.020 79.800 ;
        RECT 9.760 78.100 10.020 78.190 ;
        RECT 10.280 78.100 10.420 79.660 ;
        RECT 13.040 79.290 13.180 79.660 ;
        RECT 13.040 79.150 18.240 79.290 ;
        RECT 9.760 77.960 10.420 78.100 ;
        RECT 9.760 77.870 10.020 77.960 ;
        RECT 9.760 76.740 10.020 76.830 ;
        RECT 9.760 76.600 10.880 76.740 ;
        RECT 9.760 76.510 10.020 76.600 ;
        RECT 9.760 75.490 10.020 75.810 ;
        RECT 9.820 67.650 9.960 75.490 ;
        RECT 10.740 75.040 10.880 76.600 ;
        RECT 10.740 74.900 17.320 75.040 ;
        RECT 9.760 67.330 10.020 67.650 ;
        RECT 9.760 66.880 10.020 66.970 ;
        RECT 9.760 66.740 16.860 66.880 ;
        RECT 9.760 66.650 10.020 66.740 ;
        RECT 5.610 60.675 5.890 61.045 ;
        RECT 6.540 60.870 6.800 61.190 ;
        RECT 5.160 50.330 5.420 50.650 ;
        RECT 4.240 37.410 4.500 37.730 ;
        RECT 4.300 3.730 4.440 37.410 ;
        RECT 4.240 3.410 4.500 3.730 ;
        RECT 5.220 2.370 5.360 50.330 ;
        RECT 6.080 16.330 6.340 16.650 ;
        RECT 6.140 5.285 6.280 16.330 ;
        RECT 6.070 4.915 6.350 5.285 ;
        RECT 16.720 4.750 16.860 66.740 ;
        RECT 16.660 4.430 16.920 4.750 ;
        RECT 5.160 2.050 5.420 2.370 ;
        RECT 17.180 1.205 17.320 74.900 ;
        RECT 18.100 2.710 18.240 79.150 ;
        RECT 18.560 7.325 18.700 82.720 ;
        RECT 19.020 8.830 19.160 201.435 ;
        RECT 18.960 8.510 19.220 8.830 ;
        RECT 38.280 8.510 38.540 8.830 ;
        RECT 18.490 6.955 18.770 7.325 ;
        RECT 29.530 6.955 29.810 7.325 ;
        RECT 29.540 6.810 29.800 6.955 ;
        RECT 32.300 6.810 32.560 7.130 ;
        RECT 24.940 6.530 25.200 6.790 ;
        RECT 26.780 6.530 27.040 6.790 ;
        RECT 24.940 6.470 27.040 6.530 ;
        RECT 25.000 6.390 26.980 6.470 ;
        RECT 18.040 2.390 18.300 2.710 ;
        RECT 32.360 2.400 32.500 6.810 ;
        RECT 38.340 2.400 38.480 8.510 ;
        RECT 90.260 7.490 90.520 7.810 ;
        RECT 90.320 6.790 90.460 7.490 ;
        RECT 72.780 6.470 73.040 6.790 ;
        RECT 90.260 6.470 90.520 6.790 ;
        RECT 52.540 2.730 52.800 3.050 ;
        RECT 67.250 2.875 67.530 3.245 ;
        RECT 67.260 2.730 67.520 2.875 ;
        RECT 17.110 0.835 17.390 1.205 ;
        RECT 32.150 -4.800 32.710 2.400 ;
        RECT 38.130 -4.800 38.690 2.400 ;
        RECT 52.600 1.770 52.740 2.730 ;
        RECT 52.140 1.630 52.740 1.770 ;
        RECT 52.140 1.350 52.280 1.630 ;
        RECT 52.080 1.030 52.340 1.350 ;
        RECT 72.840 1.205 72.980 6.470 ;
        RECT 121.540 5.850 121.800 6.110 ;
        RECT 123.310 5.850 123.590 9.000 ;
        RECT 170.690 5.850 170.970 9.000 ;
        RECT 283.920 8.170 284.180 8.490 ;
        RECT 121.540 5.790 123.590 5.850 ;
        RECT 121.600 5.710 123.590 5.790 ;
        RECT 169.440 5.770 170.970 5.850 ;
        RECT 123.310 5.000 123.590 5.710 ;
        RECT 169.380 5.710 170.970 5.770 ;
        RECT 169.380 5.450 169.640 5.710 ;
        RECT 134.410 4.915 134.690 5.285 ;
        RECT 170.690 5.000 170.970 5.710 ;
        RECT 103.590 2.875 103.870 3.245 ;
        RECT 103.660 2.400 103.800 2.875 ;
        RECT 65.410 0.835 65.690 1.205 ;
        RECT 72.770 0.835 73.050 1.205 ;
        RECT 65.480 0.330 65.620 0.835 ;
        RECT 65.420 0.010 65.680 0.330 ;
        RECT 103.450 -4.800 104.010 2.400 ;
        RECT 134.480 1.690 134.620 4.915 ;
        RECT 283.980 4.750 284.120 8.170 ;
        RECT 394.320 5.450 394.580 5.770 ;
        RECT 519.900 5.450 520.160 5.770 ;
        RECT 283.920 4.430 284.180 4.750 ;
        RECT 233.320 4.090 233.580 4.410 ;
        RECT 168.520 2.990 169.580 3.130 ;
        RECT 168.520 2.565 168.660 2.990 ;
        RECT 168.450 2.195 168.730 2.565 ;
        RECT 169.440 2.400 169.580 2.990 ;
        RECT 227.860 2.990 228.920 3.130 ;
        RECT 227.860 2.565 228.000 2.990 ;
        RECT 134.420 1.370 134.680 1.690 ;
        RECT 169.230 -4.800 169.790 2.400 ;
        RECT 175.810 2.195 176.090 2.565 ;
        RECT 227.790 2.195 228.070 2.565 ;
        RECT 228.780 2.400 228.920 2.990 ;
        RECT 233.380 2.565 233.520 4.090 ;
        RECT 293.180 2.990 294.240 3.130 ;
        RECT 175.880 1.690 176.020 2.195 ;
        RECT 175.820 1.370 176.080 1.690 ;
        RECT 228.570 -4.800 229.130 2.400 ;
        RECT 233.310 2.195 233.590 2.565 ;
        RECT 249.410 2.195 249.690 2.565 ;
        RECT 249.480 1.010 249.620 2.195 ;
        RECT 293.180 1.010 293.320 2.990 ;
        RECT 294.100 2.400 294.240 2.990 ;
        RECT 249.420 0.690 249.680 1.010 ;
        RECT 293.120 0.690 293.380 1.010 ;
        RECT 293.890 -4.800 294.450 2.400 ;
        RECT 394.380 0.525 394.520 5.450 ;
        RECT 519.960 5.170 520.100 5.450 ;
        RECT 519.960 5.030 532.060 5.170 ;
        RECT 453.720 3.160 460.760 3.300 ;
        RECT 453.720 2.030 453.860 3.160 ;
        RECT 460.620 2.400 460.760 3.160 ;
        RECT 531.920 2.400 532.060 5.030 ;
        RECT 421.060 1.630 422.580 1.770 ;
        RECT 453.660 1.710 453.920 2.030 ;
        RECT 421.060 1.205 421.200 1.630 ;
        RECT 420.990 0.835 421.270 1.205 ;
        RECT 422.440 1.010 422.580 1.630 ;
        RECT 422.380 0.690 422.640 1.010 ;
        RECT 394.310 0.155 394.590 0.525 ;
        RECT 460.410 -4.800 460.970 2.400 ;
        RECT 531.710 -4.800 532.270 2.400 ;
      LAYER via2 ;
        RECT 2807.930 3402.240 2808.210 3402.520 ;
        RECT 2806.090 3401.560 2806.370 3401.840 ;
        RECT 7.910 3005.120 8.190 3005.400 ;
        RECT 7.910 2891.560 8.190 2891.840 ;
        RECT 6.530 2836.480 6.810 2836.760 ;
        RECT 7.910 2665.120 8.190 2665.400 ;
        RECT 7.910 2549.520 8.190 2549.800 ;
        RECT 6.990 2261.880 7.270 2262.160 ;
        RECT 6.530 1687.280 6.810 1687.560 ;
        RECT 15.730 1698.160 16.010 1698.440 ;
        RECT 15.730 1605.000 16.010 1605.280 ;
        RECT 6.990 1471.720 7.270 1472.000 ;
        RECT 6.990 990.960 7.270 991.240 ;
        RECT 14.350 926.360 14.630 926.640 ;
        RECT 7.450 865.160 7.730 865.440 ;
        RECT 6.990 837.960 7.270 838.240 ;
        RECT 7.910 734.600 8.190 734.880 ;
        RECT 7.450 693.120 7.730 693.400 ;
        RECT 6.070 540.800 6.350 541.080 ;
        RECT 6.070 535.360 6.350 535.640 ;
        RECT 6.530 497.960 6.810 498.240 ;
        RECT 17.570 480.280 17.850 480.560 ;
        RECT 6.070 404.120 6.350 404.400 ;
        RECT 6.530 289.880 6.810 290.160 ;
        RECT 6.530 229.360 6.810 229.640 ;
        RECT 7.450 151.160 7.730 151.440 ;
        RECT 6.070 134.840 6.350 135.120 ;
        RECT 18.950 201.480 19.230 201.760 ;
        RECT 5.610 60.720 5.890 61.000 ;
        RECT 6.070 4.960 6.350 5.240 ;
        RECT 18.490 7.000 18.770 7.280 ;
        RECT 29.530 7.000 29.810 7.280 ;
        RECT 67.250 2.920 67.530 3.200 ;
        RECT 17.110 0.880 17.390 1.160 ;
        RECT 134.410 4.960 134.690 5.240 ;
        RECT 103.590 2.920 103.870 3.200 ;
        RECT 65.410 0.880 65.690 1.160 ;
        RECT 72.770 0.880 73.050 1.160 ;
        RECT 168.450 2.240 168.730 2.520 ;
        RECT 175.810 2.240 176.090 2.520 ;
        RECT 227.790 2.240 228.070 2.520 ;
        RECT 233.310 2.240 233.590 2.520 ;
        RECT 249.410 2.240 249.690 2.520 ;
        RECT 420.990 0.880 421.270 1.160 ;
        RECT 394.310 0.200 394.590 0.480 ;
      LAYER met3 ;
        RECT 2807.905 3402.540 2808.235 3402.545 ;
        RECT 2807.905 3402.530 2808.490 3402.540 ;
        RECT 2807.680 3402.230 2808.490 3402.530 ;
        RECT 2807.905 3402.220 2808.490 3402.230 ;
        RECT 2807.905 3402.215 2808.235 3402.220 ;
        RECT 2805.350 3401.850 2805.730 3401.860 ;
        RECT 2806.065 3401.850 2806.395 3401.865 ;
        RECT 2805.350 3401.550 2806.395 3401.850 ;
        RECT 2805.350 3401.540 2805.730 3401.550 ;
        RECT 2806.065 3401.535 2806.395 3401.550 ;
        RECT 5.000 3007.920 9.000 3008.520 ;
        RECT 7.670 3005.425 7.970 3007.920 ;
        RECT 7.670 3005.110 8.215 3005.425 ;
        RECT 7.885 3005.095 8.215 3005.110 ;
        RECT 5.000 2894.360 9.000 2894.960 ;
        RECT 7.670 2891.865 7.970 2894.360 ;
        RECT 7.670 2891.550 8.215 2891.865 ;
        RECT 7.885 2891.535 8.215 2891.550 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 6.505 2836.770 6.835 2836.785 ;
        RECT -4.800 2836.470 6.835 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 6.505 2836.455 6.835 2836.470 ;
        RECT 5.000 2667.920 9.000 2668.520 ;
        RECT 7.670 2665.425 7.970 2667.920 ;
        RECT 7.670 2665.110 8.215 2665.425 ;
        RECT 7.885 2665.095 8.215 2665.110 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 7.885 2549.810 8.215 2549.825 ;
        RECT -4.800 2549.510 8.215 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 7.885 2549.495 8.215 2549.510 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 6.965 2262.170 7.295 2262.185 ;
        RECT -4.800 2261.870 7.295 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 6.965 2261.855 7.295 2261.870 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 6.505 1687.570 6.835 1687.585 ;
        RECT -4.800 1687.270 6.835 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
        RECT 6.505 1687.255 6.835 1687.270 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 6.965 1472.010 7.295 1472.025 ;
        RECT -4.800 1471.710 7.295 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 6.965 1471.695 7.295 1471.710 ;
        RECT 6.965 991.250 7.295 991.265 ;
        RECT 7.630 991.250 8.010 991.260 ;
        RECT 6.965 990.950 8.010 991.250 ;
        RECT 6.965 990.935 7.295 990.950 ;
        RECT 7.630 990.940 8.010 990.950 ;
        RECT 7.425 865.460 7.755 865.465 ;
        RECT 7.425 865.450 8.010 865.460 ;
        RECT 7.200 865.150 8.010 865.450 ;
        RECT 7.425 865.140 8.010 865.150 ;
        RECT 7.425 865.135 7.755 865.140 ;
        RECT 6.965 838.250 7.295 838.265 ;
        RECT 7.630 838.250 8.010 838.260 ;
        RECT 6.965 837.950 8.010 838.250 ;
        RECT 6.965 837.935 7.295 837.950 ;
        RECT 7.630 837.940 8.010 837.950 ;
        RECT 7.885 734.900 8.215 734.905 ;
        RECT 7.630 734.890 8.215 734.900 ;
        RECT 7.430 734.590 8.215 734.890 ;
        RECT 7.630 734.580 8.215 734.590 ;
        RECT 7.885 734.575 8.215 734.580 ;
        RECT 7.425 693.420 7.755 693.425 ;
        RECT 7.425 693.410 8.010 693.420 ;
        RECT 7.425 693.110 8.210 693.410 ;
        RECT 7.425 693.100 8.010 693.110 ;
        RECT 7.425 693.095 7.755 693.100 ;
        RECT 6.045 541.090 6.375 541.105 ;
        RECT 6.710 541.090 7.090 541.100 ;
        RECT 6.045 540.790 7.090 541.090 ;
        RECT 6.045 540.775 6.375 540.790 ;
        RECT 6.710 540.780 7.090 540.790 ;
        RECT 6.045 535.650 6.375 535.665 ;
        RECT 7.630 535.650 8.010 535.660 ;
        RECT 6.045 535.350 8.010 535.650 ;
        RECT 6.045 535.335 6.375 535.350 ;
        RECT 7.630 535.340 8.010 535.350 ;
        RECT 6.505 498.250 6.835 498.265 ;
        RECT 7.630 498.250 8.010 498.260 ;
        RECT 6.505 497.950 8.010 498.250 ;
        RECT 6.505 497.935 6.835 497.950 ;
        RECT 7.630 497.940 8.010 497.950 ;
        RECT 6.045 404.410 6.375 404.425 ;
        RECT 5.830 404.095 6.375 404.410 ;
        RECT 5.830 402.080 6.130 404.095 ;
        RECT 5.000 401.480 9.000 402.080 ;
        RECT 6.505 290.170 6.835 290.185 ;
        RECT 6.505 289.855 7.050 290.170 ;
        RECT 6.750 288.520 7.050 289.855 ;
        RECT 5.000 287.920 9.000 288.520 ;
        RECT 6.505 229.650 6.835 229.665 ;
        RECT 7.630 229.650 8.010 229.660 ;
        RECT 6.505 229.350 8.010 229.650 ;
        RECT 6.505 229.335 6.835 229.350 ;
        RECT 7.630 229.340 8.010 229.350 ;
        RECT 19.020 201.480 19.230 201.760 ;
        RECT 7.425 151.460 7.755 151.465 ;
        RECT 7.425 151.450 8.010 151.460 ;
        RECT 7.425 151.150 8.210 151.450 ;
        RECT 7.425 151.140 8.010 151.150 ;
        RECT 7.425 151.135 7.755 151.140 ;
        RECT 6.045 135.130 6.375 135.145 ;
        RECT 7.630 135.130 8.010 135.140 ;
        RECT 6.045 134.830 8.010 135.130 ;
        RECT 6.045 134.815 6.375 134.830 ;
        RECT 7.630 134.820 8.010 134.830 ;
        RECT 5.000 61.480 9.000 62.080 ;
        RECT 5.830 61.025 6.130 61.480 ;
        RECT 5.585 60.710 6.130 61.025 ;
        RECT 5.585 60.695 5.915 60.710 ;
        RECT 18.465 7.290 18.795 7.305 ;
        RECT 29.505 7.290 29.835 7.305 ;
        RECT 18.465 6.990 29.835 7.290 ;
        RECT 18.465 6.975 18.795 6.990 ;
        RECT 29.505 6.975 29.835 6.990 ;
        RECT 6.045 5.250 6.375 5.265 ;
        RECT 134.385 5.250 134.715 5.265 ;
        RECT 6.045 4.950 134.715 5.250 ;
        RECT 6.045 4.935 6.375 4.950 ;
        RECT 134.385 4.935 134.715 4.950 ;
        RECT 67.225 3.210 67.555 3.225 ;
        RECT 103.565 3.210 103.895 3.225 ;
        RECT 67.225 2.910 103.895 3.210 ;
        RECT 67.225 2.895 67.555 2.910 ;
        RECT 103.565 2.895 103.895 2.910 ;
        RECT 168.425 2.530 168.755 2.545 ;
        RECT 54.590 2.230 168.755 2.530 ;
        RECT 17.085 1.170 17.415 1.185 ;
        RECT 54.590 1.170 54.890 2.230 ;
        RECT 168.425 2.215 168.755 2.230 ;
        RECT 175.785 2.530 176.115 2.545 ;
        RECT 227.765 2.530 228.095 2.545 ;
        RECT 175.785 2.230 228.095 2.530 ;
        RECT 175.785 2.215 176.115 2.230 ;
        RECT 227.765 2.215 228.095 2.230 ;
        RECT 233.285 2.530 233.615 2.545 ;
        RECT 249.385 2.530 249.715 2.545 ;
        RECT 233.285 2.230 249.715 2.530 ;
        RECT 233.285 2.215 233.615 2.230 ;
        RECT 249.385 2.215 249.715 2.230 ;
        RECT 17.085 0.870 54.890 1.170 ;
        RECT 65.385 1.170 65.715 1.185 ;
        RECT 72.745 1.170 73.075 1.185 ;
        RECT 65.385 0.870 73.075 1.170 ;
        RECT 17.085 0.855 17.415 0.870 ;
        RECT 65.385 0.855 65.715 0.870 ;
        RECT 72.745 0.855 73.075 0.870 ;
        RECT 411.510 1.170 411.890 1.180 ;
        RECT 420.965 1.170 421.295 1.185 ;
        RECT 411.510 0.870 421.295 1.170 ;
        RECT 411.510 0.860 411.890 0.870 ;
        RECT 420.965 0.855 421.295 0.870 ;
        RECT 394.285 0.490 394.615 0.505 ;
        RECT 406.910 0.490 407.290 0.500 ;
        RECT 394.285 0.190 407.290 0.490 ;
        RECT 394.285 0.175 394.615 0.190 ;
        RECT 406.910 0.180 407.290 0.190 ;
      LAYER via3 ;
        RECT 2808.140 3402.220 2808.460 3402.540 ;
        RECT 2805.380 3401.540 2805.700 3401.860 ;
        RECT 7.660 990.940 7.980 991.260 ;
        RECT 7.660 865.140 7.980 865.460 ;
        RECT 7.660 837.940 7.980 838.260 ;
        RECT 7.660 734.580 7.980 734.900 ;
        RECT 7.660 693.100 7.980 693.420 ;
        RECT 6.740 540.780 7.060 541.100 ;
        RECT 7.660 535.340 7.980 535.660 ;
        RECT 7.660 497.940 7.980 498.260 ;
        RECT 7.660 229.340 7.980 229.660 ;
        RECT 7.660 151.140 7.980 151.460 ;
        RECT 7.660 134.820 7.980 135.140 ;
        RECT 411.540 0.860 411.860 1.180 ;
        RECT 406.940 0.180 407.260 0.500 ;
      LAYER met4 ;
        RECT 2808.135 3402.215 2808.465 3402.545 ;
        RECT 2805.375 3401.535 2805.705 3401.865 ;
        RECT 15.705 1698.450 16.035 1698.465 ;
        RECT 15.705 1698.150 17.170 1698.450 ;
        RECT 15.705 1698.135 16.035 1698.150 ;
        RECT 16.870 1671.080 17.170 1698.150 ;
        RECT 15.950 1670.780 17.170 1671.080 ;
        RECT 15.950 1633.850 16.250 1670.780 ;
        RECT 15.950 1633.550 17.170 1633.850 ;
        RECT 16.870 1620.250 17.170 1633.550 ;
        RECT 15.950 1619.950 17.170 1620.250 ;
        RECT 15.950 1616.850 16.250 1619.950 ;
        RECT 15.720 1616.550 16.250 1616.850 ;
        RECT 15.720 1605.305 16.020 1616.550 ;
        RECT 15.705 1604.975 16.035 1605.305 ;
        RECT 7.655 990.935 7.985 991.265 ;
        RECT 7.670 926.650 7.970 990.935 ;
        RECT 2805.390 987.850 2805.690 3401.535 ;
        RECT 2803.550 987.550 2805.690 987.850 ;
        RECT 2803.550 970.850 2803.850 987.550 ;
        RECT 2803.550 970.550 2805.690 970.850 ;
        RECT 14.325 926.650 14.655 926.665 ;
        RECT 7.670 926.350 14.655 926.650 ;
        RECT 14.325 926.335 14.655 926.350 ;
        RECT 7.655 865.135 7.985 865.465 ;
        RECT 7.670 838.265 7.970 865.135 ;
        RECT 7.655 837.935 7.985 838.265 ;
        RECT 7.655 734.575 7.985 734.905 ;
        RECT 7.670 693.425 7.970 734.575 ;
        RECT 7.655 693.095 7.985 693.425 ;
        RECT 6.735 540.775 7.065 541.105 ;
        RECT 6.750 481.250 7.050 540.775 ;
        RECT 7.655 535.650 7.985 535.665 ;
        RECT 7.655 535.350 15.330 535.650 ;
        RECT 7.655 535.335 7.985 535.350 ;
        RECT 7.655 498.250 7.985 498.265 ;
        RECT 15.030 498.250 15.330 535.350 ;
        RECT 7.655 497.950 15.330 498.250 ;
        RECT 7.655 497.935 7.985 497.950 ;
        RECT 6.750 480.950 17.860 481.250 ;
        RECT 17.560 480.585 17.860 480.950 ;
        RECT 17.545 480.255 17.875 480.585 ;
        RECT 7.655 229.335 7.985 229.665 ;
        RECT 7.670 219.450 7.970 229.335 ;
        RECT 7.670 219.150 19.010 219.450 ;
        RECT 18.710 201.785 19.010 219.150 ;
        RECT 18.695 201.455 19.025 201.785 ;
        RECT 2805.390 165.490 2805.690 970.550 ;
        RECT 8.150 164.310 9.330 165.490 ;
        RECT 2804.950 164.310 2806.130 165.490 ;
        RECT 2808.150 165.050 2808.450 3402.215 ;
        RECT 2808.150 164.750 2809.370 165.050 ;
        RECT 7.655 151.450 7.985 151.465 ;
        RECT 8.590 151.450 8.890 164.310 ;
        RECT 7.655 151.150 8.890 151.450 ;
        RECT 7.655 151.135 7.985 151.150 ;
        RECT 2809.070 148.490 2809.370 164.750 ;
        RECT 8.150 147.310 9.330 148.490 ;
        RECT 2808.630 147.310 2809.810 148.490 ;
        RECT 7.655 135.130 7.985 135.145 ;
        RECT 8.590 135.130 8.890 147.310 ;
        RECT 7.655 134.830 8.890 135.130 ;
        RECT 7.655 134.815 7.985 134.830 ;
        RECT 411.535 0.855 411.865 1.185 ;
        RECT 406.935 0.490 407.265 0.505 ;
        RECT 411.550 0.490 411.850 0.855 ;
        RECT 406.935 0.190 411.850 0.490 ;
        RECT 406.935 0.175 407.265 0.190 ;
      LAYER met5 ;
        RECT 7.940 164.100 2806.340 165.700 ;
        RECT 7.940 147.100 2810.020 148.700 ;
    END
  END io_in[26]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 7.045 1905.785 7.215 1935.535 ;
        RECT 9.345 1764.685 9.515 1766.215 ;
        RECT 7.505 1659.285 7.675 1680.195 ;
        RECT 9.345 1680.025 9.515 1704.335 ;
        RECT 8.885 1560.005 9.055 1659.455 ;
        RECT 7.505 1472.965 7.675 1522.095 ;
        RECT 4.285 997.305 4.455 1108.655 ;
      LAYER mcon ;
        RECT 7.045 1935.365 7.215 1935.535 ;
        RECT 9.345 1766.045 9.515 1766.215 ;
        RECT 9.345 1704.165 9.515 1704.335 ;
        RECT 7.505 1680.025 7.675 1680.195 ;
        RECT 8.885 1659.285 9.055 1659.455 ;
        RECT 7.505 1521.925 7.675 1522.095 ;
        RECT 4.285 1108.485 4.455 1108.655 ;
      LAYER met1 ;
        RECT 6.970 1935.520 7.290 1935.580 ;
        RECT 6.775 1935.380 7.290 1935.520 ;
        RECT 6.970 1935.320 7.290 1935.380 ;
        RECT 6.985 1905.940 7.275 1905.985 ;
        RECT 9.730 1905.940 10.050 1906.000 ;
        RECT 6.985 1905.800 10.050 1905.940 ;
        RECT 6.985 1905.755 7.275 1905.800 ;
        RECT 9.730 1905.740 10.050 1905.800 ;
        RECT 9.285 1766.200 9.575 1766.245 ;
        RECT 9.730 1766.200 10.050 1766.260 ;
        RECT 9.285 1766.060 10.050 1766.200 ;
        RECT 9.285 1766.015 9.575 1766.060 ;
        RECT 9.730 1766.000 10.050 1766.060 ;
        RECT 9.285 1764.840 9.575 1764.885 ;
        RECT 9.730 1764.840 10.050 1764.900 ;
        RECT 9.285 1764.700 10.050 1764.840 ;
        RECT 9.285 1764.655 9.575 1764.700 ;
        RECT 9.730 1764.640 10.050 1764.700 ;
        RECT 9.285 1704.320 9.575 1704.365 ;
        RECT 9.730 1704.320 10.050 1704.380 ;
        RECT 9.285 1704.180 10.050 1704.320 ;
        RECT 9.285 1704.135 9.575 1704.180 ;
        RECT 9.730 1704.120 10.050 1704.180 ;
        RECT 7.445 1680.180 7.735 1680.225 ;
        RECT 9.285 1680.180 9.575 1680.225 ;
        RECT 7.445 1680.040 9.575 1680.180 ;
        RECT 7.445 1679.995 7.735 1680.040 ;
        RECT 9.285 1679.995 9.575 1680.040 ;
        RECT 7.445 1659.440 7.735 1659.485 ;
        RECT 8.825 1659.440 9.115 1659.485 ;
        RECT 7.445 1659.300 9.115 1659.440 ;
        RECT 7.445 1659.255 7.735 1659.300 ;
        RECT 8.825 1659.255 9.115 1659.300 ;
        RECT 8.825 1560.160 9.115 1560.205 ;
        RECT 9.730 1560.160 10.050 1560.220 ;
        RECT 8.825 1560.020 10.050 1560.160 ;
        RECT 8.825 1559.975 9.115 1560.020 ;
        RECT 9.730 1559.960 10.050 1560.020 ;
        RECT 7.445 1522.080 7.735 1522.125 ;
        RECT 9.730 1522.080 10.050 1522.140 ;
        RECT 7.445 1521.940 10.050 1522.080 ;
        RECT 7.445 1521.895 7.735 1521.940 ;
        RECT 9.730 1521.880 10.050 1521.940 ;
        RECT 2.370 1473.120 2.690 1473.180 ;
        RECT 7.445 1473.120 7.735 1473.165 ;
        RECT 2.370 1472.980 7.735 1473.120 ;
        RECT 2.370 1472.920 2.690 1472.980 ;
        RECT 7.445 1472.935 7.735 1472.980 ;
        RECT 2.370 1208.260 2.690 1208.320 ;
        RECT 9.730 1208.260 10.050 1208.320 ;
        RECT 2.370 1208.120 10.050 1208.260 ;
        RECT 2.370 1208.060 2.690 1208.120 ;
        RECT 9.730 1208.060 10.050 1208.120 ;
        RECT 9.730 1192.280 10.050 1192.340 ;
        RECT 7.060 1192.140 10.050 1192.280 ;
        RECT 7.060 1191.260 7.200 1192.140 ;
        RECT 9.730 1192.080 10.050 1192.140 ;
        RECT 7.060 1191.120 9.960 1191.260 ;
        RECT 9.820 1190.980 9.960 1191.120 ;
        RECT 9.730 1190.720 10.050 1190.980 ;
        RECT 4.225 1108.640 4.515 1108.685 ;
        RECT 9.730 1108.640 10.050 1108.700 ;
        RECT 4.225 1108.500 10.050 1108.640 ;
        RECT 4.225 1108.455 4.515 1108.500 ;
        RECT 9.730 1108.440 10.050 1108.500 ;
        RECT 4.210 997.460 4.530 997.520 ;
        RECT 4.015 997.320 4.530 997.460 ;
        RECT 4.210 997.260 4.530 997.320 ;
        RECT 3.290 709.480 3.610 709.540 ;
        RECT 4.210 709.480 4.530 709.540 ;
        RECT 3.290 709.340 4.530 709.480 ;
        RECT 3.290 709.280 3.610 709.340 ;
        RECT 4.210 709.280 4.530 709.340 ;
        RECT 3.750 623.120 4.070 623.180 ;
        RECT 6.970 623.120 7.290 623.180 ;
        RECT 3.750 622.980 7.290 623.120 ;
        RECT 3.750 622.920 4.070 622.980 ;
        RECT 6.970 622.920 7.290 622.980 ;
      LAYER via ;
        RECT 7.000 1935.320 7.260 1935.580 ;
        RECT 9.760 1905.740 10.020 1906.000 ;
        RECT 9.760 1766.000 10.020 1766.260 ;
        RECT 9.760 1764.640 10.020 1764.900 ;
        RECT 9.760 1704.120 10.020 1704.380 ;
        RECT 9.760 1559.960 10.020 1560.220 ;
        RECT 9.760 1521.880 10.020 1522.140 ;
        RECT 2.400 1472.920 2.660 1473.180 ;
        RECT 2.400 1208.060 2.660 1208.320 ;
        RECT 9.760 1208.060 10.020 1208.320 ;
        RECT 9.760 1192.080 10.020 1192.340 ;
        RECT 9.760 1190.720 10.020 1190.980 ;
        RECT 9.760 1108.440 10.020 1108.700 ;
        RECT 4.240 997.260 4.500 997.520 ;
        RECT 3.320 709.280 3.580 709.540 ;
        RECT 4.240 709.280 4.500 709.540 ;
        RECT 3.780 622.920 4.040 623.180 ;
        RECT 7.000 622.920 7.260 623.180 ;
      LAYER met2 ;
        RECT 6.990 1974.875 7.270 1975.245 ;
        RECT 7.060 1935.610 7.200 1974.875 ;
        RECT 7.000 1935.290 7.260 1935.610 ;
        RECT 9.760 1905.770 10.020 1906.030 ;
        RECT 9.760 1905.710 12.720 1905.770 ;
        RECT 9.820 1905.630 12.720 1905.710 ;
        RECT 12.580 1847.970 12.720 1905.630 ;
        RECT 10.280 1847.830 12.720 1847.970 ;
        RECT 10.280 1810.570 10.420 1847.830 ;
        RECT 9.820 1810.430 10.420 1810.570 ;
        RECT 9.820 1766.290 9.960 1810.430 ;
        RECT 9.760 1765.970 10.020 1766.290 ;
        RECT 9.760 1764.610 10.020 1764.930 ;
        RECT 9.820 1756.850 9.960 1764.610 ;
        RECT 9.820 1756.710 10.420 1756.850 ;
        RECT 10.280 1704.490 10.420 1756.710 ;
        RECT 9.820 1704.410 10.420 1704.490 ;
        RECT 9.760 1704.350 10.420 1704.410 ;
        RECT 9.760 1704.090 10.020 1704.350 ;
        RECT 9.820 1560.250 12.260 1560.330 ;
        RECT 9.760 1560.190 12.260 1560.250 ;
        RECT 9.760 1559.930 10.020 1560.190 ;
        RECT 12.120 1522.250 12.260 1560.190 ;
        RECT 9.820 1522.170 12.260 1522.250 ;
        RECT 9.760 1522.110 12.260 1522.170 ;
        RECT 9.760 1521.850 10.020 1522.110 ;
        RECT 2.400 1472.890 2.660 1473.210 ;
        RECT 2.460 1208.350 2.600 1472.890 ;
        RECT 2.400 1208.030 2.660 1208.350 ;
        RECT 9.760 1208.260 10.020 1208.350 ;
        RECT 9.760 1208.120 10.420 1208.260 ;
        RECT 9.760 1208.030 10.020 1208.120 ;
        RECT 9.760 1192.280 10.020 1192.370 ;
        RECT 10.280 1192.280 10.420 1208.120 ;
        RECT 9.760 1192.140 10.420 1192.280 ;
        RECT 9.760 1192.050 10.020 1192.140 ;
        RECT 9.760 1190.690 10.020 1191.010 ;
        RECT 9.820 1108.730 9.960 1190.690 ;
        RECT 9.760 1108.410 10.020 1108.730 ;
        RECT 4.240 997.230 4.500 997.550 ;
        RECT 4.300 709.570 4.440 997.230 ;
        RECT 3.320 709.250 3.580 709.570 ;
        RECT 4.240 709.250 4.500 709.570 ;
        RECT 3.380 693.330 3.520 709.250 ;
        RECT 3.380 693.190 3.980 693.330 ;
        RECT 3.840 623.210 3.980 693.190 ;
        RECT 3.780 622.890 4.040 623.210 ;
        RECT 7.000 622.890 7.260 623.210 ;
        RECT 7.060 177.325 7.200 622.890 ;
        RECT 6.990 176.955 7.270 177.325 ;
      LAYER via2 ;
        RECT 6.990 1974.920 7.270 1975.200 ;
        RECT 6.990 177.000 7.270 177.280 ;
      LAYER met3 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 6.965 1975.210 7.295 1975.225 ;
        RECT -4.800 1974.910 7.295 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 6.965 1974.895 7.295 1974.910 ;
        RECT 6.965 177.290 7.295 177.305 ;
        RECT 6.750 176.975 7.295 177.290 ;
        RECT 6.750 174.960 7.050 176.975 ;
        RECT 5.000 174.360 9.000 174.960 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2873.690 552.400 2874.010 552.460 ;
        RECT 2900.830 552.400 2901.150 552.460 ;
        RECT 2873.690 552.260 2901.150 552.400 ;
        RECT 2873.690 552.200 2874.010 552.260 ;
        RECT 2900.830 552.200 2901.150 552.260 ;
      LAYER via ;
        RECT 2873.720 552.200 2873.980 552.460 ;
        RECT 2900.860 552.200 2901.120 552.460 ;
      LAYER met2 ;
        RECT 2900.850 557.075 2901.130 557.445 ;
        RECT 2900.920 552.490 2901.060 557.075 ;
        RECT 2873.720 552.170 2873.980 552.490 ;
        RECT 2900.860 552.170 2901.120 552.490 ;
        RECT 2873.780 345.285 2873.920 552.170 ;
        RECT 2873.710 344.915 2873.990 345.285 ;
      LAYER via2 ;
        RECT 2900.850 557.120 2901.130 557.400 ;
        RECT 2873.710 344.960 2873.990 345.240 ;
      LAYER met3 ;
        RECT 2900.825 557.410 2901.155 557.425 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2900.825 557.110 2924.800 557.410 ;
        RECT 2900.825 557.095 2901.155 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
        RECT 2851.000 345.250 2855.000 345.640 ;
        RECT 2873.685 345.250 2874.015 345.265 ;
        RECT 2851.000 345.040 2874.015 345.250 ;
        RECT 2854.300 344.950 2874.015 345.040 ;
        RECT 2873.685 344.935 2874.015 344.950 ;
    END
  END io_in[2]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 7.965 743.665 8.135 816.595 ;
      LAYER mcon ;
        RECT 7.965 816.425 8.135 816.595 ;
      LAYER met1 ;
        RECT 3.750 1108.300 4.070 1108.360 ;
        RECT 6.970 1108.300 7.290 1108.360 ;
        RECT 3.750 1108.160 7.290 1108.300 ;
        RECT 3.750 1108.100 4.070 1108.160 ;
        RECT 6.970 1108.100 7.290 1108.160 ;
        RECT 3.750 816.580 4.070 816.640 ;
        RECT 7.905 816.580 8.195 816.625 ;
        RECT 3.750 816.440 8.195 816.580 ;
        RECT 3.750 816.380 4.070 816.440 ;
        RECT 7.905 816.395 8.195 816.440 ;
        RECT 2.370 743.820 2.690 743.880 ;
        RECT 7.905 743.820 8.195 743.865 ;
        RECT 2.370 743.680 8.195 743.820 ;
        RECT 2.370 743.620 2.690 743.680 ;
        RECT 7.905 743.635 8.195 743.680 ;
      LAYER via ;
        RECT 3.780 1108.100 4.040 1108.360 ;
        RECT 7.000 1108.100 7.260 1108.360 ;
        RECT 3.780 816.380 4.040 816.640 ;
        RECT 2.400 743.620 2.660 743.880 ;
      LAYER met2 ;
        RECT 6.990 1256.115 7.270 1256.485 ;
        RECT 7.060 1108.390 7.200 1256.115 ;
        RECT 3.780 1108.070 4.040 1108.390 ;
        RECT 7.000 1108.070 7.260 1108.390 ;
        RECT 3.840 816.670 3.980 1108.070 ;
        RECT 3.780 816.350 4.040 816.670 ;
        RECT 2.400 743.590 2.660 743.910 ;
        RECT 2.460 517.325 2.600 743.590 ;
        RECT 2.390 516.955 2.670 517.325 ;
      LAYER via2 ;
        RECT 6.990 1256.160 7.270 1256.440 ;
        RECT 2.390 517.000 2.670 517.280 ;
      LAYER met3 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 6.965 1256.450 7.295 1256.465 ;
        RECT -4.800 1256.150 7.295 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 6.965 1256.135 7.295 1256.150 ;
        RECT 2.365 517.290 2.695 517.305 ;
        RECT 2.365 516.990 5.210 517.290 ;
        RECT 2.365 516.975 2.695 516.990 ;
        RECT 4.910 514.960 5.210 516.990 ;
        RECT 4.910 514.420 9.000 514.960 ;
        RECT 5.000 514.360 9.000 514.420 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 6.585 882.385 6.755 946.135 ;
        RECT 5.205 795.685 5.375 836.995 ;
        RECT 4.745 750.465 4.915 770.355 ;
        RECT 7.505 707.285 7.675 750.635 ;
        RECT 8.885 691.305 9.055 694.195 ;
      LAYER mcon ;
        RECT 6.585 945.965 6.755 946.135 ;
        RECT 5.205 836.825 5.375 836.995 ;
        RECT 4.745 770.185 4.915 770.355 ;
        RECT 7.505 750.465 7.675 750.635 ;
        RECT 8.885 694.025 9.055 694.195 ;
      LAYER met1 ;
        RECT 2.830 1025.340 3.150 1025.400 ;
        RECT 6.050 1025.340 6.370 1025.400 ;
        RECT 2.830 1025.200 6.370 1025.340 ;
        RECT 2.830 1025.140 3.150 1025.200 ;
        RECT 6.050 1025.140 6.370 1025.200 ;
        RECT 6.050 974.680 6.370 974.740 ;
        RECT 9.730 974.680 10.050 974.740 ;
        RECT 6.050 974.540 10.050 974.680 ;
        RECT 6.050 974.480 6.370 974.540 ;
        RECT 9.730 974.480 10.050 974.540 ;
        RECT 6.525 946.120 6.815 946.165 ;
        RECT 9.730 946.120 10.050 946.180 ;
        RECT 6.525 945.980 10.050 946.120 ;
        RECT 6.525 945.935 6.815 945.980 ;
        RECT 9.730 945.920 10.050 945.980 ;
        RECT 6.525 882.540 6.815 882.585 ;
        RECT 9.730 882.540 10.050 882.600 ;
        RECT 6.525 882.400 10.050 882.540 ;
        RECT 6.525 882.355 6.815 882.400 ;
        RECT 9.730 882.340 10.050 882.400 ;
        RECT 5.145 836.980 5.435 837.025 ;
        RECT 9.730 836.980 10.050 837.040 ;
        RECT 5.145 836.840 10.050 836.980 ;
        RECT 5.145 836.795 5.435 836.840 ;
        RECT 9.730 836.780 10.050 836.840 ;
        RECT 5.145 795.840 5.435 795.885 ;
        RECT 9.730 795.840 10.050 795.900 ;
        RECT 5.145 795.700 10.050 795.840 ;
        RECT 5.145 795.655 5.435 795.700 ;
        RECT 9.730 795.640 10.050 795.700 ;
        RECT 4.685 770.340 4.975 770.385 ;
        RECT 9.730 770.340 10.050 770.400 ;
        RECT 4.685 770.200 10.050 770.340 ;
        RECT 4.685 770.155 4.975 770.200 ;
        RECT 9.730 770.140 10.050 770.200 ;
        RECT 4.685 750.620 4.975 750.665 ;
        RECT 7.445 750.620 7.735 750.665 ;
        RECT 4.685 750.480 7.735 750.620 ;
        RECT 4.685 750.435 4.975 750.480 ;
        RECT 7.445 750.435 7.735 750.480 ;
        RECT 7.430 707.440 7.750 707.500 ;
        RECT 7.235 707.300 7.750 707.440 ;
        RECT 7.430 707.240 7.750 707.300 ;
        RECT 7.430 694.180 7.750 694.240 ;
        RECT 8.825 694.180 9.115 694.225 ;
        RECT 7.430 694.040 9.115 694.180 ;
        RECT 7.430 693.980 7.750 694.040 ;
        RECT 8.825 693.995 9.115 694.040 ;
        RECT 8.825 691.460 9.115 691.505 ;
        RECT 9.730 691.460 10.050 691.520 ;
        RECT 8.825 691.320 10.050 691.460 ;
        RECT 8.825 691.275 9.115 691.320 ;
        RECT 9.730 691.260 10.050 691.320 ;
      LAYER via ;
        RECT 2.860 1025.140 3.120 1025.400 ;
        RECT 6.080 1025.140 6.340 1025.400 ;
        RECT 6.080 974.480 6.340 974.740 ;
        RECT 9.760 974.480 10.020 974.740 ;
        RECT 9.760 945.920 10.020 946.180 ;
        RECT 9.760 882.340 10.020 882.600 ;
        RECT 9.760 836.780 10.020 837.040 ;
        RECT 9.760 795.640 10.020 795.900 ;
        RECT 9.760 770.140 10.020 770.400 ;
        RECT 7.460 707.240 7.720 707.500 ;
        RECT 7.460 693.980 7.720 694.240 ;
        RECT 9.760 691.260 10.020 691.520 ;
      LAYER met2 ;
        RECT 2.850 1040.555 3.130 1040.925 ;
        RECT 2.920 1025.430 3.060 1040.555 ;
        RECT 2.860 1025.110 3.120 1025.430 ;
        RECT 6.080 1025.110 6.340 1025.430 ;
        RECT 6.140 974.770 6.280 1025.110 ;
        RECT 6.080 974.450 6.340 974.770 ;
        RECT 9.760 974.450 10.020 974.770 ;
        RECT 9.820 974.170 9.960 974.450 ;
        RECT 9.820 974.030 11.800 974.170 ;
        RECT 11.660 947.650 11.800 974.030 ;
        RECT 10.740 947.510 11.800 947.650 ;
        RECT 9.760 946.120 10.020 946.210 ;
        RECT 10.740 946.120 10.880 947.510 ;
        RECT 9.760 945.980 10.880 946.120 ;
        RECT 9.760 945.890 10.020 945.980 ;
        RECT 9.760 882.540 10.020 882.630 ;
        RECT 9.760 882.400 11.340 882.540 ;
        RECT 9.760 882.310 10.020 882.400 ;
        RECT 11.200 881.860 11.340 882.400 ;
        RECT 11.200 881.720 11.800 881.860 ;
        RECT 11.660 837.490 11.800 881.720 ;
        RECT 9.820 837.350 11.800 837.490 ;
        RECT 9.820 837.070 9.960 837.350 ;
        RECT 9.760 836.750 10.020 837.070 ;
        RECT 9.760 795.610 10.020 795.930 ;
        RECT 9.820 770.430 9.960 795.610 ;
        RECT 9.760 770.110 10.020 770.430 ;
        RECT 7.460 707.210 7.720 707.530 ;
        RECT 7.520 694.270 7.660 707.210 ;
        RECT 7.460 693.950 7.720 694.270 ;
        RECT 9.760 691.290 10.020 691.550 ;
        RECT 9.760 691.230 10.420 691.290 ;
        RECT 9.820 691.150 10.420 691.230 ;
        RECT 10.280 666.810 10.420 691.150 ;
        RECT 8.900 666.670 10.420 666.810 ;
        RECT 8.900 660.010 9.040 666.670 ;
        RECT 7.980 659.870 9.040 660.010 ;
        RECT 7.980 632.245 8.120 659.870 ;
        RECT 7.910 631.875 8.190 632.245 ;
      LAYER via2 ;
        RECT 2.850 1040.600 3.130 1040.880 ;
        RECT 7.910 631.920 8.190 632.200 ;
      LAYER met3 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 2.825 1040.890 3.155 1040.905 ;
        RECT -4.800 1040.590 3.155 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
        RECT 2.825 1040.575 3.155 1040.590 ;
        RECT 7.885 632.210 8.215 632.225 ;
        RECT 7.670 631.895 8.215 632.210 ;
        RECT 7.670 628.520 7.970 631.895 ;
        RECT 5.000 627.920 9.000 628.520 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 6.970 781.220 7.290 781.280 ;
        RECT 7.890 781.220 8.210 781.280 ;
        RECT 6.970 781.080 8.210 781.220 ;
        RECT 6.970 781.020 7.290 781.080 ;
        RECT 7.890 781.020 8.210 781.080 ;
      LAYER via ;
        RECT 7.000 781.020 7.260 781.280 ;
        RECT 7.920 781.020 8.180 781.280 ;
      LAYER met2 ;
        RECT 6.990 824.995 7.270 825.365 ;
        RECT 7.060 781.310 7.200 824.995 ;
        RECT 7.000 780.990 7.260 781.310 ;
        RECT 7.920 780.990 8.180 781.310 ;
        RECT 7.980 743.765 8.120 780.990 ;
        RECT 7.910 743.395 8.190 743.765 ;
      LAYER via2 ;
        RECT 6.990 825.040 7.270 825.320 ;
        RECT 7.910 743.440 8.190 743.720 ;
      LAYER met3 ;
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 6.965 825.330 7.295 825.345 ;
        RECT -4.800 825.030 7.295 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
        RECT 6.965 825.015 7.295 825.030 ;
        RECT 7.885 743.730 8.215 743.745 ;
        RECT 7.670 743.415 8.215 743.730 ;
        RECT 7.670 742.080 7.970 743.415 ;
        RECT 5.000 741.480 9.000 742.080 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2.370 819.640 2.690 819.700 ;
        RECT 7.430 819.640 7.750 819.700 ;
        RECT 2.370 819.500 7.750 819.640 ;
        RECT 2.370 819.440 2.690 819.500 ;
        RECT 7.430 819.440 7.750 819.500 ;
        RECT 2.370 777.140 2.690 777.200 ;
        RECT 6.510 777.140 6.830 777.200 ;
        RECT 2.370 777.000 6.830 777.140 ;
        RECT 2.370 776.940 2.690 777.000 ;
        RECT 6.510 776.940 6.830 777.000 ;
      LAYER via ;
        RECT 2.400 819.440 2.660 819.700 ;
        RECT 7.460 819.440 7.720 819.700 ;
        RECT 2.400 776.940 2.660 777.200 ;
        RECT 6.540 776.940 6.800 777.200 ;
      LAYER met2 ;
        RECT 7.450 851.515 7.730 851.885 ;
        RECT 7.520 819.730 7.660 851.515 ;
        RECT 2.400 819.410 2.660 819.730 ;
        RECT 7.460 819.410 7.720 819.730 ;
        RECT 2.460 777.230 2.600 819.410 ;
        RECT 2.400 776.910 2.660 777.230 ;
        RECT 6.540 776.910 6.800 777.230 ;
        RECT 6.600 735.490 6.740 776.910 ;
        RECT 6.600 735.350 7.200 735.490 ;
        RECT 7.060 674.290 7.200 735.350 ;
        RECT 6.600 674.150 7.200 674.290 ;
        RECT 6.600 610.485 6.740 674.150 ;
        RECT 6.530 610.115 6.810 610.485 ;
      LAYER via2 ;
        RECT 7.450 851.560 7.730 851.840 ;
        RECT 6.530 610.160 6.810 610.440 ;
      LAYER met3 ;
        RECT 5.000 854.360 9.000 854.960 ;
        RECT 7.670 851.865 7.970 854.360 ;
        RECT 7.425 851.550 7.970 851.865 ;
        RECT 7.425 851.535 7.755 851.550 ;
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 6.505 610.450 6.835 610.465 ;
        RECT -4.800 610.150 6.835 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 6.505 610.135 6.835 610.150 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 9.345 734.655 9.515 795.515 ;
        RECT 9.345 734.485 9.975 734.655 ;
        RECT 9.805 655.775 9.975 734.485 ;
        RECT 9.345 655.605 9.975 655.775 ;
        RECT 9.345 624.665 9.515 655.605 ;
        RECT 9.345 466.225 9.515 473.875 ;
        RECT 8.425 404.685 8.595 431.715 ;
      LAYER mcon ;
        RECT 9.345 795.345 9.515 795.515 ;
        RECT 9.345 473.705 9.515 473.875 ;
        RECT 8.425 431.545 8.595 431.715 ;
      LAYER met1 ;
        RECT 3.750 808.080 4.070 808.140 ;
        RECT 6.510 808.080 6.830 808.140 ;
        RECT 3.750 807.940 6.830 808.080 ;
        RECT 3.750 807.880 4.070 807.940 ;
        RECT 6.510 807.880 6.830 807.940 ;
        RECT 3.750 795.500 4.070 795.560 ;
        RECT 9.285 795.500 9.575 795.545 ;
        RECT 3.750 795.360 9.575 795.500 ;
        RECT 3.750 795.300 4.070 795.360 ;
        RECT 9.285 795.315 9.575 795.360 ;
        RECT 9.270 624.820 9.590 624.880 ;
        RECT 9.075 624.680 9.590 624.820 ;
        RECT 9.270 624.620 9.590 624.680 ;
        RECT 9.270 473.860 9.590 473.920 ;
        RECT 9.075 473.720 9.590 473.860 ;
        RECT 9.270 473.660 9.590 473.720 ;
        RECT 9.270 466.380 9.590 466.440 ;
        RECT 9.075 466.240 9.590 466.380 ;
        RECT 9.270 466.180 9.590 466.240 ;
        RECT 8.365 431.700 8.655 431.745 ;
        RECT 9.270 431.700 9.590 431.760 ;
        RECT 8.365 431.560 9.590 431.700 ;
        RECT 8.365 431.515 8.655 431.560 ;
        RECT 9.270 431.500 9.590 431.560 ;
        RECT 2.830 404.840 3.150 404.900 ;
        RECT 8.365 404.840 8.655 404.885 ;
        RECT 2.830 404.700 8.655 404.840 ;
        RECT 2.830 404.640 3.150 404.700 ;
        RECT 8.365 404.655 8.655 404.700 ;
      LAYER via ;
        RECT 3.780 807.880 4.040 808.140 ;
        RECT 6.540 807.880 6.800 808.140 ;
        RECT 3.780 795.300 4.040 795.560 ;
        RECT 9.300 624.620 9.560 624.880 ;
        RECT 9.300 473.660 9.560 473.920 ;
        RECT 9.300 466.180 9.560 466.440 ;
        RECT 9.300 431.500 9.560 431.760 ;
        RECT 2.860 404.640 3.120 404.900 ;
      LAYER met2 ;
        RECT 6.530 965.075 6.810 965.445 ;
        RECT 6.600 808.170 6.740 965.075 ;
        RECT 3.780 807.850 4.040 808.170 ;
        RECT 6.540 807.850 6.800 808.170 ;
        RECT 3.840 795.590 3.980 807.850 ;
        RECT 3.780 795.270 4.040 795.590 ;
        RECT 9.300 624.590 9.560 624.910 ;
        RECT 9.360 473.950 9.500 624.590 ;
        RECT 9.300 473.630 9.560 473.950 ;
        RECT 9.300 466.150 9.560 466.470 ;
        RECT 9.360 431.790 9.500 466.150 ;
        RECT 9.300 431.470 9.560 431.790 ;
        RECT 2.860 404.610 3.120 404.930 ;
        RECT 2.920 394.925 3.060 404.610 ;
        RECT 2.850 394.555 3.130 394.925 ;
      LAYER via2 ;
        RECT 6.530 965.120 6.810 965.400 ;
        RECT 2.850 394.600 3.130 394.880 ;
      LAYER met3 ;
        RECT 5.000 967.920 9.000 968.520 ;
        RECT 6.750 965.425 7.050 967.920 ;
        RECT 6.505 965.110 7.050 965.425 ;
        RECT 6.505 965.095 6.835 965.110 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 2.825 394.890 3.155 394.905 ;
        RECT -4.800 394.590 3.155 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 2.825 394.575 3.155 394.590 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 0.090 1078.635 0.370 1079.005 ;
        RECT 0.160 180.725 0.300 1078.635 ;
        RECT 0.090 180.355 0.370 180.725 ;
      LAYER via2 ;
        RECT 0.090 1078.680 0.370 1078.960 ;
        RECT 0.090 180.400 0.370 180.680 ;
      LAYER met3 ;
        RECT 5.000 1081.480 9.000 1082.080 ;
        RECT 0.065 1078.970 0.395 1078.985 ;
        RECT 5.830 1078.970 6.130 1081.480 ;
        RECT 0.065 1078.670 6.130 1078.970 ;
        RECT 0.065 1078.655 0.395 1078.670 ;
        RECT 0.065 180.690 0.395 180.705 ;
        RECT 0.065 180.390 3.370 180.690 ;
        RECT 0.065 180.375 0.395 180.390 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 3.070 179.330 3.370 180.390 ;
        RECT -4.800 179.030 3.370 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2874.610 787.000 2874.930 787.060 ;
        RECT 2900.830 787.000 2901.150 787.060 ;
        RECT 2874.610 786.860 2901.150 787.000 ;
        RECT 2874.610 786.800 2874.930 786.860 ;
        RECT 2900.830 786.800 2901.150 786.860 ;
        RECT 2863.570 482.700 2863.890 482.760 ;
        RECT 2874.610 482.700 2874.930 482.760 ;
        RECT 2863.570 482.560 2874.930 482.700 ;
        RECT 2863.570 482.500 2863.890 482.560 ;
        RECT 2874.610 482.500 2874.930 482.560 ;
      LAYER via ;
        RECT 2874.640 786.800 2874.900 787.060 ;
        RECT 2900.860 786.800 2901.120 787.060 ;
        RECT 2863.600 482.500 2863.860 482.760 ;
        RECT 2874.640 482.500 2874.900 482.760 ;
      LAYER met2 ;
        RECT 2900.850 791.675 2901.130 792.045 ;
        RECT 2900.920 787.090 2901.060 791.675 ;
        RECT 2874.640 786.770 2874.900 787.090 ;
        RECT 2900.860 786.770 2901.120 787.090 ;
        RECT 2874.700 482.790 2874.840 786.770 ;
        RECT 2863.600 482.470 2863.860 482.790 ;
        RECT 2874.640 482.470 2874.900 482.790 ;
        RECT 2863.660 481.285 2863.800 482.470 ;
        RECT 2863.590 480.915 2863.870 481.285 ;
      LAYER via2 ;
        RECT 2900.850 791.720 2901.130 792.000 ;
        RECT 2863.590 480.960 2863.870 481.240 ;
      LAYER met3 ;
        RECT 2900.825 792.010 2901.155 792.025 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2900.825 791.710 2924.800 792.010 ;
        RECT 2900.825 791.695 2901.155 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
        RECT 2851.000 481.250 2855.000 481.640 ;
        RECT 2863.565 481.250 2863.895 481.265 ;
        RECT 2851.000 481.040 2863.895 481.250 ;
        RECT 2854.300 480.950 2863.895 481.040 ;
        RECT 2863.565 480.935 2863.895 480.950 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2874.150 1021.600 2874.470 1021.660 ;
        RECT 2900.830 1021.600 2901.150 1021.660 ;
        RECT 2874.150 1021.460 2901.150 1021.600 ;
        RECT 2874.150 1021.400 2874.470 1021.460 ;
        RECT 2900.830 1021.400 2901.150 1021.460 ;
        RECT 2863.570 620.400 2863.890 620.460 ;
        RECT 2874.150 620.400 2874.470 620.460 ;
        RECT 2863.570 620.260 2874.470 620.400 ;
        RECT 2863.570 620.200 2863.890 620.260 ;
        RECT 2874.150 620.200 2874.470 620.260 ;
      LAYER via ;
        RECT 2874.180 1021.400 2874.440 1021.660 ;
        RECT 2900.860 1021.400 2901.120 1021.660 ;
        RECT 2863.600 620.200 2863.860 620.460 ;
        RECT 2874.180 620.200 2874.440 620.460 ;
      LAYER met2 ;
        RECT 2900.850 1026.275 2901.130 1026.645 ;
        RECT 2900.920 1021.690 2901.060 1026.275 ;
        RECT 2874.180 1021.370 2874.440 1021.690 ;
        RECT 2900.860 1021.370 2901.120 1021.690 ;
        RECT 2874.240 620.490 2874.380 1021.370 ;
        RECT 2863.600 620.170 2863.860 620.490 ;
        RECT 2874.180 620.170 2874.440 620.490 ;
        RECT 2863.660 617.285 2863.800 620.170 ;
        RECT 2863.590 616.915 2863.870 617.285 ;
      LAYER via2 ;
        RECT 2900.850 1026.320 2901.130 1026.600 ;
        RECT 2863.590 616.960 2863.870 617.240 ;
      LAYER met3 ;
        RECT 2900.825 1026.610 2901.155 1026.625 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2900.825 1026.310 2924.800 1026.610 ;
        RECT 2900.825 1026.295 2901.155 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
        RECT 2851.000 617.250 2855.000 617.640 ;
        RECT 2863.565 617.250 2863.895 617.265 ;
        RECT 2851.000 617.040 2863.895 617.250 ;
        RECT 2854.300 616.950 2863.895 617.040 ;
        RECT 2863.565 616.935 2863.895 616.950 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2873.690 1256.200 2874.010 1256.260 ;
        RECT 2900.830 1256.200 2901.150 1256.260 ;
        RECT 2873.690 1256.060 2901.150 1256.200 ;
        RECT 2873.690 1256.000 2874.010 1256.060 ;
        RECT 2900.830 1256.000 2901.150 1256.060 ;
      LAYER via ;
        RECT 2873.720 1256.000 2873.980 1256.260 ;
        RECT 2900.860 1256.000 2901.120 1256.260 ;
      LAYER met2 ;
        RECT 2900.850 1260.875 2901.130 1261.245 ;
        RECT 2900.920 1256.290 2901.060 1260.875 ;
        RECT 2873.720 1255.970 2873.980 1256.290 ;
        RECT 2900.860 1255.970 2901.120 1256.290 ;
        RECT 2873.780 753.285 2873.920 1255.970 ;
        RECT 2873.710 752.915 2873.990 753.285 ;
      LAYER via2 ;
        RECT 2900.850 1260.920 2901.130 1261.200 ;
        RECT 2873.710 752.960 2873.990 753.240 ;
      LAYER met3 ;
        RECT 2900.825 1261.210 2901.155 1261.225 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2900.825 1260.910 2924.800 1261.210 ;
        RECT 2900.825 1260.895 2901.155 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
        RECT 2851.000 753.250 2855.000 753.640 ;
        RECT 2873.685 753.250 2874.015 753.265 ;
        RECT 2851.000 753.040 2874.015 753.250 ;
        RECT 2854.300 752.950 2874.015 753.040 ;
        RECT 2873.685 752.935 2874.015 752.950 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2875.070 1490.800 2875.390 1490.860 ;
        RECT 2900.830 1490.800 2901.150 1490.860 ;
        RECT 2875.070 1490.660 2901.150 1490.800 ;
        RECT 2875.070 1490.600 2875.390 1490.660 ;
        RECT 2900.830 1490.600 2901.150 1490.660 ;
      LAYER via ;
        RECT 2875.100 1490.600 2875.360 1490.860 ;
        RECT 2900.860 1490.600 2901.120 1490.860 ;
      LAYER met2 ;
        RECT 2900.850 1495.475 2901.130 1495.845 ;
        RECT 2900.920 1490.890 2901.060 1495.475 ;
        RECT 2875.100 1490.570 2875.360 1490.890 ;
        RECT 2900.860 1490.570 2901.120 1490.890 ;
        RECT 2875.160 889.285 2875.300 1490.570 ;
        RECT 2875.090 888.915 2875.370 889.285 ;
      LAYER via2 ;
        RECT 2900.850 1495.520 2901.130 1495.800 ;
        RECT 2875.090 888.960 2875.370 889.240 ;
      LAYER met3 ;
        RECT 2900.825 1495.810 2901.155 1495.825 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2900.825 1495.510 2924.800 1495.810 ;
        RECT 2900.825 1495.495 2901.155 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
        RECT 2851.000 889.250 2855.000 889.640 ;
        RECT 2875.065 889.250 2875.395 889.265 ;
        RECT 2851.000 889.040 2875.395 889.250 ;
        RECT 2854.300 888.950 2875.395 889.040 ;
        RECT 2875.065 888.935 2875.395 888.950 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2874.610 1725.400 2874.930 1725.460 ;
        RECT 2900.830 1725.400 2901.150 1725.460 ;
        RECT 2874.610 1725.260 2901.150 1725.400 ;
        RECT 2874.610 1725.200 2874.930 1725.260 ;
        RECT 2900.830 1725.200 2901.150 1725.260 ;
      LAYER via ;
        RECT 2874.640 1725.200 2874.900 1725.460 ;
        RECT 2900.860 1725.200 2901.120 1725.460 ;
      LAYER met2 ;
        RECT 2900.850 1730.075 2901.130 1730.445 ;
        RECT 2900.920 1725.490 2901.060 1730.075 ;
        RECT 2874.640 1725.170 2874.900 1725.490 ;
        RECT 2900.860 1725.170 2901.120 1725.490 ;
        RECT 2874.700 1025.285 2874.840 1725.170 ;
        RECT 2874.630 1024.915 2874.910 1025.285 ;
      LAYER via2 ;
        RECT 2900.850 1730.120 2901.130 1730.400 ;
        RECT 2874.630 1024.960 2874.910 1025.240 ;
      LAYER met3 ;
        RECT 2900.825 1730.410 2901.155 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2900.825 1730.110 2924.800 1730.410 ;
        RECT 2900.825 1730.095 2901.155 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
        RECT 2851.000 1025.250 2855.000 1025.640 ;
        RECT 2874.605 1025.250 2874.935 1025.265 ;
        RECT 2851.000 1025.040 2874.935 1025.250 ;
        RECT 2854.300 1024.950 2874.935 1025.040 ;
        RECT 2874.605 1024.935 2874.935 1024.950 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2874.150 1960.000 2874.470 1960.060 ;
        RECT 2900.830 1960.000 2901.150 1960.060 ;
        RECT 2874.150 1959.860 2901.150 1960.000 ;
        RECT 2874.150 1959.800 2874.470 1959.860 ;
        RECT 2900.830 1959.800 2901.150 1959.860 ;
      LAYER via ;
        RECT 2874.180 1959.800 2874.440 1960.060 ;
        RECT 2900.860 1959.800 2901.120 1960.060 ;
      LAYER met2 ;
        RECT 2900.850 1964.675 2901.130 1965.045 ;
        RECT 2900.920 1960.090 2901.060 1964.675 ;
        RECT 2874.180 1959.770 2874.440 1960.090 ;
        RECT 2900.860 1959.770 2901.120 1960.090 ;
        RECT 2874.240 1161.285 2874.380 1959.770 ;
        RECT 2874.170 1160.915 2874.450 1161.285 ;
      LAYER via2 ;
        RECT 2900.850 1964.720 2901.130 1965.000 ;
        RECT 2874.170 1160.960 2874.450 1161.240 ;
      LAYER met3 ;
        RECT 2900.825 1965.010 2901.155 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2900.825 1964.710 2924.800 1965.010 ;
        RECT 2900.825 1964.695 2901.155 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
        RECT 2851.000 1161.250 2855.000 1161.640 ;
        RECT 2874.145 1161.250 2874.475 1161.265 ;
        RECT 2851.000 1161.040 2874.475 1161.250 ;
        RECT 2854.300 1160.950 2874.475 1161.040 ;
        RECT 2874.145 1160.935 2874.475 1160.950 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2873.690 2194.600 2874.010 2194.660 ;
        RECT 2900.830 2194.600 2901.150 2194.660 ;
        RECT 2873.690 2194.460 2901.150 2194.600 ;
        RECT 2873.690 2194.400 2874.010 2194.460 ;
        RECT 2900.830 2194.400 2901.150 2194.460 ;
      LAYER via ;
        RECT 2873.720 2194.400 2873.980 2194.660 ;
        RECT 2900.860 2194.400 2901.120 2194.660 ;
      LAYER met2 ;
        RECT 2900.850 2199.275 2901.130 2199.645 ;
        RECT 2900.920 2194.690 2901.060 2199.275 ;
        RECT 2873.720 2194.370 2873.980 2194.690 ;
        RECT 2900.860 2194.370 2901.120 2194.690 ;
        RECT 2873.780 1297.285 2873.920 2194.370 ;
        RECT 2873.710 1296.915 2873.990 1297.285 ;
      LAYER via2 ;
        RECT 2900.850 2199.320 2901.130 2199.600 ;
        RECT 2873.710 1296.960 2873.990 1297.240 ;
      LAYER met3 ;
        RECT 2900.825 2199.610 2901.155 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2900.825 2199.310 2924.800 2199.610 ;
        RECT 2900.825 2199.295 2901.155 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
        RECT 2851.000 1297.250 2855.000 1297.640 ;
        RECT 2873.685 1297.250 2874.015 1297.265 ;
        RECT 2851.000 1297.040 2874.015 1297.250 ;
        RECT 2854.300 1296.950 2874.015 1297.040 ;
        RECT 2873.685 1296.935 2874.015 1296.950 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 204.420 2924.800 205.620 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2551.100 2924.800 2552.300 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2785.700 2924.800 2786.900 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3020.300 2924.800 3021.500 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3254.900 2924.800 3256.100 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3489.500 2924.800 3490.700 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 439.020 2924.800 440.220 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 3267.140 2.400 3268.340 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2979.500 2.400 2980.700 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2692.540 2.400 2693.740 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2404.900 2.400 2406.100 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2117.940 2.400 2119.140 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1830.300 2.400 1831.500 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 673.620 2924.800 674.820 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1543.340 2.400 1544.540 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1327.780 2.400 1328.980 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1112.220 2.400 1113.420 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 896.660 2.400 897.860 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 681.100 2.400 682.300 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 465.540 2.400 466.740 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 249.980 2.400 251.180 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 35.100 2.400 36.300 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 908.900 2924.800 910.100 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1143.500 2924.800 1144.700 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1378.100 2924.800 1379.300 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1612.700 2924.800 1613.900 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1847.300 2924.800 1848.500 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2081.900 2924.800 2083.100 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2316.500 2924.800 2317.700 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 145.940 2924.800 147.140 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2492.620 2924.800 2493.820 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2727.220 2924.800 2728.420 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2961.820 2924.800 2963.020 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3196.420 2924.800 3197.620 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3431.020 2924.800 3432.220 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 380.540 2924.800 381.740 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 3339.220 2.400 3340.420 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 3051.580 2.400 3052.780 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2764.620 2.400 2765.820 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2476.980 2.400 2478.180 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2189.340 2.400 2190.540 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1902.380 2.400 1903.580 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 615.140 2924.800 616.340 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1614.740 2.400 1615.940 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1399.860 2.400 1401.060 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1184.300 2.400 1185.500 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 968.740 2.400 969.940 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 753.180 2.400 754.380 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 537.620 2.400 538.820 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 322.060 2.400 323.260 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 106.500 2.400 107.700 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 849.740 2924.800 850.940 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1084.340 2924.800 1085.540 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1318.940 2924.800 1320.140 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1553.540 2924.800 1554.740 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1788.820 2924.800 1790.020 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2023.420 2924.800 2024.620 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2258.020 2924.800 2259.220 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 674.310 -4.800 674.870 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 38.915 3.130 39.285 ;
        RECT 2.920 2.400 3.060 38.915 ;
        RECT 2.710 -4.800 3.270 2.400 ;
      LAYER via2 ;
        RECT 2.850 38.960 3.130 39.240 ;
      LAYER met3 ;
        RECT 2.825 39.260 3.155 39.265 ;
        RECT 2.825 39.250 3.410 39.260 ;
        RECT 2.600 38.950 3.410 39.250 ;
        RECT 2.825 38.940 3.410 38.950 ;
        RECT 2.825 38.935 3.155 38.940 ;
      LAYER via3 ;
        RECT 3.060 38.940 3.380 39.260 ;
      LAYER met4 ;
        RECT 2.630 38.510 3.810 39.690 ;
        RECT 1128.710 31.710 1129.890 32.890 ;
      LAYER met5 ;
        RECT 69.580 41.700 108.900 43.300 ;
        RECT 69.580 39.900 71.180 41.700 ;
        RECT 2.420 38.300 71.180 39.900 ;
        RECT 107.300 39.900 108.900 41.700 ;
        RECT 192.170 41.700 304.860 43.300 ;
        RECT 192.170 39.900 193.770 41.700 ;
        RECT 107.300 38.300 193.770 39.900 ;
        RECT 303.260 39.900 304.860 41.700 ;
        RECT 398.940 41.700 421.700 43.300 ;
        RECT 398.940 39.900 400.540 41.700 ;
        RECT 303.260 38.300 324.180 39.900 ;
        RECT 322.580 36.500 324.180 38.300 ;
        RECT 364.900 38.300 400.540 39.900 ;
        RECT 364.900 36.500 366.500 38.300 ;
        RECT 322.580 34.900 366.500 36.500 ;
        RECT 420.100 36.500 421.700 41.700 ;
        RECT 485.420 41.700 559.700 43.300 ;
        RECT 485.420 36.500 487.020 41.700 ;
        RECT 420.100 34.900 487.020 36.500 ;
        RECT 558.100 36.500 559.700 41.700 ;
        RECT 605.940 41.700 636.060 43.300 ;
        RECT 605.940 39.900 607.540 41.700 ;
        RECT 571.900 38.300 607.540 39.900 ;
        RECT 634.460 39.900 636.060 41.700 ;
        RECT 678.620 41.700 835.700 43.300 ;
        RECT 678.620 39.900 680.220 41.700 ;
        RECT 634.460 38.300 643.190 39.900 ;
        RECT 571.900 36.500 573.500 38.300 ;
        RECT 558.100 34.900 573.500 36.500 ;
        RECT 641.590 36.500 643.190 38.300 ;
        RECT 675.860 38.300 680.220 39.900 ;
        RECT 834.100 39.900 835.700 41.700 ;
        RECT 896.660 41.700 946.100 43.300 ;
        RECT 896.660 39.900 898.260 41.700 ;
        RECT 834.100 38.300 850.420 39.900 ;
        RECT 675.860 36.500 677.460 38.300 ;
        RECT 641.590 34.900 677.460 36.500 ;
        RECT 848.820 36.500 850.420 38.300 ;
        RECT 882.860 38.300 898.260 39.900 ;
        RECT 882.860 36.500 884.460 38.300 ;
        RECT 848.820 34.900 884.460 36.500 ;
        RECT 944.500 36.500 946.100 41.700 ;
        RECT 1063.180 41.700 1107.100 43.300 ;
        RECT 1063.180 36.500 1064.780 41.700 ;
        RECT 1105.500 39.900 1107.100 41.700 ;
        RECT 1105.500 38.300 1130.100 39.900 ;
        RECT 944.500 34.900 1064.780 36.500 ;
        RECT 1128.500 33.090 1130.100 38.300 ;
        RECT 10.520 31.490 2849.180 33.090 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 6.585 1064.285 6.755 1107.635 ;
        RECT 8.885 703.545 9.055 731.255 ;
        RECT 4.285 630.445 4.455 703.375 ;
        RECT 2.905 8.585 3.075 51.935 ;
      LAYER mcon ;
        RECT 6.585 1107.465 6.755 1107.635 ;
        RECT 8.885 731.085 9.055 731.255 ;
        RECT 4.285 703.205 4.455 703.375 ;
        RECT 2.905 51.765 3.075 51.935 ;
      LAYER met1 ;
        RECT 6.510 1107.620 6.830 1107.680 ;
        RECT 6.315 1107.480 6.830 1107.620 ;
        RECT 6.510 1107.420 6.830 1107.480 ;
        RECT 6.525 1064.440 6.815 1064.485 ;
        RECT 9.730 1064.440 10.050 1064.500 ;
        RECT 6.525 1064.300 10.050 1064.440 ;
        RECT 6.525 1064.255 6.815 1064.300 ;
        RECT 9.730 1064.240 10.050 1064.300 ;
        RECT 9.730 1024.320 10.050 1024.380 ;
        RECT 7.060 1024.180 10.050 1024.320 ;
        RECT 7.060 1024.040 7.200 1024.180 ;
        RECT 9.730 1024.120 10.050 1024.180 ;
        RECT 6.970 1023.780 7.290 1024.040 ;
        RECT 2.830 1001.200 3.150 1001.260 ;
        RECT 6.970 1001.200 7.290 1001.260 ;
        RECT 2.830 1001.060 7.290 1001.200 ;
        RECT 2.830 1001.000 3.150 1001.060 ;
        RECT 6.970 1001.000 7.290 1001.060 ;
        RECT 2.830 731.240 3.150 731.300 ;
        RECT 8.825 731.240 9.115 731.285 ;
        RECT 2.830 731.100 9.115 731.240 ;
        RECT 2.830 731.040 3.150 731.100 ;
        RECT 8.825 731.055 9.115 731.100 ;
        RECT 8.825 703.700 9.115 703.745 ;
        RECT 4.300 703.560 9.115 703.700 ;
        RECT 4.300 703.405 4.440 703.560 ;
        RECT 8.825 703.515 9.115 703.560 ;
        RECT 4.225 703.175 4.515 703.405 ;
        RECT 1.910 630.600 2.230 630.660 ;
        RECT 4.225 630.600 4.515 630.645 ;
        RECT 1.910 630.460 4.515 630.600 ;
        RECT 1.910 630.400 2.230 630.460 ;
        RECT 4.225 630.415 4.515 630.460 ;
        RECT 1.910 490.860 2.230 490.920 ;
        RECT 6.510 490.860 6.830 490.920 ;
        RECT 1.910 490.720 6.830 490.860 ;
        RECT 1.910 490.660 2.230 490.720 ;
        RECT 6.510 490.660 6.830 490.720 ;
        RECT 6.510 417.420 6.830 417.480 ;
        RECT 9.270 417.420 9.590 417.480 ;
        RECT 6.510 417.280 9.590 417.420 ;
        RECT 6.510 417.220 6.830 417.280 ;
        RECT 9.270 417.220 9.590 417.280 ;
        RECT 2.830 363.020 3.150 363.080 ;
        RECT 9.270 363.020 9.590 363.080 ;
        RECT 2.830 362.880 9.590 363.020 ;
        RECT 2.830 362.820 3.150 362.880 ;
        RECT 9.270 362.820 9.590 362.880 ;
        RECT 2.830 51.920 3.150 51.980 ;
        RECT 2.635 51.780 3.150 51.920 ;
        RECT 2.830 51.720 3.150 51.780 ;
        RECT 2.845 8.740 3.135 8.785 ;
        RECT 8.350 8.740 8.670 8.800 ;
        RECT 2.845 8.600 8.670 8.740 ;
        RECT 2.845 8.555 3.135 8.600 ;
        RECT 8.350 8.540 8.670 8.600 ;
      LAYER via ;
        RECT 6.540 1107.420 6.800 1107.680 ;
        RECT 9.760 1064.240 10.020 1064.500 ;
        RECT 9.760 1024.120 10.020 1024.380 ;
        RECT 7.000 1023.780 7.260 1024.040 ;
        RECT 2.860 1001.000 3.120 1001.260 ;
        RECT 7.000 1001.000 7.260 1001.260 ;
        RECT 2.860 731.040 3.120 731.300 ;
        RECT 1.940 630.400 2.200 630.660 ;
        RECT 1.940 490.660 2.200 490.920 ;
        RECT 6.540 490.660 6.800 490.920 ;
        RECT 6.540 417.220 6.800 417.480 ;
        RECT 9.300 417.220 9.560 417.480 ;
        RECT 2.860 362.820 3.120 363.080 ;
        RECT 9.300 362.820 9.560 363.080 ;
        RECT 2.860 51.720 3.120 51.980 ;
        RECT 8.380 8.540 8.640 8.800 ;
      LAYER met2 ;
        RECT 6.530 1191.515 6.810 1191.885 ;
        RECT 6.600 1107.710 6.740 1191.515 ;
        RECT 6.540 1107.390 6.800 1107.710 ;
        RECT 9.760 1064.210 10.020 1064.530 ;
        RECT 9.820 1024.410 9.960 1064.210 ;
        RECT 9.760 1024.090 10.020 1024.410 ;
        RECT 7.000 1023.750 7.260 1024.070 ;
        RECT 7.060 1001.290 7.200 1023.750 ;
        RECT 2.860 1000.970 3.120 1001.290 ;
        RECT 7.000 1000.970 7.260 1001.290 ;
        RECT 2.920 731.330 3.060 1000.970 ;
        RECT 2.860 731.010 3.120 731.330 ;
        RECT 1.940 630.370 2.200 630.690 ;
        RECT 2.000 490.950 2.140 630.370 ;
        RECT 1.940 490.630 2.200 490.950 ;
        RECT 6.540 490.630 6.800 490.950 ;
        RECT 6.600 417.510 6.740 490.630 ;
        RECT 6.540 417.190 6.800 417.510 ;
        RECT 9.300 417.190 9.560 417.510 ;
        RECT 9.360 363.110 9.500 417.190 ;
        RECT 2.860 362.790 3.120 363.110 ;
        RECT 9.300 362.790 9.560 363.110 ;
        RECT 2.920 52.010 3.060 362.790 ;
        RECT 2.860 51.690 3.120 52.010 ;
        RECT 8.380 8.510 8.640 8.830 ;
        RECT 8.440 2.400 8.580 8.510 ;
        RECT 8.230 -4.800 8.790 2.400 ;
      LAYER via2 ;
        RECT 6.530 1191.560 6.810 1191.840 ;
      LAYER met3 ;
        RECT 5.000 1194.360 9.000 1194.960 ;
        RECT 6.750 1191.865 7.050 1194.360 ;
        RECT 6.505 1191.550 7.050 1191.865 ;
        RECT 6.505 1191.535 6.835 1191.550 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1453.745 8.245 1469.095 8.415 ;
        RECT 597.225 6.205 598.315 6.375 ;
        RECT 597.225 5.865 597.395 6.205 ;
        RECT 598.145 5.695 598.315 6.205 ;
        RECT 598.145 5.525 604.295 5.695 ;
        RECT 26.825 0.765 27.915 0.935 ;
        RECT 276.605 0.425 276.775 3.995 ;
        RECT 382.865 3.825 383.035 4.675 ;
        RECT 414.605 3.655 414.775 4.675 ;
        RECT 415.525 3.655 415.695 4.675 ;
        RECT 414.605 3.485 415.695 3.655 ;
        RECT 604.125 1.275 604.295 5.525 ;
        RECT 702.105 4.845 703.195 5.015 ;
        RECT 647.825 1.275 647.995 4.675 ;
        RECT 673.125 3.655 673.295 4.675 ;
        RECT 680.945 3.655 681.115 4.675 ;
        RECT 702.105 4.505 702.275 4.845 ;
        RECT 673.125 3.485 681.115 3.655 ;
        RECT 703.025 3.655 703.195 4.845 ;
        RECT 1195.225 4.165 1197.235 4.335 ;
        RECT 1208.565 4.165 1210.575 4.335 ;
        RECT 724.645 3.825 751.035 3.995 ;
        RECT 724.645 3.655 724.815 3.825 ;
        RECT 703.025 3.485 724.815 3.655 ;
        RECT 750.865 2.975 751.035 3.825 ;
        RECT 756.845 3.145 757.935 3.315 ;
        RECT 750.865 2.805 752.415 2.975 ;
        RECT 756.845 2.805 757.015 3.145 ;
        RECT 757.765 2.295 757.935 3.145 ;
        RECT 757.305 2.125 757.935 2.295 ;
        RECT 757.305 1.615 757.475 2.125 ;
        RECT 796.405 1.955 796.575 3.315 ;
        RECT 1430.745 3.145 1430.915 4.335 ;
        RECT 1448.225 2.975 1448.395 3.315 ;
        RECT 1453.745 2.975 1453.915 8.245 ;
        RECT 1468.925 7.905 1469.095 8.245 ;
        RECT 1520.905 7.565 1521.075 8.415 ;
        RECT 1573.345 8.245 1573.975 8.415 ;
        RECT 1573.805 3.825 1573.975 8.245 ;
        RECT 1587.605 4.845 1593.755 5.015 ;
        RECT 1587.605 3.825 1587.775 4.845 ;
        RECT 1782.185 3.825 1782.355 7.395 ;
        RECT 1448.225 2.805 1453.915 2.975 ;
        RECT 758.225 1.785 766.675 1.955 ;
        RECT 785.825 1.785 796.575 1.955 ;
        RECT 758.225 1.615 758.395 1.785 ;
        RECT 757.305 1.445 758.395 1.615 ;
        RECT 604.125 1.105 647.995 1.275 ;
      LAYER mcon ;
        RECT 382.865 4.505 383.035 4.675 ;
        RECT 276.605 3.825 276.775 3.995 ;
        RECT 414.605 4.505 414.775 4.675 ;
        RECT 27.745 0.765 27.915 0.935 ;
        RECT 415.525 4.505 415.695 4.675 ;
        RECT 647.825 4.505 647.995 4.675 ;
        RECT 673.125 4.505 673.295 4.675 ;
        RECT 680.945 4.505 681.115 4.675 ;
        RECT 1197.065 4.165 1197.235 4.335 ;
        RECT 1210.405 4.165 1210.575 4.335 ;
        RECT 1430.745 4.165 1430.915 4.335 ;
        RECT 752.245 2.805 752.415 2.975 ;
        RECT 796.405 3.145 796.575 3.315 ;
        RECT 1448.225 3.145 1448.395 3.315 ;
        RECT 1520.905 8.245 1521.075 8.415 ;
        RECT 1782.185 7.225 1782.355 7.395 ;
        RECT 1593.585 4.845 1593.755 5.015 ;
        RECT 766.505 1.785 766.675 1.955 ;
      LAYER met1 ;
        RECT 1520.845 8.400 1521.135 8.445 ;
        RECT 1573.285 8.400 1573.575 8.445 ;
        RECT 1520.845 8.260 1573.575 8.400 ;
        RECT 1520.845 8.215 1521.135 8.260 ;
        RECT 1573.285 8.215 1573.575 8.260 ;
        RECT 1468.865 8.060 1469.155 8.105 ;
        RECT 1468.865 7.920 1493.920 8.060 ;
        RECT 1468.865 7.875 1469.155 7.920 ;
        RECT 1493.780 7.720 1493.920 7.920 ;
        RECT 1520.845 7.720 1521.135 7.765 ;
        RECT 1493.780 7.580 1521.135 7.720 ;
        RECT 1520.845 7.535 1521.135 7.580 ;
        RECT 1782.125 7.380 1782.415 7.425 ;
        RECT 1926.550 7.380 1926.870 7.440 ;
        RECT 1782.125 7.240 1926.870 7.380 ;
        RECT 1782.125 7.195 1782.415 7.240 ;
        RECT 1926.550 7.180 1926.870 7.240 ;
        RECT 596.690 6.020 597.010 6.080 ;
        RECT 597.165 6.020 597.455 6.065 ;
        RECT 596.690 5.880 597.455 6.020 ;
        RECT 596.690 5.820 597.010 5.880 ;
        RECT 597.165 5.835 597.455 5.880 ;
        RECT 1593.525 5.000 1593.815 5.045 ;
        RECT 1597.190 5.000 1597.510 5.060 ;
        RECT 1593.525 4.860 1597.510 5.000 ;
        RECT 1593.525 4.815 1593.815 4.860 ;
        RECT 1597.190 4.800 1597.510 4.860 ;
        RECT 382.805 4.660 383.095 4.705 ;
        RECT 414.545 4.660 414.835 4.705 ;
        RECT 382.805 4.520 414.835 4.660 ;
        RECT 382.805 4.475 383.095 4.520 ;
        RECT 414.545 4.475 414.835 4.520 ;
        RECT 415.465 4.660 415.755 4.705 ;
        RECT 486.290 4.660 486.610 4.720 ;
        RECT 415.465 4.520 486.610 4.660 ;
        RECT 415.465 4.475 415.755 4.520 ;
        RECT 486.290 4.460 486.610 4.520 ;
        RECT 647.765 4.660 648.055 4.705 ;
        RECT 673.065 4.660 673.355 4.705 ;
        RECT 647.765 4.520 673.355 4.660 ;
        RECT 647.765 4.475 648.055 4.520 ;
        RECT 673.065 4.475 673.355 4.520 ;
        RECT 680.885 4.660 681.175 4.705 ;
        RECT 702.045 4.660 702.335 4.705 ;
        RECT 680.885 4.520 702.335 4.660 ;
        RECT 680.885 4.475 681.175 4.520 ;
        RECT 702.045 4.475 702.335 4.520 ;
        RECT 887.870 4.320 888.190 4.380 ;
        RECT 830.000 4.180 879.820 4.320 ;
        RECT 276.545 3.980 276.835 4.025 ;
        RECT 382.805 3.980 383.095 4.025 ;
        RECT 830.000 3.980 830.140 4.180 ;
        RECT 276.545 3.840 383.095 3.980 ;
        RECT 276.545 3.795 276.835 3.840 ;
        RECT 382.805 3.795 383.095 3.840 ;
        RECT 815.740 3.840 830.140 3.980 ;
        RECT 879.680 3.980 879.820 4.180 ;
        RECT 881.980 4.180 888.190 4.320 ;
        RECT 881.980 3.980 882.120 4.180 ;
        RECT 887.870 4.120 888.190 4.180 ;
        RECT 903.510 4.320 903.830 4.380 ;
        RECT 1195.165 4.320 1195.455 4.365 ;
        RECT 903.510 4.180 1195.455 4.320 ;
        RECT 903.510 4.120 903.830 4.180 ;
        RECT 1195.165 4.135 1195.455 4.180 ;
        RECT 1197.005 4.320 1197.295 4.365 ;
        RECT 1208.505 4.320 1208.795 4.365 ;
        RECT 1197.005 4.180 1208.795 4.320 ;
        RECT 1197.005 4.135 1197.295 4.180 ;
        RECT 1208.505 4.135 1208.795 4.180 ;
        RECT 1210.345 4.320 1210.635 4.365 ;
        RECT 1430.685 4.320 1430.975 4.365 ;
        RECT 1210.345 4.180 1430.975 4.320 ;
        RECT 1210.345 4.135 1210.635 4.180 ;
        RECT 1430.685 4.135 1430.975 4.180 ;
        RECT 879.680 3.840 882.120 3.980 ;
        RECT 1573.745 3.980 1574.035 4.025 ;
        RECT 1587.545 3.980 1587.835 4.025 ;
        RECT 1573.745 3.840 1587.835 3.980 ;
        RECT 803.690 3.640 804.010 3.700 ;
        RECT 815.740 3.640 815.880 3.840 ;
        RECT 1573.745 3.795 1574.035 3.840 ;
        RECT 1587.545 3.795 1587.835 3.840 ;
        RECT 1598.570 3.980 1598.890 4.040 ;
        RECT 1782.125 3.980 1782.415 4.025 ;
        RECT 1598.570 3.840 1782.415 3.980 ;
        RECT 1598.570 3.780 1598.890 3.840 ;
        RECT 1782.125 3.795 1782.415 3.840 ;
        RECT 803.690 3.500 815.880 3.640 ;
        RECT 803.690 3.440 804.010 3.500 ;
        RECT 796.345 3.300 796.635 3.345 ;
        RECT 797.250 3.300 797.570 3.360 ;
        RECT 796.345 3.160 797.570 3.300 ;
        RECT 796.345 3.115 796.635 3.160 ;
        RECT 797.250 3.100 797.570 3.160 ;
        RECT 1430.685 3.300 1430.975 3.345 ;
        RECT 1448.165 3.300 1448.455 3.345 ;
        RECT 1430.685 3.160 1448.455 3.300 ;
        RECT 1430.685 3.115 1430.975 3.160 ;
        RECT 1448.165 3.115 1448.455 3.160 ;
        RECT 752.185 2.960 752.475 3.005 ;
        RECT 756.785 2.960 757.075 3.005 ;
        RECT 752.185 2.820 757.075 2.960 ;
        RECT 752.185 2.775 752.475 2.820 ;
        RECT 756.785 2.775 757.075 2.820 ;
        RECT 766.445 1.940 766.735 1.985 ;
        RECT 768.730 1.940 769.050 2.000 ;
        RECT 766.445 1.800 769.050 1.940 ;
        RECT 766.445 1.755 766.735 1.800 ;
        RECT 768.730 1.740 769.050 1.800 ;
        RECT 773.330 1.940 773.650 2.000 ;
        RECT 785.765 1.940 786.055 1.985 ;
        RECT 773.330 1.800 786.055 1.940 ;
        RECT 773.330 1.740 773.650 1.800 ;
        RECT 785.765 1.755 786.055 1.800 ;
        RECT 191.890 1.260 192.210 1.320 ;
        RECT 131.260 1.120 192.210 1.260 ;
        RECT 15.250 0.920 15.570 0.980 ;
        RECT 26.765 0.920 27.055 0.965 ;
        RECT 15.250 0.780 27.055 0.920 ;
        RECT 15.250 0.720 15.570 0.780 ;
        RECT 26.765 0.735 27.055 0.780 ;
        RECT 27.685 0.920 27.975 0.965 ;
        RECT 131.260 0.920 131.400 1.120 ;
        RECT 191.890 1.060 192.210 1.120 ;
        RECT 27.685 0.780 131.400 0.920 ;
        RECT 27.685 0.735 27.975 0.780 ;
        RECT 231.450 0.580 231.770 0.640 ;
        RECT 276.545 0.580 276.835 0.625 ;
        RECT 231.450 0.440 276.835 0.580 ;
        RECT 231.450 0.380 231.770 0.440 ;
        RECT 276.545 0.395 276.835 0.440 ;
      LAYER via ;
        RECT 1926.580 7.180 1926.840 7.440 ;
        RECT 596.720 5.820 596.980 6.080 ;
        RECT 1597.220 4.800 1597.480 5.060 ;
        RECT 486.320 4.460 486.580 4.720 ;
        RECT 887.900 4.120 888.160 4.380 ;
        RECT 903.540 4.120 903.800 4.380 ;
        RECT 803.720 3.440 803.980 3.700 ;
        RECT 1598.600 3.780 1598.860 4.040 ;
        RECT 797.280 3.100 797.540 3.360 ;
        RECT 768.760 1.740 769.020 2.000 ;
        RECT 773.360 1.740 773.620 2.000 ;
        RECT 15.280 0.720 15.540 0.980 ;
        RECT 191.920 1.060 192.180 1.320 ;
        RECT 231.480 0.380 231.740 0.640 ;
      LAYER met2 ;
        RECT 1926.580 7.210 1926.840 7.470 ;
        RECT 1928.350 7.210 1928.630 9.000 ;
        RECT 1926.580 7.150 1928.630 7.210 ;
        RECT 1926.640 7.070 1928.630 7.150 ;
        RECT 584.290 6.275 584.570 6.645 ;
        RECT 584.360 6.020 584.500 6.275 ;
        RECT 596.720 6.020 596.980 6.110 ;
        RECT 584.360 5.880 596.980 6.020 ;
        RECT 596.720 5.790 596.980 5.880 ;
        RECT 486.310 4.915 486.590 5.285 ;
        RECT 486.380 4.750 486.520 4.915 ;
        RECT 1597.220 4.770 1597.480 5.090 ;
        RECT 1928.350 5.000 1928.630 7.070 ;
        RECT 486.320 4.430 486.580 4.750 ;
        RECT 1597.280 4.490 1597.420 4.770 ;
        RECT 887.900 4.090 888.160 4.410 ;
        RECT 903.540 4.090 903.800 4.410 ;
        RECT 1597.280 4.350 1598.800 4.490 ;
        RECT 191.910 3.555 192.190 3.925 ;
        RECT 231.470 3.555 231.750 3.925 ;
        RECT 887.960 3.810 888.100 4.090 ;
        RECT 803.720 3.640 803.980 3.730 ;
        RECT 887.960 3.670 890.400 3.810 ;
        RECT 14.420 2.820 15.480 2.960 ;
        RECT 14.420 2.400 14.560 2.820 ;
        RECT 14.210 -4.800 14.770 2.400 ;
        RECT 15.340 1.010 15.480 2.820 ;
        RECT 191.980 1.350 192.120 3.555 ;
        RECT 191.920 1.030 192.180 1.350 ;
        RECT 15.280 0.690 15.540 1.010 ;
        RECT 231.540 0.670 231.680 3.555 ;
        RECT 799.180 3.500 803.980 3.640 ;
        RECT 797.280 3.130 797.540 3.390 ;
        RECT 799.180 3.130 799.320 3.500 ;
        RECT 803.720 3.410 803.980 3.500 ;
        RECT 768.820 2.990 770.800 3.130 ;
        RECT 797.280 3.070 799.320 3.130 ;
        RECT 797.340 2.990 799.320 3.070 ;
        RECT 768.820 2.030 768.960 2.990 ;
        RECT 768.760 1.710 769.020 2.030 ;
        RECT 770.660 1.940 770.800 2.990 ;
        RECT 890.260 2.620 890.400 3.670 ;
        RECT 903.600 2.960 903.740 4.090 ;
        RECT 1598.660 4.070 1598.800 4.350 ;
        RECT 1598.600 3.750 1598.860 4.070 ;
        RECT 892.100 2.820 903.740 2.960 ;
        RECT 892.100 2.620 892.240 2.820 ;
        RECT 890.260 2.480 892.240 2.620 ;
        RECT 773.360 1.940 773.620 2.030 ;
        RECT 770.660 1.800 773.620 1.940 ;
        RECT 773.360 1.710 773.620 1.800 ;
        RECT 231.480 0.350 231.740 0.670 ;
      LAYER via2 ;
        RECT 584.290 6.320 584.570 6.600 ;
        RECT 486.310 4.960 486.590 5.240 ;
        RECT 191.910 3.600 192.190 3.880 ;
        RECT 231.470 3.600 231.750 3.880 ;
      LAYER met3 ;
        RECT 584.265 6.610 584.595 6.625 ;
        RECT 534.830 6.310 584.595 6.610 ;
        RECT 486.285 5.250 486.615 5.265 ;
        RECT 534.830 5.250 535.130 6.310 ;
        RECT 584.265 6.295 584.595 6.310 ;
        RECT 486.285 4.950 535.130 5.250 ;
        RECT 486.285 4.935 486.615 4.950 ;
        RECT 191.885 3.890 192.215 3.905 ;
        RECT 231.445 3.890 231.775 3.905 ;
        RECT 191.885 3.590 231.775 3.890 ;
        RECT 191.885 3.575 192.215 3.590 ;
        RECT 231.445 3.575 231.775 3.590 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 789.505 9.265 806.695 9.435 ;
        RECT 786.285 8.925 788.755 9.095 ;
        RECT 551.225 8.245 552.775 8.415 ;
        RECT 551.225 3.655 551.395 8.245 ;
        RECT 552.605 8.075 552.775 8.245 ;
        RECT 552.605 7.905 555.075 8.075 ;
        RECT 513.045 3.485 516.435 3.655 ;
        RECT 516.265 2.975 516.435 3.485 ;
        RECT 545.705 3.485 551.395 3.655 ;
        RECT 545.705 3.315 545.875 3.485 ;
        RECT 516.725 3.145 545.875 3.315 ;
        RECT 516.725 2.975 516.895 3.145 ;
        RECT 516.265 2.805 516.895 2.975 ;
        RECT 554.905 2.805 555.075 7.905 ;
        RECT 715.905 6.885 718.375 7.055 ;
        RECT 644.605 5.185 659.495 5.355 ;
        RECT 557.205 3.145 558.755 3.315 ;
        RECT 560.885 3.145 566.115 3.315 ;
        RECT 557.205 2.805 557.375 3.145 ;
        RECT 565.945 0.255 566.115 3.145 ;
        RECT 600.905 0.255 601.075 5.015 ;
        RECT 606.885 4.675 607.055 5.015 ;
        RECT 644.605 4.845 644.775 5.185 ;
        RECT 606.885 4.505 607.515 4.675 ;
        RECT 607.345 3.825 607.515 4.505 ;
        RECT 659.325 3.995 659.495 5.185 ;
        RECT 663.925 4.845 673.755 5.015 ;
        RECT 663.925 3.995 664.095 4.845 ;
        RECT 659.325 3.825 664.095 3.995 ;
        RECT 673.585 3.995 673.755 4.845 ;
        RECT 677.725 3.995 677.895 6.375 ;
        RECT 715.905 4.505 716.075 6.885 ;
        RECT 720.505 6.715 720.675 7.055 ;
        RECT 720.505 6.545 725.275 6.715 ;
        RECT 725.105 6.375 725.275 6.545 ;
        RECT 728.325 6.375 728.495 7.395 ;
        RECT 737.065 7.055 737.235 7.395 ;
        RECT 748.105 7.055 748.275 8.075 ;
        RECT 752.245 7.905 752.415 8.755 ;
        RECT 737.065 6.885 739.075 7.055 ;
        RECT 743.965 6.885 748.275 7.055 ;
        RECT 725.105 6.205 728.495 6.375 ;
        RECT 756.385 6.205 756.555 8.755 ;
        RECT 762.365 8.245 763.915 8.415 ;
        RECT 758.685 7.905 760.235 8.075 ;
        RECT 758.685 6.205 758.855 7.905 ;
        RECT 760.065 7.395 760.235 7.905 ;
        RECT 762.365 7.395 762.535 8.245 ;
        RECT 763.745 7.905 763.915 8.245 ;
        RECT 767.885 7.735 768.055 8.075 ;
        RECT 767.885 7.565 768.975 7.735 ;
        RECT 781.685 7.565 781.855 8.755 ;
        RECT 788.585 8.415 788.755 8.925 ;
        RECT 789.505 8.415 789.675 9.265 ;
        RECT 788.585 8.245 789.675 8.415 ;
        RECT 760.065 7.225 762.535 7.395 ;
        RECT 806.525 4.165 806.695 9.265 ;
        RECT 896.685 4.505 897.775 4.675 ;
        RECT 1090.345 4.505 1092.355 4.675 ;
        RECT 1209.485 4.505 1211.035 4.675 ;
        RECT 673.585 3.825 677.895 3.995 ;
        RECT 1588.065 3.825 1588.235 4.675 ;
        RECT 1597.265 3.825 1597.435 7.735 ;
        RECT 565.945 0.085 601.075 0.255 ;
      LAYER mcon ;
        RECT 752.245 8.585 752.415 8.755 ;
        RECT 748.105 7.905 748.275 8.075 ;
        RECT 756.385 8.585 756.555 8.755 ;
        RECT 728.325 7.225 728.495 7.395 ;
        RECT 718.205 6.885 718.375 7.055 ;
        RECT 720.505 6.885 720.675 7.055 ;
        RECT 677.725 6.205 677.895 6.375 ;
        RECT 600.905 4.845 601.075 5.015 ;
        RECT 558.585 3.145 558.755 3.315 ;
        RECT 606.885 4.845 607.055 5.015 ;
        RECT 737.065 7.225 737.235 7.395 ;
        RECT 738.905 6.885 739.075 7.055 ;
        RECT 781.685 8.585 781.855 8.755 ;
        RECT 767.885 7.905 768.055 8.075 ;
        RECT 768.805 7.565 768.975 7.735 ;
        RECT 1597.265 7.565 1597.435 7.735 ;
        RECT 897.605 4.505 897.775 4.675 ;
        RECT 1092.185 4.505 1092.355 4.675 ;
        RECT 1210.865 4.505 1211.035 4.675 ;
        RECT 1588.065 4.505 1588.235 4.675 ;
      LAYER met1 ;
        RECT 786.225 9.080 786.515 9.125 ;
        RECT 783.080 8.940 786.515 9.080 ;
        RECT 752.185 8.740 752.475 8.785 ;
        RECT 756.325 8.740 756.615 8.785 ;
        RECT 752.185 8.600 756.615 8.740 ;
        RECT 752.185 8.555 752.475 8.600 ;
        RECT 756.325 8.555 756.615 8.600 ;
        RECT 781.625 8.740 781.915 8.785 ;
        RECT 783.080 8.740 783.220 8.940 ;
        RECT 786.225 8.895 786.515 8.940 ;
        RECT 781.625 8.600 783.220 8.740 ;
        RECT 781.625 8.555 781.915 8.600 ;
        RECT 748.045 8.060 748.335 8.105 ;
        RECT 752.185 8.060 752.475 8.105 ;
        RECT 748.045 7.920 752.475 8.060 ;
        RECT 748.045 7.875 748.335 7.920 ;
        RECT 752.185 7.875 752.475 7.920 ;
        RECT 763.685 8.060 763.975 8.105 ;
        RECT 767.825 8.060 768.115 8.105 ;
        RECT 763.685 7.920 768.115 8.060 ;
        RECT 763.685 7.875 763.975 7.920 ;
        RECT 767.825 7.875 768.115 7.920 ;
        RECT 768.745 7.720 769.035 7.765 ;
        RECT 781.625 7.720 781.915 7.765 ;
        RECT 768.745 7.580 781.915 7.720 ;
        RECT 768.745 7.535 769.035 7.580 ;
        RECT 781.625 7.535 781.915 7.580 ;
        RECT 1597.205 7.720 1597.495 7.765 ;
        RECT 2116.990 7.720 2117.310 7.780 ;
        RECT 1597.205 7.580 2117.310 7.720 ;
        RECT 1597.205 7.535 1597.495 7.580 ;
        RECT 2116.990 7.520 2117.310 7.580 ;
        RECT 728.265 7.380 728.555 7.425 ;
        RECT 737.005 7.380 737.295 7.425 ;
        RECT 728.265 7.240 737.295 7.380 ;
        RECT 728.265 7.195 728.555 7.240 ;
        RECT 737.005 7.195 737.295 7.240 ;
        RECT 718.145 7.040 718.435 7.085 ;
        RECT 720.445 7.040 720.735 7.085 ;
        RECT 718.145 6.900 720.735 7.040 ;
        RECT 718.145 6.855 718.435 6.900 ;
        RECT 720.445 6.855 720.735 6.900 ;
        RECT 738.845 7.040 739.135 7.085 ;
        RECT 743.905 7.040 744.195 7.085 ;
        RECT 738.845 6.900 744.195 7.040 ;
        RECT 738.845 6.855 739.135 6.900 ;
        RECT 743.905 6.855 744.195 6.900 ;
        RECT 677.665 6.360 677.955 6.405 ;
        RECT 703.870 6.360 704.190 6.420 ;
        RECT 677.665 6.220 704.190 6.360 ;
        RECT 677.665 6.175 677.955 6.220 ;
        RECT 703.870 6.160 704.190 6.220 ;
        RECT 756.325 6.360 756.615 6.405 ;
        RECT 758.625 6.360 758.915 6.405 ;
        RECT 756.325 6.220 758.915 6.360 ;
        RECT 756.325 6.175 756.615 6.220 ;
        RECT 758.625 6.175 758.915 6.220 ;
        RECT 600.845 5.000 601.135 5.045 ;
        RECT 606.825 5.000 607.115 5.045 ;
        RECT 600.845 4.860 607.115 5.000 ;
        RECT 600.845 4.815 601.135 4.860 ;
        RECT 606.825 4.815 607.115 4.860 ;
        RECT 612.330 5.000 612.650 5.060 ;
        RECT 619.690 5.000 620.010 5.060 ;
        RECT 612.330 4.860 620.010 5.000 ;
        RECT 612.330 4.800 612.650 4.860 ;
        RECT 619.690 4.800 620.010 4.860 ;
        RECT 627.970 5.000 628.290 5.060 ;
        RECT 644.545 5.000 644.835 5.045 ;
        RECT 627.970 4.860 644.835 5.000 ;
        RECT 627.970 4.800 628.290 4.860 ;
        RECT 644.545 4.815 644.835 4.860 ;
        RECT 712.150 4.660 712.470 4.720 ;
        RECT 715.845 4.660 716.135 4.705 ;
        RECT 896.625 4.660 896.915 4.705 ;
        RECT 712.150 4.520 716.135 4.660 ;
        RECT 712.150 4.460 712.470 4.520 ;
        RECT 715.845 4.475 716.135 4.520 ;
        RECT 822.180 4.520 896.915 4.660 ;
        RECT 806.465 4.320 806.755 4.365 ;
        RECT 822.180 4.320 822.320 4.520 ;
        RECT 896.625 4.475 896.915 4.520 ;
        RECT 897.545 4.660 897.835 4.705 ;
        RECT 1090.285 4.660 1090.575 4.705 ;
        RECT 897.545 4.520 1090.575 4.660 ;
        RECT 897.545 4.475 897.835 4.520 ;
        RECT 1090.285 4.475 1090.575 4.520 ;
        RECT 1092.125 4.660 1092.415 4.705 ;
        RECT 1209.425 4.660 1209.715 4.705 ;
        RECT 1092.125 4.520 1209.715 4.660 ;
        RECT 1092.125 4.475 1092.415 4.520 ;
        RECT 1209.425 4.475 1209.715 4.520 ;
        RECT 1210.805 4.660 1211.095 4.705 ;
        RECT 1588.005 4.660 1588.295 4.705 ;
        RECT 1210.805 4.520 1588.295 4.660 ;
        RECT 1210.805 4.475 1211.095 4.520 ;
        RECT 1588.005 4.475 1588.295 4.520 ;
        RECT 806.465 4.180 822.320 4.320 ;
        RECT 806.465 4.135 806.755 4.180 ;
        RECT 607.285 3.980 607.575 4.025 ;
        RECT 612.330 3.980 612.650 4.040 ;
        RECT 607.285 3.840 612.650 3.980 ;
        RECT 607.285 3.795 607.575 3.840 ;
        RECT 612.330 3.780 612.650 3.840 ;
        RECT 1588.005 3.980 1588.295 4.025 ;
        RECT 1597.205 3.980 1597.495 4.025 ;
        RECT 1588.005 3.840 1597.495 3.980 ;
        RECT 1588.005 3.795 1588.295 3.840 ;
        RECT 1597.205 3.795 1597.495 3.840 ;
        RECT 512.050 3.640 512.370 3.700 ;
        RECT 512.985 3.640 513.275 3.685 ;
        RECT 512.050 3.500 513.275 3.640 ;
        RECT 512.050 3.440 512.370 3.500 ;
        RECT 512.985 3.455 513.275 3.500 ;
        RECT 558.525 3.300 558.815 3.345 ;
        RECT 560.825 3.300 561.115 3.345 ;
        RECT 558.525 3.160 561.115 3.300 ;
        RECT 558.525 3.115 558.815 3.160 ;
        RECT 560.825 3.115 561.115 3.160 ;
        RECT 554.845 2.960 555.135 3.005 ;
        RECT 557.145 2.960 557.435 3.005 ;
        RECT 554.845 2.820 557.435 2.960 ;
        RECT 554.845 2.775 555.135 2.820 ;
        RECT 557.145 2.775 557.435 2.820 ;
      LAYER via ;
        RECT 2117.020 7.520 2117.280 7.780 ;
        RECT 703.900 6.160 704.160 6.420 ;
        RECT 612.360 4.800 612.620 5.060 ;
        RECT 619.720 4.800 619.980 5.060 ;
        RECT 628.000 4.800 628.260 5.060 ;
        RECT 712.180 4.460 712.440 4.720 ;
        RECT 612.360 3.780 612.620 4.040 ;
        RECT 512.080 3.440 512.340 3.700 ;
      LAYER met2 ;
        RECT 2118.330 7.890 2118.610 9.000 ;
        RECT 2117.080 7.810 2118.610 7.890 ;
        RECT 2117.020 7.750 2118.610 7.810 ;
        RECT 2117.020 7.490 2117.280 7.750 ;
        RECT 703.900 6.360 704.160 6.450 ;
        RECT 703.900 6.220 712.380 6.360 ;
        RECT 703.900 6.130 704.160 6.220 ;
        RECT 612.360 4.770 612.620 5.090 ;
        RECT 619.720 5.000 619.980 5.090 ;
        RECT 628.000 5.000 628.260 5.090 ;
        RECT 619.720 4.860 628.260 5.000 ;
        RECT 619.720 4.770 619.980 4.860 ;
        RECT 628.000 4.770 628.260 4.860 ;
        RECT 240.670 4.235 240.950 4.605 ;
        RECT 240.740 2.400 240.880 4.235 ;
        RECT 612.420 4.070 612.560 4.770 ;
        RECT 712.240 4.750 712.380 6.220 ;
        RECT 2118.330 5.000 2118.610 7.750 ;
        RECT 712.180 4.430 712.440 4.750 ;
        RECT 458.710 3.810 458.990 3.925 ;
        RECT 460.090 3.810 460.370 3.925 ;
        RECT 458.710 3.670 460.370 3.810 ;
        RECT 458.710 3.555 458.990 3.670 ;
        RECT 460.090 3.555 460.370 3.670 ;
        RECT 511.150 3.640 511.430 3.925 ;
        RECT 612.360 3.750 612.620 4.070 ;
        RECT 512.080 3.640 512.340 3.730 ;
        RECT 511.150 3.555 512.340 3.640 ;
        RECT 511.220 3.500 512.340 3.555 ;
        RECT 512.080 3.410 512.340 3.500 ;
        RECT 240.530 -4.800 241.090 2.400 ;
      LAYER via2 ;
        RECT 240.670 4.280 240.950 4.560 ;
        RECT 458.710 3.600 458.990 3.880 ;
        RECT 460.090 3.600 460.370 3.880 ;
        RECT 511.150 3.600 511.430 3.880 ;
      LAYER met3 ;
        RECT 240.645 4.570 240.975 4.585 ;
        RECT 240.645 4.270 279.370 4.570 ;
        RECT 240.645 4.255 240.975 4.270 ;
        RECT 279.070 3.890 279.370 4.270 ;
        RECT 458.685 3.890 459.015 3.905 ;
        RECT 279.070 3.590 459.015 3.890 ;
        RECT 458.685 3.575 459.015 3.590 ;
        RECT 460.065 3.890 460.395 3.905 ;
        RECT 511.125 3.890 511.455 3.905 ;
        RECT 460.065 3.590 511.455 3.890 ;
        RECT 460.065 3.575 460.395 3.590 ;
        RECT 511.125 3.575 511.455 3.590 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1485.025 8.925 1493.475 9.095 ;
        RECT 769.265 3.655 769.435 3.995 ;
        RECT 770.645 3.655 770.815 5.695 ;
        RECT 769.265 3.485 770.815 3.655 ;
        RECT 1263.305 3.315 1263.475 8.755 ;
        RECT 1267.905 8.585 1286.015 8.755 ;
        RECT 1290.905 8.585 1291.995 8.755 ;
        RECT 1309.305 8.585 1311.775 8.755 ;
        RECT 1485.025 3.315 1485.195 8.925 ;
        RECT 1493.305 8.415 1493.475 8.925 ;
        RECT 1493.305 8.245 1500.375 8.415 ;
        RECT 1520.445 7.395 1520.615 8.415 ;
        RECT 1521.365 7.395 1521.535 7.735 ;
        RECT 1520.445 7.225 1521.535 7.395 ;
        RECT 2060.945 3.485 2061.115 8.075 ;
        RECT 1262.845 3.145 1263.475 3.315 ;
        RECT 1450.985 3.145 1453.455 3.315 ;
        RECT 1484.565 3.145 1485.195 3.315 ;
      LAYER mcon ;
        RECT 1263.305 8.585 1263.475 8.755 ;
        RECT 1285.845 8.585 1286.015 8.755 ;
        RECT 1291.825 8.585 1291.995 8.755 ;
        RECT 1311.605 8.585 1311.775 8.755 ;
        RECT 770.645 5.525 770.815 5.695 ;
        RECT 769.265 3.825 769.435 3.995 ;
        RECT 1500.205 8.245 1500.375 8.415 ;
        RECT 1520.445 8.245 1520.615 8.415 ;
        RECT 2060.945 7.905 2061.115 8.075 ;
        RECT 1521.365 7.565 1521.535 7.735 ;
        RECT 1453.285 3.145 1453.455 3.315 ;
      LAYER met1 ;
        RECT 1263.245 8.740 1263.535 8.785 ;
        RECT 1267.845 8.740 1268.135 8.785 ;
        RECT 1263.245 8.600 1268.135 8.740 ;
        RECT 1263.245 8.555 1263.535 8.600 ;
        RECT 1267.845 8.555 1268.135 8.600 ;
        RECT 1285.785 8.740 1286.075 8.785 ;
        RECT 1290.845 8.740 1291.135 8.785 ;
        RECT 1285.785 8.600 1291.135 8.740 ;
        RECT 1285.785 8.555 1286.075 8.600 ;
        RECT 1290.845 8.555 1291.135 8.600 ;
        RECT 1291.765 8.740 1292.055 8.785 ;
        RECT 1309.245 8.740 1309.535 8.785 ;
        RECT 1291.765 8.600 1309.535 8.740 ;
        RECT 1291.765 8.555 1292.055 8.600 ;
        RECT 1309.245 8.555 1309.535 8.600 ;
        RECT 1311.530 8.740 1311.850 8.800 ;
        RECT 1311.530 8.600 1312.045 8.740 ;
        RECT 1311.530 8.540 1311.850 8.600 ;
        RECT 1500.145 8.400 1500.435 8.445 ;
        RECT 1520.385 8.400 1520.675 8.445 ;
        RECT 1500.145 8.260 1520.675 8.400 ;
        RECT 1500.145 8.215 1500.435 8.260 ;
        RECT 1520.385 8.215 1520.675 8.260 ;
        RECT 2060.885 8.060 2061.175 8.105 ;
        RECT 2164.830 8.060 2165.150 8.120 ;
        RECT 2060.885 7.920 2165.150 8.060 ;
        RECT 2060.885 7.875 2061.175 7.920 ;
        RECT 2164.830 7.860 2165.150 7.920 ;
        RECT 1521.305 7.720 1521.595 7.765 ;
        RECT 1527.730 7.720 1528.050 7.780 ;
        RECT 1521.305 7.580 1528.050 7.720 ;
        RECT 1521.305 7.535 1521.595 7.580 ;
        RECT 1527.730 7.520 1528.050 7.580 ;
        RECT 1249.430 7.380 1249.750 7.440 ;
        RECT 1253.570 7.380 1253.890 7.440 ;
        RECT 1249.430 7.240 1253.890 7.380 ;
        RECT 1249.430 7.180 1249.750 7.240 ;
        RECT 1253.570 7.180 1253.890 7.240 ;
        RECT 919.610 6.020 919.930 6.080 ;
        RECT 947.210 6.020 947.530 6.080 ;
        RECT 919.610 5.880 947.530 6.020 ;
        RECT 919.610 5.820 919.930 5.880 ;
        RECT 947.210 5.820 947.530 5.880 ;
        RECT 770.585 5.680 770.875 5.725 ;
        RECT 771.030 5.680 771.350 5.740 ;
        RECT 770.585 5.540 771.350 5.680 ;
        RECT 770.585 5.495 770.875 5.540 ;
        RECT 771.030 5.480 771.350 5.540 ;
        RECT 1237.470 5.340 1237.790 5.400 ;
        RECT 1241.150 5.340 1241.470 5.400 ;
        RECT 1237.470 5.200 1241.470 5.340 ;
        RECT 1237.470 5.140 1237.790 5.200 ;
        RECT 1241.150 5.140 1241.470 5.200 ;
        RECT 1550.270 4.320 1550.590 4.380 ;
        RECT 1550.270 4.180 1597.880 4.320 ;
        RECT 1550.270 4.120 1550.590 4.180 ;
        RECT 767.350 3.980 767.670 4.040 ;
        RECT 769.205 3.980 769.495 4.025 ;
        RECT 767.350 3.840 769.495 3.980 ;
        RECT 767.350 3.780 767.670 3.840 ;
        RECT 769.205 3.795 769.495 3.840 ;
        RECT 1597.740 3.640 1597.880 4.180 ;
        RECT 2060.885 3.640 2061.175 3.685 ;
        RECT 1597.740 3.500 2061.175 3.640 ;
        RECT 2060.885 3.455 2061.175 3.500 ;
        RECT 1260.010 3.300 1260.330 3.360 ;
        RECT 1262.785 3.300 1263.075 3.345 ;
        RECT 1260.010 3.160 1263.075 3.300 ;
        RECT 1260.010 3.100 1260.330 3.160 ;
        RECT 1262.785 3.115 1263.075 3.160 ;
        RECT 1448.610 3.300 1448.930 3.360 ;
        RECT 1450.925 3.300 1451.215 3.345 ;
        RECT 1448.610 3.160 1451.215 3.300 ;
        RECT 1448.610 3.100 1448.930 3.160 ;
        RECT 1450.925 3.115 1451.215 3.160 ;
        RECT 1453.225 3.300 1453.515 3.345 ;
        RECT 1484.505 3.300 1484.795 3.345 ;
        RECT 1453.225 3.160 1484.795 3.300 ;
        RECT 1453.225 3.115 1453.515 3.160 ;
        RECT 1484.505 3.115 1484.795 3.160 ;
      LAYER via ;
        RECT 1311.560 8.540 1311.820 8.800 ;
        RECT 2164.860 7.860 2165.120 8.120 ;
        RECT 1527.760 7.520 1528.020 7.780 ;
        RECT 1249.460 7.180 1249.720 7.440 ;
        RECT 1253.600 7.180 1253.860 7.440 ;
        RECT 919.640 5.820 919.900 6.080 ;
        RECT 947.240 5.820 947.500 6.080 ;
        RECT 771.060 5.480 771.320 5.740 ;
        RECT 1237.500 5.140 1237.760 5.400 ;
        RECT 1241.180 5.140 1241.440 5.400 ;
        RECT 1550.300 4.120 1550.560 4.380 ;
        RECT 767.380 3.780 767.640 4.040 ;
        RECT 1260.040 3.100 1260.300 3.360 ;
        RECT 1448.640 3.100 1448.900 3.360 ;
      LAYER met2 ;
        RECT 1311.560 8.740 1311.820 8.830 ;
        RECT 1311.560 8.600 1312.680 8.740 ;
        RECT 1311.560 8.510 1311.820 8.600 ;
        RECT 832.300 7.580 833.820 7.720 ;
        RECT 771.060 5.680 771.320 5.770 ;
        RECT 771.060 5.540 783.220 5.680 ;
        RECT 771.060 5.450 771.320 5.540 ;
        RECT 766.910 5.170 767.190 5.285 ;
        RECT 766.910 5.030 767.580 5.170 ;
        RECT 766.910 4.915 767.190 5.030 ;
        RECT 279.770 4.235 280.050 4.605 ;
        RECT 258.220 2.990 259.280 3.130 ;
        RECT 258.220 2.400 258.360 2.990 ;
        RECT 258.010 -4.800 258.570 2.400 ;
        RECT 259.140 1.205 259.280 2.990 ;
        RECT 279.840 1.205 279.980 4.235 ;
        RECT 767.440 4.070 767.580 5.030 ;
        RECT 783.080 4.660 783.220 5.540 ;
        RECT 832.300 5.340 832.440 7.580 ;
        RECT 818.500 5.285 832.440 5.340 ;
        RECT 786.230 5.170 786.510 5.285 ;
        RECT 785.840 5.030 786.510 5.170 ;
        RECT 785.840 4.660 785.980 5.030 ;
        RECT 786.230 4.915 786.510 5.030 ;
        RECT 818.430 5.200 832.440 5.285 ;
        RECT 818.430 4.915 818.710 5.200 ;
        RECT 833.680 5.170 833.820 7.580 ;
        RECT 1249.460 7.210 1249.720 7.470 ;
        RECT 1245.840 7.150 1249.720 7.210 ;
        RECT 1253.600 7.150 1253.860 7.470 ;
        RECT 1245.840 7.070 1249.660 7.150 ;
        RECT 919.640 5.790 919.900 6.110 ;
        RECT 947.240 5.790 947.500 6.110 ;
        RECT 919.700 5.285 919.840 5.790 ;
        RECT 834.070 5.170 834.350 5.285 ;
        RECT 833.680 5.030 834.350 5.170 ;
        RECT 834.070 4.915 834.350 5.030 ;
        RECT 919.630 4.915 919.910 5.285 ;
        RECT 947.300 5.170 947.440 5.790 ;
        RECT 990.470 5.595 990.750 5.965 ;
        RECT 949.530 5.170 949.810 5.285 ;
        RECT 947.300 5.030 949.810 5.170 ;
        RECT 990.540 5.170 990.680 5.595 ;
        RECT 991.850 5.170 992.130 5.285 ;
        RECT 990.540 5.030 992.130 5.170 ;
        RECT 949.530 4.915 949.810 5.030 ;
        RECT 991.850 4.915 992.130 5.030 ;
        RECT 1237.030 5.170 1237.310 5.285 ;
        RECT 1237.500 5.170 1237.760 5.430 ;
        RECT 1237.030 5.110 1237.760 5.170 ;
        RECT 1241.180 5.340 1241.440 5.430 ;
        RECT 1245.840 5.340 1245.980 7.070 ;
        RECT 1241.180 5.200 1245.980 5.340 ;
        RECT 1253.660 5.285 1253.800 7.150 ;
        RECT 1312.540 5.285 1312.680 8.600 ;
        RECT 1529.130 7.890 1529.410 8.005 ;
        RECT 1527.760 7.490 1528.020 7.810 ;
        RECT 1528.740 7.750 1529.410 7.890 ;
        RECT 1527.820 7.210 1527.960 7.490 ;
        RECT 1528.740 7.210 1528.880 7.750 ;
        RECT 1529.130 7.635 1529.410 7.750 ;
        RECT 1535.110 7.635 1535.390 8.005 ;
        RECT 2164.860 7.890 2165.120 8.150 ;
        RECT 2166.170 7.890 2166.450 9.000 ;
        RECT 2164.860 7.830 2166.450 7.890 ;
        RECT 2164.920 7.750 2166.450 7.830 ;
        RECT 1527.820 7.070 1528.880 7.210 ;
        RECT 1438.970 5.850 1439.250 5.965 ;
        RECT 1438.120 5.710 1439.250 5.850 ;
        RECT 1241.180 5.110 1241.440 5.200 ;
        RECT 1237.030 5.030 1237.700 5.110 ;
        RECT 1237.030 4.915 1237.310 5.030 ;
        RECT 1253.590 4.915 1253.870 5.285 ;
        RECT 1258.190 4.915 1258.470 5.285 ;
        RECT 1312.470 4.915 1312.750 5.285 ;
        RECT 1428.390 5.170 1428.670 5.285 ;
        RECT 1428.390 5.030 1431.820 5.170 ;
        RECT 1428.390 4.915 1428.670 5.030 ;
        RECT 783.080 4.520 785.980 4.660 ;
        RECT 1258.260 4.490 1258.400 4.915 ;
        RECT 1258.260 4.350 1260.240 4.490 ;
        RECT 767.380 3.750 767.640 4.070 ;
        RECT 1260.100 3.390 1260.240 4.350 ;
        RECT 1431.680 3.810 1431.820 5.030 ;
        RECT 1438.120 3.810 1438.260 5.710 ;
        RECT 1438.970 5.595 1439.250 5.710 ;
        RECT 1447.710 5.595 1447.990 5.965 ;
        RECT 1431.680 3.670 1438.260 3.810 ;
        RECT 1447.780 3.810 1447.920 5.595 ;
        RECT 1535.180 5.170 1535.320 7.635 ;
        RECT 1535.570 5.170 1535.850 5.285 ;
        RECT 1535.180 5.030 1535.850 5.170 ;
        RECT 1535.570 4.915 1535.850 5.030 ;
        RECT 1546.610 4.915 1546.890 5.285 ;
        RECT 2166.170 5.000 2166.450 7.750 ;
        RECT 1546.680 3.810 1546.820 4.915 ;
        RECT 1550.300 4.090 1550.560 4.410 ;
        RECT 1550.360 3.810 1550.500 4.090 ;
        RECT 1447.780 3.670 1448.840 3.810 ;
        RECT 1546.680 3.670 1550.500 3.810 ;
        RECT 1448.700 3.390 1448.840 3.670 ;
        RECT 1260.040 3.070 1260.300 3.390 ;
        RECT 1448.640 3.070 1448.900 3.390 ;
        RECT 259.070 0.835 259.350 1.205 ;
        RECT 279.770 0.835 280.050 1.205 ;
      LAYER via2 ;
        RECT 766.910 4.960 767.190 5.240 ;
        RECT 279.770 4.280 280.050 4.560 ;
        RECT 786.230 4.960 786.510 5.240 ;
        RECT 818.430 4.960 818.710 5.240 ;
        RECT 834.070 4.960 834.350 5.240 ;
        RECT 919.630 4.960 919.910 5.240 ;
        RECT 990.470 5.640 990.750 5.920 ;
        RECT 949.530 4.960 949.810 5.240 ;
        RECT 991.850 4.960 992.130 5.240 ;
        RECT 1237.030 4.960 1237.310 5.240 ;
        RECT 1529.130 7.680 1529.410 7.960 ;
        RECT 1535.110 7.680 1535.390 7.960 ;
        RECT 1253.590 4.960 1253.870 5.240 ;
        RECT 1258.190 4.960 1258.470 5.240 ;
        RECT 1312.470 4.960 1312.750 5.240 ;
        RECT 1428.390 4.960 1428.670 5.240 ;
        RECT 1438.970 5.640 1439.250 5.920 ;
        RECT 1447.710 5.640 1447.990 5.920 ;
        RECT 1535.570 4.960 1535.850 5.240 ;
        RECT 1546.610 4.960 1546.890 5.240 ;
        RECT 259.070 0.880 259.350 1.160 ;
        RECT 279.770 0.880 280.050 1.160 ;
      LAYER met3 ;
        RECT 1529.105 7.970 1529.435 7.985 ;
        RECT 1535.085 7.970 1535.415 7.985 ;
        RECT 1529.105 7.670 1535.415 7.970 ;
        RECT 1529.105 7.655 1529.435 7.670 ;
        RECT 1535.085 7.655 1535.415 7.670 ;
        RECT 957.070 5.930 957.450 5.940 ;
        RECT 678.350 5.630 696.130 5.930 ;
        RECT 279.745 4.570 280.075 4.585 ;
        RECT 411.510 4.570 411.890 4.580 ;
        RECT 279.745 4.270 411.890 4.570 ;
        RECT 279.745 4.255 280.075 4.270 ;
        RECT 411.510 4.260 411.890 4.270 ;
        RECT 413.350 4.570 413.730 4.580 ;
        RECT 456.590 4.570 456.970 4.580 ;
        RECT 413.350 4.270 456.970 4.570 ;
        RECT 413.350 4.260 413.730 4.270 ;
        RECT 456.590 4.260 456.970 4.270 ;
        RECT 461.190 4.570 461.570 4.580 ;
        RECT 647.950 4.570 648.330 4.580 ;
        RECT 461.190 4.270 648.330 4.570 ;
        RECT 461.190 4.260 461.570 4.270 ;
        RECT 647.950 4.260 648.330 4.270 ;
        RECT 649.790 4.570 650.170 4.580 ;
        RECT 678.350 4.570 678.650 5.630 ;
        RECT 695.830 5.250 696.130 5.630 ;
        RECT 956.190 5.630 957.450 5.930 ;
        RECT 766.885 5.250 767.215 5.265 ;
        RECT 695.830 4.950 767.215 5.250 ;
        RECT 766.885 4.935 767.215 4.950 ;
        RECT 786.205 5.250 786.535 5.265 ;
        RECT 818.405 5.250 818.735 5.265 ;
        RECT 786.205 4.950 818.735 5.250 ;
        RECT 786.205 4.935 786.535 4.950 ;
        RECT 818.405 4.935 818.735 4.950 ;
        RECT 834.045 5.250 834.375 5.265 ;
        RECT 919.605 5.250 919.935 5.265 ;
        RECT 834.045 4.950 919.935 5.250 ;
        RECT 834.045 4.935 834.375 4.950 ;
        RECT 919.605 4.935 919.935 4.950 ;
        RECT 949.505 5.250 949.835 5.265 ;
        RECT 956.190 5.250 956.490 5.630 ;
        RECT 957.070 5.620 957.450 5.630 ;
        RECT 984.670 5.930 985.050 5.940 ;
        RECT 990.445 5.930 990.775 5.945 ;
        RECT 984.670 5.630 990.775 5.930 ;
        RECT 984.670 5.620 985.050 5.630 ;
        RECT 990.445 5.615 990.775 5.630 ;
        RECT 1438.945 5.930 1439.275 5.945 ;
        RECT 1447.685 5.930 1448.015 5.945 ;
        RECT 1438.945 5.630 1448.015 5.930 ;
        RECT 1438.945 5.615 1439.275 5.630 ;
        RECT 1447.685 5.615 1448.015 5.630 ;
        RECT 949.505 4.950 956.490 5.250 ;
        RECT 991.825 5.250 992.155 5.265 ;
        RECT 1237.005 5.250 1237.335 5.265 ;
        RECT 991.825 4.950 1237.335 5.250 ;
        RECT 949.505 4.935 949.835 4.950 ;
        RECT 991.825 4.935 992.155 4.950 ;
        RECT 1237.005 4.935 1237.335 4.950 ;
        RECT 1253.565 5.250 1253.895 5.265 ;
        RECT 1258.165 5.250 1258.495 5.265 ;
        RECT 1253.565 4.950 1258.495 5.250 ;
        RECT 1253.565 4.935 1253.895 4.950 ;
        RECT 1258.165 4.935 1258.495 4.950 ;
        RECT 1312.445 5.250 1312.775 5.265 ;
        RECT 1428.365 5.250 1428.695 5.265 ;
        RECT 1312.445 4.950 1428.695 5.250 ;
        RECT 1312.445 4.935 1312.775 4.950 ;
        RECT 1428.365 4.935 1428.695 4.950 ;
        RECT 1535.545 5.250 1535.875 5.265 ;
        RECT 1546.585 5.250 1546.915 5.265 ;
        RECT 1535.545 4.950 1546.915 5.250 ;
        RECT 1535.545 4.935 1535.875 4.950 ;
        RECT 1546.585 4.935 1546.915 4.950 ;
        RECT 649.790 4.270 678.650 4.570 ;
        RECT 649.790 4.260 650.170 4.270 ;
        RECT 259.045 1.170 259.375 1.185 ;
        RECT 279.745 1.170 280.075 1.185 ;
        RECT 259.045 0.870 280.075 1.170 ;
        RECT 259.045 0.855 259.375 0.870 ;
        RECT 279.745 0.855 280.075 0.870 ;
      LAYER via3 ;
        RECT 411.540 4.260 411.860 4.580 ;
        RECT 413.380 4.260 413.700 4.580 ;
        RECT 456.620 4.260 456.940 4.580 ;
        RECT 461.220 4.260 461.540 4.580 ;
        RECT 647.980 4.260 648.300 4.580 ;
        RECT 649.820 4.260 650.140 4.580 ;
        RECT 957.100 5.620 957.420 5.940 ;
        RECT 984.700 5.620 985.020 5.940 ;
      LAYER met4 ;
        RECT 456.630 6.310 461.530 6.610 ;
        RECT 411.550 4.950 413.690 5.250 ;
        RECT 411.550 4.585 411.850 4.950 ;
        RECT 413.390 4.585 413.690 4.950 ;
        RECT 456.630 4.585 456.930 6.310 ;
        RECT 461.230 4.585 461.530 6.310 ;
        RECT 957.095 5.930 957.425 5.945 ;
        RECT 984.695 5.930 985.025 5.945 ;
        RECT 957.095 5.630 985.025 5.930 ;
        RECT 957.095 5.615 957.425 5.630 ;
        RECT 984.695 5.615 985.025 5.630 ;
        RECT 411.535 4.255 411.865 4.585 ;
        RECT 413.375 4.255 413.705 4.585 ;
        RECT 456.615 4.255 456.945 4.585 ;
        RECT 461.215 4.255 461.545 4.585 ;
        RECT 647.975 4.570 648.305 4.585 ;
        RECT 649.815 4.570 650.145 4.585 ;
        RECT 647.975 4.270 650.145 4.570 ;
        RECT 647.975 4.255 648.305 4.270 ;
        RECT 649.815 4.255 650.145 4.270 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1824.045 3397.705 1824.215 3401.615 ;
        RECT 1851.185 3397.705 1851.355 3401.615 ;
        RECT 1900.405 3397.705 1900.575 3401.955 ;
        RECT 1973.545 3397.705 1973.715 3401.955 ;
        RECT 2015.865 3397.705 2016.035 3401.955 ;
        RECT 2063.705 3397.705 2063.875 3401.955 ;
        RECT 2093.145 3397.705 2093.315 3401.955 ;
        RECT 2140.985 3397.705 2141.155 3401.955 ;
        RECT 2188.825 3397.705 2188.995 3401.955 ;
        RECT 2256.905 3397.705 2257.075 3401.955 ;
        RECT 2285.885 3397.705 2286.055 3401.955 ;
        RECT 2332.805 3397.705 2332.975 3401.955 ;
        RECT 2405.945 3397.705 2406.115 3401.615 ;
        RECT 2428.945 3397.705 2429.115 3401.615 ;
        RECT 2477.245 3397.705 2477.415 3401.955 ;
        RECT 2529.685 3397.705 2529.855 3401.955 ;
        RECT 2577.065 3397.705 2577.235 3401.955 ;
        RECT 2622.145 3397.705 2622.315 3401.955 ;
        RECT 2671.825 3397.705 2671.995 3401.955 ;
        RECT 2720.125 3397.705 2720.295 3401.955 ;
        RECT 742.125 9.605 757.935 9.775 ;
        RECT 742.125 8.585 742.295 9.605 ;
        RECT 757.765 8.755 757.935 9.605 ;
        RECT 784.445 9.265 789.215 9.435 ;
        RECT 758.685 8.925 760.695 9.095 ;
        RECT 758.685 8.755 758.855 8.925 ;
        RECT 757.765 8.585 758.855 8.755 ;
        RECT 760.525 8.585 760.695 8.925 ;
        RECT 782.605 7.565 782.775 9.095 ;
        RECT 784.445 7.565 784.615 9.265 ;
        RECT 789.045 8.585 789.215 9.265 ;
        RECT 374.125 6.715 374.295 7.055 ;
        RECT 513.505 6.885 518.275 7.055 ;
        RECT 374.125 6.545 375.215 6.715 ;
        RECT 510.745 6.205 512.295 6.375 ;
        RECT 513.505 6.205 513.675 6.885 ;
        RECT 510.745 6.035 510.915 6.205 ;
        RECT 487.745 5.865 510.915 6.035 ;
        RECT 487.745 3.995 487.915 5.865 ;
        RECT 518.105 5.355 518.275 6.885 ;
        RECT 519.025 5.525 520.575 5.695 ;
        RECT 519.025 5.355 519.195 5.525 ;
        RECT 518.105 5.185 519.195 5.355 ;
        RECT 482.685 3.825 487.915 3.995 ;
        RECT 482.685 2.975 482.855 3.825 ;
        RECT 470.725 2.805 482.855 2.975 ;
        RECT 553.525 0.595 553.695 7.395 ;
        RECT 1197.525 6.205 1198.155 6.375 ;
        RECT 1193.845 5.865 1194.475 6.035 ;
        RECT 1194.305 3.995 1194.475 5.865 ;
        RECT 1197.525 3.995 1197.695 6.205 ;
        RECT 1194.305 3.825 1197.695 3.995 ;
        RECT 1396.705 3.825 1398.255 3.995 ;
        RECT 1396.705 3.485 1396.875 3.825 ;
        RECT 1398.085 3.315 1398.255 3.825 ;
        RECT 1399.005 3.315 1399.175 3.655 ;
        RECT 1398.085 3.145 1399.175 3.315 ;
        RECT 1407.285 3.315 1407.455 3.655 ;
        RECT 1407.285 3.145 1408.375 3.315 ;
        RECT 559.505 0.595 559.675 0.935 ;
        RECT 553.525 0.425 559.675 0.595 ;
      LAYER mcon ;
        RECT 1900.405 3401.785 1900.575 3401.955 ;
        RECT 1824.045 3401.445 1824.215 3401.615 ;
        RECT 1851.185 3401.445 1851.355 3401.615 ;
        RECT 1973.545 3401.785 1973.715 3401.955 ;
        RECT 2015.865 3401.785 2016.035 3401.955 ;
        RECT 2063.705 3401.785 2063.875 3401.955 ;
        RECT 2093.145 3401.785 2093.315 3401.955 ;
        RECT 2140.985 3401.785 2141.155 3401.955 ;
        RECT 2188.825 3401.785 2188.995 3401.955 ;
        RECT 2256.905 3401.785 2257.075 3401.955 ;
        RECT 2285.885 3401.785 2286.055 3401.955 ;
        RECT 2332.805 3401.785 2332.975 3401.955 ;
        RECT 2477.245 3401.785 2477.415 3401.955 ;
        RECT 2405.945 3401.445 2406.115 3401.615 ;
        RECT 2428.945 3401.445 2429.115 3401.615 ;
        RECT 2529.685 3401.785 2529.855 3401.955 ;
        RECT 2577.065 3401.785 2577.235 3401.955 ;
        RECT 2622.145 3401.785 2622.315 3401.955 ;
        RECT 2671.825 3401.785 2671.995 3401.955 ;
        RECT 2720.125 3401.785 2720.295 3401.955 ;
        RECT 782.605 8.925 782.775 9.095 ;
        RECT 553.525 7.225 553.695 7.395 ;
        RECT 374.125 6.885 374.295 7.055 ;
        RECT 375.045 6.545 375.215 6.715 ;
        RECT 512.125 6.205 512.295 6.375 ;
        RECT 520.405 5.525 520.575 5.695 ;
        RECT 1197.985 6.205 1198.155 6.375 ;
        RECT 1399.005 3.485 1399.175 3.655 ;
        RECT 1407.285 3.485 1407.455 3.655 ;
        RECT 1408.205 3.145 1408.375 3.315 ;
        RECT 559.505 0.765 559.675 0.935 ;
      LAYER met1 ;
        RECT 1429.750 3416.220 1430.070 3416.280 ;
        RECT 1476.210 3416.220 1476.530 3416.280 ;
        RECT 1429.750 3416.080 1476.530 3416.220 ;
        RECT 1429.750 3416.020 1430.070 3416.080 ;
        RECT 1476.210 3416.020 1476.530 3416.080 ;
        RECT 2787.210 3402.960 2787.530 3403.020 ;
        RECT 2816.190 3402.960 2816.510 3403.020 ;
        RECT 2787.210 3402.820 2816.510 3402.960 ;
        RECT 2787.210 3402.760 2787.530 3402.820 ;
        RECT 2816.190 3402.760 2816.510 3402.820 ;
        RECT 1900.330 3401.940 1900.650 3402.000 ;
        RECT 1973.470 3401.940 1973.790 3402.000 ;
        RECT 2015.790 3401.940 2016.110 3402.000 ;
        RECT 2063.630 3401.940 2063.950 3402.000 ;
        RECT 2093.070 3401.940 2093.390 3402.000 ;
        RECT 2140.910 3401.940 2141.230 3402.000 ;
        RECT 2188.750 3401.940 2189.070 3402.000 ;
        RECT 2256.830 3401.940 2257.150 3402.000 ;
        RECT 2285.810 3401.940 2286.130 3402.000 ;
        RECT 2332.730 3401.940 2333.050 3402.000 ;
        RECT 1900.135 3401.800 1900.650 3401.940 ;
        RECT 1973.275 3401.800 1973.790 3401.940 ;
        RECT 2015.595 3401.800 2016.110 3401.940 ;
        RECT 2063.435 3401.800 2063.950 3401.940 ;
        RECT 2092.875 3401.800 2093.390 3401.940 ;
        RECT 2140.715 3401.800 2141.230 3401.940 ;
        RECT 2188.555 3401.800 2189.070 3401.940 ;
        RECT 2256.635 3401.800 2257.150 3401.940 ;
        RECT 2285.615 3401.800 2286.130 3401.940 ;
        RECT 2332.535 3401.800 2333.050 3401.940 ;
        RECT 1900.330 3401.740 1900.650 3401.800 ;
        RECT 1973.470 3401.740 1973.790 3401.800 ;
        RECT 2015.790 3401.740 2016.110 3401.800 ;
        RECT 2063.630 3401.740 2063.950 3401.800 ;
        RECT 2093.070 3401.740 2093.390 3401.800 ;
        RECT 2140.910 3401.740 2141.230 3401.800 ;
        RECT 2188.750 3401.740 2189.070 3401.800 ;
        RECT 2256.830 3401.740 2257.150 3401.800 ;
        RECT 2285.810 3401.740 2286.130 3401.800 ;
        RECT 2332.730 3401.740 2333.050 3401.800 ;
        RECT 2477.170 3401.940 2477.490 3402.000 ;
        RECT 2529.610 3401.940 2529.930 3402.000 ;
        RECT 2576.990 3401.940 2577.310 3402.000 ;
        RECT 2477.170 3401.800 2477.685 3401.940 ;
        RECT 2529.415 3401.800 2529.930 3401.940 ;
        RECT 2576.795 3401.800 2577.310 3401.940 ;
        RECT 2477.170 3401.740 2477.490 3401.800 ;
        RECT 2529.610 3401.740 2529.930 3401.800 ;
        RECT 2576.990 3401.740 2577.310 3401.800 ;
        RECT 2622.070 3401.940 2622.390 3402.000 ;
        RECT 2671.750 3401.940 2672.070 3402.000 ;
        RECT 2720.050 3401.940 2720.370 3402.000 ;
        RECT 2622.070 3401.800 2622.585 3401.940 ;
        RECT 2671.555 3401.800 2672.070 3401.940 ;
        RECT 2719.855 3401.800 2720.370 3401.940 ;
        RECT 2622.070 3401.740 2622.390 3401.800 ;
        RECT 2671.750 3401.740 2672.070 3401.800 ;
        RECT 2720.050 3401.740 2720.370 3401.800 ;
        RECT 1476.210 3401.600 1476.530 3401.660 ;
        RECT 1483.570 3401.600 1483.890 3401.660 ;
        RECT 1823.970 3401.600 1824.290 3401.660 ;
        RECT 1851.110 3401.600 1851.430 3401.660 ;
        RECT 2405.870 3401.600 2406.190 3401.660 ;
        RECT 1476.210 3401.460 1483.890 3401.600 ;
        RECT 1823.775 3401.460 1824.290 3401.600 ;
        RECT 1850.915 3401.460 1851.430 3401.600 ;
        RECT 2405.675 3401.460 2406.190 3401.600 ;
        RECT 1476.210 3401.400 1476.530 3401.460 ;
        RECT 1483.570 3401.400 1483.890 3401.460 ;
        RECT 1823.970 3401.400 1824.290 3401.460 ;
        RECT 1851.110 3401.400 1851.430 3401.460 ;
        RECT 2405.870 3401.400 2406.190 3401.460 ;
        RECT 2428.870 3401.600 2429.190 3401.660 ;
        RECT 2428.870 3401.460 2429.385 3401.600 ;
        RECT 2428.870 3401.400 2429.190 3401.460 ;
        RECT 1823.985 3397.860 1824.275 3397.905 ;
        RECT 1851.125 3397.860 1851.415 3397.905 ;
        RECT 1823.985 3397.720 1851.415 3397.860 ;
        RECT 1823.985 3397.675 1824.275 3397.720 ;
        RECT 1851.125 3397.675 1851.415 3397.720 ;
        RECT 1900.345 3397.860 1900.635 3397.905 ;
        RECT 1973.485 3397.860 1973.775 3397.905 ;
        RECT 1900.345 3397.720 1973.775 3397.860 ;
        RECT 1900.345 3397.675 1900.635 3397.720 ;
        RECT 1973.485 3397.675 1973.775 3397.720 ;
        RECT 2015.805 3397.860 2016.095 3397.905 ;
        RECT 2063.645 3397.860 2063.935 3397.905 ;
        RECT 2015.805 3397.720 2063.935 3397.860 ;
        RECT 2015.805 3397.675 2016.095 3397.720 ;
        RECT 2063.645 3397.675 2063.935 3397.720 ;
        RECT 2093.085 3397.860 2093.375 3397.905 ;
        RECT 2140.925 3397.860 2141.215 3397.905 ;
        RECT 2093.085 3397.720 2141.215 3397.860 ;
        RECT 2093.085 3397.675 2093.375 3397.720 ;
        RECT 2140.925 3397.675 2141.215 3397.720 ;
        RECT 2188.765 3397.860 2189.055 3397.905 ;
        RECT 2256.845 3397.860 2257.135 3397.905 ;
        RECT 2188.765 3397.720 2257.135 3397.860 ;
        RECT 2188.765 3397.675 2189.055 3397.720 ;
        RECT 2256.845 3397.675 2257.135 3397.720 ;
        RECT 2285.825 3397.860 2286.115 3397.905 ;
        RECT 2332.745 3397.860 2333.035 3397.905 ;
        RECT 2285.825 3397.720 2333.035 3397.860 ;
        RECT 2285.825 3397.675 2286.115 3397.720 ;
        RECT 2332.745 3397.675 2333.035 3397.720 ;
        RECT 2405.885 3397.860 2406.175 3397.905 ;
        RECT 2428.885 3397.860 2429.175 3397.905 ;
        RECT 2405.885 3397.720 2429.175 3397.860 ;
        RECT 2405.885 3397.675 2406.175 3397.720 ;
        RECT 2428.885 3397.675 2429.175 3397.720 ;
        RECT 2477.185 3397.860 2477.475 3397.905 ;
        RECT 2529.625 3397.860 2529.915 3397.905 ;
        RECT 2477.185 3397.720 2529.915 3397.860 ;
        RECT 2477.185 3397.675 2477.475 3397.720 ;
        RECT 2529.625 3397.675 2529.915 3397.720 ;
        RECT 2577.005 3397.860 2577.295 3397.905 ;
        RECT 2622.085 3397.860 2622.375 3397.905 ;
        RECT 2577.005 3397.720 2622.375 3397.860 ;
        RECT 2577.005 3397.675 2577.295 3397.720 ;
        RECT 2622.085 3397.675 2622.375 3397.720 ;
        RECT 2671.765 3397.860 2672.055 3397.905 ;
        RECT 2720.065 3397.860 2720.355 3397.905 ;
        RECT 2671.765 3397.720 2720.355 3397.860 ;
        RECT 2671.765 3397.675 2672.055 3397.720 ;
        RECT 2720.065 3397.675 2720.355 3397.720 ;
        RECT 782.545 9.080 782.835 9.125 ;
        RECT 781.240 8.940 782.835 9.080 ;
        RECT 741.590 8.740 741.910 8.800 ;
        RECT 742.065 8.740 742.355 8.785 ;
        RECT 741.590 8.600 742.355 8.740 ;
        RECT 741.590 8.540 741.910 8.600 ;
        RECT 742.065 8.555 742.355 8.600 ;
        RECT 760.465 8.740 760.755 8.785 ;
        RECT 781.240 8.740 781.380 8.940 ;
        RECT 782.545 8.895 782.835 8.940 ;
        RECT 760.465 8.600 781.380 8.740 ;
        RECT 788.985 8.740 789.275 8.785 ;
        RECT 807.830 8.740 808.150 8.800 ;
        RECT 788.985 8.600 808.150 8.740 ;
        RECT 760.465 8.555 760.755 8.600 ;
        RECT 788.985 8.555 789.275 8.600 ;
        RECT 807.830 8.540 808.150 8.600 ;
        RECT 782.545 7.720 782.835 7.765 ;
        RECT 784.385 7.720 784.675 7.765 ;
        RECT 782.545 7.580 784.675 7.720 ;
        RECT 782.545 7.535 782.835 7.580 ;
        RECT 784.385 7.535 784.675 7.580 ;
        RECT 534.590 7.380 534.910 7.440 ;
        RECT 553.465 7.380 553.755 7.425 ;
        RECT 534.590 7.240 553.755 7.380 ;
        RECT 534.590 7.180 534.910 7.240 ;
        RECT 553.465 7.195 553.755 7.240 ;
        RECT 372.670 7.040 372.990 7.100 ;
        RECT 374.065 7.040 374.355 7.085 ;
        RECT 372.670 6.900 374.355 7.040 ;
        RECT 372.670 6.840 372.990 6.900 ;
        RECT 374.065 6.855 374.355 6.900 ;
        RECT 720.890 7.040 721.210 7.100 ;
        RECT 725.490 7.040 725.810 7.100 ;
        RECT 720.890 6.900 725.810 7.040 ;
        RECT 720.890 6.840 721.210 6.900 ;
        RECT 725.490 6.840 725.810 6.900 ;
        RECT 374.985 6.700 375.275 6.745 ;
        RECT 383.250 6.700 383.570 6.760 ;
        RECT 374.985 6.560 383.570 6.700 ;
        RECT 374.985 6.515 375.275 6.560 ;
        RECT 383.250 6.500 383.570 6.560 ;
        RECT 512.065 6.360 512.355 6.405 ;
        RECT 513.445 6.360 513.735 6.405 ;
        RECT 512.065 6.220 513.735 6.360 ;
        RECT 512.065 6.175 512.355 6.220 ;
        RECT 513.445 6.175 513.735 6.220 ;
        RECT 1197.925 6.360 1198.215 6.405 ;
        RECT 1198.830 6.360 1199.150 6.420 ;
        RECT 1197.925 6.220 1199.150 6.360 ;
        RECT 1197.925 6.175 1198.215 6.220 ;
        RECT 1198.830 6.160 1199.150 6.220 ;
        RECT 1192.850 6.020 1193.170 6.080 ;
        RECT 1193.785 6.020 1194.075 6.065 ;
        RECT 1192.850 5.880 1194.075 6.020 ;
        RECT 1192.850 5.820 1193.170 5.880 ;
        RECT 1193.785 5.835 1194.075 5.880 ;
        RECT 520.345 5.680 520.635 5.725 ;
        RECT 524.010 5.680 524.330 5.740 ;
        RECT 520.345 5.540 524.330 5.680 ;
        RECT 520.345 5.495 520.635 5.540 ;
        RECT 524.010 5.480 524.330 5.540 ;
        RECT 1089.810 5.680 1090.130 5.740 ;
        RECT 1118.790 5.680 1119.110 5.740 ;
        RECT 1089.810 5.540 1119.110 5.680 ;
        RECT 1089.810 5.480 1090.130 5.540 ;
        RECT 1118.790 5.480 1119.110 5.540 ;
        RECT 311.950 5.340 312.270 5.400 ;
        RECT 333.110 5.340 333.430 5.400 ;
        RECT 311.950 5.200 333.430 5.340 ;
        RECT 311.950 5.140 312.270 5.200 ;
        RECT 333.110 5.140 333.430 5.200 ;
        RECT 581.050 5.000 581.370 5.060 ;
        RECT 600.370 5.000 600.690 5.060 ;
        RECT 581.050 4.860 600.690 5.000 ;
        RECT 581.050 4.800 581.370 4.860 ;
        RECT 600.370 4.800 600.690 4.860 ;
        RECT 1597.650 5.000 1597.970 5.060 ;
        RECT 1638.590 5.000 1638.910 5.060 ;
        RECT 1597.650 4.860 1638.910 5.000 ;
        RECT 1597.650 4.800 1597.970 4.860 ;
        RECT 1638.590 4.800 1638.910 4.860 ;
        RECT 891.550 3.640 891.870 3.700 ;
        RECT 900.750 3.640 901.070 3.700 ;
        RECT 891.550 3.500 901.070 3.640 ;
        RECT 891.550 3.440 891.870 3.500 ;
        RECT 900.750 3.440 901.070 3.500 ;
        RECT 1366.730 3.640 1367.050 3.700 ;
        RECT 1396.645 3.640 1396.935 3.685 ;
        RECT 1366.730 3.500 1396.935 3.640 ;
        RECT 1366.730 3.440 1367.050 3.500 ;
        RECT 1396.645 3.455 1396.935 3.500 ;
        RECT 1398.945 3.640 1399.235 3.685 ;
        RECT 1407.225 3.640 1407.515 3.685 ;
        RECT 1398.945 3.500 1407.515 3.640 ;
        RECT 1398.945 3.455 1399.235 3.500 ;
        RECT 1407.225 3.455 1407.515 3.500 ;
        RECT 1122.930 3.300 1123.250 3.360 ;
        RECT 1126.610 3.300 1126.930 3.360 ;
        RECT 1122.930 3.160 1126.930 3.300 ;
        RECT 1122.930 3.100 1123.250 3.160 ;
        RECT 1126.610 3.100 1126.930 3.160 ;
        RECT 1408.145 3.300 1408.435 3.345 ;
        RECT 1430.210 3.300 1430.530 3.360 ;
        RECT 1408.145 3.160 1430.530 3.300 ;
        RECT 1408.145 3.115 1408.435 3.160 ;
        RECT 1430.210 3.100 1430.530 3.160 ;
        RECT 469.270 2.960 469.590 3.020 ;
        RECT 470.665 2.960 470.955 3.005 ;
        RECT 469.270 2.820 470.955 2.960 ;
        RECT 469.270 2.760 469.590 2.820 ;
        RECT 470.665 2.775 470.955 2.820 ;
        RECT 677.190 2.280 677.510 2.340 ;
        RECT 711.230 2.280 711.550 2.340 ;
        RECT 677.190 2.140 711.550 2.280 ;
        RECT 677.190 2.080 677.510 2.140 ;
        RECT 711.230 2.080 711.550 2.140 ;
        RECT 559.445 0.920 559.735 0.965 ;
        RECT 560.810 0.920 561.130 0.980 ;
        RECT 559.445 0.780 561.130 0.920 ;
        RECT 559.445 0.735 559.735 0.780 ;
        RECT 560.810 0.720 561.130 0.780 ;
      LAYER via ;
        RECT 1429.780 3416.020 1430.040 3416.280 ;
        RECT 1476.240 3416.020 1476.500 3416.280 ;
        RECT 2787.240 3402.760 2787.500 3403.020 ;
        RECT 2816.220 3402.760 2816.480 3403.020 ;
        RECT 1900.360 3401.740 1900.620 3402.000 ;
        RECT 1973.500 3401.740 1973.760 3402.000 ;
        RECT 2015.820 3401.740 2016.080 3402.000 ;
        RECT 2063.660 3401.740 2063.920 3402.000 ;
        RECT 2093.100 3401.740 2093.360 3402.000 ;
        RECT 2140.940 3401.740 2141.200 3402.000 ;
        RECT 2188.780 3401.740 2189.040 3402.000 ;
        RECT 2256.860 3401.740 2257.120 3402.000 ;
        RECT 2285.840 3401.740 2286.100 3402.000 ;
        RECT 2332.760 3401.740 2333.020 3402.000 ;
        RECT 2477.200 3401.740 2477.460 3402.000 ;
        RECT 2529.640 3401.740 2529.900 3402.000 ;
        RECT 2577.020 3401.740 2577.280 3402.000 ;
        RECT 2622.100 3401.740 2622.360 3402.000 ;
        RECT 2671.780 3401.740 2672.040 3402.000 ;
        RECT 2720.080 3401.740 2720.340 3402.000 ;
        RECT 1476.240 3401.400 1476.500 3401.660 ;
        RECT 1483.600 3401.400 1483.860 3401.660 ;
        RECT 1824.000 3401.400 1824.260 3401.660 ;
        RECT 1851.140 3401.400 1851.400 3401.660 ;
        RECT 2405.900 3401.400 2406.160 3401.660 ;
        RECT 2428.900 3401.400 2429.160 3401.660 ;
        RECT 741.620 8.540 741.880 8.800 ;
        RECT 807.860 8.540 808.120 8.800 ;
        RECT 534.620 7.180 534.880 7.440 ;
        RECT 372.700 6.840 372.960 7.100 ;
        RECT 720.920 6.840 721.180 7.100 ;
        RECT 725.520 6.840 725.780 7.100 ;
        RECT 383.280 6.500 383.540 6.760 ;
        RECT 1198.860 6.160 1199.120 6.420 ;
        RECT 1192.880 5.820 1193.140 6.080 ;
        RECT 524.040 5.480 524.300 5.740 ;
        RECT 1089.840 5.480 1090.100 5.740 ;
        RECT 1118.820 5.480 1119.080 5.740 ;
        RECT 311.980 5.140 312.240 5.400 ;
        RECT 333.140 5.140 333.400 5.400 ;
        RECT 581.080 4.800 581.340 5.060 ;
        RECT 600.400 4.800 600.660 5.060 ;
        RECT 1597.680 4.800 1597.940 5.060 ;
        RECT 1638.620 4.800 1638.880 5.060 ;
        RECT 891.580 3.440 891.840 3.700 ;
        RECT 900.780 3.440 901.040 3.700 ;
        RECT 1366.760 3.440 1367.020 3.700 ;
        RECT 1122.960 3.100 1123.220 3.360 ;
        RECT 1126.640 3.100 1126.900 3.360 ;
        RECT 1430.240 3.100 1430.500 3.360 ;
        RECT 469.300 2.760 469.560 3.020 ;
        RECT 677.220 2.080 677.480 2.340 ;
        RECT 711.260 2.080 711.520 2.340 ;
        RECT 560.840 0.720 561.100 0.980 ;
      LAYER met2 ;
        RECT 1429.780 3415.990 1430.040 3416.310 ;
        RECT 1476.240 3415.990 1476.500 3416.310 ;
        RECT 1429.840 3405.000 1429.980 3415.990 ;
        RECT 1429.710 3401.000 1429.990 3405.000 ;
        RECT 1476.300 3401.690 1476.440 3415.990 ;
        RECT 2787.230 3402.875 2787.510 3403.245 ;
        RECT 2787.240 3402.730 2787.500 3402.875 ;
        RECT 2816.220 3402.730 2816.480 3403.050 ;
        RECT 2816.280 3402.565 2816.420 3402.730 ;
        RECT 2816.210 3402.195 2816.490 3402.565 ;
        RECT 1900.360 3401.885 1900.620 3402.030 ;
        RECT 1973.500 3401.885 1973.760 3402.030 ;
        RECT 2015.820 3401.885 2016.080 3402.030 ;
        RECT 2063.660 3401.885 2063.920 3402.030 ;
        RECT 2093.100 3401.885 2093.360 3402.030 ;
        RECT 2140.940 3401.885 2141.200 3402.030 ;
        RECT 2188.780 3401.885 2189.040 3402.030 ;
        RECT 2256.860 3401.885 2257.120 3402.030 ;
        RECT 2285.840 3401.885 2286.100 3402.030 ;
        RECT 2332.760 3401.885 2333.020 3402.030 ;
        RECT 2477.200 3401.885 2477.460 3402.030 ;
        RECT 2529.640 3401.885 2529.900 3402.030 ;
        RECT 2577.020 3401.885 2577.280 3402.030 ;
        RECT 2622.100 3401.885 2622.360 3402.030 ;
        RECT 2671.780 3401.885 2672.040 3402.030 ;
        RECT 2720.080 3401.885 2720.340 3402.030 ;
        RECT 1476.240 3401.370 1476.500 3401.690 ;
        RECT 1483.590 3401.515 1483.870 3401.885 ;
        RECT 1823.990 3401.515 1824.270 3401.885 ;
        RECT 1851.130 3401.515 1851.410 3401.885 ;
        RECT 1900.350 3401.515 1900.630 3401.885 ;
        RECT 1973.490 3401.515 1973.770 3401.885 ;
        RECT 2015.810 3401.515 2016.090 3401.885 ;
        RECT 2063.650 3401.515 2063.930 3401.885 ;
        RECT 2093.090 3401.515 2093.370 3401.885 ;
        RECT 2140.930 3401.515 2141.210 3401.885 ;
        RECT 2188.770 3401.515 2189.050 3401.885 ;
        RECT 2256.850 3401.515 2257.130 3401.885 ;
        RECT 2285.830 3401.515 2286.110 3401.885 ;
        RECT 2332.750 3401.515 2333.030 3401.885 ;
        RECT 2405.890 3401.515 2406.170 3401.885 ;
        RECT 2428.890 3401.515 2429.170 3401.885 ;
        RECT 2477.190 3401.515 2477.470 3401.885 ;
        RECT 2529.630 3401.515 2529.910 3401.885 ;
        RECT 2577.010 3401.515 2577.290 3401.885 ;
        RECT 2622.090 3401.515 2622.370 3401.885 ;
        RECT 2671.770 3401.515 2672.050 3401.885 ;
        RECT 2720.070 3401.515 2720.350 3401.885 ;
        RECT 1483.600 3401.370 1483.860 3401.515 ;
        RECT 1824.000 3401.370 1824.260 3401.515 ;
        RECT 1851.140 3401.370 1851.400 3401.515 ;
        RECT 2405.900 3401.370 2406.160 3401.515 ;
        RECT 2428.900 3401.370 2429.160 3401.515 ;
        RECT 600.460 8.260 601.520 8.400 ;
        RECT 577.460 7.750 580.820 7.890 ;
        RECT 371.380 7.580 372.900 7.720 ;
        RECT 335.430 7.210 335.710 7.325 ;
        RECT 335.040 7.070 335.710 7.210 ;
        RECT 311.980 5.110 312.240 5.430 ;
        RECT 333.140 5.110 333.400 5.430 ;
        RECT 312.040 2.400 312.180 5.110 ;
        RECT 333.200 4.490 333.340 5.110 ;
        RECT 335.040 4.490 335.180 7.070 ;
        RECT 335.430 6.955 335.710 7.070 ;
        RECT 371.380 5.285 371.520 7.580 ;
        RECT 372.760 7.130 372.900 7.580 ;
        RECT 534.620 7.150 534.880 7.470 ;
        RECT 372.700 6.810 372.960 7.130 ;
        RECT 383.280 6.530 383.540 6.790 ;
        RECT 383.280 6.470 391.300 6.530 ;
        RECT 383.340 6.390 391.300 6.470 ;
        RECT 371.310 4.915 371.590 5.285 ;
        RECT 333.200 4.350 335.180 4.490 ;
        RECT 311.830 -4.800 312.390 2.400 ;
        RECT 391.160 1.205 391.300 6.390 ;
        RECT 524.030 5.595 524.310 5.965 ;
        RECT 534.150 5.850 534.430 5.965 ;
        RECT 534.680 5.850 534.820 7.150 ;
        RECT 534.150 5.710 534.820 5.850 ;
        RECT 534.150 5.595 534.430 5.710 ;
        RECT 524.040 5.450 524.300 5.595 ;
        RECT 577.460 5.000 577.600 7.750 ;
        RECT 580.680 7.380 580.820 7.750 ;
        RECT 580.680 7.240 581.280 7.380 ;
        RECT 581.140 5.090 581.280 7.240 ;
        RECT 600.460 5.090 600.600 8.260 ;
        RECT 601.380 7.890 601.520 8.260 ;
        RECT 713.160 8.260 715.140 8.400 ;
        RECT 725.510 8.315 725.790 8.685 ;
        RECT 728.270 8.315 728.550 8.685 ;
        RECT 741.620 8.510 741.880 8.830 ;
        RECT 807.860 8.740 808.120 8.830 ;
        RECT 807.860 8.600 831.980 8.740 ;
        RECT 807.860 8.510 808.120 8.600 ;
        RECT 601.380 7.750 606.580 7.890 ;
        RECT 606.440 5.850 606.580 7.750 ;
        RECT 610.050 6.530 610.330 6.645 ;
        RECT 609.660 6.390 610.330 6.530 ;
        RECT 609.660 5.850 609.800 6.390 ;
        RECT 610.050 6.275 610.330 6.390 ;
        RECT 656.510 6.275 656.790 6.645 ;
        RECT 606.440 5.710 609.800 5.850 ;
        RECT 561.360 4.860 577.600 5.000 ;
        RECT 412.250 4.490 412.530 4.605 ;
        RECT 410.940 4.350 412.530 4.490 ;
        RECT 410.940 1.205 411.080 4.350 ;
        RECT 412.250 4.235 412.530 4.350 ;
        RECT 469.300 2.730 469.560 3.050 ;
        RECT 561.360 2.960 561.500 4.860 ;
        RECT 581.080 4.770 581.340 5.090 ;
        RECT 600.400 4.770 600.660 5.090 ;
        RECT 656.580 3.810 656.720 6.275 ;
        RECT 656.580 3.670 676.040 3.810 ;
        RECT 560.900 2.820 561.500 2.960 ;
        RECT 391.090 0.835 391.370 1.205 ;
        RECT 410.870 0.835 411.150 1.205 ;
        RECT 469.360 0.525 469.500 2.730 ;
        RECT 560.900 1.010 561.040 2.820 ;
        RECT 675.900 2.280 676.040 3.670 ;
        RECT 677.220 2.280 677.480 2.370 ;
        RECT 675.900 2.140 677.480 2.280 ;
        RECT 677.220 2.050 677.480 2.140 ;
        RECT 711.260 2.050 711.520 2.370 ;
        RECT 711.320 1.770 711.460 2.050 ;
        RECT 713.160 1.770 713.300 8.260 ;
        RECT 715.000 7.040 715.140 8.260 ;
        RECT 725.580 7.130 725.720 8.315 ;
        RECT 728.340 7.380 728.480 8.315 ;
        RECT 728.340 7.240 739.060 7.380 ;
        RECT 720.920 7.040 721.180 7.130 ;
        RECT 715.000 6.900 721.180 7.040 ;
        RECT 720.920 6.810 721.180 6.900 ;
        RECT 725.520 6.810 725.780 7.130 ;
        RECT 738.920 4.660 739.060 7.240 ;
        RECT 741.680 4.660 741.820 8.510 ;
        RECT 831.840 5.965 831.980 8.600 ;
        RECT 1227.370 8.570 1227.650 8.685 ;
        RECT 1474.850 8.570 1475.130 8.685 ;
        RECT 1226.980 8.430 1227.650 8.570 ;
        RECT 1200.760 7.750 1209.640 7.890 ;
        RECT 891.570 6.955 891.850 7.325 ;
        RECT 845.570 6.275 845.850 6.645 ;
        RECT 831.770 5.595 832.050 5.965 ;
        RECT 843.270 5.595 843.550 5.965 ;
        RECT 843.340 5.170 843.480 5.595 ;
        RECT 845.640 5.170 845.780 6.275 ;
        RECT 843.340 5.030 845.780 5.170 ;
        RECT 738.920 4.520 741.820 4.660 ;
        RECT 891.640 3.730 891.780 6.955 ;
        RECT 900.840 6.900 905.120 7.040 ;
        RECT 900.840 3.730 900.980 6.900 ;
        RECT 904.980 5.850 905.120 6.900 ;
        RECT 1089.830 6.275 1090.110 6.645 ;
        RECT 1191.560 6.390 1193.080 6.530 ;
        RECT 914.570 5.850 914.850 5.965 ;
        RECT 904.980 5.710 914.850 5.850 ;
        RECT 1089.900 5.770 1090.040 6.275 ;
        RECT 914.570 5.595 914.850 5.710 ;
        RECT 1089.840 5.450 1090.100 5.770 ;
        RECT 1118.820 5.450 1119.080 5.770 ;
        RECT 921.470 5.170 921.750 5.285 ;
        RECT 921.470 5.030 922.600 5.170 ;
        RECT 921.470 4.915 921.750 5.030 ;
        RECT 922.460 3.810 922.600 5.030 ;
        RECT 1118.880 4.490 1119.020 5.450 ;
        RECT 1118.880 4.350 1122.700 4.490 ;
        RECT 952.290 3.810 952.570 3.925 ;
        RECT 891.580 3.410 891.840 3.730 ;
        RECT 900.780 3.410 901.040 3.730 ;
        RECT 922.460 3.670 952.570 3.810 ;
        RECT 952.290 3.555 952.570 3.670 ;
        RECT 987.710 3.810 987.990 3.925 ;
        RECT 987.710 3.670 988.380 3.810 ;
        RECT 987.710 3.555 987.990 3.670 ;
        RECT 988.240 2.565 988.380 3.670 ;
        RECT 1122.560 3.300 1122.700 4.350 ;
        RECT 1156.530 3.810 1156.810 3.925 ;
        RECT 1126.700 3.670 1156.810 3.810 ;
        RECT 1126.700 3.390 1126.840 3.670 ;
        RECT 1156.530 3.555 1156.810 3.670 ;
        RECT 1191.030 3.810 1191.310 3.925 ;
        RECT 1191.560 3.810 1191.700 6.390 ;
        RECT 1192.940 6.110 1193.080 6.390 ;
        RECT 1198.860 6.130 1199.120 6.450 ;
        RECT 1192.880 5.790 1193.140 6.110 ;
        RECT 1198.920 5.170 1199.060 6.130 ;
        RECT 1200.760 5.170 1200.900 7.750 ;
        RECT 1198.920 5.030 1200.900 5.170 ;
        RECT 1209.500 4.490 1209.640 7.750 ;
        RECT 1226.980 5.340 1227.120 8.430 ;
        RECT 1227.370 8.315 1227.650 8.430 ;
        RECT 1473.540 8.430 1475.130 8.570 ;
        RECT 1473.540 6.645 1473.680 8.430 ;
        RECT 1474.850 8.315 1475.130 8.430 ;
        RECT 1597.670 7.635 1597.950 8.005 ;
        RECT 1448.170 6.530 1448.450 6.645 ;
        RECT 1446.860 6.390 1448.450 6.530 ;
        RECT 1346.050 5.850 1346.330 5.965 ;
        RECT 1217.320 5.200 1227.120 5.340 ;
        RECT 1345.200 5.710 1346.330 5.850 ;
        RECT 1209.500 4.350 1210.100 4.490 ;
        RECT 1209.960 3.980 1210.100 4.350 ;
        RECT 1209.960 3.840 1210.560 3.980 ;
        RECT 1191.030 3.670 1191.700 3.810 ;
        RECT 1210.420 3.810 1210.560 3.840 ;
        RECT 1217.320 3.810 1217.460 5.200 ;
        RECT 1345.200 3.810 1345.340 5.710 ;
        RECT 1346.050 5.595 1346.330 5.710 ;
        RECT 1366.290 5.850 1366.570 5.965 ;
        RECT 1366.290 5.710 1366.960 5.850 ;
        RECT 1366.290 5.595 1366.570 5.710 ;
        RECT 1210.420 3.670 1217.460 3.810 ;
        RECT 1334.160 3.670 1345.340 3.810 ;
        RECT 1366.820 3.730 1366.960 5.710 ;
        RECT 1191.030 3.555 1191.310 3.670 ;
        RECT 1122.960 3.300 1123.220 3.390 ;
        RECT 1122.560 3.160 1123.220 3.300 ;
        RECT 1122.960 3.070 1123.220 3.160 ;
        RECT 1126.640 3.070 1126.900 3.390 ;
        RECT 1334.160 3.245 1334.300 3.670 ;
        RECT 1366.760 3.410 1367.020 3.730 ;
        RECT 1334.090 2.875 1334.370 3.245 ;
        RECT 1430.240 3.130 1430.500 3.390 ;
        RECT 1430.240 3.070 1442.860 3.130 ;
        RECT 1430.300 2.990 1442.860 3.070 ;
        RECT 988.170 2.195 988.450 2.565 ;
        RECT 711.320 1.630 713.300 1.770 ;
        RECT 1442.720 1.090 1442.860 2.990 ;
        RECT 1446.860 1.090 1447.000 6.390 ;
        RECT 1448.170 6.275 1448.450 6.390 ;
        RECT 1473.470 6.275 1473.750 6.645 ;
        RECT 1597.740 5.090 1597.880 7.635 ;
        RECT 1638.610 6.275 1638.890 6.645 ;
        RECT 1638.680 5.090 1638.820 6.275 ;
        RECT 1597.680 4.770 1597.940 5.090 ;
        RECT 1638.620 4.770 1638.880 5.090 ;
        RECT 560.840 0.690 561.100 1.010 ;
        RECT 1442.720 0.950 1447.000 1.090 ;
        RECT 469.290 0.155 469.570 0.525 ;
      LAYER via2 ;
        RECT 2787.230 3402.920 2787.510 3403.200 ;
        RECT 2816.210 3402.240 2816.490 3402.520 ;
        RECT 1483.590 3401.560 1483.870 3401.840 ;
        RECT 1823.990 3401.560 1824.270 3401.840 ;
        RECT 1851.130 3401.560 1851.410 3401.840 ;
        RECT 1900.350 3401.560 1900.630 3401.840 ;
        RECT 1973.490 3401.560 1973.770 3401.840 ;
        RECT 2015.810 3401.560 2016.090 3401.840 ;
        RECT 2063.650 3401.560 2063.930 3401.840 ;
        RECT 2093.090 3401.560 2093.370 3401.840 ;
        RECT 2140.930 3401.560 2141.210 3401.840 ;
        RECT 2188.770 3401.560 2189.050 3401.840 ;
        RECT 2256.850 3401.560 2257.130 3401.840 ;
        RECT 2285.830 3401.560 2286.110 3401.840 ;
        RECT 2332.750 3401.560 2333.030 3401.840 ;
        RECT 2405.890 3401.560 2406.170 3401.840 ;
        RECT 2428.890 3401.560 2429.170 3401.840 ;
        RECT 2477.190 3401.560 2477.470 3401.840 ;
        RECT 2529.630 3401.560 2529.910 3401.840 ;
        RECT 2577.010 3401.560 2577.290 3401.840 ;
        RECT 2622.090 3401.560 2622.370 3401.840 ;
        RECT 2671.770 3401.560 2672.050 3401.840 ;
        RECT 2720.070 3401.560 2720.350 3401.840 ;
        RECT 335.430 7.000 335.710 7.280 ;
        RECT 371.310 4.960 371.590 5.240 ;
        RECT 524.030 5.640 524.310 5.920 ;
        RECT 534.150 5.640 534.430 5.920 ;
        RECT 725.510 8.360 725.790 8.640 ;
        RECT 728.270 8.360 728.550 8.640 ;
        RECT 610.050 6.320 610.330 6.600 ;
        RECT 656.510 6.320 656.790 6.600 ;
        RECT 412.250 4.280 412.530 4.560 ;
        RECT 391.090 0.880 391.370 1.160 ;
        RECT 410.870 0.880 411.150 1.160 ;
        RECT 891.570 7.000 891.850 7.280 ;
        RECT 845.570 6.320 845.850 6.600 ;
        RECT 831.770 5.640 832.050 5.920 ;
        RECT 843.270 5.640 843.550 5.920 ;
        RECT 1089.830 6.320 1090.110 6.600 ;
        RECT 914.570 5.640 914.850 5.920 ;
        RECT 921.470 4.960 921.750 5.240 ;
        RECT 952.290 3.600 952.570 3.880 ;
        RECT 987.710 3.600 987.990 3.880 ;
        RECT 1156.530 3.600 1156.810 3.880 ;
        RECT 1191.030 3.600 1191.310 3.880 ;
        RECT 1227.370 8.360 1227.650 8.640 ;
        RECT 1474.850 8.360 1475.130 8.640 ;
        RECT 1597.670 7.680 1597.950 7.960 ;
        RECT 1346.050 5.640 1346.330 5.920 ;
        RECT 1366.290 5.640 1366.570 5.920 ;
        RECT 1334.090 2.920 1334.370 3.200 ;
        RECT 988.170 2.240 988.450 2.520 ;
        RECT 1448.170 6.320 1448.450 6.600 ;
        RECT 1473.470 6.320 1473.750 6.600 ;
        RECT 1638.610 6.320 1638.890 6.600 ;
        RECT 469.290 0.200 469.570 0.480 ;
      LAYER met3 ;
        RECT 2787.205 3403.210 2787.535 3403.225 ;
        RECT 2769.510 3402.910 2787.535 3403.210 ;
        RECT 1483.565 3401.850 1483.895 3401.865 ;
        RECT 1823.965 3401.850 1824.295 3401.865 ;
        RECT 1483.565 3401.550 1824.295 3401.850 ;
        RECT 1483.565 3401.535 1483.895 3401.550 ;
        RECT 1823.965 3401.535 1824.295 3401.550 ;
        RECT 1851.105 3401.850 1851.435 3401.865 ;
        RECT 1900.325 3401.850 1900.655 3401.865 ;
        RECT 1851.105 3401.550 1900.655 3401.850 ;
        RECT 1851.105 3401.535 1851.435 3401.550 ;
        RECT 1900.325 3401.535 1900.655 3401.550 ;
        RECT 1973.465 3401.850 1973.795 3401.865 ;
        RECT 2015.785 3401.850 2016.115 3401.865 ;
        RECT 1973.465 3401.550 2016.115 3401.850 ;
        RECT 1973.465 3401.535 1973.795 3401.550 ;
        RECT 2015.785 3401.535 2016.115 3401.550 ;
        RECT 2063.625 3401.850 2063.955 3401.865 ;
        RECT 2093.065 3401.850 2093.395 3401.865 ;
        RECT 2063.625 3401.550 2093.395 3401.850 ;
        RECT 2063.625 3401.535 2063.955 3401.550 ;
        RECT 2093.065 3401.535 2093.395 3401.550 ;
        RECT 2140.905 3401.850 2141.235 3401.865 ;
        RECT 2188.745 3401.850 2189.075 3401.865 ;
        RECT 2140.905 3401.550 2189.075 3401.850 ;
        RECT 2140.905 3401.535 2141.235 3401.550 ;
        RECT 2188.745 3401.535 2189.075 3401.550 ;
        RECT 2256.825 3401.850 2257.155 3401.865 ;
        RECT 2285.805 3401.850 2286.135 3401.865 ;
        RECT 2256.825 3401.550 2286.135 3401.850 ;
        RECT 2256.825 3401.535 2257.155 3401.550 ;
        RECT 2285.805 3401.535 2286.135 3401.550 ;
        RECT 2332.725 3401.850 2333.055 3401.865 ;
        RECT 2405.865 3401.850 2406.195 3401.865 ;
        RECT 2332.725 3401.550 2406.195 3401.850 ;
        RECT 2332.725 3401.535 2333.055 3401.550 ;
        RECT 2405.865 3401.535 2406.195 3401.550 ;
        RECT 2428.865 3401.850 2429.195 3401.865 ;
        RECT 2477.165 3401.850 2477.495 3401.865 ;
        RECT 2428.865 3401.550 2477.495 3401.850 ;
        RECT 2428.865 3401.535 2429.195 3401.550 ;
        RECT 2477.165 3401.535 2477.495 3401.550 ;
        RECT 2529.605 3401.850 2529.935 3401.865 ;
        RECT 2576.985 3401.850 2577.315 3401.865 ;
        RECT 2529.605 3401.550 2577.315 3401.850 ;
        RECT 2529.605 3401.535 2529.935 3401.550 ;
        RECT 2576.985 3401.535 2577.315 3401.550 ;
        RECT 2622.065 3401.850 2622.395 3401.865 ;
        RECT 2671.745 3401.850 2672.075 3401.865 ;
        RECT 2622.065 3401.550 2672.075 3401.850 ;
        RECT 2622.065 3401.535 2622.395 3401.550 ;
        RECT 2671.745 3401.535 2672.075 3401.550 ;
        RECT 2720.045 3401.850 2720.375 3401.865 ;
        RECT 2769.510 3401.850 2769.810 3402.910 ;
        RECT 2787.205 3402.895 2787.535 3402.910 ;
        RECT 2816.185 3402.530 2816.515 3402.545 ;
        RECT 2822.830 3402.530 2823.210 3402.540 ;
        RECT 2816.185 3402.230 2823.210 3402.530 ;
        RECT 2816.185 3402.215 2816.515 3402.230 ;
        RECT 2822.830 3402.220 2823.210 3402.230 ;
        RECT 2720.045 3401.550 2769.810 3401.850 ;
        RECT 2720.045 3401.535 2720.375 3401.550 ;
        RECT 725.485 8.650 725.815 8.665 ;
        RECT 728.245 8.650 728.575 8.665 ;
        RECT 725.485 8.350 728.575 8.650 ;
        RECT 725.485 8.335 725.815 8.350 ;
        RECT 728.245 8.335 728.575 8.350 ;
        RECT 849.430 8.650 849.810 8.660 ;
        RECT 878.870 8.650 879.250 8.660 ;
        RECT 849.430 8.350 879.250 8.650 ;
        RECT 849.430 8.340 849.810 8.350 ;
        RECT 878.870 8.340 879.250 8.350 ;
        RECT 1227.345 8.650 1227.675 8.665 ;
        RECT 1237.670 8.650 1238.050 8.660 ;
        RECT 1227.345 8.350 1238.050 8.650 ;
        RECT 1227.345 8.335 1227.675 8.350 ;
        RECT 1237.670 8.340 1238.050 8.350 ;
        RECT 1474.825 8.650 1475.155 8.665 ;
        RECT 1474.825 8.350 1548.970 8.650 ;
        RECT 1474.825 8.335 1475.155 8.350 ;
        RECT 1548.670 7.970 1548.970 8.350 ;
        RECT 1597.645 7.970 1597.975 7.985 ;
        RECT 1548.670 7.670 1597.975 7.970 ;
        RECT 1597.645 7.655 1597.975 7.670 ;
        RECT 335.405 7.290 335.735 7.305 ;
        RECT 367.350 7.290 367.730 7.300 ;
        RECT 335.405 6.990 367.730 7.290 ;
        RECT 335.405 6.975 335.735 6.990 ;
        RECT 367.350 6.980 367.730 6.990 ;
        RECT 889.910 7.290 890.290 7.300 ;
        RECT 891.545 7.290 891.875 7.305 ;
        RECT 889.910 6.990 891.875 7.290 ;
        RECT 889.910 6.980 890.290 6.990 ;
        RECT 891.545 6.975 891.875 6.990 ;
        RECT 610.025 6.610 610.355 6.625 ;
        RECT 656.485 6.610 656.815 6.625 ;
        RECT 610.025 6.310 656.815 6.610 ;
        RECT 610.025 6.295 610.355 6.310 ;
        RECT 656.485 6.295 656.815 6.310 ;
        RECT 845.545 6.610 845.875 6.625 ;
        RECT 849.430 6.610 849.810 6.620 ;
        RECT 845.545 6.310 849.810 6.610 ;
        RECT 845.545 6.295 845.875 6.310 ;
        RECT 849.430 6.300 849.810 6.310 ;
        RECT 1087.710 6.610 1088.090 6.620 ;
        RECT 1089.805 6.610 1090.135 6.625 ;
        RECT 1087.710 6.310 1090.135 6.610 ;
        RECT 1087.710 6.300 1088.090 6.310 ;
        RECT 1089.805 6.295 1090.135 6.310 ;
        RECT 1448.145 6.610 1448.475 6.625 ;
        RECT 1473.445 6.610 1473.775 6.625 ;
        RECT 1638.585 6.620 1638.915 6.625 ;
        RECT 1638.585 6.610 1639.170 6.620 ;
        RECT 1448.145 6.310 1473.775 6.610 ;
        RECT 1638.360 6.310 1639.170 6.610 ;
        RECT 1448.145 6.295 1448.475 6.310 ;
        RECT 1473.445 6.295 1473.775 6.310 ;
        RECT 1638.585 6.300 1639.170 6.310 ;
        RECT 1638.585 6.295 1638.915 6.300 ;
        RECT 524.005 5.930 524.335 5.945 ;
        RECT 534.125 5.930 534.455 5.945 ;
        RECT 524.005 5.630 534.455 5.930 ;
        RECT 524.005 5.615 524.335 5.630 ;
        RECT 534.125 5.615 534.455 5.630 ;
        RECT 831.745 5.930 832.075 5.945 ;
        RECT 843.245 5.930 843.575 5.945 ;
        RECT 831.745 5.630 843.575 5.930 ;
        RECT 831.745 5.615 832.075 5.630 ;
        RECT 843.245 5.615 843.575 5.630 ;
        RECT 914.545 5.930 914.875 5.945 ;
        RECT 1346.025 5.930 1346.355 5.945 ;
        RECT 1366.265 5.930 1366.595 5.945 ;
        RECT 914.545 5.630 920.610 5.930 ;
        RECT 914.545 5.615 914.875 5.630 ;
        RECT 367.350 5.250 367.730 5.260 ;
        RECT 371.285 5.250 371.615 5.265 ;
        RECT 416.110 5.250 416.490 5.260 ;
        RECT 367.350 4.950 371.615 5.250 ;
        RECT 367.350 4.940 367.730 4.950 ;
        RECT 371.285 4.935 371.615 4.950 ;
        RECT 412.470 4.950 416.490 5.250 ;
        RECT 920.310 5.250 920.610 5.630 ;
        RECT 1346.025 5.630 1366.595 5.930 ;
        RECT 1346.025 5.615 1346.355 5.630 ;
        RECT 1366.265 5.615 1366.595 5.630 ;
        RECT 921.445 5.250 921.775 5.265 ;
        RECT 920.310 4.950 921.775 5.250 ;
        RECT 412.470 4.585 412.770 4.950 ;
        RECT 416.110 4.940 416.490 4.950 ;
        RECT 921.445 4.935 921.775 4.950 ;
        RECT 412.225 4.270 412.770 4.585 ;
        RECT 1790.590 4.570 1790.970 4.580 ;
        RECT 2822.830 4.570 2823.210 4.580 ;
        RECT 1790.590 4.270 2823.210 4.570 ;
        RECT 412.225 4.255 412.555 4.270 ;
        RECT 1790.590 4.260 1790.970 4.270 ;
        RECT 2822.830 4.260 2823.210 4.270 ;
        RECT 952.265 3.890 952.595 3.905 ;
        RECT 987.685 3.890 988.015 3.905 ;
        RECT 952.265 3.590 988.015 3.890 ;
        RECT 952.265 3.575 952.595 3.590 ;
        RECT 987.685 3.575 988.015 3.590 ;
        RECT 1156.505 3.890 1156.835 3.905 ;
        RECT 1191.005 3.890 1191.335 3.905 ;
        RECT 1156.505 3.590 1191.335 3.890 ;
        RECT 1156.505 3.575 1156.835 3.590 ;
        RECT 1191.005 3.575 1191.335 3.590 ;
        RECT 1324.150 3.210 1324.530 3.220 ;
        RECT 1334.065 3.210 1334.395 3.225 ;
        RECT 1324.150 2.910 1334.395 3.210 ;
        RECT 1324.150 2.900 1324.530 2.910 ;
        RECT 1334.065 2.895 1334.395 2.910 ;
        RECT 1693.990 3.210 1694.370 3.220 ;
        RECT 1713.310 3.210 1713.690 3.220 ;
        RECT 1693.990 2.910 1713.690 3.210 ;
        RECT 1693.990 2.900 1694.370 2.910 ;
        RECT 1713.310 2.900 1713.690 2.910 ;
        RECT 988.145 2.530 988.475 2.545 ;
        RECT 989.270 2.530 989.650 2.540 ;
        RECT 988.145 2.230 989.650 2.530 ;
        RECT 988.145 2.215 988.475 2.230 ;
        RECT 989.270 2.220 989.650 2.230 ;
        RECT 391.065 1.170 391.395 1.185 ;
        RECT 410.845 1.170 411.175 1.185 ;
        RECT 391.065 0.870 411.175 1.170 ;
        RECT 391.065 0.855 391.395 0.870 ;
        RECT 410.845 0.855 411.175 0.870 ;
        RECT 421.630 0.490 422.010 0.500 ;
        RECT 448.310 0.490 448.690 0.500 ;
        RECT 421.630 0.190 448.690 0.490 ;
        RECT 421.630 0.180 422.010 0.190 ;
        RECT 448.310 0.180 448.690 0.190 ;
        RECT 463.030 0.490 463.410 0.500 ;
        RECT 469.265 0.490 469.595 0.505 ;
        RECT 463.030 0.190 469.595 0.490 ;
        RECT 463.030 0.180 463.410 0.190 ;
        RECT 469.265 0.175 469.595 0.190 ;
      LAYER via3 ;
        RECT 2822.860 3402.220 2823.180 3402.540 ;
        RECT 849.460 8.340 849.780 8.660 ;
        RECT 878.900 8.340 879.220 8.660 ;
        RECT 1237.700 8.340 1238.020 8.660 ;
        RECT 367.380 6.980 367.700 7.300 ;
        RECT 889.940 6.980 890.260 7.300 ;
        RECT 849.460 6.300 849.780 6.620 ;
        RECT 1087.740 6.300 1088.060 6.620 ;
        RECT 1638.820 6.300 1639.140 6.620 ;
        RECT 367.380 4.940 367.700 5.260 ;
        RECT 416.140 4.940 416.460 5.260 ;
        RECT 1790.620 4.260 1790.940 4.580 ;
        RECT 2822.860 4.260 2823.180 4.580 ;
        RECT 1324.180 2.900 1324.500 3.220 ;
        RECT 1694.020 2.900 1694.340 3.220 ;
        RECT 1713.340 2.900 1713.660 3.220 ;
        RECT 989.300 2.220 989.620 2.540 ;
        RECT 421.660 0.180 421.980 0.500 ;
        RECT 448.340 0.180 448.660 0.500 ;
        RECT 463.060 0.180 463.380 0.500 ;
      LAYER met4 ;
        RECT 2822.855 3402.215 2823.185 3402.545 ;
        RECT 878.910 9.030 881.050 9.330 ;
        RECT 878.910 8.665 879.210 9.030 ;
        RECT 849.455 8.335 849.785 8.665 ;
        RECT 878.895 8.335 879.225 8.665 ;
        RECT 880.750 8.650 881.050 9.030 ;
        RECT 1237.695 8.650 1238.025 8.665 ;
        RECT 880.750 8.350 886.570 8.650 ;
        RECT 367.375 6.975 367.705 7.305 ;
        RECT 367.390 5.265 367.690 6.975 ;
        RECT 849.470 6.625 849.770 8.335 ;
        RECT 886.270 7.290 886.570 8.350 ;
        RECT 1237.695 8.350 1240.770 8.650 ;
        RECT 1237.695 8.335 1238.025 8.350 ;
        RECT 889.935 7.290 890.265 7.305 ;
        RECT 886.270 6.990 890.265 7.290 ;
        RECT 889.935 6.975 890.265 6.990 ;
        RECT 849.455 6.295 849.785 6.625 ;
        RECT 1087.735 6.295 1088.065 6.625 ;
        RECT 367.375 4.935 367.705 5.265 ;
        RECT 416.135 4.935 416.465 5.265 ;
        RECT 1087.750 5.250 1088.050 6.295 ;
        RECT 1087.750 4.950 1088.970 5.250 ;
        RECT 416.150 0.490 416.450 4.935 ;
        RECT 1088.670 3.210 1088.970 4.950 ;
        RECT 1088.670 2.910 1089.200 3.210 ;
        RECT 989.295 2.290 989.625 2.545 ;
        RECT 1088.900 2.290 1089.200 2.910 ;
        RECT 1240.470 2.290 1240.770 8.350 ;
        RECT 1638.815 6.295 1639.145 6.625 ;
        RECT 1638.830 5.690 1639.130 6.295 ;
        RECT 1638.390 4.510 1639.570 5.690 ;
        RECT 1693.590 4.510 1694.770 5.690 ;
        RECT 2822.870 4.585 2823.170 3402.215 ;
        RECT 1694.030 3.225 1694.330 4.510 ;
        RECT 1790.615 4.255 1790.945 4.585 ;
        RECT 2822.855 4.255 2823.185 4.585 ;
        RECT 1324.175 2.895 1324.505 3.225 ;
        RECT 1694.015 2.895 1694.345 3.225 ;
        RECT 1713.335 2.895 1713.665 3.225 ;
        RECT 1324.190 2.290 1324.490 2.895 ;
        RECT 988.870 1.110 990.050 2.290 ;
        RECT 1088.230 1.110 1089.410 2.290 ;
        RECT 1240.030 1.110 1241.210 2.290 ;
        RECT 1323.750 1.110 1324.930 2.290 ;
        RECT 1713.350 1.850 1713.650 2.895 ;
        RECT 1790.630 2.290 1790.930 4.255 ;
        RECT 1717.510 1.850 1718.690 2.290 ;
        RECT 1713.350 1.550 1718.690 1.850 ;
        RECT 1717.510 1.110 1718.690 1.550 ;
        RECT 1790.190 1.110 1791.370 2.290 ;
        RECT 421.655 0.490 421.985 0.505 ;
        RECT 416.150 0.190 421.985 0.490 ;
        RECT 421.655 0.175 421.985 0.190 ;
        RECT 448.335 0.490 448.665 0.505 ;
        RECT 463.055 0.490 463.385 0.505 ;
        RECT 448.335 0.190 463.385 0.490 ;
        RECT 448.335 0.175 448.665 0.190 ;
        RECT 463.055 0.175 463.385 0.190 ;
      LAYER met5 ;
        RECT 1638.180 4.300 1694.980 5.900 ;
        RECT 988.660 0.900 1089.620 2.500 ;
        RECT 1239.820 0.900 1325.140 2.500 ;
        RECT 1717.300 0.900 1791.580 2.500 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 9.345 1419.585 9.515 1479.935 ;
        RECT 7.965 879.665 8.135 990.335 ;
        RECT 9.805 990.165 9.975 1106.955 ;
        RECT 9.805 817.615 9.975 845.495 ;
        RECT 9.345 817.445 9.975 817.615 ;
        RECT 7.045 707.115 7.215 796.195 ;
        RECT 9.345 796.025 9.515 817.445 ;
        RECT 7.045 706.945 8.135 707.115 ;
        RECT 7.965 655.605 8.135 706.945 ;
        RECT 9.805 624.665 9.975 655.435 ;
        RECT 9.805 535.245 9.975 590.155 ;
        RECT 8.885 456.025 9.055 492.235 ;
        RECT 9.805 332.265 9.975 432.055 ;
        RECT 0.145 174.845 0.315 252.195 ;
        RECT 9.345 252.025 9.515 323.935 ;
        RECT 18.545 8.415 18.715 8.755 ;
        RECT 18.545 8.245 21.015 8.415 ;
        RECT 26.365 8.075 26.535 8.415 ;
        RECT 26.365 7.905 27.915 8.075 ;
        RECT 27.745 4.335 27.915 7.905 ;
        RECT 27.745 4.165 28.375 4.335 ;
        RECT 128.945 4.165 129.115 8.415 ;
        RECT 190.585 0.765 190.755 3.995 ;
        RECT 198.405 0.765 198.575 9.095 ;
        RECT 254.065 8.585 255.155 8.755 ;
        RECT 283.045 7.735 283.215 8.415 ;
        RECT 283.045 7.565 283.675 7.735 ;
      LAYER mcon ;
        RECT 9.345 1479.765 9.515 1479.935 ;
        RECT 9.805 1106.785 9.975 1106.955 ;
        RECT 7.965 990.165 8.135 990.335 ;
        RECT 9.805 845.325 9.975 845.495 ;
        RECT 7.045 796.025 7.215 796.195 ;
        RECT 9.805 655.265 9.975 655.435 ;
        RECT 9.805 589.985 9.975 590.155 ;
        RECT 8.885 492.065 9.055 492.235 ;
        RECT 9.805 431.885 9.975 432.055 ;
        RECT 9.345 323.765 9.515 323.935 ;
        RECT 0.145 252.025 0.315 252.195 ;
        RECT 198.405 8.925 198.575 9.095 ;
        RECT 18.545 8.585 18.715 8.755 ;
        RECT 20.845 8.245 21.015 8.415 ;
        RECT 26.365 8.245 26.535 8.415 ;
        RECT 128.945 8.245 129.115 8.415 ;
        RECT 28.205 4.165 28.375 4.335 ;
        RECT 190.585 3.825 190.755 3.995 ;
        RECT 254.985 8.585 255.155 8.755 ;
        RECT 283.045 8.245 283.215 8.415 ;
        RECT 283.505 7.565 283.675 7.735 ;
      LAYER met1 ;
        RECT 6.970 1479.920 7.290 1479.980 ;
        RECT 9.285 1479.920 9.575 1479.965 ;
        RECT 6.970 1479.780 9.575 1479.920 ;
        RECT 6.970 1479.720 7.290 1479.780 ;
        RECT 9.285 1479.735 9.575 1479.780 ;
        RECT 9.285 1419.740 9.575 1419.785 ;
        RECT 9.730 1419.740 10.050 1419.800 ;
        RECT 9.285 1419.600 10.050 1419.740 ;
        RECT 9.285 1419.555 9.575 1419.600 ;
        RECT 9.730 1419.540 10.050 1419.600 ;
        RECT 1.910 1321.480 2.230 1321.540 ;
        RECT 9.730 1321.480 10.050 1321.540 ;
        RECT 1.910 1321.340 10.050 1321.480 ;
        RECT 1.910 1321.280 2.230 1321.340 ;
        RECT 9.730 1321.280 10.050 1321.340 ;
        RECT 1.910 1106.940 2.230 1107.000 ;
        RECT 9.745 1106.940 10.035 1106.985 ;
        RECT 1.910 1106.800 10.035 1106.940 ;
        RECT 1.910 1106.740 2.230 1106.800 ;
        RECT 9.745 1106.755 10.035 1106.800 ;
        RECT 7.905 990.320 8.195 990.365 ;
        RECT 9.745 990.320 10.035 990.365 ;
        RECT 7.905 990.180 10.035 990.320 ;
        RECT 7.905 990.135 8.195 990.180 ;
        RECT 9.745 990.135 10.035 990.180 ;
        RECT 7.905 879.820 8.195 879.865 ;
        RECT 9.730 879.820 10.050 879.880 ;
        RECT 7.905 879.680 10.050 879.820 ;
        RECT 7.905 879.635 8.195 879.680 ;
        RECT 9.730 879.620 10.050 879.680 ;
        RECT 9.730 845.480 10.050 845.540 ;
        RECT 9.730 845.340 10.245 845.480 ;
        RECT 9.730 845.280 10.050 845.340 ;
        RECT 6.985 796.180 7.275 796.225 ;
        RECT 9.285 796.180 9.575 796.225 ;
        RECT 6.985 796.040 9.575 796.180 ;
        RECT 6.985 795.995 7.275 796.040 ;
        RECT 9.285 795.995 9.575 796.040 ;
        RECT 7.905 655.760 8.195 655.805 ;
        RECT 7.905 655.620 9.500 655.760 ;
        RECT 7.905 655.575 8.195 655.620 ;
        RECT 9.360 655.420 9.500 655.620 ;
        RECT 9.745 655.420 10.035 655.465 ;
        RECT 9.360 655.280 10.035 655.420 ;
        RECT 9.745 655.235 10.035 655.280 ;
        RECT 9.730 624.820 10.050 624.880 ;
        RECT 9.730 624.680 10.245 624.820 ;
        RECT 9.730 624.620 10.050 624.680 ;
        RECT 9.730 590.140 10.050 590.200 ;
        RECT 9.535 590.000 10.050 590.140 ;
        RECT 9.730 589.940 10.050 590.000 ;
        RECT 9.730 535.400 10.050 535.460 ;
        RECT 9.535 535.260 10.050 535.400 ;
        RECT 9.730 535.200 10.050 535.260 ;
        RECT 8.825 492.220 9.115 492.265 ;
        RECT 9.730 492.220 10.050 492.280 ;
        RECT 8.825 492.080 10.050 492.220 ;
        RECT 8.825 492.035 9.115 492.080 ;
        RECT 9.730 492.020 10.050 492.080 ;
        RECT 8.825 456.180 9.115 456.225 ;
        RECT 9.730 456.180 10.050 456.240 ;
        RECT 8.825 456.040 10.050 456.180 ;
        RECT 8.825 455.995 9.115 456.040 ;
        RECT 9.730 455.980 10.050 456.040 ;
        RECT 9.730 432.040 10.050 432.100 ;
        RECT 9.535 431.900 10.050 432.040 ;
        RECT 9.730 431.840 10.050 431.900 ;
        RECT 9.730 332.420 10.050 332.480 ;
        RECT 9.535 332.280 10.050 332.420 ;
        RECT 9.730 332.220 10.050 332.280 ;
        RECT 9.285 323.920 9.575 323.965 ;
        RECT 9.730 323.920 10.050 323.980 ;
        RECT 9.285 323.780 10.050 323.920 ;
        RECT 9.285 323.735 9.575 323.780 ;
        RECT 9.730 323.720 10.050 323.780 ;
        RECT 0.085 252.180 0.375 252.225 ;
        RECT 9.285 252.180 9.575 252.225 ;
        RECT 0.085 252.040 9.575 252.180 ;
        RECT 0.085 251.995 0.375 252.040 ;
        RECT 9.285 251.995 9.575 252.040 ;
        RECT 0.070 175.000 0.390 175.060 ;
        RECT 0.070 174.860 0.585 175.000 ;
        RECT 0.070 174.800 0.390 174.860 ;
        RECT 198.345 9.080 198.635 9.125 ;
        RECT 198.345 8.940 244.560 9.080 ;
        RECT 198.345 8.895 198.635 8.940 ;
        RECT 244.420 8.800 244.560 8.940 ;
        RECT 18.485 8.740 18.775 8.785 ;
        RECT 8.900 8.600 18.775 8.740 ;
        RECT 0.070 8.060 0.390 8.120 ;
        RECT 8.900 8.060 9.040 8.600 ;
        RECT 18.485 8.555 18.775 8.600 ;
        RECT 244.330 8.540 244.650 8.800 ;
        RECT 253.990 8.740 254.310 8.800 ;
        RECT 253.795 8.600 254.310 8.740 ;
        RECT 253.990 8.540 254.310 8.600 ;
        RECT 254.925 8.740 255.215 8.785 ;
        RECT 254.925 8.600 281.820 8.740 ;
        RECT 254.925 8.555 255.215 8.600 ;
        RECT 20.785 8.400 21.075 8.445 ;
        RECT 26.305 8.400 26.595 8.445 ;
        RECT 20.785 8.260 26.595 8.400 ;
        RECT 20.785 8.215 21.075 8.260 ;
        RECT 26.305 8.215 26.595 8.260 ;
        RECT 128.885 8.400 129.175 8.445 ;
        RECT 133.010 8.400 133.330 8.460 ;
        RECT 128.885 8.260 133.330 8.400 ;
        RECT 281.680 8.400 281.820 8.600 ;
        RECT 282.985 8.400 283.275 8.445 ;
        RECT 281.680 8.260 283.275 8.400 ;
        RECT 128.885 8.215 129.175 8.260 ;
        RECT 133.010 8.200 133.330 8.260 ;
        RECT 282.985 8.215 283.275 8.260 ;
        RECT 0.070 7.920 9.040 8.060 ;
        RECT 0.070 7.860 0.390 7.920 ;
        RECT 283.445 7.720 283.735 7.765 ;
        RECT 290.330 7.720 290.650 7.780 ;
        RECT 283.445 7.580 290.650 7.720 ;
        RECT 283.445 7.535 283.735 7.580 ;
        RECT 290.330 7.520 290.650 7.580 ;
        RECT 290.330 4.660 290.650 4.720 ;
        RECT 305.970 4.660 306.290 4.720 ;
        RECT 290.330 4.520 306.290 4.660 ;
        RECT 290.330 4.460 290.650 4.520 ;
        RECT 305.970 4.460 306.290 4.520 ;
        RECT 28.145 4.320 28.435 4.365 ;
        RECT 128.885 4.320 129.175 4.365 ;
        RECT 28.145 4.180 129.175 4.320 ;
        RECT 28.145 4.135 28.435 4.180 ;
        RECT 128.885 4.135 129.175 4.180 ;
        RECT 148.650 3.980 148.970 4.040 ;
        RECT 190.525 3.980 190.815 4.025 ;
        RECT 148.650 3.840 190.815 3.980 ;
        RECT 148.650 3.780 148.970 3.840 ;
        RECT 190.525 3.795 190.815 3.840 ;
        RECT 190.525 0.920 190.815 0.965 ;
        RECT 198.345 0.920 198.635 0.965 ;
        RECT 190.525 0.780 198.635 0.920 ;
        RECT 190.525 0.735 190.815 0.780 ;
        RECT 198.345 0.735 198.635 0.780 ;
      LAYER via ;
        RECT 7.000 1479.720 7.260 1479.980 ;
        RECT 9.760 1419.540 10.020 1419.800 ;
        RECT 1.940 1321.280 2.200 1321.540 ;
        RECT 9.760 1321.280 10.020 1321.540 ;
        RECT 1.940 1106.740 2.200 1107.000 ;
        RECT 9.760 879.620 10.020 879.880 ;
        RECT 9.760 845.280 10.020 845.540 ;
        RECT 9.760 624.620 10.020 624.880 ;
        RECT 9.760 589.940 10.020 590.200 ;
        RECT 9.760 535.200 10.020 535.460 ;
        RECT 9.760 492.020 10.020 492.280 ;
        RECT 9.760 455.980 10.020 456.240 ;
        RECT 9.760 431.840 10.020 432.100 ;
        RECT 9.760 332.220 10.020 332.480 ;
        RECT 9.760 323.720 10.020 323.980 ;
        RECT 0.100 174.800 0.360 175.060 ;
        RECT 0.100 7.860 0.360 8.120 ;
        RECT 244.360 8.540 244.620 8.800 ;
        RECT 254.020 8.540 254.280 8.800 ;
        RECT 133.040 8.200 133.300 8.460 ;
        RECT 290.360 7.520 290.620 7.780 ;
        RECT 290.360 4.460 290.620 4.720 ;
        RECT 306.000 4.460 306.260 4.720 ;
        RECT 148.680 3.780 148.940 4.040 ;
      LAYER met2 ;
        RECT 6.990 1531.515 7.270 1531.885 ;
        RECT 7.060 1480.010 7.200 1531.515 ;
        RECT 7.000 1479.690 7.260 1480.010 ;
        RECT 9.760 1419.740 10.020 1419.830 ;
        RECT 9.760 1419.600 10.880 1419.740 ;
        RECT 9.760 1419.510 10.020 1419.600 ;
        RECT 10.740 1366.530 10.880 1419.600 ;
        RECT 10.740 1366.390 13.180 1366.530 ;
        RECT 13.040 1322.330 13.180 1366.390 ;
        RECT 9.820 1322.190 13.180 1322.330 ;
        RECT 9.820 1321.570 9.960 1322.190 ;
        RECT 1.940 1321.250 2.200 1321.570 ;
        RECT 9.760 1321.250 10.020 1321.570 ;
        RECT 2.000 1107.030 2.140 1321.250 ;
        RECT 1.940 1106.710 2.200 1107.030 ;
        RECT 9.760 879.590 10.020 879.910 ;
        RECT 9.820 845.570 9.960 879.590 ;
        RECT 9.760 845.250 10.020 845.570 ;
        RECT 9.760 624.590 10.020 624.910 ;
        RECT 9.820 590.230 9.960 624.590 ;
        RECT 9.760 589.910 10.020 590.230 ;
        RECT 9.760 535.170 10.020 535.490 ;
        RECT 9.820 492.310 9.960 535.170 ;
        RECT 9.760 491.990 10.020 492.310 ;
        RECT 9.760 455.950 10.020 456.270 ;
        RECT 9.820 432.130 9.960 455.950 ;
        RECT 9.760 431.810 10.020 432.130 ;
        RECT 9.760 332.190 10.020 332.510 ;
        RECT 9.820 324.010 9.960 332.190 ;
        RECT 9.760 323.690 10.020 324.010 ;
        RECT 0.100 174.770 0.360 175.090 ;
        RECT 0.160 8.150 0.300 174.770 ;
        RECT 244.360 8.570 244.620 8.830 ;
        RECT 244.360 8.510 245.480 8.570 ;
        RECT 254.020 8.510 254.280 8.830 ;
        RECT 133.040 8.170 133.300 8.490 ;
        RECT 244.420 8.430 245.480 8.510 ;
        RECT 0.100 7.830 0.360 8.150 ;
        RECT 133.100 8.005 133.240 8.170 ;
        RECT 133.030 7.635 133.310 8.005 ;
        RECT 148.670 7.635 148.950 8.005 ;
        RECT 245.340 7.890 245.480 8.430 ;
        RECT 254.080 8.005 254.220 8.510 ;
        RECT 246.650 7.890 246.930 8.005 ;
        RECT 245.340 7.750 246.930 7.890 ;
        RECT 246.650 7.635 246.930 7.750 ;
        RECT 254.010 7.635 254.290 8.005 ;
        RECT 148.740 4.070 148.880 7.635 ;
        RECT 290.360 7.490 290.620 7.810 ;
        RECT 305.990 7.635 306.270 8.005 ;
        RECT 322.550 7.635 322.830 8.005 ;
        RECT 290.420 4.750 290.560 7.490 ;
        RECT 306.060 4.750 306.200 7.635 ;
        RECT 322.620 6.700 322.760 7.635 ;
        RECT 322.620 6.560 323.680 6.700 ;
        RECT 323.540 6.360 323.680 6.560 ;
        RECT 323.540 6.220 325.520 6.360 ;
        RECT 290.360 4.430 290.620 4.750 ;
        RECT 306.000 4.430 306.260 4.750 ;
        RECT 325.380 4.320 325.520 6.220 ;
        RECT 325.380 4.180 330.120 4.320 ;
        RECT 148.680 3.750 148.940 4.070 ;
        RECT 329.980 2.400 330.120 4.180 ;
        RECT 329.770 -4.800 330.330 2.400 ;
      LAYER via2 ;
        RECT 6.990 1531.560 7.270 1531.840 ;
        RECT 133.030 7.680 133.310 7.960 ;
        RECT 148.670 7.680 148.950 7.960 ;
        RECT 246.650 7.680 246.930 7.960 ;
        RECT 254.010 7.680 254.290 7.960 ;
        RECT 305.990 7.680 306.270 7.960 ;
        RECT 322.550 7.680 322.830 7.960 ;
      LAYER met3 ;
        RECT 5.000 1534.360 9.000 1534.960 ;
        RECT 6.750 1531.865 7.050 1534.360 ;
        RECT 6.750 1531.550 7.295 1531.865 ;
        RECT 6.965 1531.535 7.295 1531.550 ;
        RECT 133.005 7.970 133.335 7.985 ;
        RECT 148.645 7.970 148.975 7.985 ;
        RECT 133.005 7.670 148.975 7.970 ;
        RECT 133.005 7.655 133.335 7.670 ;
        RECT 148.645 7.655 148.975 7.670 ;
        RECT 246.625 7.970 246.955 7.985 ;
        RECT 253.985 7.970 254.315 7.985 ;
        RECT 246.625 7.670 254.315 7.970 ;
        RECT 246.625 7.655 246.955 7.670 ;
        RECT 253.985 7.655 254.315 7.670 ;
        RECT 305.965 7.970 306.295 7.985 ;
        RECT 322.525 7.970 322.855 7.985 ;
        RECT 305.965 7.670 322.855 7.970 ;
        RECT 305.965 7.655 306.295 7.670 ;
        RECT 322.525 7.655 322.855 7.670 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 9.345 932.365 9.515 975.715 ;
        RECT 9.805 881.025 9.975 888.335 ;
        RECT 1.525 728.025 1.695 839.035 ;
        RECT 295.465 1.445 295.635 6.715 ;
        RECT 304.205 0.765 304.375 1.615 ;
      LAYER mcon ;
        RECT 9.345 975.545 9.515 975.715 ;
        RECT 9.805 888.165 9.975 888.335 ;
        RECT 1.525 838.865 1.695 839.035 ;
        RECT 295.465 6.545 295.635 6.715 ;
        RECT 304.205 1.445 304.375 1.615 ;
      LAYER met1 ;
        RECT 3.290 975.700 3.610 975.760 ;
        RECT 9.285 975.700 9.575 975.745 ;
        RECT 3.290 975.560 9.575 975.700 ;
        RECT 3.290 975.500 3.610 975.560 ;
        RECT 9.285 975.515 9.575 975.560 ;
        RECT 9.285 932.520 9.575 932.565 ;
        RECT 9.730 932.520 10.050 932.580 ;
        RECT 9.285 932.380 10.050 932.520 ;
        RECT 9.285 932.335 9.575 932.380 ;
        RECT 9.730 932.320 10.050 932.380 ;
        RECT 9.730 888.320 10.050 888.380 ;
        RECT 9.535 888.180 10.050 888.320 ;
        RECT 9.730 888.120 10.050 888.180 ;
        RECT 9.730 881.180 10.050 881.240 ;
        RECT 9.535 881.040 10.050 881.180 ;
        RECT 9.730 880.980 10.050 881.040 ;
        RECT 1.465 839.020 1.755 839.065 ;
        RECT 9.730 839.020 10.050 839.080 ;
        RECT 1.465 838.880 10.050 839.020 ;
        RECT 1.465 838.835 1.755 838.880 ;
        RECT 9.730 838.820 10.050 838.880 ;
        RECT 1.450 728.180 1.770 728.240 ;
        RECT 1.255 728.040 1.770 728.180 ;
        RECT 1.450 727.980 1.770 728.040 ;
        RECT 291.250 6.700 291.570 6.760 ;
        RECT 295.405 6.700 295.695 6.745 ;
        RECT 291.250 6.560 295.695 6.700 ;
        RECT 291.250 6.500 291.570 6.560 ;
        RECT 295.405 6.515 295.695 6.560 ;
        RECT 295.405 1.600 295.695 1.645 ;
        RECT 304.145 1.600 304.435 1.645 ;
        RECT 295.405 1.460 304.435 1.600 ;
        RECT 295.405 1.415 295.695 1.460 ;
        RECT 304.145 1.415 304.435 1.460 ;
        RECT 304.145 0.920 304.435 0.965 ;
        RECT 346.450 0.920 346.770 0.980 ;
        RECT 304.145 0.780 346.770 0.920 ;
        RECT 304.145 0.735 304.435 0.780 ;
        RECT 346.450 0.720 346.770 0.780 ;
      LAYER via ;
        RECT 3.320 975.500 3.580 975.760 ;
        RECT 9.760 932.320 10.020 932.580 ;
        RECT 9.760 888.120 10.020 888.380 ;
        RECT 9.760 880.980 10.020 881.240 ;
        RECT 9.760 838.820 10.020 839.080 ;
        RECT 1.480 727.980 1.740 728.240 ;
        RECT 291.280 6.500 291.540 6.760 ;
        RECT 346.480 0.720 346.740 0.980 ;
      LAYER met2 ;
        RECT 3.310 1645.075 3.590 1645.445 ;
        RECT 3.380 975.790 3.520 1645.075 ;
        RECT 3.320 975.470 3.580 975.790 ;
        RECT 9.760 932.290 10.020 932.610 ;
        RECT 9.820 888.410 9.960 932.290 ;
        RECT 9.760 888.090 10.020 888.410 ;
        RECT 9.760 881.180 10.020 881.270 ;
        RECT 9.760 881.040 10.420 881.180 ;
        RECT 9.760 880.950 10.020 881.040 ;
        RECT 10.280 880.500 10.420 881.040 ;
        RECT 10.280 880.360 10.880 880.500 ;
        RECT 9.760 839.020 10.020 839.110 ;
        RECT 10.740 839.020 10.880 880.360 ;
        RECT 9.760 838.880 10.880 839.020 ;
        RECT 9.760 838.790 10.020 838.880 ;
        RECT 1.480 727.950 1.740 728.270 ;
        RECT 1.540 1.885 1.680 727.950 ;
        RECT 196.510 6.955 196.790 7.325 ;
        RECT 211.230 6.955 211.510 7.325 ;
        RECT 196.580 5.965 196.720 6.955 ;
        RECT 211.300 5.965 211.440 6.955 ;
        RECT 291.280 6.470 291.540 6.790 ;
        RECT 196.510 5.595 196.790 5.965 ;
        RECT 211.230 5.595 211.510 5.965 ;
        RECT 290.810 5.850 291.090 5.965 ;
        RECT 291.340 5.850 291.480 6.470 ;
        RECT 290.810 5.710 291.480 5.850 ;
        RECT 290.810 5.595 291.090 5.710 ;
        RECT 346.540 2.990 347.600 3.130 ;
        RECT 1.470 1.515 1.750 1.885 ;
        RECT 346.540 1.010 346.680 2.990 ;
        RECT 347.460 2.400 347.600 2.990 ;
        RECT 346.480 0.690 346.740 1.010 ;
        RECT 347.250 -4.800 347.810 2.400 ;
      LAYER via2 ;
        RECT 3.310 1645.120 3.590 1645.400 ;
        RECT 196.510 7.000 196.790 7.280 ;
        RECT 211.230 7.000 211.510 7.280 ;
        RECT 196.510 5.640 196.790 5.920 ;
        RECT 211.230 5.640 211.510 5.920 ;
        RECT 290.810 5.640 291.090 5.920 ;
        RECT 1.470 1.560 1.750 1.840 ;
      LAYER met3 ;
        RECT 5.000 1647.920 9.000 1648.520 ;
        RECT 3.285 1645.410 3.615 1645.425 ;
        RECT 5.830 1645.410 6.130 1647.920 ;
        RECT 3.285 1645.110 6.130 1645.410 ;
        RECT 3.285 1645.095 3.615 1645.110 ;
        RECT 196.485 7.290 196.815 7.305 ;
        RECT 211.205 7.290 211.535 7.305 ;
        RECT 196.485 6.990 211.535 7.290 ;
        RECT 196.485 6.975 196.815 6.990 ;
        RECT 211.205 6.975 211.535 6.990 ;
        RECT 54.550 5.930 54.930 5.940 ;
        RECT 196.485 5.930 196.815 5.945 ;
        RECT 54.550 5.630 196.815 5.930 ;
        RECT 54.550 5.620 54.930 5.630 ;
        RECT 196.485 5.615 196.815 5.630 ;
        RECT 211.205 5.930 211.535 5.945 ;
        RECT 290.785 5.930 291.115 5.945 ;
        RECT 211.205 5.630 291.115 5.930 ;
        RECT 211.205 5.615 211.535 5.630 ;
        RECT 290.785 5.615 291.115 5.630 ;
        RECT 1.445 1.850 1.775 1.865 ;
        RECT 2.110 1.850 2.490 1.860 ;
        RECT 1.445 1.550 2.490 1.850 ;
        RECT 1.445 1.535 1.775 1.550 ;
        RECT 2.110 1.540 2.490 1.550 ;
      LAYER via3 ;
        RECT 54.580 5.620 54.900 5.940 ;
        RECT 2.140 1.540 2.460 1.860 ;
      LAYER met4 ;
        RECT 54.575 5.615 54.905 5.945 ;
        RECT 54.590 2.290 54.890 5.615 ;
        RECT 1.710 1.110 2.890 2.290 ;
        RECT 54.150 1.110 55.330 2.290 ;
      LAYER met5 ;
        RECT 1.500 0.900 55.540 2.500 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 967.450 2.280 967.770 2.340 ;
        RECT 991.830 2.280 992.150 2.340 ;
        RECT 967.450 2.140 992.150 2.280 ;
        RECT 967.450 2.080 967.770 2.140 ;
        RECT 991.830 2.080 992.150 2.140 ;
      LAYER via ;
        RECT 967.480 2.080 967.740 2.340 ;
        RECT 991.860 2.080 992.120 2.340 ;
      LAYER met2 ;
        RECT 2213.550 5.000 2213.830 9.000 ;
        RECT 401.280 2.990 402.340 3.130 ;
        RECT 401.280 2.400 401.420 2.990 ;
        RECT 402.200 2.565 402.340 2.990 ;
        RECT 953.280 2.990 955.260 3.130 ;
        RECT 953.280 2.565 953.420 2.990 ;
        RECT 401.070 -4.800 401.630 2.400 ;
        RECT 402.130 2.195 402.410 2.565 ;
        RECT 646.390 2.450 646.670 2.565 ;
        RECT 649.610 2.450 649.890 2.565 ;
        RECT 646.390 2.310 649.890 2.450 ;
        RECT 646.390 2.195 646.670 2.310 ;
        RECT 649.610 2.195 649.890 2.310 ;
        RECT 784.390 2.450 784.670 2.565 ;
        RECT 785.770 2.450 786.050 2.565 ;
        RECT 784.390 2.310 786.050 2.450 ;
        RECT 784.390 2.195 784.670 2.310 ;
        RECT 785.770 2.195 786.050 2.310 ;
        RECT 953.210 2.195 953.490 2.565 ;
        RECT 955.120 1.260 955.260 2.990 ;
        RECT 959.260 2.990 967.220 3.130 ;
        RECT 959.260 1.260 959.400 2.990 ;
        RECT 967.080 2.280 967.220 2.990 ;
        RECT 2213.680 2.565 2213.820 5.000 ;
        RECT 967.480 2.280 967.740 2.370 ;
        RECT 967.080 2.140 967.740 2.280 ;
        RECT 991.850 2.195 992.130 2.565 ;
        RECT 2213.610 2.195 2213.890 2.565 ;
        RECT 967.480 2.050 967.740 2.140 ;
        RECT 991.860 2.050 992.120 2.195 ;
        RECT 955.120 1.120 959.400 1.260 ;
      LAYER via2 ;
        RECT 402.130 2.240 402.410 2.520 ;
        RECT 646.390 2.240 646.670 2.520 ;
        RECT 649.610 2.240 649.890 2.520 ;
        RECT 784.390 2.240 784.670 2.520 ;
        RECT 785.770 2.240 786.050 2.520 ;
        RECT 953.210 2.240 953.490 2.520 ;
        RECT 991.850 2.240 992.130 2.520 ;
        RECT 2213.610 2.240 2213.890 2.520 ;
      LAYER met3 ;
        RECT 752.870 2.910 755.010 3.210 ;
        RECT 402.105 2.530 402.435 2.545 ;
        RECT 512.710 2.530 513.090 2.540 ;
        RECT 402.105 2.230 513.090 2.530 ;
        RECT 402.105 2.215 402.435 2.230 ;
        RECT 512.710 2.220 513.090 2.230 ;
        RECT 516.390 2.530 516.770 2.540 ;
        RECT 558.710 2.530 559.090 2.540 ;
        RECT 516.390 2.230 559.090 2.530 ;
        RECT 516.390 2.220 516.770 2.230 ;
        RECT 558.710 2.220 559.090 2.230 ;
        RECT 561.470 2.530 561.850 2.540 ;
        RECT 646.365 2.530 646.695 2.545 ;
        RECT 561.470 2.230 614.250 2.530 ;
        RECT 561.470 2.220 561.850 2.230 ;
        RECT 613.950 1.850 614.250 2.230 ;
        RECT 615.790 2.230 646.695 2.530 ;
        RECT 615.790 1.850 616.090 2.230 ;
        RECT 646.365 2.215 646.695 2.230 ;
        RECT 649.585 2.530 649.915 2.545 ;
        RECT 752.870 2.530 753.170 2.910 ;
        RECT 649.585 2.230 753.170 2.530 ;
        RECT 754.710 2.530 755.010 2.910 ;
        RECT 784.365 2.530 784.695 2.545 ;
        RECT 754.710 2.230 784.695 2.530 ;
        RECT 649.585 2.215 649.915 2.230 ;
        RECT 784.365 2.215 784.695 2.230 ;
        RECT 785.745 2.530 786.075 2.545 ;
        RECT 953.185 2.530 953.515 2.545 ;
        RECT 785.745 2.230 953.515 2.530 ;
        RECT 785.745 2.215 786.075 2.230 ;
        RECT 953.185 2.215 953.515 2.230 ;
        RECT 991.825 2.530 992.155 2.545 ;
        RECT 2213.585 2.530 2213.915 2.545 ;
        RECT 991.825 2.230 2213.915 2.530 ;
        RECT 991.825 2.215 992.155 2.230 ;
        RECT 2213.585 2.215 2213.915 2.230 ;
        RECT 613.950 1.550 616.090 1.850 ;
      LAYER via3 ;
        RECT 512.740 2.220 513.060 2.540 ;
        RECT 516.420 2.220 516.740 2.540 ;
        RECT 558.740 2.220 559.060 2.540 ;
        RECT 561.500 2.220 561.820 2.540 ;
      LAYER met4 ;
        RECT 512.750 2.910 516.730 3.210 ;
        RECT 512.750 2.545 513.050 2.910 ;
        RECT 516.430 2.545 516.730 2.910 ;
        RECT 512.735 2.215 513.065 2.545 ;
        RECT 516.415 2.215 516.745 2.545 ;
        RECT 558.735 2.530 559.065 2.545 ;
        RECT 561.495 2.530 561.825 2.545 ;
        RECT 558.735 2.230 561.825 2.530 ;
        RECT 558.735 2.215 559.065 2.230 ;
        RECT 561.495 2.215 561.825 2.230 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1491.925 8.585 1493.015 8.755 ;
        RECT 584.805 7.565 600.615 7.735 ;
        RECT 191.505 4.165 191.675 5.015 ;
        RECT 414.145 3.315 414.315 5.015 ;
        RECT 417.825 3.655 417.995 5.015 ;
        RECT 580.665 4.335 580.835 5.015 ;
        RECT 584.805 4.335 584.975 7.565 ;
        RECT 600.445 7.395 600.615 7.565 ;
        RECT 600.445 7.225 602.915 7.395 ;
        RECT 602.745 6.035 602.915 7.225 ;
        RECT 602.745 5.865 605.215 6.035 ;
        RECT 580.665 4.165 584.975 4.335 ;
        RECT 415.985 3.485 417.995 3.655 ;
        RECT 415.985 3.315 416.155 3.485 ;
        RECT 414.145 3.145 416.155 3.315 ;
        RECT 605.045 1.615 605.215 5.865 ;
        RECT 1484.565 5.015 1484.735 8.415 ;
        RECT 1491.925 8.245 1492.095 8.585 ;
        RECT 1492.845 8.075 1493.015 8.585 ;
        RECT 1492.845 7.905 1494.395 8.075 ;
        RECT 647.365 4.845 659.035 5.015 ;
        RECT 703.485 4.845 704.575 5.015 ;
        RECT 727.865 4.845 728.955 5.015 ;
        RECT 647.365 1.615 647.535 4.845 ;
        RECT 728.785 4.505 728.955 4.845 ;
        RECT 760.065 4.675 760.235 5.015 ;
        RECT 761.445 4.675 761.615 5.015 ;
        RECT 896.225 4.845 897.315 5.015 ;
        RECT 1091.725 4.845 1092.815 5.015 ;
        RECT 1209.025 4.845 1210.575 5.015 ;
        RECT 1484.105 4.845 1484.735 5.015 ;
        RECT 760.065 4.505 761.615 4.675 ;
        RECT 605.045 1.445 647.535 1.615 ;
      LAYER mcon ;
        RECT 1484.565 8.245 1484.735 8.415 ;
        RECT 191.505 4.845 191.675 5.015 ;
        RECT 414.145 4.845 414.315 5.015 ;
        RECT 417.825 4.845 417.995 5.015 ;
        RECT 580.665 4.845 580.835 5.015 ;
        RECT 1494.225 7.905 1494.395 8.075 ;
        RECT 658.865 4.845 659.035 5.015 ;
        RECT 704.405 4.845 704.575 5.015 ;
        RECT 760.065 4.845 760.235 5.015 ;
        RECT 761.445 4.845 761.615 5.015 ;
        RECT 897.145 4.845 897.315 5.015 ;
        RECT 1092.645 4.845 1092.815 5.015 ;
        RECT 1210.405 4.845 1210.575 5.015 ;
      LAYER met1 ;
        RECT 1484.505 8.400 1484.795 8.445 ;
        RECT 1491.865 8.400 1492.155 8.445 ;
        RECT 1484.505 8.260 1492.155 8.400 ;
        RECT 1484.505 8.215 1484.795 8.260 ;
        RECT 1491.865 8.215 1492.155 8.260 ;
        RECT 1494.165 8.060 1494.455 8.105 ;
        RECT 1974.390 8.060 1974.710 8.120 ;
        RECT 1494.165 7.920 1974.710 8.060 ;
        RECT 1494.165 7.875 1494.455 7.920 ;
        RECT 1974.390 7.860 1974.710 7.920 ;
        RECT 191.445 5.000 191.735 5.045 ;
        RECT 414.085 5.000 414.375 5.045 ;
        RECT 191.445 4.860 414.375 5.000 ;
        RECT 191.445 4.815 191.735 4.860 ;
        RECT 414.085 4.815 414.375 4.860 ;
        RECT 417.765 5.000 418.055 5.045 ;
        RECT 580.605 5.000 580.895 5.045 ;
        RECT 417.765 4.860 580.895 5.000 ;
        RECT 417.765 4.815 418.055 4.860 ;
        RECT 580.605 4.815 580.895 4.860 ;
        RECT 658.805 5.000 659.095 5.045 ;
        RECT 703.425 5.000 703.715 5.045 ;
        RECT 658.805 4.860 703.715 5.000 ;
        RECT 658.805 4.815 659.095 4.860 ;
        RECT 703.425 4.815 703.715 4.860 ;
        RECT 704.345 5.000 704.635 5.045 ;
        RECT 727.805 5.000 728.095 5.045 ;
        RECT 760.005 5.000 760.295 5.045 ;
        RECT 704.345 4.860 728.095 5.000 ;
        RECT 704.345 4.815 704.635 4.860 ;
        RECT 727.805 4.815 728.095 4.860 ;
        RECT 731.100 4.860 760.295 5.000 ;
        RECT 728.725 4.660 729.015 4.705 ;
        RECT 731.100 4.660 731.240 4.860 ;
        RECT 760.005 4.815 760.295 4.860 ;
        RECT 761.385 5.000 761.675 5.045 ;
        RECT 896.165 5.000 896.455 5.045 ;
        RECT 761.385 4.860 804.840 5.000 ;
        RECT 761.385 4.815 761.675 4.860 ;
        RECT 728.725 4.520 731.240 4.660 ;
        RECT 804.700 4.660 804.840 4.860 ;
        RECT 805.620 4.860 896.455 5.000 ;
        RECT 805.620 4.660 805.760 4.860 ;
        RECT 896.165 4.815 896.455 4.860 ;
        RECT 897.085 5.000 897.375 5.045 ;
        RECT 1091.665 5.000 1091.955 5.045 ;
        RECT 897.085 4.860 1091.955 5.000 ;
        RECT 897.085 4.815 897.375 4.860 ;
        RECT 1091.665 4.815 1091.955 4.860 ;
        RECT 1092.585 5.000 1092.875 5.045 ;
        RECT 1208.965 5.000 1209.255 5.045 ;
        RECT 1092.585 4.860 1209.255 5.000 ;
        RECT 1092.585 4.815 1092.875 4.860 ;
        RECT 1208.965 4.815 1209.255 4.860 ;
        RECT 1210.345 5.000 1210.635 5.045 ;
        RECT 1484.045 5.000 1484.335 5.045 ;
        RECT 1210.345 4.860 1484.335 5.000 ;
        RECT 1210.345 4.815 1210.635 4.860 ;
        RECT 1484.045 4.815 1484.335 4.860 ;
        RECT 804.700 4.520 805.760 4.660 ;
        RECT 728.725 4.475 729.015 4.520 ;
        RECT 141.290 4.320 141.610 4.380 ;
        RECT 191.445 4.320 191.735 4.365 ;
        RECT 141.290 4.180 191.735 4.320 ;
        RECT 141.290 4.120 141.610 4.180 ;
        RECT 191.445 4.135 191.735 4.180 ;
      LAYER via ;
        RECT 1974.420 7.860 1974.680 8.120 ;
        RECT 141.320 4.120 141.580 4.380 ;
      LAYER met2 ;
        RECT 1974.420 7.890 1974.680 8.150 ;
        RECT 1975.730 7.890 1976.010 9.000 ;
        RECT 1974.420 7.830 1976.010 7.890 ;
        RECT 1974.480 7.750 1976.010 7.830 ;
        RECT 73.230 6.955 73.510 7.325 ;
        RECT 141.310 6.955 141.590 7.325 ;
        RECT 62.260 2.990 63.320 3.130 ;
        RECT 62.260 2.400 62.400 2.990 ;
        RECT 62.050 -4.800 62.610 2.400 ;
        RECT 63.180 1.885 63.320 2.990 ;
        RECT 73.300 1.885 73.440 6.955 ;
        RECT 141.380 4.410 141.520 6.955 ;
        RECT 1975.730 5.000 1976.010 7.750 ;
        RECT 141.320 4.090 141.580 4.410 ;
        RECT 63.110 1.515 63.390 1.885 ;
        RECT 73.230 1.515 73.510 1.885 ;
      LAYER via2 ;
        RECT 73.230 7.000 73.510 7.280 ;
        RECT 141.310 7.000 141.590 7.280 ;
        RECT 63.110 1.560 63.390 1.840 ;
        RECT 73.230 1.560 73.510 1.840 ;
      LAYER met3 ;
        RECT 73.205 7.290 73.535 7.305 ;
        RECT 141.285 7.290 141.615 7.305 ;
        RECT 73.205 6.990 141.615 7.290 ;
        RECT 73.205 6.975 73.535 6.990 ;
        RECT 141.285 6.975 141.615 6.990 ;
        RECT 63.085 1.850 63.415 1.865 ;
        RECT 73.205 1.850 73.535 1.865 ;
        RECT 63.085 1.550 73.535 1.850 ;
        RECT 63.085 1.535 63.415 1.550 ;
        RECT 73.205 1.535 73.535 1.550 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 870.925 9.265 891.335 9.435 ;
        RECT 870.925 8.585 871.095 9.265 ;
        RECT 804.225 8.245 805.315 8.415 ;
        RECT 804.225 7.905 804.395 8.245 ;
        RECT 891.165 8.075 891.335 9.265 ;
        RECT 891.165 7.905 894.095 8.075 ;
        RECT 516.265 6.205 516.895 6.375 ;
        RECT 516.725 3.655 516.895 6.205 ;
        RECT 545.245 3.655 545.415 3.995 ;
        RECT 516.725 3.485 545.415 3.655 ;
        RECT 555.365 3.655 555.535 3.995 ;
        RECT 556.745 3.655 556.915 7.055 ;
        RECT 555.365 3.485 556.915 3.655 ;
        RECT 984.545 1.785 991.615 1.955 ;
      LAYER mcon ;
        RECT 805.145 8.245 805.315 8.415 ;
        RECT 893.925 7.905 894.095 8.075 ;
        RECT 556.745 6.885 556.915 7.055 ;
        RECT 545.245 3.825 545.415 3.995 ;
        RECT 555.365 3.825 555.535 3.995 ;
        RECT 991.445 1.785 991.615 1.955 ;
      LAYER met1 ;
        RECT 1897.110 3402.960 1897.430 3403.020 ;
        RECT 1908.150 3402.960 1908.470 3403.020 ;
        RECT 1897.110 3402.820 1908.470 3402.960 ;
        RECT 1897.110 3402.760 1897.430 3402.820 ;
        RECT 1908.150 3402.760 1908.470 3402.820 ;
        RECT 2318.930 3402.280 2319.250 3402.340 ;
        RECT 2333.190 3402.280 2333.510 3402.340 ;
        RECT 2318.930 3402.140 2333.510 3402.280 ;
        RECT 2318.930 3402.080 2319.250 3402.140 ;
        RECT 2333.190 3402.080 2333.510 3402.140 ;
        RECT 731.010 8.740 731.330 8.800 ;
        RECT 735.150 8.740 735.470 8.800 ;
        RECT 731.010 8.600 735.470 8.740 ;
        RECT 731.010 8.540 731.330 8.600 ;
        RECT 735.150 8.540 735.470 8.600 ;
        RECT 855.210 8.740 855.530 8.800 ;
        RECT 870.865 8.740 871.155 8.785 ;
        RECT 855.210 8.600 871.155 8.740 ;
        RECT 855.210 8.540 855.530 8.600 ;
        RECT 870.865 8.555 871.155 8.600 ;
        RECT 2374.590 8.740 2374.910 8.800 ;
        RECT 2406.330 8.740 2406.650 8.800 ;
        RECT 2374.590 8.600 2406.650 8.740 ;
        RECT 2374.590 8.540 2374.910 8.600 ;
        RECT 2406.330 8.540 2406.650 8.600 ;
        RECT 2444.970 8.740 2445.290 8.800 ;
        RECT 2508.910 8.740 2509.230 8.800 ;
        RECT 2444.970 8.600 2509.230 8.740 ;
        RECT 2444.970 8.540 2445.290 8.600 ;
        RECT 2508.910 8.540 2509.230 8.600 ;
        RECT 2561.810 8.740 2562.130 8.800 ;
        RECT 2646.910 8.740 2647.230 8.800 ;
        RECT 2561.810 8.600 2647.230 8.740 ;
        RECT 2561.810 8.540 2562.130 8.600 ;
        RECT 2646.910 8.540 2647.230 8.600 ;
        RECT 805.085 8.400 805.375 8.445 ;
        RECT 845.550 8.400 845.870 8.460 ;
        RECT 805.085 8.260 845.870 8.400 ;
        RECT 805.085 8.215 805.375 8.260 ;
        RECT 845.550 8.200 845.870 8.260 ;
        RECT 2078.350 8.400 2078.670 8.460 ;
        RECT 2093.990 8.400 2094.310 8.460 ;
        RECT 2078.350 8.260 2094.310 8.400 ;
        RECT 2078.350 8.200 2078.670 8.260 ;
        RECT 2093.990 8.200 2094.310 8.260 ;
        RECT 2161.610 8.400 2161.930 8.460 ;
        RECT 2218.190 8.400 2218.510 8.460 ;
        RECT 2161.610 8.260 2218.510 8.400 ;
        RECT 2161.610 8.200 2161.930 8.260 ;
        RECT 2218.190 8.200 2218.510 8.260 ;
        RECT 2266.490 8.400 2266.810 8.460 ;
        RECT 2314.330 8.400 2314.650 8.460 ;
        RECT 2266.490 8.260 2314.650 8.400 ;
        RECT 2266.490 8.200 2266.810 8.260 ;
        RECT 2314.330 8.200 2314.650 8.260 ;
        RECT 796.790 8.060 797.110 8.120 ;
        RECT 804.165 8.060 804.455 8.105 ;
        RECT 796.790 7.920 804.455 8.060 ;
        RECT 796.790 7.860 797.110 7.920 ;
        RECT 804.165 7.875 804.455 7.920 ;
        RECT 893.850 8.060 894.170 8.120 ;
        RECT 1977.150 8.060 1977.470 8.120 ;
        RECT 1993.250 8.060 1993.570 8.120 ;
        RECT 893.850 7.920 894.365 8.060 ;
        RECT 1977.150 7.920 1993.570 8.060 ;
        RECT 893.850 7.860 894.170 7.920 ;
        RECT 1977.150 7.860 1977.470 7.920 ;
        RECT 1993.250 7.860 1993.570 7.920 ;
        RECT 1997.850 8.060 1998.170 8.120 ;
        RECT 2018.550 8.060 2018.870 8.120 ;
        RECT 1997.850 7.920 2018.870 8.060 ;
        RECT 1997.850 7.860 1998.170 7.920 ;
        RECT 2018.550 7.860 2018.870 7.920 ;
        RECT 556.685 7.040 556.975 7.085 ;
        RECT 557.130 7.040 557.450 7.100 ;
        RECT 556.685 6.900 557.450 7.040 ;
        RECT 556.685 6.855 556.975 6.900 ;
        RECT 557.130 6.840 557.450 6.900 ;
        RECT 513.890 6.360 514.210 6.420 ;
        RECT 516.205 6.360 516.495 6.405 ;
        RECT 513.890 6.220 516.495 6.360 ;
        RECT 513.890 6.160 514.210 6.220 ;
        RECT 516.205 6.175 516.495 6.220 ;
        RECT 1120.170 5.680 1120.490 5.740 ;
        RECT 1125.230 5.680 1125.550 5.740 ;
        RECT 1120.170 5.540 1125.550 5.680 ;
        RECT 1120.170 5.480 1120.490 5.540 ;
        RECT 1125.230 5.480 1125.550 5.540 ;
        RECT 545.185 3.980 545.475 4.025 ;
        RECT 555.305 3.980 555.595 4.025 ;
        RECT 545.185 3.840 555.595 3.980 ;
        RECT 545.185 3.795 545.475 3.840 ;
        RECT 555.305 3.795 555.595 3.840 ;
        RECT 983.090 1.940 983.410 2.000 ;
        RECT 984.485 1.940 984.775 1.985 ;
        RECT 983.090 1.800 984.775 1.940 ;
        RECT 983.090 1.740 983.410 1.800 ;
        RECT 984.485 1.755 984.775 1.800 ;
        RECT 991.370 1.940 991.690 2.000 ;
        RECT 991.370 1.800 991.885 1.940 ;
        RECT 991.370 1.740 991.690 1.800 ;
      LAYER via ;
        RECT 1897.140 3402.760 1897.400 3403.020 ;
        RECT 1908.180 3402.760 1908.440 3403.020 ;
        RECT 2318.960 3402.080 2319.220 3402.340 ;
        RECT 2333.220 3402.080 2333.480 3402.340 ;
        RECT 731.040 8.540 731.300 8.800 ;
        RECT 735.180 8.540 735.440 8.800 ;
        RECT 855.240 8.540 855.500 8.800 ;
        RECT 2374.620 8.540 2374.880 8.800 ;
        RECT 2406.360 8.540 2406.620 8.800 ;
        RECT 2445.000 8.540 2445.260 8.800 ;
        RECT 2508.940 8.540 2509.200 8.800 ;
        RECT 2561.840 8.540 2562.100 8.800 ;
        RECT 2646.940 8.540 2647.200 8.800 ;
        RECT 845.580 8.200 845.840 8.460 ;
        RECT 2078.380 8.200 2078.640 8.460 ;
        RECT 2094.020 8.200 2094.280 8.460 ;
        RECT 2161.640 8.200 2161.900 8.460 ;
        RECT 2218.220 8.200 2218.480 8.460 ;
        RECT 2266.520 8.200 2266.780 8.460 ;
        RECT 2314.360 8.200 2314.620 8.460 ;
        RECT 796.820 7.860 797.080 8.120 ;
        RECT 893.880 7.860 894.140 8.120 ;
        RECT 1977.180 7.860 1977.440 8.120 ;
        RECT 1993.280 7.860 1993.540 8.120 ;
        RECT 1997.880 7.860 1998.140 8.120 ;
        RECT 2018.580 7.860 2018.840 8.120 ;
        RECT 557.160 6.840 557.420 7.100 ;
        RECT 513.920 6.160 514.180 6.420 ;
        RECT 1120.200 5.480 1120.460 5.740 ;
        RECT 1125.260 5.480 1125.520 5.740 ;
        RECT 983.120 1.740 983.380 2.000 ;
        RECT 991.400 1.740 991.660 2.000 ;
      LAYER met2 ;
        RECT 1626.130 3402.450 1626.410 3405.000 ;
        RECT 2823.570 3404.915 2823.850 3405.285 ;
        RECT 2197.510 3404.235 2197.790 3404.605 ;
        RECT 1897.130 3402.875 1897.410 3403.245 ;
        RECT 1897.140 3402.730 1897.400 3402.875 ;
        RECT 1908.180 3402.730 1908.440 3403.050 ;
        RECT 1628.030 3402.450 1628.310 3402.565 ;
        RECT 1626.130 3402.310 1628.310 3402.450 ;
        RECT 1626.130 3401.000 1626.410 3402.310 ;
        RECT 1628.030 3402.195 1628.310 3402.310 ;
        RECT 1908.240 3401.885 1908.380 3402.730 ;
        RECT 2197.580 3401.885 2197.720 3404.235 ;
        RECT 2719.150 3402.875 2719.430 3403.245 ;
        RECT 2318.960 3402.050 2319.220 3402.370 ;
        RECT 2333.210 3402.195 2333.490 3402.565 ;
        RECT 2333.220 3402.050 2333.480 3402.195 ;
        RECT 1908.170 3401.515 1908.450 3401.885 ;
        RECT 2197.510 3401.515 2197.790 3401.885 ;
        RECT 2318.490 3401.770 2318.770 3401.885 ;
        RECT 2319.020 3401.770 2319.160 3402.050 ;
        RECT 2719.220 3401.885 2719.360 3402.875 ;
        RECT 2823.640 3402.565 2823.780 3404.915 ;
        RECT 2823.570 3402.195 2823.850 3402.565 ;
        RECT 2318.490 3401.630 2319.160 3401.770 ;
        RECT 2318.490 3401.515 2318.770 3401.630 ;
        RECT 2719.150 3401.515 2719.430 3401.885 ;
        RECT 731.040 8.685 731.300 8.830 ;
        RECT 735.180 8.740 735.440 8.830 ;
        RECT 731.030 8.315 731.310 8.685 ;
        RECT 735.180 8.600 739.520 8.740 ;
        RECT 735.180 8.510 735.440 8.600 ;
        RECT 557.150 6.955 557.430 7.325 ;
        RECT 557.160 6.810 557.420 6.955 ;
        RECT 739.380 6.645 739.520 8.600 ;
        RECT 845.570 8.315 845.850 8.685 ;
        RECT 855.240 8.510 855.500 8.830 ;
        RECT 2374.620 8.685 2374.880 8.830 ;
        RECT 2406.360 8.685 2406.620 8.830 ;
        RECT 2445.000 8.685 2445.260 8.830 ;
        RECT 2508.940 8.685 2509.200 8.830 ;
        RECT 2561.840 8.685 2562.100 8.830 ;
        RECT 2646.940 8.685 2647.200 8.830 ;
        RECT 845.580 8.170 845.840 8.315 ;
        RECT 761.920 8.005 769.880 8.060 ;
        RECT 761.920 7.920 769.950 8.005 ;
        RECT 761.920 6.645 762.060 7.920 ;
        RECT 769.670 7.635 769.950 7.920 ;
        RECT 796.820 7.830 797.080 8.150 ;
        RECT 855.300 8.005 855.440 8.510 ;
        RECT 893.870 8.315 894.150 8.685 ;
        RECT 953.210 8.570 953.490 8.685 ;
        RECT 1428.850 8.570 1429.130 8.685 ;
        RECT 953.210 8.430 953.880 8.570 ;
        RECT 953.210 8.315 953.490 8.430 ;
        RECT 893.940 8.150 894.080 8.315 ;
        RECT 796.880 6.645 797.020 7.830 ;
        RECT 855.230 7.635 855.510 8.005 ;
        RECT 893.880 7.830 894.140 8.150 ;
        RECT 658.350 6.530 658.630 6.645 ;
        RECT 513.920 6.360 514.180 6.450 ;
        RECT 513.520 6.220 514.180 6.360 ;
        RECT 513.520 4.660 513.660 6.220 ;
        RECT 513.920 6.130 514.180 6.220 ;
        RECT 657.960 6.390 658.630 6.530 ;
        RECT 657.430 5.170 657.710 5.285 ;
        RECT 657.960 5.170 658.100 6.390 ;
        RECT 658.350 6.275 658.630 6.390 ;
        RECT 739.310 6.275 739.590 6.645 ;
        RECT 760.010 6.275 760.290 6.645 ;
        RECT 761.850 6.275 762.130 6.645 ;
        RECT 796.810 6.275 797.090 6.645 ;
        RECT 657.430 5.030 658.100 5.170 ;
        RECT 657.430 4.915 657.710 5.030 ;
        RECT 508.920 4.520 513.660 4.660 ;
        RECT 436.700 2.990 437.760 3.130 ;
        RECT 436.700 2.400 436.840 2.990 ;
        RECT 436.490 -4.800 437.050 2.400 ;
        RECT 437.620 1.205 437.760 2.990 ;
        RECT 437.550 0.835 437.830 1.205 ;
        RECT 508.920 0.525 509.060 4.520 ;
        RECT 755.870 4.490 756.150 4.605 ;
        RECT 760.080 4.490 760.220 6.275 ;
        RECT 755.870 4.350 760.220 4.490 ;
        RECT 953.740 4.490 953.880 8.430 ;
        RECT 1407.760 8.430 1429.130 8.570 ;
        RECT 1037.390 7.890 1037.670 8.005 ;
        RECT 959.720 7.750 961.240 7.890 ;
        RECT 959.720 4.490 959.860 7.750 ;
        RECT 953.740 4.350 959.860 4.490 ;
        RECT 755.870 4.235 756.150 4.350 ;
        RECT 961.100 3.980 961.240 7.750 ;
        RECT 1037.390 7.750 1039.440 7.890 ;
        RECT 1037.390 7.635 1037.670 7.750 ;
        RECT 1039.300 3.980 1039.440 7.750 ;
        RECT 1407.760 7.325 1407.900 8.430 ;
        RECT 1428.850 8.315 1429.130 8.430 ;
        RECT 1741.650 8.315 1741.930 8.685 ;
        RECT 1868.610 8.315 1868.890 8.685 ;
        RECT 1945.430 8.315 1945.710 8.685 ;
        RECT 1977.170 8.315 1977.450 8.685 ;
        RECT 1993.270 8.315 1993.550 8.685 ;
        RECT 1997.870 8.315 1998.150 8.685 ;
        RECT 2018.570 8.315 2018.850 8.685 ;
        RECT 2078.370 8.315 2078.650 8.685 ;
        RECT 2094.010 8.315 2094.290 8.685 ;
        RECT 2161.630 8.315 2161.910 8.685 ;
        RECT 2218.210 8.315 2218.490 8.685 ;
        RECT 2266.510 8.315 2266.790 8.685 ;
        RECT 2314.350 8.315 2314.630 8.685 ;
        RECT 2374.610 8.315 2374.890 8.685 ;
        RECT 2406.350 8.315 2406.630 8.685 ;
        RECT 2444.990 8.315 2445.270 8.685 ;
        RECT 2508.930 8.315 2509.210 8.685 ;
        RECT 2561.830 8.315 2562.110 8.685 ;
        RECT 2646.930 8.315 2647.210 8.685 ;
        RECT 1119.730 6.955 1120.010 7.325 ;
        RECT 1407.690 6.955 1407.970 7.325 ;
        RECT 1119.800 5.680 1119.940 6.955 ;
        RECT 1741.720 5.965 1741.860 8.315 ;
        RECT 1868.680 5.965 1868.820 8.315 ;
        RECT 1945.500 5.965 1945.640 8.315 ;
        RECT 1977.240 8.150 1977.380 8.315 ;
        RECT 1993.340 8.150 1993.480 8.315 ;
        RECT 1997.940 8.150 1998.080 8.315 ;
        RECT 2018.640 8.150 2018.780 8.315 ;
        RECT 2078.380 8.170 2078.640 8.315 ;
        RECT 2094.020 8.170 2094.280 8.315 ;
        RECT 2161.640 8.170 2161.900 8.315 ;
        RECT 2218.220 8.170 2218.480 8.315 ;
        RECT 2266.520 8.170 2266.780 8.315 ;
        RECT 2314.360 8.170 2314.620 8.315 ;
        RECT 1977.180 7.830 1977.440 8.150 ;
        RECT 1993.280 7.830 1993.540 8.150 ;
        RECT 1997.880 7.830 1998.140 8.150 ;
        RECT 2018.580 7.830 2018.840 8.150 ;
        RECT 1125.710 5.850 1125.990 5.965 ;
        RECT 1125.320 5.770 1125.990 5.850 ;
        RECT 1120.200 5.680 1120.460 5.770 ;
        RECT 1119.800 5.540 1120.460 5.680 ;
        RECT 1120.200 5.450 1120.460 5.540 ;
        RECT 1125.260 5.710 1125.990 5.770 ;
        RECT 1125.260 5.450 1125.520 5.710 ;
        RECT 1125.710 5.595 1125.990 5.710 ;
        RECT 1680.010 5.595 1680.290 5.965 ;
        RECT 1741.650 5.595 1741.930 5.965 ;
        RECT 1868.610 5.595 1868.890 5.965 ;
        RECT 1945.430 5.595 1945.710 5.965 ;
        RECT 1680.080 4.605 1680.220 5.595 ;
        RECT 1642.750 4.235 1643.030 4.605 ;
        RECT 1649.190 4.235 1649.470 4.605 ;
        RECT 1680.010 4.235 1680.290 4.605 ;
        RECT 961.100 3.840 968.600 3.980 ;
        RECT 968.460 3.810 968.600 3.840 ;
        RECT 1023.200 3.840 1039.440 3.980 ;
        RECT 968.460 3.670 973.200 3.810 ;
        RECT 973.060 3.300 973.200 3.670 ;
        RECT 973.060 3.160 979.180 3.300 ;
        RECT 979.040 1.940 979.180 3.160 ;
        RECT 994.220 2.990 1014.600 3.130 ;
        RECT 983.120 1.940 983.380 2.030 ;
        RECT 979.040 1.800 983.380 1.940 ;
        RECT 983.120 1.710 983.380 1.800 ;
        RECT 991.400 1.710 991.660 2.030 ;
        RECT 508.850 0.155 509.130 0.525 ;
        RECT 991.460 0.410 991.600 1.710 ;
        RECT 994.220 0.410 994.360 2.990 ;
        RECT 1014.460 1.770 1014.600 2.990 ;
        RECT 1016.300 2.990 1020.580 3.130 ;
        RECT 1016.300 1.770 1016.440 2.990 ;
        RECT 1020.440 2.450 1020.580 2.990 ;
        RECT 1023.200 2.450 1023.340 3.840 ;
        RECT 1642.820 3.810 1642.960 4.235 ;
        RECT 1649.260 3.810 1649.400 4.235 ;
        RECT 1642.820 3.670 1649.400 3.810 ;
        RECT 1020.440 2.310 1023.340 2.450 ;
        RECT 1014.460 1.630 1016.440 1.770 ;
        RECT 991.460 0.270 994.360 0.410 ;
      LAYER via2 ;
        RECT 2823.570 3404.960 2823.850 3405.240 ;
        RECT 2197.510 3404.280 2197.790 3404.560 ;
        RECT 1897.130 3402.920 1897.410 3403.200 ;
        RECT 1628.030 3402.240 1628.310 3402.520 ;
        RECT 2719.150 3402.920 2719.430 3403.200 ;
        RECT 2333.210 3402.240 2333.490 3402.520 ;
        RECT 1908.170 3401.560 1908.450 3401.840 ;
        RECT 2197.510 3401.560 2197.790 3401.840 ;
        RECT 2318.490 3401.560 2318.770 3401.840 ;
        RECT 2823.570 3402.240 2823.850 3402.520 ;
        RECT 2719.150 3401.560 2719.430 3401.840 ;
        RECT 731.030 8.360 731.310 8.640 ;
        RECT 557.150 7.000 557.430 7.280 ;
        RECT 845.570 8.360 845.850 8.640 ;
        RECT 769.670 7.680 769.950 7.960 ;
        RECT 893.870 8.360 894.150 8.640 ;
        RECT 953.210 8.360 953.490 8.640 ;
        RECT 855.230 7.680 855.510 7.960 ;
        RECT 657.430 4.960 657.710 5.240 ;
        RECT 658.350 6.320 658.630 6.600 ;
        RECT 739.310 6.320 739.590 6.600 ;
        RECT 760.010 6.320 760.290 6.600 ;
        RECT 761.850 6.320 762.130 6.600 ;
        RECT 796.810 6.320 797.090 6.600 ;
        RECT 437.550 0.880 437.830 1.160 ;
        RECT 755.870 4.280 756.150 4.560 ;
        RECT 1037.390 7.680 1037.670 7.960 ;
        RECT 1428.850 8.360 1429.130 8.640 ;
        RECT 1741.650 8.360 1741.930 8.640 ;
        RECT 1868.610 8.360 1868.890 8.640 ;
        RECT 1945.430 8.360 1945.710 8.640 ;
        RECT 1977.170 8.360 1977.450 8.640 ;
        RECT 1993.270 8.360 1993.550 8.640 ;
        RECT 1997.870 8.360 1998.150 8.640 ;
        RECT 2018.570 8.360 2018.850 8.640 ;
        RECT 2078.370 8.360 2078.650 8.640 ;
        RECT 2094.010 8.360 2094.290 8.640 ;
        RECT 2161.630 8.360 2161.910 8.640 ;
        RECT 2218.210 8.360 2218.490 8.640 ;
        RECT 2266.510 8.360 2266.790 8.640 ;
        RECT 2314.350 8.360 2314.630 8.640 ;
        RECT 2374.610 8.360 2374.890 8.640 ;
        RECT 2406.350 8.360 2406.630 8.640 ;
        RECT 2444.990 8.360 2445.270 8.640 ;
        RECT 2508.930 8.360 2509.210 8.640 ;
        RECT 2561.830 8.360 2562.110 8.640 ;
        RECT 2646.930 8.360 2647.210 8.640 ;
        RECT 1119.730 7.000 1120.010 7.280 ;
        RECT 1407.690 7.000 1407.970 7.280 ;
        RECT 1125.710 5.640 1125.990 5.920 ;
        RECT 1680.010 5.640 1680.290 5.920 ;
        RECT 1741.650 5.640 1741.930 5.920 ;
        RECT 1868.610 5.640 1868.890 5.920 ;
        RECT 1945.430 5.640 1945.710 5.920 ;
        RECT 1642.750 4.280 1643.030 4.560 ;
        RECT 1649.190 4.280 1649.470 4.560 ;
        RECT 1680.010 4.280 1680.290 4.560 ;
        RECT 508.850 0.200 509.130 0.480 ;
      LAYER met3 ;
        RECT 2752.910 3405.250 2753.290 3405.260 ;
        RECT 2823.545 3405.250 2823.875 3405.265 ;
        RECT 2752.910 3404.950 2823.875 3405.250 ;
        RECT 2752.910 3404.940 2753.290 3404.950 ;
        RECT 2823.545 3404.935 2823.875 3404.950 ;
        RECT 2173.310 3404.570 2173.690 3404.580 ;
        RECT 2197.485 3404.570 2197.815 3404.585 ;
        RECT 2173.310 3404.270 2197.815 3404.570 ;
        RECT 2173.310 3404.260 2173.690 3404.270 ;
        RECT 2197.485 3404.255 2197.815 3404.270 ;
        RECT 1821.910 3403.590 1830.490 3403.890 ;
        RECT 1628.005 3402.530 1628.335 3402.545 ;
        RECT 1821.910 3402.530 1822.210 3403.590 ;
        RECT 1628.005 3402.230 1822.210 3402.530 ;
        RECT 1628.005 3402.215 1628.335 3402.230 ;
        RECT 1830.190 3401.850 1830.490 3403.590 ;
        RECT 2090.550 3403.590 2098.210 3403.890 ;
        RECT 1897.105 3403.210 1897.435 3403.225 ;
        RECT 1849.510 3402.910 1897.435 3403.210 ;
        RECT 1849.510 3401.850 1849.810 3402.910 ;
        RECT 1897.105 3402.895 1897.435 3402.910 ;
        RECT 2090.550 3402.530 2090.850 3403.590 ;
        RECT 1967.270 3402.230 2017.250 3402.530 ;
        RECT 1830.190 3401.550 1849.810 3401.850 ;
        RECT 1908.145 3401.850 1908.475 3401.865 ;
        RECT 1967.270 3401.850 1967.570 3402.230 ;
        RECT 1908.145 3401.550 1967.570 3401.850 ;
        RECT 2016.950 3401.850 2017.250 3402.230 ;
        RECT 2062.950 3402.230 2090.850 3402.530 ;
        RECT 2062.950 3401.850 2063.250 3402.230 ;
        RECT 2016.950 3401.550 2063.250 3401.850 ;
        RECT 2097.910 3401.850 2098.210 3403.590 ;
        RECT 2283.750 3403.590 2291.410 3403.890 ;
        RECT 2173.310 3403.210 2173.690 3403.220 ;
        RECT 2139.310 3402.910 2173.690 3403.210 ;
        RECT 2139.310 3401.850 2139.610 3402.910 ;
        RECT 2173.310 3402.900 2173.690 3402.910 ;
        RECT 2283.750 3402.530 2284.050 3403.590 ;
        RECT 2256.150 3402.230 2284.050 3402.530 ;
        RECT 2097.910 3401.550 2139.610 3401.850 ;
        RECT 2197.485 3401.850 2197.815 3401.865 ;
        RECT 2256.150 3401.850 2256.450 3402.230 ;
        RECT 2197.485 3401.550 2256.450 3401.850 ;
        RECT 2291.110 3401.850 2291.410 3403.590 ;
        RECT 2670.150 3403.590 2677.810 3403.890 ;
        RECT 2333.185 3402.530 2333.515 3402.545 ;
        RECT 2670.150 3402.530 2670.450 3403.590 ;
        RECT 2333.185 3402.230 2479.090 3402.530 ;
        RECT 2333.185 3402.215 2333.515 3402.230 ;
        RECT 2318.465 3401.850 2318.795 3401.865 ;
        RECT 2291.110 3401.550 2318.795 3401.850 ;
        RECT 2478.790 3401.850 2479.090 3402.230 ;
        RECT 2525.710 3402.230 2670.450 3402.530 ;
        RECT 2525.710 3401.850 2526.010 3402.230 ;
        RECT 2478.790 3401.550 2526.010 3401.850 ;
        RECT 2677.510 3401.850 2677.810 3403.590 ;
        RECT 2719.125 3403.210 2719.455 3403.225 ;
        RECT 2752.910 3403.210 2753.290 3403.220 ;
        RECT 2719.125 3402.910 2753.290 3403.210 ;
        RECT 2719.125 3402.895 2719.455 3402.910 ;
        RECT 2752.910 3402.900 2753.290 3402.910 ;
        RECT 2823.545 3402.530 2823.875 3402.545 ;
        RECT 2835.710 3402.530 2836.090 3402.540 ;
        RECT 2823.545 3402.230 2836.090 3402.530 ;
        RECT 2823.545 3402.215 2823.875 3402.230 ;
        RECT 2835.710 3402.220 2836.090 3402.230 ;
        RECT 2719.125 3401.850 2719.455 3401.865 ;
        RECT 2677.510 3401.550 2719.455 3401.850 ;
        RECT 1908.145 3401.535 1908.475 3401.550 ;
        RECT 2197.485 3401.535 2197.815 3401.550 ;
        RECT 2318.465 3401.535 2318.795 3401.550 ;
        RECT 2719.125 3401.535 2719.455 3401.550 ;
        RECT 731.005 8.660 731.335 8.665 ;
        RECT 730.750 8.650 731.335 8.660 ;
        RECT 730.550 8.350 731.335 8.650 ;
        RECT 730.750 8.340 731.335 8.350 ;
        RECT 731.005 8.335 731.335 8.340 ;
        RECT 845.545 8.650 845.875 8.665 ;
        RECT 893.845 8.650 894.175 8.665 ;
        RECT 894.510 8.650 894.890 8.660 ;
        RECT 845.545 8.350 847.930 8.650 ;
        RECT 845.545 8.335 845.875 8.350 ;
        RECT 769.645 7.970 769.975 7.985 ;
        RECT 847.630 7.970 847.930 8.350 ;
        RECT 893.845 8.350 894.890 8.650 ;
        RECT 893.845 8.335 894.175 8.350 ;
        RECT 894.510 8.340 894.890 8.350 ;
        RECT 924.870 8.650 925.250 8.660 ;
        RECT 953.185 8.650 953.515 8.665 ;
        RECT 1039.870 8.650 1040.250 8.660 ;
        RECT 924.870 8.350 953.515 8.650 ;
        RECT 924.870 8.340 925.250 8.350 ;
        RECT 953.185 8.335 953.515 8.350 ;
        RECT 1037.380 8.350 1040.250 8.650 ;
        RECT 1037.380 7.985 1037.680 8.350 ;
        RECT 1039.870 8.340 1040.250 8.350 ;
        RECT 1360.950 8.650 1361.330 8.660 ;
        RECT 1394.990 8.650 1395.370 8.660 ;
        RECT 1360.950 8.350 1395.370 8.650 ;
        RECT 1360.950 8.340 1361.330 8.350 ;
        RECT 1394.990 8.340 1395.370 8.350 ;
        RECT 1428.825 8.650 1429.155 8.665 ;
        RECT 1470.430 8.650 1470.810 8.830 ;
        RECT 1428.825 8.510 1470.810 8.650 ;
        RECT 1741.625 8.650 1741.955 8.665 ;
        RECT 1868.585 8.650 1868.915 8.665 ;
        RECT 1428.825 8.350 1470.770 8.510 ;
        RECT 1741.625 8.350 1868.915 8.650 ;
        RECT 1428.825 8.335 1429.155 8.350 ;
        RECT 1741.625 8.335 1741.955 8.350 ;
        RECT 1868.585 8.335 1868.915 8.350 ;
        RECT 1945.405 8.650 1945.735 8.665 ;
        RECT 1977.145 8.650 1977.475 8.665 ;
        RECT 1945.405 8.350 1977.475 8.650 ;
        RECT 1945.405 8.335 1945.735 8.350 ;
        RECT 1977.145 8.335 1977.475 8.350 ;
        RECT 1993.245 8.650 1993.575 8.665 ;
        RECT 1997.845 8.650 1998.175 8.665 ;
        RECT 1993.245 8.350 1998.175 8.650 ;
        RECT 1993.245 8.335 1993.575 8.350 ;
        RECT 1997.845 8.335 1998.175 8.350 ;
        RECT 2018.545 8.650 2018.875 8.665 ;
        RECT 2078.345 8.650 2078.675 8.665 ;
        RECT 2018.545 8.350 2078.675 8.650 ;
        RECT 2018.545 8.335 2018.875 8.350 ;
        RECT 2078.345 8.335 2078.675 8.350 ;
        RECT 2093.985 8.650 2094.315 8.665 ;
        RECT 2161.605 8.650 2161.935 8.665 ;
        RECT 2093.985 8.350 2161.935 8.650 ;
        RECT 2093.985 8.335 2094.315 8.350 ;
        RECT 2161.605 8.335 2161.935 8.350 ;
        RECT 2218.185 8.650 2218.515 8.665 ;
        RECT 2266.485 8.650 2266.815 8.665 ;
        RECT 2218.185 8.350 2266.815 8.650 ;
        RECT 2218.185 8.335 2218.515 8.350 ;
        RECT 2266.485 8.335 2266.815 8.350 ;
        RECT 2314.325 8.650 2314.655 8.665 ;
        RECT 2374.585 8.650 2374.915 8.665 ;
        RECT 2314.325 8.350 2374.915 8.650 ;
        RECT 2314.325 8.335 2314.655 8.350 ;
        RECT 2374.585 8.335 2374.915 8.350 ;
        RECT 2406.325 8.650 2406.655 8.665 ;
        RECT 2444.965 8.650 2445.295 8.665 ;
        RECT 2406.325 8.350 2445.295 8.650 ;
        RECT 2406.325 8.335 2406.655 8.350 ;
        RECT 2444.965 8.335 2445.295 8.350 ;
        RECT 2508.905 8.650 2509.235 8.665 ;
        RECT 2561.805 8.650 2562.135 8.665 ;
        RECT 2508.905 8.350 2562.135 8.650 ;
        RECT 2508.905 8.335 2509.235 8.350 ;
        RECT 2561.805 8.335 2562.135 8.350 ;
        RECT 2646.905 8.650 2647.235 8.665 ;
        RECT 2835.710 8.650 2836.090 8.660 ;
        RECT 2646.905 8.350 2836.090 8.650 ;
        RECT 2646.905 8.335 2647.235 8.350 ;
        RECT 2835.710 8.340 2836.090 8.350 ;
        RECT 855.205 7.970 855.535 7.985 ;
        RECT 769.645 7.670 789.050 7.970 ;
        RECT 847.630 7.670 855.535 7.970 ;
        RECT 769.645 7.655 769.975 7.670 ;
        RECT 557.125 7.290 557.455 7.305 ;
        RECT 558.710 7.290 559.090 7.300 ;
        RECT 557.125 6.990 559.090 7.290 ;
        RECT 557.125 6.975 557.455 6.990 ;
        RECT 558.710 6.980 559.090 6.990 ;
        RECT 658.325 6.610 658.655 6.625 ;
        RECT 671.870 6.610 672.250 6.620 ;
        RECT 658.325 6.310 672.250 6.610 ;
        RECT 658.325 6.295 658.655 6.310 ;
        RECT 671.870 6.300 672.250 6.310 ;
        RECT 739.285 6.610 739.615 6.625 ;
        RECT 739.950 6.610 740.330 6.620 ;
        RECT 739.285 6.310 740.330 6.610 ;
        RECT 739.285 6.295 739.615 6.310 ;
        RECT 739.950 6.300 740.330 6.310 ;
        RECT 759.985 6.610 760.315 6.625 ;
        RECT 761.825 6.610 762.155 6.625 ;
        RECT 759.985 6.310 762.155 6.610 ;
        RECT 788.750 6.610 789.050 7.670 ;
        RECT 855.205 7.655 855.535 7.670 ;
        RECT 1037.365 7.655 1037.695 7.985 ;
        RECT 1050.910 7.970 1051.290 7.980 ;
        RECT 1291.950 7.970 1292.330 7.980 ;
        RECT 1309.430 7.970 1309.810 7.980 ;
        RECT 1050.910 7.670 1055.850 7.970 ;
        RECT 1050.910 7.660 1051.290 7.670 ;
        RECT 1055.550 7.290 1055.850 7.670 ;
        RECT 1291.950 7.670 1309.810 7.970 ;
        RECT 1291.950 7.660 1292.330 7.670 ;
        RECT 1309.430 7.660 1309.810 7.670 ;
        RECT 1060.110 7.290 1060.490 7.300 ;
        RECT 1055.550 6.990 1060.490 7.290 ;
        RECT 1060.110 6.980 1060.490 6.990 ;
        RECT 1091.390 7.290 1091.770 7.300 ;
        RECT 1119.705 7.290 1120.035 7.305 ;
        RECT 1091.390 6.990 1120.035 7.290 ;
        RECT 1091.390 6.980 1091.770 6.990 ;
        RECT 1119.705 6.975 1120.035 6.990 ;
        RECT 1233.990 7.290 1234.370 7.300 ;
        RECT 1244.110 7.290 1244.490 7.300 ;
        RECT 1233.990 6.990 1244.490 7.290 ;
        RECT 1233.990 6.980 1234.370 6.990 ;
        RECT 1244.110 6.980 1244.490 6.990 ;
        RECT 1406.950 7.290 1407.330 7.300 ;
        RECT 1407.665 7.290 1407.995 7.305 ;
        RECT 1406.950 6.990 1407.995 7.290 ;
        RECT 1406.950 6.980 1407.330 6.990 ;
        RECT 1407.665 6.975 1407.995 6.990 ;
        RECT 796.785 6.610 797.115 6.625 ;
        RECT 788.750 6.310 797.115 6.610 ;
        RECT 759.985 6.295 760.315 6.310 ;
        RECT 761.825 6.295 762.155 6.310 ;
        RECT 796.785 6.295 797.115 6.310 ;
        RECT 1125.685 5.940 1126.015 5.945 ;
        RECT 1060.110 5.930 1060.490 5.940 ;
        RECT 1088.630 5.930 1089.010 5.940 ;
        RECT 1060.110 5.630 1089.010 5.930 ;
        RECT 1060.110 5.620 1060.490 5.630 ;
        RECT 1088.630 5.620 1089.010 5.630 ;
        RECT 1125.430 5.930 1126.015 5.940 ;
        RECT 1484.230 5.930 1484.610 5.940 ;
        RECT 1544.030 5.930 1544.410 5.940 ;
        RECT 1125.430 5.630 1126.240 5.930 ;
        RECT 1484.230 5.630 1544.410 5.930 ;
        RECT 1125.430 5.620 1126.015 5.630 ;
        RECT 1484.230 5.620 1484.610 5.630 ;
        RECT 1544.030 5.620 1544.410 5.630 ;
        RECT 1679.985 5.930 1680.315 5.945 ;
        RECT 1741.625 5.930 1741.955 5.945 ;
        RECT 1679.985 5.630 1741.955 5.930 ;
        RECT 1125.685 5.615 1126.015 5.620 ;
        RECT 1679.985 5.615 1680.315 5.630 ;
        RECT 1741.625 5.615 1741.955 5.630 ;
        RECT 1868.585 5.930 1868.915 5.945 ;
        RECT 1945.405 5.930 1945.735 5.945 ;
        RECT 1868.585 5.630 1945.735 5.930 ;
        RECT 1868.585 5.615 1868.915 5.630 ;
        RECT 1945.405 5.615 1945.735 5.630 ;
        RECT 620.350 5.250 620.730 5.260 ;
        RECT 643.350 5.250 643.730 5.260 ;
        RECT 620.350 4.950 643.730 5.250 ;
        RECT 620.350 4.940 620.730 4.950 ;
        RECT 643.350 4.940 643.730 4.950 ;
        RECT 649.790 5.250 650.170 5.260 ;
        RECT 657.405 5.250 657.735 5.265 ;
        RECT 649.790 4.950 657.735 5.250 ;
        RECT 649.790 4.940 650.170 4.950 ;
        RECT 657.405 4.935 657.735 4.950 ;
        RECT 754.670 4.570 755.050 4.580 ;
        RECT 755.845 4.570 756.175 4.585 ;
        RECT 1642.725 4.580 1643.055 4.585 ;
        RECT 754.670 4.270 756.175 4.570 ;
        RECT 754.670 4.260 755.050 4.270 ;
        RECT 755.845 4.255 756.175 4.270 ;
        RECT 1574.390 4.570 1574.770 4.580 ;
        RECT 1641.550 4.570 1641.930 4.580 ;
        RECT 1574.390 4.270 1641.930 4.570 ;
        RECT 1574.390 4.260 1574.770 4.270 ;
        RECT 1641.550 4.260 1641.930 4.270 ;
        RECT 1642.700 4.570 1643.080 4.580 ;
        RECT 1649.165 4.570 1649.495 4.585 ;
        RECT 1679.985 4.570 1680.315 4.585 ;
        RECT 1642.700 4.270 1643.510 4.570 ;
        RECT 1649.165 4.270 1680.315 4.570 ;
        RECT 1642.700 4.260 1643.080 4.270 ;
        RECT 1642.725 4.255 1643.055 4.260 ;
        RECT 1649.165 4.255 1649.495 4.270 ;
        RECT 1679.985 4.255 1680.315 4.270 ;
        RECT 437.525 1.170 437.855 1.185 ;
        RECT 464.870 1.170 465.250 1.180 ;
        RECT 437.525 0.870 465.250 1.170 ;
        RECT 437.525 0.855 437.855 0.870 ;
        RECT 464.870 0.860 465.250 0.870 ;
        RECT 507.190 0.490 507.570 0.500 ;
        RECT 508.825 0.490 509.155 0.505 ;
        RECT 507.190 0.190 509.155 0.490 ;
        RECT 507.190 0.180 507.570 0.190 ;
        RECT 508.825 0.175 509.155 0.190 ;
      LAYER via3 ;
        RECT 2752.940 3404.940 2753.260 3405.260 ;
        RECT 2173.340 3404.260 2173.660 3404.580 ;
        RECT 2173.340 3402.900 2173.660 3403.220 ;
        RECT 2752.940 3402.900 2753.260 3403.220 ;
        RECT 2835.740 3402.220 2836.060 3402.540 ;
        RECT 730.780 8.340 731.100 8.660 ;
        RECT 894.540 8.340 894.860 8.660 ;
        RECT 924.900 8.340 925.220 8.660 ;
        RECT 1039.900 8.340 1040.220 8.660 ;
        RECT 1360.980 8.340 1361.300 8.660 ;
        RECT 1395.020 8.340 1395.340 8.660 ;
        RECT 1470.460 8.510 1470.780 8.830 ;
        RECT 2835.740 8.340 2836.060 8.660 ;
        RECT 558.740 6.980 559.060 7.300 ;
        RECT 671.900 6.300 672.220 6.620 ;
        RECT 739.980 6.300 740.300 6.620 ;
        RECT 1050.940 7.660 1051.260 7.980 ;
        RECT 1291.980 7.660 1292.300 7.980 ;
        RECT 1309.460 7.660 1309.780 7.980 ;
        RECT 1060.140 6.980 1060.460 7.300 ;
        RECT 1091.420 6.980 1091.740 7.300 ;
        RECT 1234.020 6.980 1234.340 7.300 ;
        RECT 1244.140 6.980 1244.460 7.300 ;
        RECT 1406.980 6.980 1407.300 7.300 ;
        RECT 1060.140 5.620 1060.460 5.940 ;
        RECT 1088.660 5.620 1088.980 5.940 ;
        RECT 1125.460 5.620 1125.780 5.940 ;
        RECT 1484.260 5.620 1484.580 5.940 ;
        RECT 1544.060 5.620 1544.380 5.940 ;
        RECT 620.380 4.940 620.700 5.260 ;
        RECT 643.380 4.940 643.700 5.260 ;
        RECT 649.820 4.940 650.140 5.260 ;
        RECT 754.700 4.260 755.020 4.580 ;
        RECT 1574.420 4.260 1574.740 4.580 ;
        RECT 1641.580 4.260 1641.900 4.580 ;
        RECT 1642.730 4.260 1643.050 4.580 ;
        RECT 464.900 0.860 465.220 1.180 ;
        RECT 507.220 0.180 507.540 0.500 ;
      LAYER met4 ;
        RECT 2752.935 3404.935 2753.265 3405.265 ;
        RECT 2173.335 3404.255 2173.665 3404.585 ;
        RECT 2173.350 3403.225 2173.650 3404.255 ;
        RECT 2752.950 3403.225 2753.250 3404.935 ;
        RECT 2173.335 3402.895 2173.665 3403.225 ;
        RECT 2752.935 3402.895 2753.265 3403.225 ;
        RECT 2835.735 3402.215 2836.065 3402.545 ;
        RECT 697.670 11.750 727.410 12.050 ;
        RECT 681.110 9.030 683.250 9.330 ;
        RECT 558.735 7.290 559.065 7.305 ;
        RECT 681.110 7.290 681.410 9.030 ;
        RECT 682.950 8.650 683.250 9.030 ;
        RECT 682.950 8.350 684.170 8.650 ;
        RECT 558.735 6.990 559.970 7.290 ;
        RECT 558.735 6.975 559.065 6.990 ;
        RECT 559.670 5.250 559.970 6.990 ;
        RECT 676.510 6.990 681.410 7.290 ;
        RECT 671.895 6.610 672.225 6.625 ;
        RECT 676.510 6.610 676.810 6.990 ;
        RECT 671.895 6.310 676.810 6.610 ;
        RECT 671.895 6.295 672.225 6.310 ;
        RECT 683.870 5.930 684.170 8.350 ;
        RECT 697.670 6.610 697.970 11.750 ;
        RECT 727.110 9.330 727.410 11.750 ;
        RECT 1395.030 11.750 1402.690 12.050 ;
        RECT 727.110 9.030 730.170 9.330 ;
        RECT 729.870 8.650 730.170 9.030 ;
        RECT 1311.310 9.030 1332.770 9.330 ;
        RECT 730.775 8.650 731.105 8.665 ;
        RECT 729.870 8.350 731.105 8.650 ;
        RECT 730.775 8.335 731.105 8.350 ;
        RECT 894.535 8.650 894.865 8.665 ;
        RECT 924.895 8.650 925.225 8.665 ;
        RECT 894.535 8.350 925.225 8.650 ;
        RECT 894.535 8.335 894.865 8.350 ;
        RECT 924.895 8.335 925.225 8.350 ;
        RECT 1039.895 8.335 1040.225 8.665 ;
        RECT 1039.910 7.970 1040.210 8.335 ;
        RECT 1050.935 7.970 1051.265 7.985 ;
        RECT 1291.975 7.970 1292.305 7.985 ;
        RECT 1039.910 7.670 1051.265 7.970 ;
        RECT 1050.935 7.655 1051.265 7.670 ;
        RECT 1226.670 7.670 1234.330 7.970 ;
        RECT 1060.135 6.975 1060.465 7.305 ;
        RECT 1091.415 6.975 1091.745 7.305 ;
        RECT 696.750 6.310 697.970 6.610 ;
        RECT 696.750 5.930 697.050 6.310 ;
        RECT 739.975 6.295 740.305 6.625 ;
        RECT 683.870 5.630 697.050 5.930 ;
        RECT 739.990 5.690 740.290 6.295 ;
        RECT 1060.150 5.945 1060.450 6.975 ;
        RECT 1091.430 6.610 1091.730 6.975 ;
        RECT 1226.670 6.610 1226.970 7.670 ;
        RECT 1234.030 7.305 1234.330 7.670 ;
        RECT 1269.910 7.670 1292.305 7.970 ;
        RECT 1234.015 6.975 1234.345 7.305 ;
        RECT 1244.135 6.975 1244.465 7.305 ;
        RECT 1088.670 6.310 1091.730 6.610 ;
        RECT 1157.670 6.310 1168.090 6.610 ;
        RECT 1088.670 5.945 1088.970 6.310 ;
        RECT 620.375 5.250 620.705 5.265 ;
        RECT 559.670 4.950 562.730 5.250 ;
        RECT 562.430 3.890 562.730 4.950 ;
        RECT 587.270 4.950 617.930 5.250 ;
        RECT 587.270 3.890 587.570 4.950 ;
        RECT 617.630 4.570 617.930 4.950 ;
        RECT 619.470 4.950 620.705 5.250 ;
        RECT 619.470 4.570 619.770 4.950 ;
        RECT 620.375 4.935 620.705 4.950 ;
        RECT 643.375 5.250 643.705 5.265 ;
        RECT 649.815 5.250 650.145 5.265 ;
        RECT 643.375 4.950 650.145 5.250 ;
        RECT 643.375 4.935 643.705 4.950 ;
        RECT 649.815 4.935 650.145 4.950 ;
        RECT 617.630 4.270 619.770 4.570 ;
        RECT 739.550 4.510 740.730 5.690 ;
        RECT 751.510 4.510 752.690 5.690 ;
        RECT 1060.135 5.615 1060.465 5.945 ;
        RECT 1088.655 5.615 1088.985 5.945 ;
        RECT 1125.455 5.615 1125.785 5.945 ;
        RECT 562.430 3.590 587.570 3.890 ;
        RECT 751.950 3.890 752.250 4.510 ;
        RECT 754.695 4.255 755.025 4.585 ;
        RECT 754.710 3.890 755.010 4.255 ;
        RECT 751.950 3.590 755.010 3.890 ;
        RECT 1125.470 3.210 1125.770 5.615 ;
        RECT 1157.670 3.210 1157.970 6.310 ;
        RECT 1167.790 3.890 1168.090 6.310 ;
        RECT 1170.550 6.310 1226.970 6.610 ;
        RECT 1170.550 3.890 1170.850 6.310 ;
        RECT 1167.790 3.590 1170.850 3.890 ;
        RECT 1125.470 2.910 1157.970 3.210 ;
        RECT 1244.150 3.210 1244.450 6.975 ;
        RECT 1269.910 3.890 1270.210 7.670 ;
        RECT 1291.975 7.655 1292.305 7.670 ;
        RECT 1309.455 7.970 1309.785 7.985 ;
        RECT 1311.310 7.970 1311.610 9.030 ;
        RECT 1332.470 8.650 1332.770 9.030 ;
        RECT 1338.910 9.030 1361.290 9.330 ;
        RECT 1338.910 8.650 1339.210 9.030 ;
        RECT 1360.990 8.665 1361.290 9.030 ;
        RECT 1395.030 8.665 1395.330 11.750 ;
        RECT 1402.390 9.330 1402.690 11.750 ;
        RECT 1402.390 9.030 1406.370 9.330 ;
        RECT 1332.470 8.350 1339.210 8.650 ;
        RECT 1360.975 8.335 1361.305 8.665 ;
        RECT 1395.015 8.335 1395.345 8.665 ;
        RECT 1309.455 7.670 1311.610 7.970 ;
        RECT 1309.455 7.655 1309.785 7.670 ;
        RECT 1406.070 7.290 1406.370 9.030 ;
        RECT 1470.455 8.505 1470.785 8.835 ;
        RECT 2835.750 8.665 2836.050 3402.215 ;
        RECT 1470.470 7.970 1470.770 8.505 ;
        RECT 2835.735 8.335 2836.065 8.665 ;
        RECT 1470.470 7.670 1479.050 7.970 ;
        RECT 1406.975 7.290 1407.305 7.305 ;
        RECT 1406.070 6.990 1407.305 7.290 ;
        RECT 1406.975 6.975 1407.305 6.990 ;
        RECT 1478.750 5.930 1479.050 7.670 ;
        RECT 1484.255 5.930 1484.585 5.945 ;
        RECT 1478.750 5.630 1484.585 5.930 ;
        RECT 1484.255 5.615 1484.585 5.630 ;
        RECT 1544.055 5.930 1544.385 5.945 ;
        RECT 1544.055 5.630 1550.810 5.930 ;
        RECT 1544.055 5.615 1544.385 5.630 ;
        RECT 1550.510 4.570 1550.810 5.630 ;
        RECT 1574.415 4.570 1574.745 4.585 ;
        RECT 1550.510 4.270 1574.745 4.570 ;
        RECT 1574.415 4.255 1574.745 4.270 ;
        RECT 1641.575 4.255 1641.905 4.585 ;
        RECT 1642.725 4.255 1643.055 4.585 ;
        RECT 1263.470 3.590 1270.210 3.890 ;
        RECT 1263.470 3.210 1263.770 3.590 ;
        RECT 1244.150 2.910 1263.770 3.210 ;
        RECT 1641.590 3.210 1641.890 4.255 ;
        RECT 1642.740 3.210 1643.040 4.255 ;
        RECT 1641.590 2.910 1643.040 3.210 ;
        RECT 464.895 0.855 465.225 1.185 ;
        RECT 464.910 0.490 465.210 0.855 ;
        RECT 507.215 0.490 507.545 0.505 ;
        RECT 464.910 0.190 507.545 0.490 ;
        RECT 507.215 0.175 507.545 0.190 ;
      LAYER met5 ;
        RECT 739.340 4.300 752.900 5.900 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 585.265 6.885 602.455 7.055 ;
        RECT 604.585 6.885 606.595 7.055 ;
        RECT 488.205 5.525 504.935 5.695 ;
        RECT 472.105 2.465 484.235 2.635 ;
        RECT 463.365 1.615 463.535 1.955 ;
        RECT 472.105 1.615 472.275 2.465 ;
        RECT 484.065 1.955 484.235 2.465 ;
        RECT 488.205 1.955 488.375 5.525 ;
        RECT 504.765 5.185 504.935 5.525 ;
        RECT 559.045 5.185 560.595 5.355 ;
        RECT 582.045 4.675 582.215 5.355 ;
        RECT 582.045 4.505 583.595 4.675 ;
        RECT 585.265 4.505 585.435 6.885 ;
        RECT 606.425 5.185 606.595 6.885 ;
        RECT 618.385 5.525 619.475 5.695 ;
        RECT 615.165 5.015 615.335 5.355 ;
        RECT 618.385 5.015 618.555 5.525 ;
        RECT 615.165 4.845 618.555 5.015 ;
        RECT 619.305 5.015 619.475 5.525 ;
        RECT 700.265 5.185 703.195 5.355 ;
        RECT 619.305 4.845 620.395 5.015 ;
        RECT 737.065 4.505 737.235 5.355 ;
        RECT 747.185 4.505 747.355 5.355 ;
        RECT 896.685 5.185 898.235 5.355 ;
        RECT 1124.845 5.015 1125.015 5.355 ;
        RECT 1127.145 5.015 1127.315 5.355 ;
        RECT 1124.845 4.845 1127.315 5.015 ;
        RECT 1195.225 5.015 1195.395 5.355 ;
        RECT 1196.605 5.015 1196.775 5.355 ;
        RECT 1227.425 5.185 1241.855 5.355 ;
        RECT 1710.885 5.185 1716.115 5.355 ;
        RECT 1195.225 4.845 1196.775 5.015 ;
        RECT 1715.945 4.505 1716.115 5.185 ;
        RECT 1821.285 4.505 1821.455 5.355 ;
        RECT 1892.125 4.165 1892.295 5.355 ;
        RECT 1968.025 5.185 1968.195 7.395 ;
        RECT 484.065 1.785 488.375 1.955 ;
        RECT 463.365 1.445 472.275 1.615 ;
      LAYER mcon ;
        RECT 1968.025 7.225 1968.195 7.395 ;
        RECT 602.285 6.885 602.455 7.055 ;
        RECT 463.365 1.785 463.535 1.955 ;
        RECT 560.425 5.185 560.595 5.355 ;
        RECT 582.045 5.185 582.215 5.355 ;
        RECT 615.165 5.185 615.335 5.355 ;
        RECT 703.025 5.185 703.195 5.355 ;
        RECT 737.065 5.185 737.235 5.355 ;
        RECT 620.225 4.845 620.395 5.015 ;
        RECT 583.425 4.505 583.595 4.675 ;
        RECT 747.185 5.185 747.355 5.355 ;
        RECT 898.065 5.185 898.235 5.355 ;
        RECT 1124.845 5.185 1125.015 5.355 ;
        RECT 1127.145 5.185 1127.315 5.355 ;
        RECT 1195.225 5.185 1195.395 5.355 ;
        RECT 1196.605 5.185 1196.775 5.355 ;
        RECT 1241.685 5.185 1241.855 5.355 ;
        RECT 1821.285 5.185 1821.455 5.355 ;
        RECT 1892.125 5.185 1892.295 5.355 ;
      LAYER met1 ;
        RECT 1967.965 7.380 1968.255 7.425 ;
        RECT 2259.590 7.380 2259.910 7.440 ;
        RECT 1967.965 7.240 2259.910 7.380 ;
        RECT 1967.965 7.195 1968.255 7.240 ;
        RECT 2259.590 7.180 2259.910 7.240 ;
        RECT 602.225 7.040 602.515 7.085 ;
        RECT 604.525 7.040 604.815 7.085 ;
        RECT 602.225 6.900 604.815 7.040 ;
        RECT 602.225 6.855 602.515 6.900 ;
        RECT 604.525 6.855 604.815 6.900 ;
        RECT 504.705 5.340 504.995 5.385 ;
        RECT 558.985 5.340 559.275 5.385 ;
        RECT 504.705 5.200 559.275 5.340 ;
        RECT 504.705 5.155 504.995 5.200 ;
        RECT 558.985 5.155 559.275 5.200 ;
        RECT 560.365 5.340 560.655 5.385 ;
        RECT 581.985 5.340 582.275 5.385 ;
        RECT 560.365 5.200 582.275 5.340 ;
        RECT 560.365 5.155 560.655 5.200 ;
        RECT 581.985 5.155 582.275 5.200 ;
        RECT 606.365 5.340 606.655 5.385 ;
        RECT 615.105 5.340 615.395 5.385 ;
        RECT 700.205 5.340 700.495 5.385 ;
        RECT 606.365 5.200 615.395 5.340 ;
        RECT 606.365 5.155 606.655 5.200 ;
        RECT 615.105 5.155 615.395 5.200 ;
        RECT 621.160 5.200 700.495 5.340 ;
        RECT 620.165 5.000 620.455 5.045 ;
        RECT 621.160 5.000 621.300 5.200 ;
        RECT 700.205 5.155 700.495 5.200 ;
        RECT 702.965 5.340 703.255 5.385 ;
        RECT 737.005 5.340 737.295 5.385 ;
        RECT 702.965 5.200 737.295 5.340 ;
        RECT 702.965 5.155 703.255 5.200 ;
        RECT 737.005 5.155 737.295 5.200 ;
        RECT 747.125 5.340 747.415 5.385 ;
        RECT 896.625 5.340 896.915 5.385 ;
        RECT 747.125 5.200 896.915 5.340 ;
        RECT 747.125 5.155 747.415 5.200 ;
        RECT 896.625 5.155 896.915 5.200 ;
        RECT 898.005 5.340 898.295 5.385 ;
        RECT 1124.785 5.340 1125.075 5.385 ;
        RECT 898.005 5.200 1125.075 5.340 ;
        RECT 898.005 5.155 898.295 5.200 ;
        RECT 1124.785 5.155 1125.075 5.200 ;
        RECT 1127.085 5.340 1127.375 5.385 ;
        RECT 1195.165 5.340 1195.455 5.385 ;
        RECT 1127.085 5.200 1195.455 5.340 ;
        RECT 1127.085 5.155 1127.375 5.200 ;
        RECT 1195.165 5.155 1195.455 5.200 ;
        RECT 1196.545 5.340 1196.835 5.385 ;
        RECT 1227.365 5.340 1227.655 5.385 ;
        RECT 1196.545 5.200 1227.655 5.340 ;
        RECT 1196.545 5.155 1196.835 5.200 ;
        RECT 1227.365 5.155 1227.655 5.200 ;
        RECT 1241.625 5.340 1241.915 5.385 ;
        RECT 1710.825 5.340 1711.115 5.385 ;
        RECT 1760.950 5.340 1761.270 5.400 ;
        RECT 1241.625 5.200 1711.115 5.340 ;
        RECT 1241.625 5.155 1241.915 5.200 ;
        RECT 1710.825 5.155 1711.115 5.200 ;
        RECT 1728.380 5.200 1761.270 5.340 ;
        RECT 620.165 4.860 621.300 5.000 ;
        RECT 620.165 4.815 620.455 4.860 ;
        RECT 583.365 4.660 583.655 4.705 ;
        RECT 585.205 4.660 585.495 4.705 ;
        RECT 583.365 4.520 585.495 4.660 ;
        RECT 583.365 4.475 583.655 4.520 ;
        RECT 585.205 4.475 585.495 4.520 ;
        RECT 737.005 4.660 737.295 4.705 ;
        RECT 747.125 4.660 747.415 4.705 ;
        RECT 737.005 4.520 747.415 4.660 ;
        RECT 737.005 4.475 737.295 4.520 ;
        RECT 747.125 4.475 747.415 4.520 ;
        RECT 1715.885 4.660 1716.175 4.705 ;
        RECT 1728.380 4.660 1728.520 5.200 ;
        RECT 1760.950 5.140 1761.270 5.200 ;
        RECT 1821.225 5.340 1821.515 5.385 ;
        RECT 1863.990 5.340 1864.310 5.400 ;
        RECT 1821.225 5.200 1864.310 5.340 ;
        RECT 1821.225 5.155 1821.515 5.200 ;
        RECT 1863.990 5.140 1864.310 5.200 ;
        RECT 1892.065 5.340 1892.355 5.385 ;
        RECT 1967.965 5.340 1968.255 5.385 ;
        RECT 1892.065 5.200 1968.255 5.340 ;
        RECT 1892.065 5.155 1892.355 5.200 ;
        RECT 1967.965 5.155 1968.255 5.200 ;
        RECT 1715.885 4.520 1728.520 4.660 ;
        RECT 1781.190 4.660 1781.510 4.720 ;
        RECT 1821.225 4.660 1821.515 4.705 ;
        RECT 1781.190 4.520 1821.515 4.660 ;
        RECT 1715.885 4.475 1716.175 4.520 ;
        RECT 1781.190 4.460 1781.510 4.520 ;
        RECT 1821.225 4.475 1821.515 4.520 ;
        RECT 1865.370 4.320 1865.690 4.380 ;
        RECT 1892.065 4.320 1892.355 4.365 ;
        RECT 1865.370 4.180 1892.355 4.320 ;
        RECT 1865.370 4.120 1865.690 4.180 ;
        RECT 1892.065 4.135 1892.355 4.180 ;
        RECT 455.470 1.940 455.790 2.000 ;
        RECT 463.305 1.940 463.595 1.985 ;
        RECT 455.470 1.800 463.595 1.940 ;
        RECT 455.470 1.740 455.790 1.800 ;
        RECT 463.305 1.755 463.595 1.800 ;
      LAYER via ;
        RECT 2259.620 7.180 2259.880 7.440 ;
        RECT 1760.980 5.140 1761.240 5.400 ;
        RECT 1864.020 5.140 1864.280 5.400 ;
        RECT 1781.220 4.460 1781.480 4.720 ;
        RECT 1865.400 4.120 1865.660 4.380 ;
        RECT 455.500 1.740 455.760 2.000 ;
      LAYER met2 ;
        RECT 2259.620 7.210 2259.880 7.470 ;
        RECT 2260.930 7.210 2261.210 9.000 ;
        RECT 2259.620 7.150 2261.210 7.210 ;
        RECT 2259.680 7.070 2261.210 7.150 ;
        RECT 1760.980 5.110 1761.240 5.430 ;
        RECT 1864.020 5.170 1864.280 5.430 ;
        RECT 1864.020 5.110 1865.600 5.170 ;
        RECT 1761.040 4.605 1761.180 5.110 ;
        RECT 1864.080 5.030 1865.600 5.110 ;
        RECT 1781.220 4.605 1781.480 4.750 ;
        RECT 1760.970 4.235 1761.250 4.605 ;
        RECT 1781.210 4.235 1781.490 4.605 ;
        RECT 1865.460 4.410 1865.600 5.030 ;
        RECT 2260.930 5.000 2261.210 7.070 ;
        RECT 1865.400 4.090 1865.660 4.410 ;
        RECT 454.640 2.820 455.700 2.960 ;
        RECT 454.640 2.400 454.780 2.820 ;
        RECT 454.430 -4.800 454.990 2.400 ;
        RECT 455.560 2.030 455.700 2.820 ;
        RECT 455.500 1.710 455.760 2.030 ;
      LAYER via2 ;
        RECT 1760.970 4.280 1761.250 4.560 ;
        RECT 1781.210 4.280 1781.490 4.560 ;
      LAYER met3 ;
        RECT 1760.945 4.570 1761.275 4.585 ;
        RECT 1781.185 4.570 1781.515 4.585 ;
        RECT 1760.945 4.270 1781.515 4.570 ;
        RECT 1760.945 4.255 1761.275 4.270 ;
        RECT 1781.185 4.255 1781.515 4.270 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 7.045 990.165 7.215 1084.175 ;
        RECT 5.665 480.165 5.835 693.515 ;
        RECT 7.965 361.505 8.135 480.335 ;
        RECT 8.885 238.085 9.055 361.675 ;
        RECT 4.285 51.425 4.455 85.595 ;
        RECT 8.425 85.425 8.595 217.515 ;
        RECT 9.805 217.345 9.975 238.255 ;
        RECT 7.965 5.865 8.135 51.595 ;
        RECT 25.905 5.865 26.995 6.035 ;
        RECT 34.645 5.865 34.815 7.395 ;
        RECT 462.905 3.825 463.995 3.995 ;
        RECT 463.825 1.955 463.995 3.825 ;
        RECT 463.825 1.785 464.455 1.955 ;
      LAYER mcon ;
        RECT 7.045 1084.005 7.215 1084.175 ;
        RECT 5.665 693.345 5.835 693.515 ;
        RECT 7.965 480.165 8.135 480.335 ;
        RECT 8.885 361.505 9.055 361.675 ;
        RECT 9.805 238.085 9.975 238.255 ;
        RECT 8.425 217.345 8.595 217.515 ;
        RECT 4.285 85.425 4.455 85.595 ;
        RECT 7.965 51.425 8.135 51.595 ;
        RECT 34.645 7.225 34.815 7.395 ;
        RECT 26.825 5.865 26.995 6.035 ;
        RECT 464.285 1.785 464.455 1.955 ;
      LAYER met1 ;
        RECT 0.530 1084.160 0.850 1084.220 ;
        RECT 6.985 1084.160 7.275 1084.205 ;
        RECT 0.530 1084.020 7.275 1084.160 ;
        RECT 0.530 1083.960 0.850 1084.020 ;
        RECT 6.985 1083.975 7.275 1084.020 ;
        RECT 6.970 990.320 7.290 990.380 ;
        RECT 6.970 990.180 7.485 990.320 ;
        RECT 6.970 990.120 7.290 990.180 ;
        RECT 6.050 859.760 6.370 859.820 ;
        RECT 6.970 859.760 7.290 859.820 ;
        RECT 6.050 859.620 7.290 859.760 ;
        RECT 6.050 859.560 6.370 859.620 ;
        RECT 6.970 859.560 7.290 859.620 ;
        RECT 5.605 693.500 5.895 693.545 ;
        RECT 6.510 693.500 6.830 693.560 ;
        RECT 5.605 693.360 6.830 693.500 ;
        RECT 5.605 693.315 5.895 693.360 ;
        RECT 6.510 693.300 6.830 693.360 ;
        RECT 5.605 480.320 5.895 480.365 ;
        RECT 7.905 480.320 8.195 480.365 ;
        RECT 5.605 480.180 8.195 480.320 ;
        RECT 5.605 480.135 5.895 480.180 ;
        RECT 7.905 480.135 8.195 480.180 ;
        RECT 7.905 361.660 8.195 361.705 ;
        RECT 8.825 361.660 9.115 361.705 ;
        RECT 7.905 361.520 9.115 361.660 ;
        RECT 7.905 361.475 8.195 361.520 ;
        RECT 8.825 361.475 9.115 361.520 ;
        RECT 8.825 238.240 9.115 238.285 ;
        RECT 9.745 238.240 10.035 238.285 ;
        RECT 8.825 238.100 10.035 238.240 ;
        RECT 8.825 238.055 9.115 238.100 ;
        RECT 9.745 238.055 10.035 238.100 ;
        RECT 8.365 217.500 8.655 217.545 ;
        RECT 9.745 217.500 10.035 217.545 ;
        RECT 8.365 217.360 10.035 217.500 ;
        RECT 8.365 217.315 8.655 217.360 ;
        RECT 9.745 217.315 10.035 217.360 ;
        RECT 4.225 85.580 4.515 85.625 ;
        RECT 8.365 85.580 8.655 85.625 ;
        RECT 4.225 85.440 8.655 85.580 ;
        RECT 4.225 85.395 4.515 85.440 ;
        RECT 8.365 85.395 8.655 85.440 ;
        RECT 4.225 51.580 4.515 51.625 ;
        RECT 7.905 51.580 8.195 51.625 ;
        RECT 4.225 51.440 8.195 51.580 ;
        RECT 4.225 51.395 4.515 51.440 ;
        RECT 7.905 51.395 8.195 51.440 ;
        RECT 89.770 7.720 90.090 7.780 ;
        RECT 52.140 7.580 90.090 7.720 ;
        RECT 34.585 7.380 34.875 7.425 ;
        RECT 52.140 7.380 52.280 7.580 ;
        RECT 89.770 7.520 90.090 7.580 ;
        RECT 34.585 7.240 52.280 7.380 ;
        RECT 34.585 7.195 34.875 7.240 ;
        RECT 7.905 6.020 8.195 6.065 ;
        RECT 25.845 6.020 26.135 6.065 ;
        RECT 7.905 5.880 26.135 6.020 ;
        RECT 7.905 5.835 8.195 5.880 ;
        RECT 25.845 5.835 26.135 5.880 ;
        RECT 26.765 6.020 27.055 6.065 ;
        RECT 34.585 6.020 34.875 6.065 ;
        RECT 26.765 5.880 34.875 6.020 ;
        RECT 26.765 5.835 27.055 5.880 ;
        RECT 34.585 5.835 34.875 5.880 ;
        RECT 462.845 3.980 463.135 4.025 ;
        RECT 418.760 3.840 463.135 3.980 ;
        RECT 89.770 3.640 90.090 3.700 ;
        RECT 418.760 3.640 418.900 3.840 ;
        RECT 462.845 3.795 463.135 3.840 ;
        RECT 89.770 3.500 418.900 3.640 ;
        RECT 89.770 3.440 90.090 3.500 ;
        RECT 464.225 1.940 464.515 1.985 ;
        RECT 471.110 1.940 471.430 2.000 ;
        RECT 464.225 1.800 471.430 1.940 ;
        RECT 464.225 1.755 464.515 1.800 ;
        RECT 471.110 1.740 471.430 1.800 ;
      LAYER via ;
        RECT 0.560 1083.960 0.820 1084.220 ;
        RECT 7.000 990.120 7.260 990.380 ;
        RECT 6.080 859.560 6.340 859.820 ;
        RECT 7.000 859.560 7.260 859.820 ;
        RECT 6.540 693.300 6.800 693.560 ;
        RECT 89.800 7.520 90.060 7.780 ;
        RECT 89.800 3.440 90.060 3.700 ;
        RECT 471.140 1.740 471.400 2.000 ;
      LAYER met2 ;
        RECT 0.550 1760.675 0.830 1761.045 ;
        RECT 0.620 1084.250 0.760 1760.675 ;
        RECT 0.560 1083.930 0.820 1084.250 ;
        RECT 7.000 990.090 7.260 990.410 ;
        RECT 7.060 859.850 7.200 990.090 ;
        RECT 6.080 859.530 6.340 859.850 ;
        RECT 7.000 859.530 7.260 859.850 ;
        RECT 6.140 734.810 6.280 859.530 ;
        RECT 6.140 734.670 6.740 734.810 ;
        RECT 6.600 693.590 6.740 734.670 ;
        RECT 6.540 693.270 6.800 693.590 ;
        RECT 89.800 7.490 90.060 7.810 ;
        RECT 89.860 3.730 90.000 7.490 ;
        RECT 89.800 3.410 90.060 3.730 ;
        RECT 471.200 2.820 472.720 2.960 ;
        RECT 471.200 2.030 471.340 2.820 ;
        RECT 472.580 2.400 472.720 2.820 ;
        RECT 471.140 1.710 471.400 2.030 ;
        RECT 472.370 -4.800 472.930 2.400 ;
      LAYER via2 ;
        RECT 0.550 1760.720 0.830 1761.000 ;
      LAYER met3 ;
        RECT 5.000 1761.480 9.000 1762.080 ;
        RECT 0.525 1761.010 0.855 1761.025 ;
        RECT 5.830 1761.010 6.130 1761.480 ;
        RECT 0.525 1760.710 6.130 1761.010 ;
        RECT 0.525 1760.695 0.855 1760.710 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 756.770 1.260 757.090 1.320 ;
        RECT 758.610 1.260 758.930 1.320 ;
        RECT 756.770 1.120 758.930 1.260 ;
        RECT 756.770 1.060 757.090 1.120 ;
        RECT 758.610 1.060 758.930 1.120 ;
      LAYER via ;
        RECT 756.800 1.060 757.060 1.320 ;
        RECT 758.640 1.060 758.900 1.320 ;
      LAYER met2 ;
        RECT 2308.310 5.000 2308.590 9.000 ;
        RECT 490.520 2.820 491.580 2.960 ;
        RECT 490.520 2.400 490.660 2.820 ;
        RECT 490.310 -4.800 490.870 2.400 ;
        RECT 491.440 1.205 491.580 2.820 ;
        RECT 491.370 0.835 491.650 1.205 ;
        RECT 582.910 1.090 583.190 1.205 ;
        RECT 584.290 1.090 584.570 1.205 ;
        RECT 582.910 0.950 584.570 1.090 ;
        RECT 582.910 0.835 583.190 0.950 ;
        RECT 584.290 0.835 584.570 0.950 ;
        RECT 754.950 1.090 755.230 1.205 ;
        RECT 756.800 1.090 757.060 1.350 ;
        RECT 754.950 1.030 757.060 1.090 ;
        RECT 758.640 1.090 758.900 1.350 ;
        RECT 2308.440 1.205 2308.580 5.000 ;
        RECT 759.090 1.090 759.370 1.205 ;
        RECT 758.640 1.030 759.370 1.090 ;
        RECT 754.950 0.950 757.000 1.030 ;
        RECT 758.700 0.950 759.370 1.030 ;
        RECT 754.950 0.835 755.230 0.950 ;
        RECT 759.090 0.835 759.370 0.950 ;
        RECT 991.850 1.090 992.130 1.205 ;
        RECT 992.770 1.090 993.050 1.205 ;
        RECT 991.850 0.950 993.050 1.090 ;
        RECT 991.850 0.835 992.130 0.950 ;
        RECT 992.770 0.835 993.050 0.950 ;
        RECT 1242.090 1.090 1242.370 1.205 ;
        RECT 1243.470 1.090 1243.750 1.205 ;
        RECT 1242.090 0.950 1243.750 1.090 ;
        RECT 1242.090 0.835 1242.370 0.950 ;
        RECT 1243.470 0.835 1243.750 0.950 ;
        RECT 1325.350 0.835 1325.630 1.205 ;
        RECT 1328.110 0.835 1328.390 1.205 ;
        RECT 2308.370 0.835 2308.650 1.205 ;
        RECT 1325.420 0.410 1325.560 0.835 ;
        RECT 1328.180 0.410 1328.320 0.835 ;
        RECT 1325.420 0.270 1328.320 0.410 ;
      LAYER via2 ;
        RECT 491.370 0.880 491.650 1.160 ;
        RECT 582.910 0.880 583.190 1.160 ;
        RECT 584.290 0.880 584.570 1.160 ;
        RECT 754.950 0.880 755.230 1.160 ;
        RECT 759.090 0.880 759.370 1.160 ;
        RECT 991.850 0.880 992.130 1.160 ;
        RECT 992.770 0.880 993.050 1.160 ;
        RECT 1242.090 0.880 1242.370 1.160 ;
        RECT 1243.470 0.880 1243.750 1.160 ;
        RECT 1325.350 0.880 1325.630 1.160 ;
        RECT 1328.110 0.880 1328.390 1.160 ;
        RECT 2308.370 0.880 2308.650 1.160 ;
      LAYER met3 ;
        RECT 491.345 1.170 491.675 1.185 ;
        RECT 582.885 1.170 583.215 1.185 ;
        RECT 491.345 0.870 544.330 1.170 ;
        RECT 491.345 0.855 491.675 0.870 ;
        RECT 544.030 0.490 544.330 0.870 ;
        RECT 559.440 0.870 583.215 1.170 ;
        RECT 559.440 0.490 559.740 0.870 ;
        RECT 582.885 0.855 583.215 0.870 ;
        RECT 584.265 1.170 584.595 1.185 ;
        RECT 754.925 1.170 755.255 1.185 ;
        RECT 584.265 0.870 755.255 1.170 ;
        RECT 584.265 0.855 584.595 0.870 ;
        RECT 754.925 0.855 755.255 0.870 ;
        RECT 759.065 1.170 759.395 1.185 ;
        RECT 991.825 1.170 992.155 1.185 ;
        RECT 759.065 0.870 992.155 1.170 ;
        RECT 759.065 0.855 759.395 0.870 ;
        RECT 991.825 0.855 992.155 0.870 ;
        RECT 992.745 1.170 993.075 1.185 ;
        RECT 1242.065 1.170 1242.395 1.185 ;
        RECT 992.745 0.870 1242.395 1.170 ;
        RECT 992.745 0.855 993.075 0.870 ;
        RECT 1242.065 0.855 1242.395 0.870 ;
        RECT 1243.445 1.170 1243.775 1.185 ;
        RECT 1325.325 1.170 1325.655 1.185 ;
        RECT 1243.445 0.870 1325.655 1.170 ;
        RECT 1243.445 0.855 1243.775 0.870 ;
        RECT 1325.325 0.855 1325.655 0.870 ;
        RECT 1328.085 1.170 1328.415 1.185 ;
        RECT 2308.345 1.170 2308.675 1.185 ;
        RECT 1328.085 0.870 2308.675 1.170 ;
        RECT 1328.085 0.855 1328.415 0.870 ;
        RECT 2308.345 0.855 2308.675 0.870 ;
        RECT 544.030 0.190 559.740 0.490 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 7.505 1191.445 7.675 1251.455 ;
        RECT 1.525 997.305 1.695 1105.255 ;
        RECT 1.525 854.845 1.695 914.175 ;
        RECT 8.885 195.925 9.055 237.575 ;
        RECT 6.585 105.995 6.755 178.415 ;
        RECT 6.585 105.825 7.215 105.995 ;
        RECT 7.045 63.835 7.215 105.825 ;
        RECT 7.045 63.665 7.675 63.835 ;
        RECT 7.505 1.785 7.675 63.665 ;
        RECT 504.305 3.825 504.475 5.355 ;
        RECT 27.745 2.125 29.295 2.295 ;
        RECT 27.745 1.955 27.915 2.125 ;
        RECT 26.825 1.785 27.915 1.955 ;
        RECT 29.125 1.785 29.295 2.125 ;
      LAYER mcon ;
        RECT 7.505 1251.285 7.675 1251.455 ;
        RECT 1.525 1105.085 1.695 1105.255 ;
        RECT 1.525 914.005 1.695 914.175 ;
        RECT 8.885 237.405 9.055 237.575 ;
        RECT 6.585 178.245 6.755 178.415 ;
        RECT 504.305 5.185 504.475 5.355 ;
      LAYER met1 ;
        RECT 2.830 1286.460 3.150 1286.520 ;
        RECT 9.730 1286.460 10.050 1286.520 ;
        RECT 2.830 1286.320 10.050 1286.460 ;
        RECT 2.830 1286.260 3.150 1286.320 ;
        RECT 9.730 1286.260 10.050 1286.320 ;
        RECT 7.445 1251.440 7.735 1251.485 ;
        RECT 9.730 1251.440 10.050 1251.500 ;
        RECT 7.445 1251.300 10.050 1251.440 ;
        RECT 7.445 1251.255 7.735 1251.300 ;
        RECT 9.730 1251.240 10.050 1251.300 ;
        RECT 7.445 1191.600 7.735 1191.645 ;
        RECT 9.730 1191.600 10.050 1191.660 ;
        RECT 7.445 1191.460 10.050 1191.600 ;
        RECT 7.445 1191.415 7.735 1191.460 ;
        RECT 9.730 1191.400 10.050 1191.460 ;
        RECT 1.465 1105.240 1.755 1105.285 ;
        RECT 9.730 1105.240 10.050 1105.300 ;
        RECT 1.465 1105.100 10.050 1105.240 ;
        RECT 1.465 1105.055 1.755 1105.100 ;
        RECT 9.730 1105.040 10.050 1105.100 ;
        RECT 1.450 997.460 1.770 997.520 ;
        RECT 1.255 997.320 1.770 997.460 ;
        RECT 1.450 997.260 1.770 997.320 ;
        RECT 1.450 914.160 1.770 914.220 ;
        RECT 1.255 914.020 1.770 914.160 ;
        RECT 1.450 913.960 1.770 914.020 ;
        RECT 0.530 855.000 0.850 855.060 ;
        RECT 1.465 855.000 1.755 855.045 ;
        RECT 0.530 854.860 1.755 855.000 ;
        RECT 0.530 854.800 0.850 854.860 ;
        RECT 1.465 854.815 1.755 854.860 ;
        RECT 0.530 760.140 0.850 760.200 ;
        RECT 1.910 760.140 2.230 760.200 ;
        RECT 0.530 760.000 2.230 760.140 ;
        RECT 0.530 759.940 0.850 760.000 ;
        RECT 1.910 759.940 2.230 760.000 ;
        RECT 0.530 735.660 0.850 735.720 ;
        RECT 1.910 735.660 2.230 735.720 ;
        RECT 0.530 735.520 2.230 735.660 ;
        RECT 0.530 735.460 0.850 735.520 ;
        RECT 1.910 735.460 2.230 735.520 ;
        RECT 0.530 237.560 0.850 237.620 ;
        RECT 8.825 237.560 9.115 237.605 ;
        RECT 0.530 237.420 9.115 237.560 ;
        RECT 0.530 237.360 0.850 237.420 ;
        RECT 8.825 237.375 9.115 237.420 ;
        RECT 8.825 196.080 9.115 196.125 ;
        RECT 9.730 196.080 10.050 196.140 ;
        RECT 8.825 195.940 10.050 196.080 ;
        RECT 8.825 195.895 9.115 195.940 ;
        RECT 9.730 195.880 10.050 195.940 ;
        RECT 6.525 178.400 6.815 178.445 ;
        RECT 9.730 178.400 10.050 178.460 ;
        RECT 6.525 178.260 10.050 178.400 ;
        RECT 6.525 178.215 6.815 178.260 ;
        RECT 9.730 178.200 10.050 178.260 ;
        RECT 464.210 5.340 464.530 5.400 ;
        RECT 504.245 5.340 504.535 5.385 ;
        RECT 464.210 5.200 504.535 5.340 ;
        RECT 464.210 5.140 464.530 5.200 ;
        RECT 504.245 5.155 504.535 5.200 ;
        RECT 463.290 3.980 463.610 4.040 ;
        RECT 464.210 3.980 464.530 4.040 ;
        RECT 463.290 3.840 464.530 3.980 ;
        RECT 463.290 3.780 463.610 3.840 ;
        RECT 464.210 3.780 464.530 3.840 ;
        RECT 504.245 3.980 504.535 4.025 ;
        RECT 506.990 3.980 507.310 4.040 ;
        RECT 504.245 3.840 507.310 3.980 ;
        RECT 504.245 3.795 504.535 3.840 ;
        RECT 506.990 3.780 507.310 3.840 ;
        RECT 462.830 2.280 463.150 2.340 ;
        RECT 51.680 2.140 370.140 2.280 ;
        RECT 7.445 1.940 7.735 1.985 ;
        RECT 26.765 1.940 27.055 1.985 ;
        RECT 7.445 1.800 27.055 1.940 ;
        RECT 7.445 1.755 7.735 1.800 ;
        RECT 26.765 1.755 27.055 1.800 ;
        RECT 29.065 1.940 29.355 1.985 ;
        RECT 51.680 1.940 51.820 2.140 ;
        RECT 29.065 1.800 51.820 1.940 ;
        RECT 370.000 1.940 370.140 2.140 ;
        RECT 371.380 2.140 463.150 2.280 ;
        RECT 371.380 1.940 371.520 2.140 ;
        RECT 462.830 2.080 463.150 2.140 ;
        RECT 370.000 1.800 371.520 1.940 ;
        RECT 29.065 1.755 29.355 1.800 ;
      LAYER via ;
        RECT 2.860 1286.260 3.120 1286.520 ;
        RECT 9.760 1286.260 10.020 1286.520 ;
        RECT 9.760 1251.240 10.020 1251.500 ;
        RECT 9.760 1191.400 10.020 1191.660 ;
        RECT 9.760 1105.040 10.020 1105.300 ;
        RECT 1.480 997.260 1.740 997.520 ;
        RECT 1.480 913.960 1.740 914.220 ;
        RECT 0.560 854.800 0.820 855.060 ;
        RECT 0.560 759.940 0.820 760.200 ;
        RECT 1.940 759.940 2.200 760.200 ;
        RECT 0.560 735.460 0.820 735.720 ;
        RECT 1.940 735.460 2.200 735.720 ;
        RECT 0.560 237.360 0.820 237.620 ;
        RECT 9.760 195.880 10.020 196.140 ;
        RECT 9.760 178.200 10.020 178.460 ;
        RECT 464.240 5.140 464.500 5.400 ;
        RECT 463.320 3.780 463.580 4.040 ;
        RECT 464.240 3.780 464.500 4.040 ;
        RECT 507.020 3.780 507.280 4.040 ;
        RECT 462.860 2.080 463.120 2.340 ;
      LAYER met2 ;
        RECT 2.850 1871.515 3.130 1871.885 ;
        RECT 2.920 1286.550 3.060 1871.515 ;
        RECT 2.860 1286.230 3.120 1286.550 ;
        RECT 9.760 1286.290 10.020 1286.550 ;
        RECT 9.760 1286.230 10.420 1286.290 ;
        RECT 9.820 1286.150 10.420 1286.230 ;
        RECT 10.280 1284.930 10.420 1286.150 ;
        RECT 10.280 1284.790 11.340 1284.930 ;
        RECT 11.200 1259.770 11.340 1284.790 ;
        RECT 10.280 1259.630 11.340 1259.770 ;
        RECT 10.280 1251.610 10.420 1259.630 ;
        RECT 9.820 1251.530 10.420 1251.610 ;
        RECT 9.760 1251.470 10.420 1251.530 ;
        RECT 9.760 1251.210 10.020 1251.470 ;
        RECT 9.760 1191.600 10.020 1191.690 ;
        RECT 9.760 1191.460 11.340 1191.600 ;
        RECT 9.760 1191.370 10.020 1191.460 ;
        RECT 11.200 1130.570 11.340 1191.460 ;
        RECT 10.740 1130.430 11.340 1130.570 ;
        RECT 10.740 1105.410 10.880 1130.430 ;
        RECT 9.820 1105.330 10.880 1105.410 ;
        RECT 9.760 1105.270 10.880 1105.330 ;
        RECT 9.760 1105.010 10.020 1105.270 ;
        RECT 1.480 997.230 1.740 997.550 ;
        RECT 1.540 914.250 1.680 997.230 ;
        RECT 1.480 913.930 1.740 914.250 ;
        RECT 0.560 854.770 0.820 855.090 ;
        RECT 0.620 760.230 0.760 854.770 ;
        RECT 0.560 759.910 0.820 760.230 ;
        RECT 1.940 759.910 2.200 760.230 ;
        RECT 2.000 735.750 2.140 759.910 ;
        RECT 0.560 735.430 0.820 735.750 ;
        RECT 1.940 735.430 2.200 735.750 ;
        RECT 0.620 237.650 0.760 735.430 ;
        RECT 0.560 237.330 0.820 237.650 ;
        RECT 9.760 195.850 10.020 196.170 ;
        RECT 9.820 195.570 9.960 195.850 ;
        RECT 9.820 195.430 12.260 195.570 ;
        RECT 12.120 178.570 12.260 195.430 ;
        RECT 9.820 178.490 12.260 178.570 ;
        RECT 9.760 178.430 12.260 178.490 ;
        RECT 9.760 178.170 10.020 178.430 ;
        RECT 464.240 5.110 464.500 5.430 ;
        RECT 464.300 4.070 464.440 5.110 ;
        RECT 463.320 3.750 463.580 4.070 ;
        RECT 464.240 3.750 464.500 4.070 ;
        RECT 507.020 3.750 507.280 4.070 ;
        RECT 462.860 2.280 463.120 2.370 ;
        RECT 463.380 2.280 463.520 3.750 ;
        RECT 507.080 2.960 507.220 3.750 ;
        RECT 507.080 2.820 508.140 2.960 ;
        RECT 508.000 2.400 508.140 2.820 ;
        RECT 462.860 2.140 463.520 2.280 ;
        RECT 462.860 2.050 463.120 2.140 ;
        RECT 507.790 -4.800 508.350 2.400 ;
      LAYER via2 ;
        RECT 2.850 1871.560 3.130 1871.840 ;
      LAYER met3 ;
        RECT 5.000 1874.360 9.000 1874.960 ;
        RECT 2.825 1871.850 3.155 1871.865 ;
        RECT 5.830 1871.850 6.130 1874.360 ;
        RECT 2.825 1871.550 6.130 1871.850 ;
        RECT 2.825 1871.535 3.155 1871.550 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 4.745 979.625 4.915 988.295 ;
        RECT 4.285 796.365 4.455 834.615 ;
        RECT 9.345 715.445 9.515 729.555 ;
        RECT 4.745 673.115 4.915 693.855 ;
        RECT 7.045 693.685 7.215 706.435 ;
        RECT 4.745 672.945 5.375 673.115 ;
        RECT 5.205 633.165 5.375 672.945 ;
        RECT 9.345 481.185 9.515 589.135 ;
        RECT 3.825 18.445 3.995 52.275 ;
        RECT 7.965 52.105 8.135 91.375 ;
        RECT 505.685 4.505 506.775 4.675 ;
        RECT 505.685 4.165 505.855 4.505 ;
      LAYER mcon ;
        RECT 4.745 988.125 4.915 988.295 ;
        RECT 4.285 834.445 4.455 834.615 ;
        RECT 9.345 729.385 9.515 729.555 ;
        RECT 7.045 706.265 7.215 706.435 ;
        RECT 4.745 693.685 4.915 693.855 ;
        RECT 9.345 588.965 9.515 589.135 ;
        RECT 7.965 91.205 8.135 91.375 ;
        RECT 3.825 52.105 3.995 52.275 ;
        RECT 506.605 4.505 506.775 4.675 ;
      LAYER met1 ;
        RECT 4.670 988.280 4.990 988.340 ;
        RECT 4.475 988.140 4.990 988.280 ;
        RECT 4.670 988.080 4.990 988.140 ;
        RECT 4.685 979.780 4.975 979.825 ;
        RECT 9.730 979.780 10.050 979.840 ;
        RECT 4.685 979.640 10.050 979.780 ;
        RECT 4.685 979.595 4.975 979.640 ;
        RECT 9.730 979.580 10.050 979.640 ;
        RECT 4.225 834.600 4.515 834.645 ;
        RECT 9.730 834.600 10.050 834.660 ;
        RECT 4.225 834.460 10.050 834.600 ;
        RECT 4.225 834.415 4.515 834.460 ;
        RECT 9.730 834.400 10.050 834.460 ;
        RECT 4.225 796.520 4.515 796.565 ;
        RECT 9.730 796.520 10.050 796.580 ;
        RECT 4.225 796.380 10.050 796.520 ;
        RECT 4.225 796.335 4.515 796.380 ;
        RECT 9.730 796.320 10.050 796.380 ;
        RECT 9.270 729.540 9.590 729.600 ;
        RECT 9.075 729.400 9.590 729.540 ;
        RECT 9.270 729.340 9.590 729.400 ;
        RECT 9.270 715.600 9.590 715.660 ;
        RECT 9.075 715.460 9.590 715.600 ;
        RECT 9.270 715.400 9.590 715.460 ;
        RECT 6.985 706.420 7.275 706.465 ;
        RECT 9.270 706.420 9.590 706.480 ;
        RECT 6.985 706.280 9.590 706.420 ;
        RECT 6.985 706.235 7.275 706.280 ;
        RECT 9.270 706.220 9.590 706.280 ;
        RECT 4.685 693.840 4.975 693.885 ;
        RECT 6.985 693.840 7.275 693.885 ;
        RECT 4.685 693.700 7.275 693.840 ;
        RECT 4.685 693.655 4.975 693.700 ;
        RECT 6.985 693.655 7.275 693.700 ;
        RECT 5.145 633.320 5.435 633.365 ;
        RECT 8.810 633.320 9.130 633.380 ;
        RECT 5.145 633.180 9.130 633.320 ;
        RECT 5.145 633.135 5.435 633.180 ;
        RECT 8.810 633.120 9.130 633.180 ;
        RECT 9.285 589.120 9.575 589.165 ;
        RECT 9.730 589.120 10.050 589.180 ;
        RECT 9.285 588.980 10.050 589.120 ;
        RECT 9.285 588.935 9.575 588.980 ;
        RECT 9.730 588.920 10.050 588.980 ;
        RECT 2.370 481.340 2.690 481.400 ;
        RECT 9.285 481.340 9.575 481.385 ;
        RECT 2.370 481.200 9.575 481.340 ;
        RECT 2.370 481.140 2.690 481.200 ;
        RECT 9.285 481.155 9.575 481.200 ;
        RECT 2.370 91.360 2.690 91.420 ;
        RECT 7.905 91.360 8.195 91.405 ;
        RECT 2.370 91.220 8.195 91.360 ;
        RECT 2.370 91.160 2.690 91.220 ;
        RECT 7.905 91.175 8.195 91.220 ;
        RECT 3.765 52.260 4.055 52.305 ;
        RECT 7.905 52.260 8.195 52.305 ;
        RECT 3.765 52.120 8.195 52.260 ;
        RECT 3.765 52.075 4.055 52.120 ;
        RECT 7.905 52.075 8.195 52.120 ;
        RECT 3.750 18.600 4.070 18.660 ;
        RECT 3.555 18.460 4.070 18.600 ;
        RECT 3.750 18.400 4.070 18.460 ;
        RECT 506.545 4.660 506.835 4.705 ;
        RECT 506.545 4.520 508.140 4.660 ;
        RECT 506.545 4.475 506.835 4.520 ;
        RECT 485.370 4.320 485.690 4.380 ;
        RECT 505.625 4.320 505.915 4.365 ;
        RECT 485.370 4.180 505.915 4.320 ;
        RECT 508.000 4.320 508.140 4.520 ;
        RECT 517.110 4.320 517.430 4.380 ;
        RECT 508.000 4.180 517.430 4.320 ;
        RECT 485.370 4.120 485.690 4.180 ;
        RECT 505.625 4.135 505.915 4.180 ;
        RECT 517.110 4.120 517.430 4.180 ;
      LAYER via ;
        RECT 4.700 988.080 4.960 988.340 ;
        RECT 9.760 979.580 10.020 979.840 ;
        RECT 9.760 834.400 10.020 834.660 ;
        RECT 9.760 796.320 10.020 796.580 ;
        RECT 9.300 729.340 9.560 729.600 ;
        RECT 9.300 715.400 9.560 715.660 ;
        RECT 9.300 706.220 9.560 706.480 ;
        RECT 8.840 633.120 9.100 633.380 ;
        RECT 9.760 588.920 10.020 589.180 ;
        RECT 2.400 481.140 2.660 481.400 ;
        RECT 2.400 91.160 2.660 91.420 ;
        RECT 3.780 18.400 4.040 18.660 ;
        RECT 485.400 4.120 485.660 4.380 ;
        RECT 517.140 4.120 517.400 4.380 ;
      LAYER met2 ;
        RECT 4.690 1986.435 4.970 1986.805 ;
        RECT 4.760 988.370 4.900 1986.435 ;
        RECT 4.700 988.050 4.960 988.370 ;
        RECT 9.760 979.610 10.020 979.870 ;
        RECT 9.760 979.550 13.180 979.610 ;
        RECT 9.820 979.470 13.180 979.550 ;
        RECT 13.040 944.760 13.180 979.470 ;
        RECT 12.580 944.620 13.180 944.760 ;
        RECT 12.580 931.330 12.720 944.620 ;
        RECT 11.200 931.190 12.720 931.330 ;
        RECT 11.200 885.090 11.340 931.190 ;
        RECT 11.200 884.950 13.180 885.090 ;
        RECT 13.040 834.770 13.180 884.950 ;
        RECT 9.820 834.690 13.180 834.770 ;
        RECT 9.760 834.630 13.180 834.690 ;
        RECT 9.760 834.370 10.020 834.630 ;
        RECT 9.760 796.520 10.020 796.610 ;
        RECT 9.760 796.380 10.420 796.520 ;
        RECT 9.760 796.290 10.020 796.380 ;
        RECT 10.280 755.890 10.420 796.380 ;
        RECT 9.360 755.750 10.420 755.890 ;
        RECT 9.360 729.630 9.500 755.750 ;
        RECT 9.300 729.310 9.560 729.630 ;
        RECT 9.300 715.370 9.560 715.690 ;
        RECT 9.360 706.510 9.500 715.370 ;
        RECT 9.300 706.190 9.560 706.510 ;
        RECT 8.840 633.090 9.100 633.410 ;
        RECT 8.900 630.090 9.040 633.090 ;
        RECT 8.900 629.950 10.420 630.090 ;
        RECT 10.280 589.290 10.420 629.950 ;
        RECT 9.820 589.210 10.420 589.290 ;
        RECT 9.760 589.150 10.420 589.210 ;
        RECT 9.760 588.890 10.020 589.150 ;
        RECT 2.400 481.110 2.660 481.430 ;
        RECT 2.460 91.450 2.600 481.110 ;
        RECT 2.400 91.130 2.660 91.450 ;
        RECT 3.780 18.370 4.040 18.690 ;
        RECT 3.840 6.645 3.980 18.370 ;
        RECT 315.260 6.900 319.080 7.040 ;
        RECT 315.260 6.645 315.400 6.900 ;
        RECT 318.940 6.645 319.080 6.900 ;
        RECT 3.770 6.275 4.050 6.645 ;
        RECT 301.390 6.275 301.670 6.645 ;
        RECT 304.150 6.275 304.430 6.645 ;
        RECT 315.190 6.275 315.470 6.645 ;
        RECT 318.870 6.275 319.150 6.645 ;
        RECT 301.460 5.340 301.600 6.275 ;
        RECT 304.220 5.340 304.360 6.275 ;
        RECT 301.460 5.200 304.360 5.340 ;
        RECT 485.390 4.915 485.670 5.285 ;
        RECT 485.460 4.410 485.600 4.915 ;
        RECT 485.400 4.090 485.660 4.410 ;
        RECT 517.140 4.090 517.400 4.410 ;
        RECT 519.500 4.180 526.080 4.320 ;
        RECT 517.200 3.130 517.340 4.090 ;
        RECT 519.500 3.130 519.640 4.180 ;
        RECT 517.200 2.990 519.640 3.130 ;
        RECT 525.940 2.400 526.080 4.180 ;
        RECT 525.730 -4.800 526.290 2.400 ;
      LAYER via2 ;
        RECT 4.690 1986.480 4.970 1986.760 ;
        RECT 3.770 6.320 4.050 6.600 ;
        RECT 301.390 6.320 301.670 6.600 ;
        RECT 304.150 6.320 304.430 6.600 ;
        RECT 315.190 6.320 315.470 6.600 ;
        RECT 318.870 6.320 319.150 6.600 ;
        RECT 485.390 4.960 485.670 5.240 ;
      LAYER met3 ;
        RECT 5.000 1987.920 9.000 1988.520 ;
        RECT 4.665 1986.770 4.995 1986.785 ;
        RECT 5.830 1986.770 6.130 1987.920 ;
        RECT 4.665 1986.470 6.130 1986.770 ;
        RECT 4.665 1986.455 4.995 1986.470 ;
        RECT 3.745 6.610 4.075 6.625 ;
        RECT 301.365 6.610 301.695 6.625 ;
        RECT 3.745 6.310 301.695 6.610 ;
        RECT 3.745 6.295 4.075 6.310 ;
        RECT 301.365 6.295 301.695 6.310 ;
        RECT 304.125 6.610 304.455 6.625 ;
        RECT 315.165 6.610 315.495 6.625 ;
        RECT 304.125 6.310 315.495 6.610 ;
        RECT 304.125 6.295 304.455 6.310 ;
        RECT 315.165 6.295 315.495 6.310 ;
        RECT 318.845 6.610 319.175 6.625 ;
        RECT 415.190 6.610 415.570 6.620 ;
        RECT 318.845 6.310 415.570 6.610 ;
        RECT 318.845 6.295 319.175 6.310 ;
        RECT 415.190 6.300 415.570 6.310 ;
        RECT 417.030 5.250 417.410 5.260 ;
        RECT 485.365 5.250 485.695 5.265 ;
        RECT 417.030 4.950 485.695 5.250 ;
        RECT 417.030 4.940 417.410 4.950 ;
        RECT 485.365 4.935 485.695 4.950 ;
      LAYER via3 ;
        RECT 415.220 6.300 415.540 6.620 ;
        RECT 417.060 4.940 417.380 5.260 ;
      LAYER met4 ;
        RECT 415.215 6.295 415.545 6.625 ;
        RECT 415.230 5.930 415.530 6.295 ;
        RECT 415.230 5.630 417.370 5.930 ;
        RECT 417.070 5.265 417.370 5.630 ;
        RECT 417.055 4.935 417.385 5.265 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 8.425 1838.805 8.595 1852.575 ;
        RECT 8.425 624.325 8.595 672.775 ;
        RECT 8.425 323.765 8.595 329.375 ;
        RECT 17.625 9.265 30.675 9.435 ;
        RECT 17.625 7.395 17.795 9.265 ;
        RECT 17.165 7.225 17.795 7.395 ;
        RECT 30.505 2.465 30.675 9.265 ;
        RECT 481.765 4.505 486.995 4.675 ;
        RECT 481.765 4.165 481.935 4.505 ;
        RECT 505.225 3.995 505.395 4.675 ;
        RECT 506.145 3.995 506.315 4.335 ;
        RECT 505.225 3.825 506.315 3.995 ;
      LAYER mcon ;
        RECT 8.425 1852.405 8.595 1852.575 ;
        RECT 8.425 672.605 8.595 672.775 ;
        RECT 8.425 329.205 8.595 329.375 ;
        RECT 486.825 4.505 486.995 4.675 ;
        RECT 505.225 4.505 505.395 4.675 ;
        RECT 506.145 4.165 506.315 4.335 ;
      LAYER met1 ;
        RECT 6.970 2073.220 7.290 2073.280 ;
        RECT 8.350 2073.220 8.670 2073.280 ;
        RECT 6.970 2073.080 8.670 2073.220 ;
        RECT 6.970 2073.020 7.290 2073.080 ;
        RECT 8.350 2073.020 8.670 2073.080 ;
        RECT 8.350 1852.560 8.670 1852.620 ;
        RECT 8.155 1852.420 8.670 1852.560 ;
        RECT 8.350 1852.360 8.670 1852.420 ;
        RECT 8.350 1838.960 8.670 1839.020 ;
        RECT 8.155 1838.820 8.670 1838.960 ;
        RECT 8.350 1838.760 8.670 1838.820 ;
        RECT 8.350 672.760 8.670 672.820 ;
        RECT 8.155 672.620 8.670 672.760 ;
        RECT 8.350 672.560 8.670 672.620 ;
        RECT 8.350 624.480 8.670 624.540 ;
        RECT 8.155 624.340 8.670 624.480 ;
        RECT 8.350 624.280 8.670 624.340 ;
        RECT 8.350 329.360 8.670 329.420 ;
        RECT 8.155 329.220 8.670 329.360 ;
        RECT 8.350 329.160 8.670 329.220 ;
        RECT 8.350 323.920 8.670 323.980 ;
        RECT 8.155 323.780 8.670 323.920 ;
        RECT 8.350 323.720 8.670 323.780 ;
        RECT 7.890 7.380 8.210 7.440 ;
        RECT 17.105 7.380 17.395 7.425 ;
        RECT 7.890 7.240 17.395 7.380 ;
        RECT 7.890 7.180 8.210 7.240 ;
        RECT 17.105 7.195 17.395 7.240 ;
        RECT 486.765 4.660 487.055 4.705 ;
        RECT 505.165 4.660 505.455 4.705 ;
        RECT 486.765 4.520 505.455 4.660 ;
        RECT 486.765 4.475 487.055 4.520 ;
        RECT 505.165 4.475 505.455 4.520 ;
        RECT 470.190 4.320 470.510 4.380 ;
        RECT 481.705 4.320 481.995 4.365 ;
        RECT 470.190 4.180 481.995 4.320 ;
        RECT 470.190 4.120 470.510 4.180 ;
        RECT 481.705 4.135 481.995 4.180 ;
        RECT 506.085 4.320 506.375 4.365 ;
        RECT 506.085 4.180 507.680 4.320 ;
        RECT 506.085 4.135 506.375 4.180 ;
        RECT 507.540 3.980 507.680 4.180 ;
        RECT 509.750 3.980 510.070 4.040 ;
        RECT 507.540 3.840 510.070 3.980 ;
        RECT 509.750 3.780 510.070 3.840 ;
        RECT 30.445 2.620 30.735 2.665 ;
        RECT 366.230 2.620 366.550 2.680 ;
        RECT 30.445 2.480 366.550 2.620 ;
        RECT 30.445 2.435 30.735 2.480 ;
        RECT 366.230 2.420 366.550 2.480 ;
      LAYER via ;
        RECT 7.000 2073.020 7.260 2073.280 ;
        RECT 8.380 2073.020 8.640 2073.280 ;
        RECT 8.380 1852.360 8.640 1852.620 ;
        RECT 8.380 1838.760 8.640 1839.020 ;
        RECT 8.380 672.560 8.640 672.820 ;
        RECT 8.380 624.280 8.640 624.540 ;
        RECT 8.380 329.160 8.640 329.420 ;
        RECT 8.380 323.720 8.640 323.980 ;
        RECT 7.920 7.180 8.180 7.440 ;
        RECT 470.220 4.120 470.480 4.380 ;
        RECT 509.780 3.780 510.040 4.040 ;
        RECT 366.260 2.420 366.520 2.680 ;
      LAYER met2 ;
        RECT 6.990 2098.635 7.270 2099.005 ;
        RECT 7.060 2073.310 7.200 2098.635 ;
        RECT 7.000 2072.990 7.260 2073.310 ;
        RECT 8.380 2072.990 8.640 2073.310 ;
        RECT 8.440 1852.650 8.580 2072.990 ;
        RECT 8.380 1852.330 8.640 1852.650 ;
        RECT 8.380 1838.730 8.640 1839.050 ;
        RECT 8.440 672.850 8.580 1838.730 ;
        RECT 8.380 672.530 8.640 672.850 ;
        RECT 8.380 624.250 8.640 624.570 ;
        RECT 8.440 329.450 8.580 624.250 ;
        RECT 8.380 329.130 8.640 329.450 ;
        RECT 8.380 323.690 8.640 324.010 ;
        RECT 8.440 25.570 8.580 323.690 ;
        RECT 7.980 25.430 8.580 25.570 ;
        RECT 7.980 7.470 8.120 25.430 ;
        RECT 7.920 7.150 8.180 7.470 ;
        RECT 470.220 4.320 470.480 4.410 ;
        RECT 467.980 4.180 470.480 4.320 ;
        RECT 366.260 2.450 366.520 2.710 ;
        RECT 366.260 2.390 369.680 2.450 ;
        RECT 366.320 2.310 369.680 2.390 ;
        RECT 369.540 0.525 369.680 2.310 ;
        RECT 467.980 1.205 468.120 4.180 ;
        RECT 470.220 4.090 470.480 4.180 ;
        RECT 509.780 3.750 510.040 4.070 ;
        RECT 467.910 0.835 468.190 1.205 ;
        RECT 509.840 0.525 509.980 3.750 ;
        RECT 542.960 2.990 544.020 3.130 ;
        RECT 542.960 0.525 543.100 2.990 ;
        RECT 543.880 2.400 544.020 2.990 ;
        RECT 369.470 0.155 369.750 0.525 ;
        RECT 509.770 0.155 510.050 0.525 ;
        RECT 542.890 0.155 543.170 0.525 ;
        RECT 543.670 -4.800 544.230 2.400 ;
      LAYER via2 ;
        RECT 6.990 2098.680 7.270 2098.960 ;
        RECT 467.910 0.880 468.190 1.160 ;
        RECT 369.470 0.200 369.750 0.480 ;
        RECT 509.770 0.200 510.050 0.480 ;
        RECT 542.890 0.200 543.170 0.480 ;
      LAYER met3 ;
        RECT 5.000 2101.480 9.000 2102.080 ;
        RECT 6.750 2098.985 7.050 2101.480 ;
        RECT 6.750 2098.670 7.295 2098.985 ;
        RECT 6.965 2098.655 7.295 2098.670 ;
        RECT 465.790 1.170 466.170 1.180 ;
        RECT 467.885 1.170 468.215 1.185 ;
        RECT 465.790 0.870 468.215 1.170 ;
        RECT 465.790 0.860 466.170 0.870 ;
        RECT 467.885 0.855 468.215 0.870 ;
        RECT 369.445 0.490 369.775 0.505 ;
        RECT 371.030 0.490 371.410 0.500 ;
        RECT 369.445 0.190 371.410 0.490 ;
        RECT 369.445 0.175 369.775 0.190 ;
        RECT 371.030 0.180 371.410 0.190 ;
        RECT 509.745 0.490 510.075 0.505 ;
        RECT 542.865 0.490 543.195 0.505 ;
        RECT 509.745 0.190 543.195 0.490 ;
        RECT 509.745 0.175 510.075 0.190 ;
        RECT 542.865 0.175 543.195 0.190 ;
      LAYER via3 ;
        RECT 465.820 0.860 466.140 1.180 ;
        RECT 371.060 0.180 371.380 0.500 ;
      LAYER met4 ;
        RECT 372.470 1.110 373.650 2.290 ;
        RECT 462.630 1.850 463.810 2.290 ;
        RECT 462.630 1.550 466.130 1.850 ;
        RECT 462.630 1.110 463.810 1.550 ;
        RECT 465.830 1.185 466.130 1.550 ;
        RECT 371.055 0.490 371.385 0.505 ;
        RECT 372.910 0.490 373.210 1.110 ;
        RECT 465.815 0.855 466.145 1.185 ;
        RECT 371.055 0.190 373.210 0.490 ;
        RECT 371.055 0.175 371.385 0.190 ;
      LAYER met5 ;
        RECT 372.260 0.900 464.020 2.500 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 950.505 9.265 957.115 9.435 ;
        RECT 877.825 8.925 879.375 9.095 ;
        RECT 846.545 8.585 848.555 8.755 ;
        RECT 846.545 8.075 846.715 8.585 ;
        RECT 824.925 7.905 846.715 8.075 ;
        RECT 605.045 6.545 606.135 6.715 ;
        RECT 605.045 6.205 605.215 6.545 ;
        RECT 605.965 4.335 606.135 6.545 ;
        RECT 824.925 6.035 825.095 7.905 ;
        RECT 879.205 7.565 879.375 8.925 ;
        RECT 882.885 6.885 883.055 7.735 ;
        RECT 948.665 7.225 949.755 7.395 ;
        RECT 948.665 6.205 948.835 7.225 ;
        RECT 949.585 6.715 949.755 7.225 ;
        RECT 950.505 6.715 950.675 9.265 ;
        RECT 956.945 8.415 957.115 9.265 ;
        RECT 949.585 6.545 950.675 6.715 ;
        RECT 956.485 8.245 957.115 8.415 ;
        RECT 1259.165 9.265 1264.855 9.435 ;
        RECT 956.485 6.205 956.655 8.245 ;
        RECT 1182.805 7.565 1183.895 7.735 ;
        RECT 1123.465 6.545 1125.015 6.715 ;
        RECT 1123.465 6.375 1123.635 6.545 ;
        RECT 1122.085 6.205 1123.635 6.375 ;
        RECT 1124.845 6.205 1125.015 6.545 ;
        RECT 815.265 5.865 825.095 6.035 ;
        RECT 605.965 4.165 607.055 4.335 ;
        RECT 766.505 4.165 769.895 4.335 ;
        RECT 769.725 3.825 769.895 4.165 ;
        RECT 771.565 3.825 771.735 5.695 ;
        RECT 787.205 4.165 787.375 5.695 ;
        RECT 805.145 3.145 805.315 4.335 ;
        RECT 811.125 3.485 812.215 3.655 ;
        RECT 811.125 3.145 811.295 3.485 ;
        RECT 812.045 1.275 812.215 3.485 ;
        RECT 813.425 1.275 813.595 4.675 ;
        RECT 815.265 4.505 815.435 5.865 ;
        RECT 1161.185 5.695 1161.355 6.375 ;
        RECT 1166.245 5.695 1166.415 7.395 ;
        RECT 1182.805 7.225 1182.975 7.565 ;
        RECT 1183.725 5.865 1183.895 7.565 ;
        RECT 1189.705 7.225 1195.395 7.395 ;
        RECT 1189.705 5.865 1189.875 7.225 ;
        RECT 1257.325 6.035 1257.495 6.375 ;
        RECT 1259.165 6.035 1259.335 9.265 ;
        RECT 1264.685 6.715 1264.855 9.265 ;
        RECT 1469.385 7.735 1469.555 8.755 ;
        RECT 1454.665 7.565 1469.555 7.735 ;
        RECT 1292.285 6.715 1292.455 7.055 ;
        RECT 1264.685 6.545 1292.455 6.715 ;
        RECT 1353.465 6.205 1361.915 6.375 ;
        RECT 1369.105 6.205 1400.095 6.375 ;
        RECT 1454.665 6.205 1454.835 7.565 ;
        RECT 1475.825 7.055 1475.995 8.755 ;
        RECT 1548.505 8.585 1575.355 8.755 ;
        RECT 1475.825 6.885 1476.915 7.055 ;
        RECT 1257.325 5.865 1259.335 6.035 ;
        RECT 1476.745 5.865 1476.915 6.885 ;
        RECT 1547.125 6.375 1547.295 7.055 ;
        RECT 1548.505 6.885 1548.675 8.585 ;
        RECT 1546.205 6.205 1547.295 6.375 ;
        RECT 1575.185 6.375 1575.355 8.585 ;
        RECT 1575.185 6.205 1593.295 6.375 ;
        RECT 1161.185 5.525 1166.415 5.695 ;
        RECT 1687.885 2.465 1688.055 6.375 ;
        RECT 1726.985 5.185 1727.155 6.375 ;
        RECT 1789.545 5.185 1789.715 6.375 ;
        RECT 1820.825 5.525 1821.915 5.695 ;
        RECT 1820.825 5.185 1820.995 5.525 ;
        RECT 1693.865 2.465 1694.035 5.015 ;
        RECT 1821.745 4.505 1821.915 5.525 ;
        RECT 1842.445 4.505 1842.615 7.055 ;
        RECT 1873.265 6.205 1873.435 7.055 ;
        RECT 1932.145 4.335 1932.315 6.375 ;
        RECT 1932.145 4.165 1932.775 4.335 ;
        RECT 2021.385 4.165 2021.555 6.375 ;
        RECT 2161.225 6.205 2161.395 7.735 ;
        RECT 2297.845 6.205 2298.015 7.395 ;
        RECT 2365.925 6.205 2366.095 7.395 ;
        RECT 2366.845 5.185 2367.015 6.375 ;
        RECT 2504.845 6.205 2505.015 7.735 ;
        RECT 2547.625 6.205 2547.795 7.735 ;
        RECT 2780.845 6.205 2781.015 8.075 ;
        RECT 2583.965 4.505 2584.135 5.355 ;
        RECT 812.045 1.105 813.595 1.275 ;
      LAYER mcon ;
        RECT 848.385 8.585 848.555 8.755 ;
        RECT 882.885 7.565 883.055 7.735 ;
        RECT 1166.245 7.225 1166.415 7.395 ;
        RECT 1161.185 6.205 1161.355 6.375 ;
        RECT 771.565 5.525 771.735 5.695 ;
        RECT 606.885 4.165 607.055 4.335 ;
        RECT 787.205 5.525 787.375 5.695 ;
        RECT 1195.225 7.225 1195.395 7.395 ;
        RECT 1257.325 6.205 1257.495 6.375 ;
        RECT 1469.385 8.585 1469.555 8.755 ;
        RECT 1475.825 8.585 1475.995 8.755 ;
        RECT 1292.285 6.885 1292.455 7.055 ;
        RECT 1361.745 6.205 1361.915 6.375 ;
        RECT 1399.925 6.205 1400.095 6.375 ;
        RECT 1547.125 6.885 1547.295 7.055 ;
        RECT 2780.845 7.905 2781.015 8.075 ;
        RECT 2161.225 7.565 2161.395 7.735 ;
        RECT 1842.445 6.885 1842.615 7.055 ;
        RECT 1593.125 6.205 1593.295 6.375 ;
        RECT 1687.885 6.205 1688.055 6.375 ;
        RECT 813.425 4.505 813.595 4.675 ;
        RECT 805.145 4.165 805.315 4.335 ;
        RECT 1726.985 6.205 1727.155 6.375 ;
        RECT 1789.545 6.205 1789.715 6.375 ;
        RECT 1693.865 4.845 1694.035 5.015 ;
        RECT 1873.265 6.885 1873.435 7.055 ;
        RECT 2504.845 7.565 2505.015 7.735 ;
        RECT 1932.145 6.205 1932.315 6.375 ;
        RECT 2021.385 6.205 2021.555 6.375 ;
        RECT 2297.845 7.225 2298.015 7.395 ;
        RECT 2365.925 7.225 2366.095 7.395 ;
        RECT 2366.845 6.205 2367.015 6.375 ;
        RECT 2547.625 7.565 2547.795 7.735 ;
        RECT 2583.965 5.185 2584.135 5.355 ;
        RECT 1932.605 4.165 1932.775 4.335 ;
      LAYER met1 ;
        RECT 877.765 9.080 878.055 9.125 ;
        RECT 850.700 8.940 878.055 9.080 ;
        RECT 848.325 8.740 848.615 8.785 ;
        RECT 850.700 8.740 850.840 8.940 ;
        RECT 877.765 8.895 878.055 8.940 ;
        RECT 848.325 8.600 850.840 8.740 ;
        RECT 1469.325 8.740 1469.615 8.785 ;
        RECT 1475.765 8.740 1476.055 8.785 ;
        RECT 1469.325 8.600 1476.055 8.740 ;
        RECT 848.325 8.555 848.615 8.600 ;
        RECT 1469.325 8.555 1469.615 8.600 ;
        RECT 1475.765 8.555 1476.055 8.600 ;
        RECT 2746.270 8.060 2746.590 8.120 ;
        RECT 2780.785 8.060 2781.075 8.105 ;
        RECT 2746.270 7.920 2781.075 8.060 ;
        RECT 2746.270 7.860 2746.590 7.920 ;
        RECT 2780.785 7.875 2781.075 7.920 ;
        RECT 879.145 7.720 879.435 7.765 ;
        RECT 882.825 7.720 883.115 7.765 ;
        RECT 879.145 7.580 883.115 7.720 ;
        RECT 879.145 7.535 879.435 7.580 ;
        RECT 882.825 7.535 883.115 7.580 ;
        RECT 2125.270 7.720 2125.590 7.780 ;
        RECT 2161.165 7.720 2161.455 7.765 ;
        RECT 2125.270 7.580 2161.455 7.720 ;
        RECT 2125.270 7.520 2125.590 7.580 ;
        RECT 2161.165 7.535 2161.455 7.580 ;
        RECT 2504.785 7.720 2505.075 7.765 ;
        RECT 2547.565 7.720 2547.855 7.765 ;
        RECT 2504.785 7.580 2547.855 7.720 ;
        RECT 2504.785 7.535 2505.075 7.580 ;
        RECT 2547.565 7.535 2547.855 7.580 ;
        RECT 889.250 7.380 889.570 7.440 ;
        RECT 883.820 7.240 889.570 7.380 ;
        RECT 882.825 7.040 883.115 7.085 ;
        RECT 883.820 7.040 883.960 7.240 ;
        RECT 889.250 7.180 889.570 7.240 ;
        RECT 1166.185 7.380 1166.475 7.425 ;
        RECT 1182.745 7.380 1183.035 7.425 ;
        RECT 1166.185 7.240 1183.035 7.380 ;
        RECT 1166.185 7.195 1166.475 7.240 ;
        RECT 1182.745 7.195 1183.035 7.240 ;
        RECT 1195.165 7.380 1195.455 7.425 ;
        RECT 1206.650 7.380 1206.970 7.440 ;
        RECT 1195.165 7.240 1206.970 7.380 ;
        RECT 1195.165 7.195 1195.455 7.240 ;
        RECT 1206.650 7.180 1206.970 7.240 ;
        RECT 1361.670 7.380 1361.990 7.440 ;
        RECT 1369.030 7.380 1369.350 7.440 ;
        RECT 1361.670 7.240 1369.350 7.380 ;
        RECT 1361.670 7.180 1361.990 7.240 ;
        RECT 1369.030 7.180 1369.350 7.240 ;
        RECT 2297.785 7.380 2298.075 7.425 ;
        RECT 2365.865 7.380 2366.155 7.425 ;
        RECT 2297.785 7.240 2366.155 7.380 ;
        RECT 2297.785 7.195 2298.075 7.240 ;
        RECT 2365.865 7.195 2366.155 7.240 ;
        RECT 882.825 6.900 883.960 7.040 ;
        RECT 1292.225 7.040 1292.515 7.085 ;
        RECT 1295.430 7.040 1295.750 7.100 ;
        RECT 1292.225 6.900 1295.750 7.040 ;
        RECT 882.825 6.855 883.115 6.900 ;
        RECT 1292.225 6.855 1292.515 6.900 ;
        RECT 1295.430 6.840 1295.750 6.900 ;
        RECT 1547.065 7.040 1547.355 7.085 ;
        RECT 1548.445 7.040 1548.735 7.085 ;
        RECT 1547.065 6.900 1548.735 7.040 ;
        RECT 1547.065 6.855 1547.355 6.900 ;
        RECT 1548.445 6.855 1548.735 6.900 ;
        RECT 1842.385 7.040 1842.675 7.085 ;
        RECT 1873.205 7.040 1873.495 7.085 ;
        RECT 1842.385 6.900 1873.495 7.040 ;
        RECT 1842.385 6.855 1842.675 6.900 ;
        RECT 1873.205 6.855 1873.495 6.900 ;
        RECT 583.810 6.360 584.130 6.420 ;
        RECT 604.985 6.360 605.275 6.405 ;
        RECT 583.810 6.220 605.275 6.360 ;
        RECT 583.810 6.160 584.130 6.220 ;
        RECT 604.985 6.175 605.275 6.220 ;
        RECT 890.630 6.360 890.950 6.420 ;
        RECT 948.605 6.360 948.895 6.405 ;
        RECT 890.630 6.220 948.895 6.360 ;
        RECT 890.630 6.160 890.950 6.220 ;
        RECT 948.605 6.175 948.895 6.220 ;
        RECT 956.425 6.360 956.715 6.405 ;
        RECT 1122.025 6.360 1122.315 6.405 ;
        RECT 956.425 6.220 1122.315 6.360 ;
        RECT 956.425 6.175 956.715 6.220 ;
        RECT 1122.025 6.175 1122.315 6.220 ;
        RECT 1124.785 6.360 1125.075 6.405 ;
        RECT 1161.125 6.360 1161.415 6.405 ;
        RECT 1124.785 6.220 1161.415 6.360 ;
        RECT 1124.785 6.175 1125.075 6.220 ;
        RECT 1161.125 6.175 1161.415 6.220 ;
        RECT 1206.650 6.360 1206.970 6.420 ;
        RECT 1257.265 6.360 1257.555 6.405 ;
        RECT 1206.650 6.220 1257.555 6.360 ;
        RECT 1206.650 6.160 1206.970 6.220 ;
        RECT 1257.265 6.175 1257.555 6.220 ;
        RECT 1302.330 6.360 1302.650 6.420 ;
        RECT 1353.405 6.360 1353.695 6.405 ;
        RECT 1361.670 6.360 1361.990 6.420 ;
        RECT 1369.030 6.360 1369.350 6.420 ;
        RECT 1302.330 6.220 1353.695 6.360 ;
        RECT 1361.475 6.220 1361.990 6.360 ;
        RECT 1368.835 6.220 1369.350 6.360 ;
        RECT 1302.330 6.160 1302.650 6.220 ;
        RECT 1353.405 6.175 1353.695 6.220 ;
        RECT 1361.670 6.160 1361.990 6.220 ;
        RECT 1369.030 6.160 1369.350 6.220 ;
        RECT 1399.865 6.360 1400.155 6.405 ;
        RECT 1454.605 6.360 1454.895 6.405 ;
        RECT 1546.145 6.360 1546.435 6.405 ;
        RECT 1399.865 6.220 1454.895 6.360 ;
        RECT 1399.865 6.175 1400.155 6.220 ;
        RECT 1454.605 6.175 1454.895 6.220 ;
        RECT 1490.100 6.220 1546.435 6.360 ;
        RECT 1183.665 6.020 1183.955 6.065 ;
        RECT 1189.645 6.020 1189.935 6.065 ;
        RECT 1183.665 5.880 1189.935 6.020 ;
        RECT 1183.665 5.835 1183.955 5.880 ;
        RECT 1189.645 5.835 1189.935 5.880 ;
        RECT 1476.685 6.020 1476.975 6.065 ;
        RECT 1490.100 6.020 1490.240 6.220 ;
        RECT 1546.145 6.175 1546.435 6.220 ;
        RECT 1593.065 6.360 1593.355 6.405 ;
        RECT 1687.825 6.360 1688.115 6.405 ;
        RECT 1593.065 6.220 1635.140 6.360 ;
        RECT 1593.065 6.175 1593.355 6.220 ;
        RECT 1476.685 5.880 1490.240 6.020 ;
        RECT 1635.000 6.020 1635.140 6.220 ;
        RECT 1679.620 6.220 1688.115 6.360 ;
        RECT 1679.620 6.020 1679.760 6.220 ;
        RECT 1687.825 6.175 1688.115 6.220 ;
        RECT 1726.925 6.360 1727.215 6.405 ;
        RECT 1789.485 6.360 1789.775 6.405 ;
        RECT 1726.925 6.220 1789.775 6.360 ;
        RECT 1726.925 6.175 1727.215 6.220 ;
        RECT 1789.485 6.175 1789.775 6.220 ;
        RECT 1873.205 6.360 1873.495 6.405 ;
        RECT 1932.085 6.360 1932.375 6.405 ;
        RECT 1873.205 6.220 1932.375 6.360 ;
        RECT 1873.205 6.175 1873.495 6.220 ;
        RECT 1932.085 6.175 1932.375 6.220 ;
        RECT 2021.325 6.360 2021.615 6.405 ;
        RECT 2124.810 6.360 2125.130 6.420 ;
        RECT 2021.325 6.220 2125.130 6.360 ;
        RECT 2021.325 6.175 2021.615 6.220 ;
        RECT 2124.810 6.160 2125.130 6.220 ;
        RECT 2161.165 6.360 2161.455 6.405 ;
        RECT 2297.785 6.360 2298.075 6.405 ;
        RECT 2161.165 6.220 2298.075 6.360 ;
        RECT 2161.165 6.175 2161.455 6.220 ;
        RECT 2297.785 6.175 2298.075 6.220 ;
        RECT 2365.865 6.360 2366.155 6.405 ;
        RECT 2366.785 6.360 2367.075 6.405 ;
        RECT 2365.865 6.220 2367.075 6.360 ;
        RECT 2365.865 6.175 2366.155 6.220 ;
        RECT 2366.785 6.175 2367.075 6.220 ;
        RECT 2400.810 6.360 2401.130 6.420 ;
        RECT 2462.450 6.360 2462.770 6.420 ;
        RECT 2400.810 6.220 2462.770 6.360 ;
        RECT 2400.810 6.160 2401.130 6.220 ;
        RECT 2462.450 6.160 2462.770 6.220 ;
        RECT 2463.370 6.360 2463.690 6.420 ;
        RECT 2504.785 6.360 2505.075 6.405 ;
        RECT 2463.370 6.220 2505.075 6.360 ;
        RECT 2463.370 6.160 2463.690 6.220 ;
        RECT 2504.785 6.175 2505.075 6.220 ;
        RECT 2547.565 6.360 2547.855 6.405 ;
        RECT 2559.970 6.360 2560.290 6.420 ;
        RECT 2547.565 6.220 2560.290 6.360 ;
        RECT 2547.565 6.175 2547.855 6.220 ;
        RECT 2559.970 6.160 2560.290 6.220 ;
        RECT 2676.810 6.360 2677.130 6.420 ;
        RECT 2745.810 6.360 2746.130 6.420 ;
        RECT 2676.810 6.220 2746.130 6.360 ;
        RECT 2676.810 6.160 2677.130 6.220 ;
        RECT 2745.810 6.160 2746.130 6.220 ;
        RECT 2780.785 6.360 2781.075 6.405 ;
        RECT 2822.170 6.360 2822.490 6.420 ;
        RECT 2780.785 6.220 2822.490 6.360 ;
        RECT 2780.785 6.175 2781.075 6.220 ;
        RECT 2822.170 6.160 2822.490 6.220 ;
        RECT 1635.000 5.880 1679.760 6.020 ;
        RECT 1476.685 5.835 1476.975 5.880 ;
        RECT 771.505 5.680 771.795 5.725 ;
        RECT 787.145 5.680 787.435 5.725 ;
        RECT 771.505 5.540 787.435 5.680 ;
        RECT 771.505 5.495 771.795 5.540 ;
        RECT 787.145 5.495 787.435 5.540 ;
        RECT 1726.925 5.340 1727.215 5.385 ;
        RECT 1711.360 5.200 1727.215 5.340 ;
        RECT 1693.805 5.000 1694.095 5.045 ;
        RECT 1711.360 5.000 1711.500 5.200 ;
        RECT 1726.925 5.155 1727.215 5.200 ;
        RECT 1789.485 5.340 1789.775 5.385 ;
        RECT 1820.765 5.340 1821.055 5.385 ;
        RECT 1789.485 5.200 1821.055 5.340 ;
        RECT 1789.485 5.155 1789.775 5.200 ;
        RECT 1820.765 5.155 1821.055 5.200 ;
        RECT 2366.785 5.340 2367.075 5.385 ;
        RECT 2400.810 5.340 2401.130 5.400 ;
        RECT 2366.785 5.200 2401.130 5.340 ;
        RECT 2366.785 5.155 2367.075 5.200 ;
        RECT 2400.810 5.140 2401.130 5.200 ;
        RECT 2583.905 5.340 2584.195 5.385 ;
        RECT 2676.810 5.340 2677.130 5.400 ;
        RECT 2583.905 5.200 2677.130 5.340 ;
        RECT 2583.905 5.155 2584.195 5.200 ;
        RECT 2676.810 5.140 2677.130 5.200 ;
        RECT 1693.805 4.860 1711.500 5.000 ;
        RECT 1693.805 4.815 1694.095 4.860 ;
        RECT 813.365 4.660 813.655 4.705 ;
        RECT 815.205 4.660 815.495 4.705 ;
        RECT 813.365 4.520 815.495 4.660 ;
        RECT 813.365 4.475 813.655 4.520 ;
        RECT 815.205 4.475 815.495 4.520 ;
        RECT 1821.685 4.660 1821.975 4.705 ;
        RECT 1842.385 4.660 1842.675 4.705 ;
        RECT 1821.685 4.520 1842.675 4.660 ;
        RECT 1821.685 4.475 1821.975 4.520 ;
        RECT 1842.385 4.475 1842.675 4.520 ;
        RECT 2559.970 4.660 2560.290 4.720 ;
        RECT 2583.905 4.660 2584.195 4.705 ;
        RECT 2559.970 4.520 2584.195 4.660 ;
        RECT 2559.970 4.460 2560.290 4.520 ;
        RECT 2583.905 4.475 2584.195 4.520 ;
        RECT 606.825 4.320 607.115 4.365 ;
        RECT 766.445 4.320 766.735 4.365 ;
        RECT 606.825 4.180 766.735 4.320 ;
        RECT 606.825 4.135 607.115 4.180 ;
        RECT 766.445 4.135 766.735 4.180 ;
        RECT 787.145 4.320 787.435 4.365 ;
        RECT 805.085 4.320 805.375 4.365 ;
        RECT 787.145 4.180 805.375 4.320 ;
        RECT 787.145 4.135 787.435 4.180 ;
        RECT 805.085 4.135 805.375 4.180 ;
        RECT 1932.545 4.320 1932.835 4.365 ;
        RECT 2021.325 4.320 2021.615 4.365 ;
        RECT 1932.545 4.180 2021.615 4.320 ;
        RECT 1932.545 4.135 1932.835 4.180 ;
        RECT 2021.325 4.135 2021.615 4.180 ;
        RECT 769.665 3.980 769.955 4.025 ;
        RECT 771.505 3.980 771.795 4.025 ;
        RECT 769.665 3.840 771.795 3.980 ;
        RECT 769.665 3.795 769.955 3.840 ;
        RECT 771.505 3.795 771.795 3.840 ;
        RECT 805.085 3.300 805.375 3.345 ;
        RECT 811.065 3.300 811.355 3.345 ;
        RECT 805.085 3.160 811.355 3.300 ;
        RECT 805.085 3.115 805.375 3.160 ;
        RECT 811.065 3.115 811.355 3.160 ;
        RECT 1687.825 2.620 1688.115 2.665 ;
        RECT 1693.805 2.620 1694.095 2.665 ;
        RECT 1687.825 2.480 1694.095 2.620 ;
        RECT 1687.825 2.435 1688.115 2.480 ;
        RECT 1693.805 2.435 1694.095 2.480 ;
      LAYER via ;
        RECT 2746.300 7.860 2746.560 8.120 ;
        RECT 2125.300 7.520 2125.560 7.780 ;
        RECT 889.280 7.180 889.540 7.440 ;
        RECT 1206.680 7.180 1206.940 7.440 ;
        RECT 1361.700 7.180 1361.960 7.440 ;
        RECT 1369.060 7.180 1369.320 7.440 ;
        RECT 1295.460 6.840 1295.720 7.100 ;
        RECT 583.840 6.160 584.100 6.420 ;
        RECT 890.660 6.160 890.920 6.420 ;
        RECT 1206.680 6.160 1206.940 6.420 ;
        RECT 1302.360 6.160 1302.620 6.420 ;
        RECT 1361.700 6.160 1361.960 6.420 ;
        RECT 1369.060 6.160 1369.320 6.420 ;
        RECT 2124.840 6.160 2125.100 6.420 ;
        RECT 2400.840 6.160 2401.100 6.420 ;
        RECT 2462.480 6.160 2462.740 6.420 ;
        RECT 2463.400 6.160 2463.660 6.420 ;
        RECT 2560.000 6.160 2560.260 6.420 ;
        RECT 2676.840 6.160 2677.100 6.420 ;
        RECT 2745.840 6.160 2746.100 6.420 ;
        RECT 2822.200 6.160 2822.460 6.420 ;
        RECT 2400.840 5.140 2401.100 5.400 ;
        RECT 2676.840 5.140 2677.100 5.400 ;
        RECT 2560.000 4.460 2560.260 4.720 ;
      LAYER met2 ;
        RECT 1724.570 3403.130 1724.850 3405.000 ;
        RECT 1725.090 3403.130 1725.370 3403.245 ;
        RECT 1724.570 3402.990 1725.370 3403.130 ;
        RECT 1724.570 3401.000 1724.850 3402.990 ;
        RECT 1725.090 3402.875 1725.370 3402.990 ;
        RECT 2746.300 7.830 2746.560 8.150 ;
        RECT 2125.300 7.490 2125.560 7.810 ;
        RECT 889.280 7.380 889.540 7.470 ;
        RECT 889.280 7.240 890.860 7.380 ;
        RECT 889.280 7.150 889.540 7.240 ;
        RECT 890.720 6.450 890.860 7.240 ;
        RECT 1206.680 7.150 1206.940 7.470 ;
        RECT 1206.740 6.450 1206.880 7.150 ;
        RECT 1295.450 6.955 1295.730 7.325 ;
        RECT 1302.350 6.955 1302.630 7.325 ;
        RECT 1361.700 7.150 1361.960 7.470 ;
        RECT 1369.060 7.150 1369.320 7.470 ;
        RECT 1295.460 6.810 1295.720 6.955 ;
        RECT 1302.420 6.450 1302.560 6.955 ;
        RECT 1361.760 6.450 1361.900 7.150 ;
        RECT 1369.120 6.450 1369.260 7.150 ;
        RECT 2125.360 6.530 2125.500 7.490 ;
        RECT 2746.360 6.530 2746.500 7.830 ;
        RECT 2124.900 6.450 2125.500 6.530 ;
        RECT 2745.900 6.450 2746.500 6.530 ;
        RECT 583.840 6.130 584.100 6.450 ;
        RECT 890.660 6.130 890.920 6.450 ;
        RECT 1206.680 6.130 1206.940 6.450 ;
        RECT 1302.360 6.130 1302.620 6.450 ;
        RECT 1361.700 6.130 1361.960 6.450 ;
        RECT 1369.060 6.130 1369.320 6.450 ;
        RECT 2124.840 6.390 2125.500 6.450 ;
        RECT 2124.840 6.130 2125.100 6.390 ;
        RECT 2400.840 6.130 2401.100 6.450 ;
        RECT 2462.480 6.130 2462.740 6.450 ;
        RECT 2463.400 6.130 2463.660 6.450 ;
        RECT 2560.000 6.130 2560.260 6.450 ;
        RECT 2676.840 6.130 2677.100 6.450 ;
        RECT 2745.840 6.390 2746.500 6.450 ;
        RECT 2745.840 6.130 2746.100 6.390 ;
        RECT 2822.190 6.275 2822.470 6.645 ;
        RECT 2822.200 6.130 2822.460 6.275 ;
        RECT 583.900 5.850 584.040 6.130 ;
        RECT 582.060 5.710 584.040 5.850 ;
        RECT 582.060 3.925 582.200 5.710 ;
        RECT 2400.900 5.430 2401.040 6.130 ;
        RECT 2400.840 5.110 2401.100 5.430 ;
        RECT 2462.540 5.340 2462.680 6.130 ;
        RECT 2463.460 5.340 2463.600 6.130 ;
        RECT 2462.540 5.200 2463.600 5.340 ;
        RECT 2560.060 4.750 2560.200 6.130 ;
        RECT 2676.900 5.430 2677.040 6.130 ;
        RECT 2676.840 5.110 2677.100 5.430 ;
        RECT 2560.000 4.430 2560.260 4.750 ;
        RECT 581.990 3.555 582.270 3.925 ;
        RECT 561.750 2.875 562.030 3.245 ;
        RECT 561.820 2.400 561.960 2.875 ;
        RECT 561.610 -4.800 562.170 2.400 ;
      LAYER via2 ;
        RECT 1725.090 3402.920 1725.370 3403.200 ;
        RECT 1295.450 7.000 1295.730 7.280 ;
        RECT 1302.350 7.000 1302.630 7.280 ;
        RECT 2822.190 6.320 2822.470 6.600 ;
        RECT 581.990 3.600 582.270 3.880 ;
        RECT 561.750 2.920 562.030 3.200 ;
      LAYER met3 ;
        RECT 1724.350 3403.210 1724.730 3403.220 ;
        RECT 1725.065 3403.210 1725.395 3403.225 ;
        RECT 1724.350 3402.910 1725.395 3403.210 ;
        RECT 1724.350 3402.900 1724.730 3402.910 ;
        RECT 1725.065 3402.895 1725.395 3402.910 ;
        RECT 1295.425 7.290 1295.755 7.305 ;
        RECT 1302.325 7.290 1302.655 7.305 ;
        RECT 1295.425 6.990 1302.655 7.290 ;
        RECT 1295.425 6.975 1295.755 6.990 ;
        RECT 1302.325 6.975 1302.655 6.990 ;
        RECT 2822.165 6.610 2822.495 6.625 ;
        RECT 2824.670 6.610 2825.050 6.620 ;
        RECT 2822.165 6.310 2825.050 6.610 ;
        RECT 2822.165 6.295 2822.495 6.310 ;
        RECT 2824.670 6.300 2825.050 6.310 ;
        RECT 581.965 3.890 582.295 3.905 ;
        RECT 569.790 3.590 582.295 3.890 ;
        RECT 561.725 3.210 562.055 3.225 ;
        RECT 569.790 3.210 570.090 3.590 ;
        RECT 581.965 3.575 582.295 3.590 ;
        RECT 561.725 2.910 570.090 3.210 ;
        RECT 561.725 2.895 562.055 2.910 ;
      LAYER via3 ;
        RECT 1724.380 3402.900 1724.700 3403.220 ;
        RECT 2824.700 6.300 2825.020 6.620 ;
      LAYER met4 ;
        RECT 1724.375 3402.895 1724.705 3403.225 ;
        RECT 1724.390 3402.290 1724.690 3402.895 ;
        RECT 1723.950 3401.110 1725.130 3402.290 ;
        RECT 2824.270 3401.110 2825.450 3402.290 ;
        RECT 2824.710 6.625 2825.010 3401.110 ;
        RECT 2824.695 6.295 2825.025 6.625 ;
      LAYER met5 ;
        RECT 1821.260 3407.700 1850.460 3409.300 ;
        RECT 1821.260 3402.500 1822.860 3407.700 ;
        RECT 1848.860 3405.900 1850.460 3407.700 ;
        RECT 2330.940 3407.700 2336.220 3409.300 ;
        RECT 2330.940 3405.900 2332.540 3407.700 ;
        RECT 1848.860 3404.300 1897.380 3405.900 ;
        RECT 1723.740 3400.900 1822.860 3402.500 ;
        RECT 1895.780 3402.500 1897.380 3404.300 ;
        RECT 2283.100 3404.300 2332.540 3405.900 ;
        RECT 2334.620 3405.900 2336.220 3407.700 ;
        RECT 2379.700 3407.700 2432.820 3409.300 ;
        RECT 2379.700 3405.900 2381.300 3407.700 ;
        RECT 2334.620 3404.300 2381.300 3405.900 ;
        RECT 2431.220 3405.900 2432.820 3407.700 ;
        RECT 2476.300 3407.700 2528.500 3409.300 ;
        RECT 2476.300 3405.900 2477.900 3407.700 ;
        RECT 2431.220 3404.300 2477.900 3405.900 ;
        RECT 2526.900 3405.900 2528.500 3407.700 ;
        RECT 2526.900 3404.300 2573.580 3405.900 ;
        RECT 2283.100 3402.500 2284.700 3404.300 ;
        RECT 1895.780 3400.900 2284.700 3402.500 ;
        RECT 2571.980 3402.500 2573.580 3404.300 ;
        RECT 2571.980 3400.900 2825.660 3402.500 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2405.025 3401.445 2405.655 3401.615 ;
        RECT 2405.485 3399.745 2405.655 3401.445 ;
        RECT 2448.725 3399.745 2448.895 3401.615 ;
        RECT 2767.505 3399.065 2767.675 3401.615 ;
        RECT 2808.905 3399.065 2809.075 3401.615 ;
        RECT 640.465 10.285 648.915 10.455 ;
        RECT 507.065 9.265 530.695 9.435 ;
        RECT 290.405 7.565 291.495 7.735 ;
        RECT 507.065 7.565 507.235 9.265 ;
        RECT 530.525 8.925 530.695 9.265 ;
        RECT 534.205 8.925 550.015 9.095 ;
        RECT 290.405 6.545 290.575 7.565 ;
        RECT 379.185 2.975 379.355 3.315 ;
        RECT 383.325 2.975 383.495 3.995 ;
        RECT 394.825 3.825 394.995 5.695 ;
        RECT 413.685 5.525 413.855 7.395 ;
        RECT 415.985 7.225 417.075 7.395 ;
        RECT 549.845 6.885 550.015 8.925 ;
        RECT 582.045 8.585 607.975 8.755 ;
        RECT 640.465 8.585 640.635 10.285 ;
        RECT 648.745 10.115 648.915 10.285 ;
        RECT 648.745 9.945 672.835 10.115 ;
        RECT 672.665 9.775 672.835 9.945 ;
        RECT 1070.565 9.945 1110.755 10.115 ;
        RECT 672.665 9.605 694.455 9.775 ;
        RECT 694.285 9.095 694.455 9.605 ;
        RECT 695.665 9.605 709.175 9.775 ;
        RECT 695.665 9.095 695.835 9.605 ;
        RECT 694.285 8.925 695.835 9.095 ;
        RECT 709.005 8.755 709.175 9.605 ;
        RECT 724.645 9.265 734.015 9.435 ;
        RECT 673.585 8.585 693.075 8.755 ;
        RECT 709.005 8.585 722.975 8.755 ;
        RECT 555.825 3.825 555.995 7.055 ;
        RECT 574.225 4.165 574.395 7.395 ;
        RECT 582.045 5.695 582.215 8.585 ;
        RECT 580.665 5.525 582.215 5.695 ;
        RECT 580.665 5.355 580.835 5.525 ;
        RECT 580.205 5.185 580.835 5.355 ;
        RECT 580.205 4.675 580.375 5.185 ;
        RECT 609.645 4.845 609.815 7.055 ;
        RECT 645.065 6.545 647.075 6.715 ;
        RECT 645.065 5.695 645.235 6.545 ;
        RECT 646.905 6.205 647.075 6.545 ;
        RECT 672.205 6.205 672.375 7.055 ;
        RECT 673.585 6.885 673.755 8.585 ;
        RECT 692.905 8.245 693.075 8.585 ;
        RECT 722.805 7.735 722.975 8.585 ;
        RECT 724.645 7.735 724.815 9.265 ;
        RECT 733.845 8.755 734.015 9.265 ;
        RECT 760.985 9.265 767.135 9.435 ;
        RECT 740.285 8.755 740.455 9.095 ;
        RECT 733.845 8.585 740.455 8.755 ;
        RECT 722.805 7.565 724.815 7.735 ;
        RECT 742.585 7.735 742.755 9.095 ;
        RECT 745.345 8.755 745.515 9.095 ;
        RECT 746.265 8.925 751.035 9.095 ;
        RECT 746.265 8.755 746.435 8.925 ;
        RECT 745.345 8.585 746.435 8.755 ;
        RECT 744.885 8.245 745.975 8.415 ;
        RECT 744.885 7.735 745.055 8.245 ;
        RECT 745.805 7.905 745.975 8.245 ;
        RECT 742.585 7.565 745.055 7.735 ;
        RECT 747.645 7.225 747.815 8.075 ;
        RECT 750.865 7.055 751.035 8.925 ;
        RECT 755.465 8.925 757.015 9.095 ;
        RECT 750.865 6.885 751.495 7.055 ;
        RECT 629.885 5.525 645.235 5.695 ;
        RECT 629.885 5.015 630.055 5.525 ;
        RECT 576.065 4.505 580.375 4.675 ;
        RECT 611.945 4.675 612.115 5.015 ;
        RECT 621.145 4.845 621.775 5.015 ;
        RECT 627.585 4.845 630.055 5.015 ;
        RECT 611.945 4.505 613.495 4.675 ;
        RECT 558.585 3.825 559.215 3.995 ;
        RECT 559.045 3.655 559.215 3.825 ;
        RECT 576.065 3.655 576.235 4.505 ;
        RECT 621.145 4.335 621.315 4.845 ;
        RECT 610.565 4.165 621.315 4.335 ;
        RECT 751.325 4.335 751.495 6.885 ;
        RECT 752.245 6.205 752.415 7.395 ;
        RECT 755.465 6.205 755.635 8.925 ;
        RECT 756.845 8.585 757.015 8.925 ;
        RECT 760.065 8.415 760.235 8.755 ;
        RECT 760.985 8.415 761.155 9.265 ;
        RECT 766.965 8.925 767.135 9.265 ;
        RECT 760.065 8.245 761.155 8.415 ;
        RECT 771.105 8.415 771.275 9.095 ;
        RECT 794.105 8.585 802.555 8.755 ;
        RECT 771.105 8.245 776.335 8.415 ;
        RECT 764.665 6.545 765.755 6.715 ;
        RECT 764.665 4.675 764.835 6.545 ;
        RECT 762.825 4.505 764.835 4.675 ;
        RECT 762.825 4.335 762.995 4.505 ;
        RECT 751.325 4.165 762.995 4.335 ;
        RECT 559.045 3.485 576.235 3.655 ;
        RECT 606.425 3.655 606.595 3.995 ;
        RECT 606.425 3.485 607.975 3.655 ;
        RECT 607.805 3.145 607.975 3.485 ;
        RECT 610.565 3.145 610.735 4.165 ;
        RECT 379.185 2.805 383.495 2.975 ;
        RECT 765.585 2.975 765.755 6.545 ;
        RECT 776.165 4.505 776.335 8.245 ;
        RECT 794.105 6.035 794.275 8.585 ;
        RECT 802.385 8.245 802.555 8.585 ;
        RECT 823.085 8.245 846.255 8.415 ;
        RECT 796.405 7.905 798.415 8.075 ;
        RECT 789.045 5.865 794.275 6.035 ;
        RECT 789.045 3.825 789.215 5.865 ;
        RECT 798.245 5.355 798.415 7.905 ;
        RECT 823.085 7.225 823.255 8.245 ;
        RECT 878.745 7.565 878.915 8.755 ;
        RECT 798.245 5.185 800.255 5.355 ;
        RECT 800.085 3.485 800.255 5.185 ;
        RECT 812.965 4.845 814.055 5.015 ;
        RECT 812.965 3.995 813.135 4.845 ;
        RECT 807.905 3.825 813.135 3.995 ;
        RECT 765.585 2.805 769.895 2.975 ;
        RECT 769.725 0.595 769.895 2.805 ;
        RECT 803.305 2.295 803.475 3.655 ;
        RECT 807.905 2.295 808.075 3.825 ;
        RECT 803.305 2.125 808.075 2.295 ;
        RECT 813.885 0.935 814.055 4.845 ;
        RECT 814.805 2.635 814.975 7.055 ;
        RECT 888.865 6.375 889.035 8.755 ;
        RECT 889.325 8.245 890.415 8.415 ;
        RECT 889.325 7.905 889.495 8.245 ;
        RECT 890.245 7.225 890.415 8.245 ;
        RECT 894.845 7.225 895.015 8.075 ;
        RECT 951.885 7.905 954.355 8.075 ;
        RECT 1070.565 7.905 1070.735 9.945 ;
        RECT 1110.585 7.905 1110.755 9.945 ;
        RECT 1123.005 8.075 1123.175 8.415 ;
        RECT 1123.005 7.905 1125.015 8.075 ;
        RECT 1163.025 7.905 1163.195 9.095 ;
        RECT 1169.925 7.905 1170.095 8.755 ;
        RECT 951.885 7.225 952.055 7.905 ;
        RECT 888.865 6.205 889.495 6.375 ;
        RECT 1021.345 3.485 1022.895 3.655 ;
        RECT 1040.665 3.315 1040.835 3.655 ;
        RECT 1042.045 3.485 1044.055 3.655 ;
        RECT 1069.645 3.485 1071.655 3.655 ;
        RECT 1042.045 3.315 1042.215 3.485 ;
        RECT 1040.665 3.145 1042.215 3.315 ;
        RECT 1306.545 2.975 1306.715 3.655 ;
        RECT 1316.205 2.975 1316.375 9.095 ;
        RECT 1401.305 8.925 1409.755 9.095 ;
        RECT 1399.925 8.415 1400.095 8.755 ;
        RECT 1401.305 8.415 1401.475 8.925 ;
        RECT 1399.925 8.245 1401.475 8.415 ;
        RECT 1409.585 7.225 1409.755 8.925 ;
        RECT 1306.545 2.805 1316.375 2.975 ;
        RECT 814.805 2.465 815.895 2.635 ;
        RECT 1617.045 2.465 1617.215 4.675 ;
        RECT 812.045 0.765 814.515 0.935 ;
        RECT 812.045 0.595 812.215 0.765 ;
        RECT 769.725 0.425 812.215 0.595 ;
        RECT 813.885 0.255 814.055 0.765 ;
        RECT 814.345 0.595 814.515 0.765 ;
        RECT 815.725 0.595 815.895 2.465 ;
        RECT 852.525 2.125 856.375 2.295 ;
        RECT 852.525 1.615 852.695 2.125 ;
        RECT 814.345 0.425 815.895 0.595 ;
        RECT 820.785 1.445 852.695 1.615 ;
        RECT 856.205 1.615 856.375 2.125 ;
        RECT 856.205 1.445 876.615 1.615 ;
        RECT 820.785 0.255 820.955 1.445 ;
        RECT 876.445 0.935 876.615 1.445 ;
        RECT 876.445 0.765 918.935 0.935 ;
        RECT 813.885 0.085 820.955 0.255 ;
      LAYER mcon ;
        RECT 2448.725 3401.445 2448.895 3401.615 ;
        RECT 2767.505 3401.445 2767.675 3401.615 ;
        RECT 2808.905 3401.445 2809.075 3401.615 ;
        RECT 291.325 7.565 291.495 7.735 ;
        RECT 413.685 7.225 413.855 7.395 ;
        RECT 416.905 7.225 417.075 7.395 ;
        RECT 607.805 8.585 607.975 8.755 ;
        RECT 574.225 7.225 574.395 7.395 ;
        RECT 555.825 6.885 555.995 7.055 ;
        RECT 394.825 5.525 394.995 5.695 ;
        RECT 383.325 3.825 383.495 3.995 ;
        RECT 740.285 8.925 740.455 9.095 ;
        RECT 742.585 8.925 742.755 9.095 ;
        RECT 745.345 8.925 745.515 9.095 ;
        RECT 747.645 7.905 747.815 8.075 ;
        RECT 609.645 6.885 609.815 7.055 ;
        RECT 672.205 6.885 672.375 7.055 ;
        RECT 752.245 7.225 752.415 7.395 ;
        RECT 611.945 4.845 612.115 5.015 ;
        RECT 621.605 4.845 621.775 5.015 ;
        RECT 613.325 4.505 613.495 4.675 ;
        RECT 379.185 3.145 379.355 3.315 ;
        RECT 760.065 8.585 760.235 8.755 ;
        RECT 771.105 8.925 771.275 9.095 ;
        RECT 606.425 3.825 606.595 3.995 ;
        RECT 878.745 8.585 878.915 8.755 ;
        RECT 846.085 8.245 846.255 8.415 ;
        RECT 888.865 8.585 889.035 8.755 ;
        RECT 814.805 6.885 814.975 7.055 ;
        RECT 803.305 3.485 803.475 3.655 ;
        RECT 894.845 7.905 895.015 8.075 ;
        RECT 954.185 7.905 954.355 8.075 ;
        RECT 1163.025 8.925 1163.195 9.095 ;
        RECT 1123.005 8.245 1123.175 8.415 ;
        RECT 1316.205 8.925 1316.375 9.095 ;
        RECT 1124.845 7.905 1125.015 8.075 ;
        RECT 1169.925 8.585 1170.095 8.755 ;
        RECT 889.325 6.205 889.495 6.375 ;
        RECT 1022.725 3.485 1022.895 3.655 ;
        RECT 1040.665 3.485 1040.835 3.655 ;
        RECT 1043.885 3.485 1044.055 3.655 ;
        RECT 1071.485 3.485 1071.655 3.655 ;
        RECT 1306.545 3.485 1306.715 3.655 ;
        RECT 1399.925 8.585 1400.095 8.755 ;
        RECT 1617.045 4.505 1617.215 4.675 ;
        RECT 918.765 0.765 918.935 0.935 ;
      LAYER met1 ;
        RECT 1822.590 3416.220 1822.910 3416.280 ;
        RECT 1876.870 3416.220 1877.190 3416.280 ;
        RECT 1822.590 3416.080 1877.190 3416.220 ;
        RECT 1822.590 3416.020 1822.910 3416.080 ;
        RECT 1876.870 3416.020 1877.190 3416.080 ;
        RECT 2041.640 3402.140 2042.700 3402.280 ;
        RECT 1876.870 3401.600 1877.190 3401.660 ;
        RECT 2041.640 3401.600 2041.780 3402.140 ;
        RECT 1876.870 3401.460 2041.780 3401.600 ;
        RECT 2042.560 3401.600 2042.700 3402.140 ;
        RECT 2404.965 3401.600 2405.255 3401.645 ;
        RECT 2042.560 3401.460 2405.255 3401.600 ;
        RECT 1876.870 3401.400 1877.190 3401.460 ;
        RECT 2404.965 3401.415 2405.255 3401.460 ;
        RECT 2448.665 3401.600 2448.955 3401.645 ;
        RECT 2767.445 3401.600 2767.735 3401.645 ;
        RECT 2808.830 3401.600 2809.150 3401.660 ;
        RECT 2448.665 3401.460 2767.735 3401.600 ;
        RECT 2808.635 3401.460 2809.150 3401.600 ;
        RECT 2448.665 3401.415 2448.955 3401.460 ;
        RECT 2767.445 3401.415 2767.735 3401.460 ;
        RECT 2808.830 3401.400 2809.150 3401.460 ;
        RECT 2405.425 3399.900 2405.715 3399.945 ;
        RECT 2448.665 3399.900 2448.955 3399.945 ;
        RECT 2405.425 3399.760 2448.955 3399.900 ;
        RECT 2405.425 3399.715 2405.715 3399.760 ;
        RECT 2448.665 3399.715 2448.955 3399.760 ;
        RECT 2767.445 3399.220 2767.735 3399.265 ;
        RECT 2808.845 3399.220 2809.135 3399.265 ;
        RECT 2767.445 3399.080 2809.135 3399.220 ;
        RECT 2767.445 3399.035 2767.735 3399.080 ;
        RECT 2808.845 3399.035 2809.135 3399.080 ;
        RECT 530.465 9.080 530.755 9.125 ;
        RECT 534.145 9.080 534.435 9.125 ;
        RECT 530.465 8.940 534.435 9.080 ;
        RECT 530.465 8.895 530.755 8.940 ;
        RECT 534.145 8.895 534.435 8.940 ;
        RECT 740.225 9.080 740.515 9.125 ;
        RECT 742.525 9.080 742.815 9.125 ;
        RECT 745.285 9.080 745.575 9.125 ;
        RECT 740.225 8.940 742.815 9.080 ;
        RECT 740.225 8.895 740.515 8.940 ;
        RECT 742.525 8.895 742.815 8.940 ;
        RECT 743.060 8.940 745.575 9.080 ;
        RECT 743.060 8.800 743.200 8.940 ;
        RECT 745.285 8.895 745.575 8.940 ;
        RECT 766.905 9.080 767.195 9.125 ;
        RECT 771.045 9.080 771.335 9.125 ;
        RECT 1162.965 9.080 1163.255 9.125 ;
        RECT 766.905 8.940 771.335 9.080 ;
        RECT 766.905 8.895 767.195 8.940 ;
        RECT 771.045 8.895 771.335 8.940 ;
        RECT 1161.200 8.940 1163.255 9.080 ;
        RECT 607.745 8.740 608.035 8.785 ;
        RECT 640.405 8.740 640.695 8.785 ;
        RECT 607.745 8.600 640.695 8.740 ;
        RECT 607.745 8.555 608.035 8.600 ;
        RECT 640.405 8.555 640.695 8.600 ;
        RECT 742.970 8.540 743.290 8.800 ;
        RECT 756.785 8.740 757.075 8.785 ;
        RECT 760.005 8.740 760.295 8.785 ;
        RECT 756.785 8.600 760.295 8.740 ;
        RECT 756.785 8.555 757.075 8.600 ;
        RECT 760.005 8.555 760.295 8.600 ;
        RECT 878.685 8.740 878.975 8.785 ;
        RECT 888.805 8.740 889.095 8.785 ;
        RECT 1161.200 8.740 1161.340 8.940 ;
        RECT 1162.965 8.895 1163.255 8.940 ;
        RECT 1316.145 9.080 1316.435 9.125 ;
        RECT 1316.145 8.940 1344.420 9.080 ;
        RECT 1316.145 8.895 1316.435 8.940 ;
        RECT 878.685 8.600 889.095 8.740 ;
        RECT 878.685 8.555 878.975 8.600 ;
        RECT 888.805 8.555 889.095 8.600 ;
        RECT 1159.820 8.600 1161.340 8.740 ;
        RECT 1169.865 8.740 1170.155 8.785 ;
        RECT 1182.730 8.740 1183.050 8.800 ;
        RECT 1169.865 8.600 1183.050 8.740 ;
        RECT 1344.280 8.740 1344.420 8.940 ;
        RECT 1399.865 8.740 1400.155 8.785 ;
        RECT 1344.280 8.600 1400.155 8.740 ;
        RECT 692.845 8.400 693.135 8.445 ;
        RECT 693.750 8.400 694.070 8.460 ;
        RECT 692.845 8.260 694.070 8.400 ;
        RECT 692.845 8.215 693.135 8.260 ;
        RECT 693.750 8.200 694.070 8.260 ;
        RECT 802.325 8.400 802.615 8.445 ;
        RECT 846.025 8.400 846.315 8.445 ;
        RECT 847.850 8.400 848.170 8.460 ;
        RECT 1122.945 8.400 1123.235 8.445 ;
        RECT 802.325 8.260 804.840 8.400 ;
        RECT 802.325 8.215 802.615 8.260 ;
        RECT 745.745 8.060 746.035 8.105 ;
        RECT 747.585 8.060 747.875 8.105 ;
        RECT 745.745 7.920 747.875 8.060 ;
        RECT 745.745 7.875 746.035 7.920 ;
        RECT 747.585 7.875 747.875 7.920 ;
        RECT 794.030 8.060 794.350 8.120 ;
        RECT 796.345 8.060 796.635 8.105 ;
        RECT 794.030 7.920 796.635 8.060 ;
        RECT 804.700 8.060 804.840 8.260 ;
        RECT 846.025 8.260 848.170 8.400 ;
        RECT 846.025 8.215 846.315 8.260 ;
        RECT 847.850 8.200 848.170 8.260 ;
        RECT 1120.720 8.260 1123.235 8.400 ;
        RECT 889.265 8.060 889.555 8.105 ;
        RECT 804.700 7.920 805.300 8.060 ;
        RECT 794.030 7.860 794.350 7.920 ;
        RECT 796.345 7.875 796.635 7.920 ;
        RECT 291.265 7.720 291.555 7.765 ;
        RECT 296.310 7.720 296.630 7.780 ;
        RECT 507.005 7.720 507.295 7.765 ;
        RECT 291.265 7.580 296.630 7.720 ;
        RECT 291.265 7.535 291.555 7.580 ;
        RECT 296.310 7.520 296.630 7.580 ;
        RECT 438.080 7.580 507.295 7.720 ;
        RECT 413.625 7.380 413.915 7.425 ;
        RECT 415.925 7.380 416.215 7.425 ;
        RECT 413.625 7.240 416.215 7.380 ;
        RECT 413.625 7.195 413.915 7.240 ;
        RECT 415.925 7.195 416.215 7.240 ;
        RECT 416.845 7.380 417.135 7.425 ;
        RECT 438.080 7.380 438.220 7.580 ;
        RECT 507.005 7.535 507.295 7.580 ;
        RECT 508.370 7.720 508.690 7.780 ;
        RECT 511.130 7.720 511.450 7.780 ;
        RECT 508.370 7.580 511.450 7.720 ;
        RECT 805.160 7.720 805.300 7.920 ;
        RECT 848.860 7.920 889.555 8.060 ;
        RECT 848.860 7.720 849.000 7.920 ;
        RECT 889.265 7.875 889.555 7.920 ;
        RECT 894.785 8.060 895.075 8.105 ;
        RECT 919.610 8.060 919.930 8.120 ;
        RECT 894.785 7.920 919.930 8.060 ;
        RECT 894.785 7.875 895.075 7.920 ;
        RECT 919.610 7.860 919.930 7.920 ;
        RECT 954.125 8.060 954.415 8.105 ;
        RECT 1070.505 8.060 1070.795 8.105 ;
        RECT 954.125 7.920 1070.795 8.060 ;
        RECT 954.125 7.875 954.415 7.920 ;
        RECT 1070.505 7.875 1070.795 7.920 ;
        RECT 1110.525 8.060 1110.815 8.105 ;
        RECT 1120.720 8.060 1120.860 8.260 ;
        RECT 1122.945 8.215 1123.235 8.260 ;
        RECT 1110.525 7.920 1120.860 8.060 ;
        RECT 1124.785 8.060 1125.075 8.105 ;
        RECT 1159.820 8.060 1159.960 8.600 ;
        RECT 1169.865 8.555 1170.155 8.600 ;
        RECT 1182.730 8.540 1183.050 8.600 ;
        RECT 1399.865 8.555 1400.155 8.600 ;
        RECT 1124.785 7.920 1159.960 8.060 ;
        RECT 1162.965 8.060 1163.255 8.105 ;
        RECT 1169.865 8.060 1170.155 8.105 ;
        RECT 1162.965 7.920 1170.155 8.060 ;
        RECT 1110.525 7.875 1110.815 7.920 ;
        RECT 1124.785 7.875 1125.075 7.920 ;
        RECT 1162.965 7.875 1163.255 7.920 ;
        RECT 1169.865 7.875 1170.155 7.920 ;
        RECT 805.160 7.580 849.000 7.720 ;
        RECT 849.230 7.720 849.550 7.780 ;
        RECT 878.685 7.720 878.975 7.765 ;
        RECT 849.230 7.580 878.975 7.720 ;
        RECT 508.370 7.520 508.690 7.580 ;
        RECT 511.130 7.520 511.450 7.580 ;
        RECT 849.230 7.520 849.550 7.580 ;
        RECT 878.685 7.535 878.975 7.580 ;
        RECT 416.845 7.240 438.220 7.380 ;
        RECT 556.210 7.380 556.530 7.440 ;
        RECT 574.165 7.380 574.455 7.425 ;
        RECT 556.210 7.240 574.455 7.380 ;
        RECT 416.845 7.195 417.135 7.240 ;
        RECT 556.210 7.180 556.530 7.240 ;
        RECT 574.165 7.195 574.455 7.240 ;
        RECT 747.585 7.380 747.875 7.425 ;
        RECT 752.185 7.380 752.475 7.425 ;
        RECT 747.585 7.240 752.475 7.380 ;
        RECT 747.585 7.195 747.875 7.240 ;
        RECT 752.185 7.195 752.475 7.240 ;
        RECT 823.025 7.195 823.315 7.425 ;
        RECT 890.185 7.380 890.475 7.425 ;
        RECT 894.785 7.380 895.075 7.425 ;
        RECT 951.810 7.380 952.130 7.440 ;
        RECT 890.185 7.240 895.075 7.380 ;
        RECT 951.615 7.240 952.130 7.380 ;
        RECT 890.185 7.195 890.475 7.240 ;
        RECT 894.785 7.195 895.075 7.240 ;
        RECT 549.785 7.040 550.075 7.085 ;
        RECT 555.765 7.040 556.055 7.085 ;
        RECT 549.785 6.900 556.055 7.040 ;
        RECT 549.785 6.855 550.075 6.900 ;
        RECT 555.765 6.855 556.055 6.900 ;
        RECT 604.970 7.040 605.290 7.100 ;
        RECT 609.585 7.040 609.875 7.085 ;
        RECT 604.970 6.900 609.875 7.040 ;
        RECT 604.970 6.840 605.290 6.900 ;
        RECT 609.585 6.855 609.875 6.900 ;
        RECT 672.145 7.040 672.435 7.085 ;
        RECT 673.525 7.040 673.815 7.085 ;
        RECT 672.145 6.900 673.815 7.040 ;
        RECT 672.145 6.855 672.435 6.900 ;
        RECT 673.525 6.855 673.815 6.900 ;
        RECT 673.970 7.040 674.290 7.100 ;
        RECT 679.030 7.040 679.350 7.100 ;
        RECT 673.970 6.900 679.350 7.040 ;
        RECT 673.970 6.840 674.290 6.900 ;
        RECT 679.030 6.840 679.350 6.900 ;
        RECT 693.750 7.040 694.070 7.100 ;
        RECT 695.590 7.040 695.910 7.100 ;
        RECT 693.750 6.900 695.910 7.040 ;
        RECT 693.750 6.840 694.070 6.900 ;
        RECT 695.590 6.840 695.910 6.900 ;
        RECT 814.745 7.040 815.035 7.085 ;
        RECT 823.100 7.040 823.240 7.195 ;
        RECT 951.810 7.180 952.130 7.240 ;
        RECT 1409.525 7.380 1409.815 7.425 ;
        RECT 1410.430 7.380 1410.750 7.440 ;
        RECT 1409.525 7.240 1410.750 7.380 ;
        RECT 1409.525 7.195 1409.815 7.240 ;
        RECT 1410.430 7.180 1410.750 7.240 ;
        RECT 814.745 6.900 823.240 7.040 ;
        RECT 814.745 6.855 815.035 6.900 ;
        RECT 275.150 6.700 275.470 6.760 ;
        RECT 290.345 6.700 290.635 6.745 ;
        RECT 275.150 6.560 290.635 6.700 ;
        RECT 275.150 6.500 275.470 6.560 ;
        RECT 290.345 6.515 290.635 6.560 ;
        RECT 646.845 6.360 647.135 6.405 ;
        RECT 672.145 6.360 672.435 6.405 ;
        RECT 646.845 6.220 672.435 6.360 ;
        RECT 646.845 6.175 647.135 6.220 ;
        RECT 672.145 6.175 672.435 6.220 ;
        RECT 752.185 6.360 752.475 6.405 ;
        RECT 755.405 6.360 755.695 6.405 ;
        RECT 752.185 6.220 755.695 6.360 ;
        RECT 752.185 6.175 752.475 6.220 ;
        RECT 755.405 6.175 755.695 6.220 ;
        RECT 889.265 6.360 889.555 6.405 ;
        RECT 890.170 6.360 890.490 6.420 ;
        RECT 889.265 6.220 890.490 6.360 ;
        RECT 889.265 6.175 889.555 6.220 ;
        RECT 890.170 6.160 890.490 6.220 ;
        RECT 394.765 5.680 395.055 5.725 ;
        RECT 413.625 5.680 413.915 5.725 ;
        RECT 394.765 5.540 413.915 5.680 ;
        RECT 394.765 5.495 395.055 5.540 ;
        RECT 413.625 5.495 413.915 5.540 ;
        RECT 2068.230 5.340 2068.550 5.400 ;
        RECT 2266.490 5.340 2266.810 5.400 ;
        RECT 2068.230 5.200 2266.810 5.340 ;
        RECT 2068.230 5.140 2068.550 5.200 ;
        RECT 2266.490 5.140 2266.810 5.200 ;
        RECT 609.585 5.000 609.875 5.045 ;
        RECT 611.885 5.000 612.175 5.045 ;
        RECT 609.585 4.860 612.175 5.000 ;
        RECT 609.585 4.815 609.875 4.860 ;
        RECT 611.885 4.815 612.175 4.860 ;
        RECT 621.545 5.000 621.835 5.045 ;
        RECT 627.525 5.000 627.815 5.045 ;
        RECT 621.545 4.860 627.815 5.000 ;
        RECT 621.545 4.815 621.835 4.860 ;
        RECT 627.525 4.815 627.815 4.860 ;
        RECT 613.265 4.660 613.555 4.705 ;
        RECT 617.390 4.660 617.710 4.720 ;
        RECT 613.265 4.520 617.710 4.660 ;
        RECT 613.265 4.475 613.555 4.520 ;
        RECT 617.390 4.460 617.710 4.520 ;
        RECT 776.105 4.660 776.395 4.705 ;
        RECT 1588.450 4.660 1588.770 4.720 ;
        RECT 1616.985 4.660 1617.275 4.705 ;
        RECT 776.105 4.520 785.520 4.660 ;
        RECT 776.105 4.475 776.395 4.520 ;
        RECT 574.165 4.320 574.455 4.365 ;
        RECT 574.165 4.180 606.580 4.320 ;
        RECT 574.165 4.135 574.455 4.180 ;
        RECT 606.440 4.025 606.580 4.180 ;
        RECT 383.265 3.980 383.555 4.025 ;
        RECT 394.765 3.980 395.055 4.025 ;
        RECT 383.265 3.840 395.055 3.980 ;
        RECT 383.265 3.795 383.555 3.840 ;
        RECT 394.765 3.795 395.055 3.840 ;
        RECT 555.765 3.980 556.055 4.025 ;
        RECT 558.525 3.980 558.815 4.025 ;
        RECT 555.765 3.840 558.815 3.980 ;
        RECT 555.765 3.795 556.055 3.840 ;
        RECT 558.525 3.795 558.815 3.840 ;
        RECT 606.365 3.795 606.655 4.025 ;
        RECT 785.380 3.980 785.520 4.520 ;
        RECT 1588.450 4.520 1617.275 4.660 ;
        RECT 1588.450 4.460 1588.770 4.520 ;
        RECT 1616.985 4.475 1617.275 4.520 ;
        RECT 788.985 3.980 789.275 4.025 ;
        RECT 785.380 3.840 789.275 3.980 ;
        RECT 788.985 3.795 789.275 3.840 ;
        RECT 1164.790 3.980 1165.110 4.040 ;
        RECT 1164.790 3.840 1166.860 3.980 ;
        RECT 1164.790 3.780 1165.110 3.840 ;
        RECT 800.025 3.640 800.315 3.685 ;
        RECT 803.245 3.640 803.535 3.685 ;
        RECT 800.025 3.500 803.535 3.640 ;
        RECT 800.025 3.455 800.315 3.500 ;
        RECT 803.245 3.455 803.535 3.500 ;
        RECT 920.070 3.640 920.390 3.700 ;
        RECT 1021.285 3.640 1021.575 3.685 ;
        RECT 920.070 3.500 1021.575 3.640 ;
        RECT 920.070 3.440 920.390 3.500 ;
        RECT 1021.285 3.455 1021.575 3.500 ;
        RECT 1022.665 3.640 1022.955 3.685 ;
        RECT 1040.605 3.640 1040.895 3.685 ;
        RECT 1022.665 3.500 1040.895 3.640 ;
        RECT 1022.665 3.455 1022.955 3.500 ;
        RECT 1040.605 3.455 1040.895 3.500 ;
        RECT 1043.825 3.640 1044.115 3.685 ;
        RECT 1069.585 3.640 1069.875 3.685 ;
        RECT 1043.825 3.500 1069.875 3.640 ;
        RECT 1043.825 3.455 1044.115 3.500 ;
        RECT 1069.585 3.455 1069.875 3.500 ;
        RECT 1071.425 3.640 1071.715 3.685 ;
        RECT 1106.830 3.640 1107.150 3.700 ;
        RECT 1071.425 3.500 1107.150 3.640 ;
        RECT 1166.720 3.640 1166.860 3.840 ;
        RECT 1306.485 3.640 1306.775 3.685 ;
        RECT 1166.720 3.500 1306.775 3.640 ;
        RECT 1071.425 3.455 1071.715 3.500 ;
        RECT 1106.830 3.440 1107.150 3.500 ;
        RECT 1306.485 3.455 1306.775 3.500 ;
        RECT 1451.830 3.640 1452.150 3.700 ;
        RECT 1475.750 3.640 1476.070 3.700 ;
        RECT 1451.830 3.500 1476.070 3.640 ;
        RECT 1451.830 3.440 1452.150 3.500 ;
        RECT 1475.750 3.440 1476.070 3.500 ;
        RECT 378.190 3.300 378.510 3.360 ;
        RECT 379.125 3.300 379.415 3.345 ;
        RECT 378.190 3.160 379.415 3.300 ;
        RECT 378.190 3.100 378.510 3.160 ;
        RECT 379.125 3.115 379.415 3.160 ;
        RECT 607.745 3.300 608.035 3.345 ;
        RECT 610.505 3.300 610.795 3.345 ;
        RECT 607.745 3.160 610.795 3.300 ;
        RECT 607.745 3.115 608.035 3.160 ;
        RECT 610.505 3.115 610.795 3.160 ;
        RECT 1616.985 2.620 1617.275 2.665 ;
        RECT 1639.510 2.620 1639.830 2.680 ;
        RECT 1616.985 2.480 1639.830 2.620 ;
        RECT 1616.985 2.435 1617.275 2.480 ;
        RECT 1639.510 2.420 1639.830 2.480 ;
        RECT 918.705 0.920 918.995 0.965 ;
        RECT 919.610 0.920 919.930 0.980 ;
        RECT 918.705 0.780 919.930 0.920 ;
        RECT 918.705 0.735 918.995 0.780 ;
        RECT 919.610 0.720 919.930 0.780 ;
      LAYER via ;
        RECT 1822.620 3416.020 1822.880 3416.280 ;
        RECT 1876.900 3416.020 1877.160 3416.280 ;
        RECT 1876.900 3401.400 1877.160 3401.660 ;
        RECT 2808.860 3401.400 2809.120 3401.660 ;
        RECT 743.000 8.540 743.260 8.800 ;
        RECT 693.780 8.200 694.040 8.460 ;
        RECT 794.060 7.860 794.320 8.120 ;
        RECT 847.880 8.200 848.140 8.460 ;
        RECT 296.340 7.520 296.600 7.780 ;
        RECT 508.400 7.520 508.660 7.780 ;
        RECT 511.160 7.520 511.420 7.780 ;
        RECT 919.640 7.860 919.900 8.120 ;
        RECT 1182.760 8.540 1183.020 8.800 ;
        RECT 849.260 7.520 849.520 7.780 ;
        RECT 556.240 7.180 556.500 7.440 ;
        RECT 605.000 6.840 605.260 7.100 ;
        RECT 674.000 6.840 674.260 7.100 ;
        RECT 679.060 6.840 679.320 7.100 ;
        RECT 693.780 6.840 694.040 7.100 ;
        RECT 695.620 6.840 695.880 7.100 ;
        RECT 951.840 7.180 952.100 7.440 ;
        RECT 1410.460 7.180 1410.720 7.440 ;
        RECT 275.180 6.500 275.440 6.760 ;
        RECT 890.200 6.160 890.460 6.420 ;
        RECT 2068.260 5.140 2068.520 5.400 ;
        RECT 2266.520 5.140 2266.780 5.400 ;
        RECT 617.420 4.460 617.680 4.720 ;
        RECT 1588.480 4.460 1588.740 4.720 ;
        RECT 1164.820 3.780 1165.080 4.040 ;
        RECT 920.100 3.440 920.360 3.700 ;
        RECT 1106.860 3.440 1107.120 3.700 ;
        RECT 1451.860 3.440 1452.120 3.700 ;
        RECT 1475.780 3.440 1476.040 3.700 ;
        RECT 378.220 3.100 378.480 3.360 ;
        RECT 1639.540 2.420 1639.800 2.680 ;
        RECT 919.640 0.720 919.900 0.980 ;
      LAYER met2 ;
        RECT 1822.620 3415.990 1822.880 3416.310 ;
        RECT 1876.900 3415.990 1877.160 3416.310 ;
        RECT 1822.680 3405.000 1822.820 3415.990 ;
        RECT 1822.550 3401.000 1822.830 3405.000 ;
        RECT 1876.960 3401.690 1877.100 3415.990 ;
        RECT 2808.850 3402.195 2809.130 3402.565 ;
        RECT 2808.920 3401.690 2809.060 3402.195 ;
        RECT 1876.900 3401.370 1877.160 3401.690 ;
        RECT 2808.860 3401.370 2809.120 3401.690 ;
        RECT 296.330 8.315 296.610 8.685 ;
        RECT 324.390 8.570 324.670 8.685 ;
        RECT 681.350 8.570 681.630 8.685 ;
        RECT 697.060 8.600 703.640 8.740 ;
        RECT 697.060 8.570 697.200 8.600 ;
        RECT 324.390 8.430 326.440 8.570 ;
        RECT 324.390 8.315 324.670 8.430 ;
        RECT 296.400 7.810 296.540 8.315 ;
        RECT 326.300 7.890 326.440 8.430 ;
        RECT 462.920 8.430 484.680 8.570 ;
        RECT 462.920 8.005 463.060 8.430 ;
        RECT 326.690 7.890 326.970 8.005 ;
        RECT 296.340 7.490 296.600 7.810 ;
        RECT 326.300 7.750 326.970 7.890 ;
        RECT 326.690 7.635 326.970 7.750 ;
        RECT 462.850 7.635 463.130 8.005 ;
        RECT 484.540 7.890 484.680 8.430 ;
        RECT 681.350 8.430 685.240 8.570 ;
        RECT 681.350 8.315 681.630 8.430 ;
        RECT 484.930 7.890 485.210 8.005 ;
        RECT 484.540 7.750 485.210 7.890 ;
        RECT 484.930 7.635 485.210 7.750 ;
        RECT 508.390 7.635 508.670 8.005 ;
        RECT 511.680 7.920 515.960 8.060 ;
        RECT 511.160 7.720 511.420 7.810 ;
        RECT 511.680 7.720 511.820 7.920 ;
        RECT 508.400 7.490 508.660 7.635 ;
        RECT 511.160 7.580 511.820 7.720 ;
        RECT 511.160 7.490 511.420 7.580 ;
        RECT 275.180 6.700 275.440 6.790 ;
        RECT 270.180 6.560 275.440 6.700 ;
        RECT 270.180 2.400 270.320 6.560 ;
        RECT 275.180 6.470 275.440 6.560 ;
        RECT 515.820 5.850 515.960 7.920 ;
        RECT 517.130 7.635 517.410 8.005 ;
        RECT 517.200 5.850 517.340 7.635 ;
        RECT 556.240 7.325 556.500 7.470 ;
        RECT 556.230 6.955 556.510 7.325 ;
        RECT 605.000 6.810 605.260 7.130 ;
        RECT 645.010 6.955 645.290 7.325 ;
        RECT 673.990 6.955 674.270 7.325 ;
        RECT 515.820 5.710 517.340 5.850 ;
        RECT 378.220 3.130 378.480 3.390 ;
        RECT 605.060 3.300 605.200 6.810 ;
        RECT 617.420 4.430 617.680 4.750 ;
        RECT 604.600 3.245 605.200 3.300 ;
        RECT 377.360 3.070 378.480 3.130 ;
        RECT 377.360 2.990 378.420 3.070 ;
        RECT 377.360 2.400 377.500 2.990 ;
        RECT 579.690 2.875 579.970 3.245 ;
        RECT 604.530 3.160 605.200 3.245 ;
        RECT 604.530 2.875 604.810 3.160 ;
        RECT 579.760 2.400 579.900 2.875 ;
        RECT 269.970 -4.800 270.530 2.400 ;
        RECT 377.150 -4.800 377.710 2.400 ;
        RECT 579.550 -4.800 580.110 2.400 ;
        RECT 617.480 1.090 617.620 4.430 ;
        RECT 645.080 4.320 645.220 6.955 ;
        RECT 674.000 6.810 674.260 6.955 ;
        RECT 679.060 6.810 679.320 7.130 ;
        RECT 679.120 6.020 679.260 6.810 ;
        RECT 685.100 6.020 685.240 8.430 ;
        RECT 693.780 8.170 694.040 8.490 ;
        RECT 696.600 8.430 697.200 8.570 ;
        RECT 693.840 7.130 693.980 8.170 ;
        RECT 693.780 6.810 694.040 7.130 ;
        RECT 695.620 6.810 695.880 7.130 ;
        RECT 695.680 6.530 695.820 6.810 ;
        RECT 696.600 6.530 696.740 8.430 ;
        RECT 703.500 7.380 703.640 8.600 ;
        RECT 743.000 8.510 743.260 8.830 ;
        RECT 704.810 7.890 705.090 8.005 ;
        RECT 704.420 7.750 705.090 7.890 ;
        RECT 704.420 7.380 704.560 7.750 ;
        RECT 704.810 7.635 705.090 7.750 ;
        RECT 703.500 7.240 704.560 7.380 ;
        RECT 695.680 6.390 696.740 6.530 ;
        RECT 679.120 5.880 685.240 6.020 ;
        RECT 743.060 5.965 743.200 8.510 ;
        RECT 794.050 8.315 794.330 8.685 ;
        RECT 794.120 8.150 794.260 8.315 ;
        RECT 847.880 8.170 848.140 8.490 ;
        RECT 921.540 8.260 923.980 8.400 ;
        RECT 794.060 7.830 794.320 8.150 ;
        RECT 847.940 7.720 848.080 8.170 ;
        RECT 919.640 7.830 919.900 8.150 ;
        RECT 849.260 7.720 849.520 7.810 ;
        RECT 847.940 7.580 849.520 7.720 ;
        RECT 849.260 7.490 849.520 7.580 ;
        RECT 919.700 7.380 919.840 7.830 ;
        RECT 921.540 7.380 921.680 8.260 ;
        RECT 919.700 7.240 921.680 7.380 ;
        RECT 890.190 6.275 890.470 6.645 ;
        RECT 913.190 6.530 913.470 6.645 ;
        RECT 913.190 6.390 920.300 6.530 ;
        RECT 913.190 6.275 913.470 6.390 ;
        RECT 890.200 6.130 890.460 6.275 ;
        RECT 742.990 5.595 743.270 5.965 ;
        RECT 920.160 5.850 920.300 6.390 ;
        RECT 923.840 6.360 923.980 8.260 ;
        RECT 931.070 6.360 931.350 9.000 ;
        RECT 1182.760 8.740 1183.020 8.830 ;
        RECT 1182.760 8.600 1191.240 8.740 ;
        RECT 1182.760 8.510 1183.020 8.600 ;
        RECT 951.840 7.150 952.100 7.470 ;
        RECT 1191.100 7.210 1191.240 8.600 ;
        RECT 1193.330 7.210 1193.610 7.325 ;
        RECT 923.840 6.220 931.800 6.360 ;
        RECT 921.010 5.850 921.290 5.965 ;
        RECT 920.160 5.710 921.290 5.850 ;
        RECT 921.010 5.595 921.290 5.710 ;
        RECT 929.290 5.850 929.570 5.965 ;
        RECT 931.070 5.850 931.350 6.220 ;
        RECT 929.290 5.710 931.350 5.850 ;
        RECT 931.660 5.850 931.800 6.220 ;
        RECT 951.900 5.965 952.040 7.150 ;
        RECT 1191.100 7.070 1193.610 7.210 ;
        RECT 1193.330 6.955 1193.610 7.070 ;
        RECT 1214.490 7.210 1214.770 7.325 ;
        RECT 1215.810 7.210 1216.090 9.000 ;
        RECT 1214.490 7.070 1216.090 7.210 ;
        RECT 1410.460 7.150 1410.720 7.470 ;
        RECT 1214.490 6.955 1214.770 7.070 ;
        RECT 932.510 5.850 932.790 5.965 ;
        RECT 931.660 5.710 932.790 5.850 ;
        RECT 929.290 5.595 929.570 5.710 ;
        RECT 931.070 5.000 931.350 5.710 ;
        RECT 932.510 5.595 932.790 5.710 ;
        RECT 951.830 5.595 952.110 5.965 ;
        RECT 1215.810 5.000 1216.090 7.070 ;
        RECT 1410.520 6.530 1410.660 7.150 ;
        RECT 1410.520 6.390 1427.220 6.530 ;
        RECT 644.620 4.180 645.220 4.320 ;
        RECT 644.620 3.810 644.760 4.180 ;
        RECT 620.240 3.670 644.760 3.810 ;
        RECT 1164.820 3.750 1165.080 4.070 ;
        RECT 1427.080 3.810 1427.220 6.390 ;
        RECT 1475.770 6.275 1476.050 6.645 ;
        RECT 1588.470 6.275 1588.750 6.645 ;
        RECT 1639.530 6.275 1639.810 6.645 ;
        RECT 1823.530 6.275 1823.810 6.645 ;
        RECT 1866.770 6.275 1867.050 6.645 ;
        RECT 2033.290 6.275 2033.570 6.645 ;
        RECT 2266.510 6.275 2266.790 6.645 ;
        RECT 2302.850 6.275 2303.130 6.645 ;
        RECT 2382.890 6.275 2383.170 6.645 ;
        RECT 2410.950 6.275 2411.230 6.645 ;
        RECT 2520.890 6.275 2521.170 6.645 ;
        RECT 2583.450 6.275 2583.730 6.645 ;
        RECT 2797.810 6.275 2798.090 6.645 ;
        RECT 1428.850 3.810 1429.130 3.925 ;
        RECT 620.240 1.090 620.380 3.670 ;
        RECT 920.100 3.640 920.360 3.730 ;
        RECT 617.480 0.950 620.380 1.090 ;
        RECT 919.700 3.500 920.360 3.640 ;
        RECT 919.700 1.010 919.840 3.500 ;
        RECT 920.100 3.410 920.360 3.500 ;
        RECT 1106.860 3.410 1107.120 3.730 ;
        RECT 1106.920 3.245 1107.060 3.410 ;
        RECT 1164.880 3.245 1165.020 3.750 ;
        RECT 1427.080 3.670 1429.130 3.810 ;
        RECT 1428.850 3.555 1429.130 3.670 ;
        RECT 1451.850 3.555 1452.130 3.925 ;
        RECT 1475.840 3.730 1475.980 6.275 ;
        RECT 1588.540 4.750 1588.680 6.275 ;
        RECT 1588.480 4.430 1588.740 4.750 ;
        RECT 1451.860 3.410 1452.120 3.555 ;
        RECT 1475.780 3.410 1476.040 3.730 ;
        RECT 1106.850 2.875 1107.130 3.245 ;
        RECT 1164.810 2.875 1165.090 3.245 ;
        RECT 1639.600 2.710 1639.740 6.275 ;
        RECT 1823.600 3.925 1823.740 6.275 ;
        RECT 1866.840 3.925 1866.980 6.275 ;
        RECT 1823.530 3.555 1823.810 3.925 ;
        RECT 1866.770 3.555 1867.050 3.925 ;
        RECT 1639.540 2.390 1639.800 2.710 ;
        RECT 2033.360 1.885 2033.500 6.275 ;
        RECT 2266.580 5.430 2266.720 6.275 ;
        RECT 2068.260 5.110 2068.520 5.430 ;
        RECT 2266.520 5.110 2266.780 5.430 ;
        RECT 2068.320 1.885 2068.460 5.110 ;
        RECT 2302.920 3.925 2303.060 6.275 ;
        RECT 2382.960 3.925 2383.100 6.275 ;
        RECT 2411.020 3.925 2411.160 6.275 ;
        RECT 2520.960 3.925 2521.100 6.275 ;
        RECT 2583.520 3.925 2583.660 6.275 ;
        RECT 2658.890 5.595 2659.170 5.965 ;
        RECT 2658.960 3.925 2659.100 5.595 ;
        RECT 2797.880 3.925 2798.020 6.275 ;
        RECT 2302.850 3.555 2303.130 3.925 ;
        RECT 2382.890 3.555 2383.170 3.925 ;
        RECT 2410.950 3.555 2411.230 3.925 ;
        RECT 2520.890 3.555 2521.170 3.925 ;
        RECT 2583.450 3.555 2583.730 3.925 ;
        RECT 2658.890 3.555 2659.170 3.925 ;
        RECT 2797.810 3.555 2798.090 3.925 ;
        RECT 2033.290 1.515 2033.570 1.885 ;
        RECT 2068.250 1.515 2068.530 1.885 ;
        RECT 919.640 0.690 919.900 1.010 ;
      LAYER via2 ;
        RECT 2808.850 3402.240 2809.130 3402.520 ;
        RECT 296.330 8.360 296.610 8.640 ;
        RECT 324.390 8.360 324.670 8.640 ;
        RECT 326.690 7.680 326.970 7.960 ;
        RECT 462.850 7.680 463.130 7.960 ;
        RECT 681.350 8.360 681.630 8.640 ;
        RECT 484.930 7.680 485.210 7.960 ;
        RECT 508.390 7.680 508.670 7.960 ;
        RECT 517.130 7.680 517.410 7.960 ;
        RECT 556.230 7.000 556.510 7.280 ;
        RECT 645.010 7.000 645.290 7.280 ;
        RECT 673.990 7.000 674.270 7.280 ;
        RECT 579.690 2.920 579.970 3.200 ;
        RECT 604.530 2.920 604.810 3.200 ;
        RECT 704.810 7.680 705.090 7.960 ;
        RECT 794.050 8.360 794.330 8.640 ;
        RECT 890.190 6.320 890.470 6.600 ;
        RECT 913.190 6.320 913.470 6.600 ;
        RECT 742.990 5.640 743.270 5.920 ;
        RECT 921.010 5.640 921.290 5.920 ;
        RECT 929.290 5.640 929.570 5.920 ;
        RECT 1193.330 7.000 1193.610 7.280 ;
        RECT 1214.490 7.000 1214.770 7.280 ;
        RECT 932.510 5.640 932.790 5.920 ;
        RECT 951.830 5.640 952.110 5.920 ;
        RECT 1475.770 6.320 1476.050 6.600 ;
        RECT 1588.470 6.320 1588.750 6.600 ;
        RECT 1639.530 6.320 1639.810 6.600 ;
        RECT 1823.530 6.320 1823.810 6.600 ;
        RECT 1866.770 6.320 1867.050 6.600 ;
        RECT 2033.290 6.320 2033.570 6.600 ;
        RECT 2266.510 6.320 2266.790 6.600 ;
        RECT 2302.850 6.320 2303.130 6.600 ;
        RECT 2382.890 6.320 2383.170 6.600 ;
        RECT 2410.950 6.320 2411.230 6.600 ;
        RECT 2520.890 6.320 2521.170 6.600 ;
        RECT 2583.450 6.320 2583.730 6.600 ;
        RECT 2797.810 6.320 2798.090 6.600 ;
        RECT 1428.850 3.600 1429.130 3.880 ;
        RECT 1451.850 3.600 1452.130 3.880 ;
        RECT 1106.850 2.920 1107.130 3.200 ;
        RECT 1164.810 2.920 1165.090 3.200 ;
        RECT 1823.530 3.600 1823.810 3.880 ;
        RECT 1866.770 3.600 1867.050 3.880 ;
        RECT 2658.890 5.640 2659.170 5.920 ;
        RECT 2302.850 3.600 2303.130 3.880 ;
        RECT 2382.890 3.600 2383.170 3.880 ;
        RECT 2410.950 3.600 2411.230 3.880 ;
        RECT 2520.890 3.600 2521.170 3.880 ;
        RECT 2583.450 3.600 2583.730 3.880 ;
        RECT 2658.890 3.600 2659.170 3.880 ;
        RECT 2797.810 3.600 2798.090 3.880 ;
        RECT 2033.290 1.560 2033.570 1.840 ;
        RECT 2068.250 1.560 2068.530 1.840 ;
      LAYER met3 ;
        RECT 2808.825 3402.530 2809.155 3402.545 ;
        RECT 2815.470 3402.530 2815.850 3402.540 ;
        RECT 2808.825 3402.230 2815.850 3402.530 ;
        RECT 2808.825 3402.215 2809.155 3402.230 ;
        RECT 2815.470 3402.220 2815.850 3402.230 ;
        RECT 296.305 8.650 296.635 8.665 ;
        RECT 324.365 8.650 324.695 8.665 ;
        RECT 296.305 8.350 324.695 8.650 ;
        RECT 296.305 8.335 296.635 8.350 ;
        RECT 324.365 8.335 324.695 8.350 ;
        RECT 440.950 8.650 441.330 8.660 ;
        RECT 680.380 8.650 680.760 8.660 ;
        RECT 681.325 8.650 681.655 8.665 ;
        RECT 440.950 8.350 457.620 8.650 ;
        RECT 440.950 8.340 441.330 8.350 ;
        RECT 326.665 7.970 326.995 7.985 ;
        RECT 333.310 7.970 333.690 7.980 ;
        RECT 326.665 7.670 333.690 7.970 ;
        RECT 457.320 7.970 457.620 8.350 ;
        RECT 680.380 8.350 681.655 8.650 ;
        RECT 680.380 8.340 680.760 8.350 ;
        RECT 681.325 8.335 681.655 8.350 ;
        RECT 792.390 8.650 792.770 8.660 ;
        RECT 794.025 8.650 794.355 8.665 ;
        RECT 792.390 8.350 794.355 8.650 ;
        RECT 792.390 8.340 792.770 8.350 ;
        RECT 794.025 8.335 794.355 8.350 ;
        RECT 462.825 7.970 463.155 7.985 ;
        RECT 457.320 7.670 463.155 7.970 ;
        RECT 326.665 7.655 326.995 7.670 ;
        RECT 333.310 7.660 333.690 7.670 ;
        RECT 462.825 7.655 463.155 7.670 ;
        RECT 484.905 7.970 485.235 7.985 ;
        RECT 508.365 7.970 508.695 7.985 ;
        RECT 484.905 7.670 508.695 7.970 ;
        RECT 484.905 7.655 485.235 7.670 ;
        RECT 508.365 7.655 508.695 7.670 ;
        RECT 517.105 7.970 517.435 7.985 ;
        RECT 704.785 7.970 705.115 7.985 ;
        RECT 517.105 7.670 555.600 7.970 ;
        RECT 517.105 7.655 517.435 7.670 ;
        RECT 555.300 7.290 555.600 7.670 ;
        RECT 704.785 7.670 707.170 7.970 ;
        RECT 704.785 7.655 705.115 7.670 ;
        RECT 556.205 7.290 556.535 7.305 ;
        RECT 555.300 6.990 556.535 7.290 ;
        RECT 556.205 6.975 556.535 6.990 ;
        RECT 644.985 7.290 645.315 7.305 ;
        RECT 673.965 7.290 674.295 7.305 ;
        RECT 644.985 6.990 674.295 7.290 ;
        RECT 644.985 6.975 645.315 6.990 ;
        RECT 673.965 6.975 674.295 6.990 ;
        RECT 706.870 6.610 707.170 7.670 ;
        RECT 1193.305 7.290 1193.635 7.305 ;
        RECT 1214.465 7.290 1214.795 7.305 ;
        RECT 1193.305 6.990 1214.795 7.290 ;
        RECT 1193.305 6.975 1193.635 6.990 ;
        RECT 1214.465 6.975 1214.795 6.990 ;
        RECT 890.165 6.610 890.495 6.625 ;
        RECT 897.270 6.610 897.650 6.620 ;
        RECT 706.870 6.310 738.450 6.610 ;
        RECT 738.150 5.930 738.450 6.310 ;
        RECT 890.165 6.310 897.650 6.610 ;
        RECT 890.165 6.295 890.495 6.310 ;
        RECT 897.270 6.300 897.650 6.310 ;
        RECT 901.870 6.610 902.250 6.620 ;
        RECT 913.165 6.610 913.495 6.625 ;
        RECT 901.870 6.310 913.495 6.610 ;
        RECT 901.870 6.300 902.250 6.310 ;
        RECT 913.165 6.295 913.495 6.310 ;
        RECT 1475.745 6.610 1476.075 6.625 ;
        RECT 1588.445 6.610 1588.775 6.625 ;
        RECT 1475.745 6.310 1588.775 6.610 ;
        RECT 1475.745 6.295 1476.075 6.310 ;
        RECT 1588.445 6.295 1588.775 6.310 ;
        RECT 1639.505 6.610 1639.835 6.625 ;
        RECT 1823.505 6.610 1823.835 6.625 ;
        RECT 1639.505 6.310 1823.835 6.610 ;
        RECT 1639.505 6.295 1639.835 6.310 ;
        RECT 1823.505 6.295 1823.835 6.310 ;
        RECT 1866.745 6.610 1867.075 6.625 ;
        RECT 2033.265 6.610 2033.595 6.625 ;
        RECT 1866.745 6.310 2033.595 6.610 ;
        RECT 1866.745 6.295 1867.075 6.310 ;
        RECT 2033.265 6.295 2033.595 6.310 ;
        RECT 2266.485 6.610 2266.815 6.625 ;
        RECT 2302.825 6.610 2303.155 6.625 ;
        RECT 2266.485 6.310 2303.155 6.610 ;
        RECT 2266.485 6.295 2266.815 6.310 ;
        RECT 2302.825 6.295 2303.155 6.310 ;
        RECT 2382.865 6.610 2383.195 6.625 ;
        RECT 2410.925 6.610 2411.255 6.625 ;
        RECT 2382.865 6.310 2411.255 6.610 ;
        RECT 2382.865 6.295 2383.195 6.310 ;
        RECT 2410.925 6.295 2411.255 6.310 ;
        RECT 2520.865 6.610 2521.195 6.625 ;
        RECT 2583.425 6.610 2583.755 6.625 ;
        RECT 2797.785 6.610 2798.115 6.625 ;
        RECT 2520.865 6.310 2583.755 6.610 ;
        RECT 2520.865 6.295 2521.195 6.310 ;
        RECT 2583.425 6.295 2583.755 6.310 ;
        RECT 2763.070 6.310 2798.115 6.610 ;
        RECT 742.965 5.930 743.295 5.945 ;
        RECT 738.150 5.630 743.295 5.930 ;
        RECT 742.965 5.615 743.295 5.630 ;
        RECT 920.985 5.930 921.315 5.945 ;
        RECT 929.265 5.930 929.595 5.945 ;
        RECT 920.985 5.630 929.595 5.930 ;
        RECT 920.985 5.615 921.315 5.630 ;
        RECT 929.265 5.615 929.595 5.630 ;
        RECT 932.485 5.930 932.815 5.945 ;
        RECT 951.805 5.930 952.135 5.945 ;
        RECT 932.485 5.630 952.135 5.930 ;
        RECT 932.485 5.615 932.815 5.630 ;
        RECT 951.805 5.615 952.135 5.630 ;
        RECT 2658.865 5.930 2659.195 5.945 ;
        RECT 2763.070 5.930 2763.370 6.310 ;
        RECT 2797.785 6.295 2798.115 6.310 ;
        RECT 2658.865 5.630 2763.370 5.930 ;
        RECT 2658.865 5.615 2659.195 5.630 ;
        RECT 1428.825 3.890 1429.155 3.905 ;
        RECT 1451.825 3.890 1452.155 3.905 ;
        RECT 1428.825 3.590 1452.155 3.890 ;
        RECT 1428.825 3.575 1429.155 3.590 ;
        RECT 1451.825 3.575 1452.155 3.590 ;
        RECT 1823.505 3.890 1823.835 3.905 ;
        RECT 1866.745 3.890 1867.075 3.905 ;
        RECT 1823.505 3.590 1867.075 3.890 ;
        RECT 1823.505 3.575 1823.835 3.590 ;
        RECT 1866.745 3.575 1867.075 3.590 ;
        RECT 2302.825 3.890 2303.155 3.905 ;
        RECT 2382.865 3.890 2383.195 3.905 ;
        RECT 2302.825 3.590 2383.195 3.890 ;
        RECT 2302.825 3.575 2303.155 3.590 ;
        RECT 2382.865 3.575 2383.195 3.590 ;
        RECT 2410.925 3.890 2411.255 3.905 ;
        RECT 2520.865 3.890 2521.195 3.905 ;
        RECT 2410.925 3.590 2521.195 3.890 ;
        RECT 2410.925 3.575 2411.255 3.590 ;
        RECT 2520.865 3.575 2521.195 3.590 ;
        RECT 2583.425 3.890 2583.755 3.905 ;
        RECT 2658.865 3.890 2659.195 3.905 ;
        RECT 2583.425 3.590 2659.195 3.890 ;
        RECT 2583.425 3.575 2583.755 3.590 ;
        RECT 2658.865 3.575 2659.195 3.590 ;
        RECT 2797.785 3.890 2798.115 3.905 ;
        RECT 2815.470 3.890 2815.850 3.900 ;
        RECT 2797.785 3.590 2815.850 3.890 ;
        RECT 2797.785 3.575 2798.115 3.590 ;
        RECT 2815.470 3.580 2815.850 3.590 ;
        RECT 579.665 3.210 579.995 3.225 ;
        RECT 604.505 3.210 604.835 3.225 ;
        RECT 579.665 2.910 604.835 3.210 ;
        RECT 579.665 2.895 579.995 2.910 ;
        RECT 604.505 2.895 604.835 2.910 ;
        RECT 1106.825 3.210 1107.155 3.225 ;
        RECT 1164.785 3.210 1165.115 3.225 ;
        RECT 1106.825 2.910 1165.115 3.210 ;
        RECT 1106.825 2.895 1107.155 2.910 ;
        RECT 1164.785 2.895 1165.115 2.910 ;
        RECT 2033.265 1.850 2033.595 1.865 ;
        RECT 2068.225 1.850 2068.555 1.865 ;
        RECT 2033.265 1.550 2068.555 1.850 ;
        RECT 2033.265 1.535 2033.595 1.550 ;
        RECT 2068.225 1.535 2068.555 1.550 ;
      LAYER via3 ;
        RECT 2815.500 3402.220 2815.820 3402.540 ;
        RECT 440.980 8.340 441.300 8.660 ;
        RECT 333.340 7.660 333.660 7.980 ;
        RECT 680.410 8.340 680.730 8.660 ;
        RECT 792.420 8.340 792.740 8.660 ;
        RECT 897.300 6.300 897.620 6.620 ;
        RECT 901.900 6.300 902.220 6.620 ;
        RECT 2815.500 3.580 2815.820 3.900 ;
      LAYER met4 ;
        RECT 2815.495 3402.215 2815.825 3402.545 ;
        RECT 682.510 14.710 683.690 15.890 ;
        RECT 729.430 14.710 730.610 15.890 ;
        RECT 682.950 12.050 683.250 14.710 ;
        RECT 680.190 11.750 683.250 12.050 ;
        RECT 729.870 12.050 730.170 14.710 ;
        RECT 729.870 11.750 733.850 12.050 ;
        RECT 680.190 8.665 680.490 11.750 ;
        RECT 333.350 8.350 336.410 8.650 ;
        RECT 333.350 7.985 333.650 8.350 ;
        RECT 333.335 7.655 333.665 7.985 ;
        RECT 336.110 5.250 336.410 8.350 ;
        RECT 440.975 8.335 441.305 8.665 ;
        RECT 680.190 8.350 680.735 8.665 ;
        RECT 680.405 8.335 680.735 8.350 ;
        RECT 440.990 5.690 441.290 8.335 ;
        RECT 733.550 5.930 733.850 11.750 ;
        RECT 792.415 8.335 792.745 8.665 ;
        RECT 741.830 7.670 761.450 7.970 ;
        RECT 344.870 5.250 346.050 5.690 ;
        RECT 336.110 4.950 346.050 5.250 ;
        RECT 344.870 4.510 346.050 4.950 ;
        RECT 440.550 4.510 441.730 5.690 ;
        RECT 733.550 5.630 736.610 5.930 ;
        RECT 736.310 3.890 736.610 5.630 ;
        RECT 741.830 3.890 742.130 7.670 ;
        RECT 761.150 5.930 761.450 7.670 ;
        RECT 792.430 5.930 792.730 8.335 ;
        RECT 897.295 6.610 897.625 6.625 ;
        RECT 901.895 6.610 902.225 6.625 ;
        RECT 897.295 6.310 902.225 6.610 ;
        RECT 897.295 6.295 897.625 6.310 ;
        RECT 901.895 6.295 902.225 6.310 ;
        RECT 761.150 5.630 792.730 5.930 ;
        RECT 2815.510 3.905 2815.810 3402.215 ;
        RECT 736.310 3.590 742.130 3.890 ;
        RECT 2815.495 3.575 2815.825 3.905 ;
      LAYER met5 ;
        RECT 682.300 14.500 730.820 16.100 ;
        RECT 344.660 4.300 441.940 5.900 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2849.845 2090.745 2850.015 2162.655 ;
        RECT 2849.845 1968.855 2850.015 1997.755 ;
        RECT 2849.385 1968.685 2850.015 1968.855 ;
        RECT 2849.385 1913.265 2849.555 1968.685 ;
        RECT 2850.305 1882.665 2850.475 1909.355 ;
        RECT 2850.765 1738.505 2850.935 1848.835 ;
        RECT 2849.385 1521.245 2850.015 1521.415 ;
        RECT 2849.385 1463.955 2849.555 1521.245 ;
        RECT 2849.385 1463.785 2850.015 1463.955 ;
        RECT 2849.845 1426.895 2850.015 1427.575 ;
        RECT 2849.385 1426.725 2850.015 1426.895 ;
        RECT 2849.385 1370.115 2849.555 1426.725 ;
        RECT 2849.385 1369.945 2850.015 1370.115 ;
        RECT 2850.305 1348.865 2850.475 1369.435 ;
        RECT 2849.845 1299.225 2850.015 1336.455 ;
        RECT 2850.305 1027.225 2850.475 1134.495 ;
        RECT 2851.225 1022.125 2851.395 1027.395 ;
        RECT 2852.145 957.525 2852.315 963.815 ;
        RECT 2849.385 886.465 2850.015 886.635 ;
        RECT 2849.385 817.615 2849.555 886.465 ;
        RECT 2849.385 817.445 2850.015 817.615 ;
        RECT 2849.845 746.385 2850.015 789.395 ;
        RECT 2851.685 665.465 2851.855 742.475 ;
        RECT 2852.605 282.965 2852.775 330.055 ;
        RECT 2852.605 195.245 2852.775 216.495 ;
      LAYER mcon ;
        RECT 2849.845 2162.485 2850.015 2162.655 ;
        RECT 2849.845 1997.585 2850.015 1997.755 ;
        RECT 2850.305 1909.185 2850.475 1909.355 ;
        RECT 2850.765 1848.665 2850.935 1848.835 ;
        RECT 2849.845 1521.245 2850.015 1521.415 ;
        RECT 2849.845 1463.785 2850.015 1463.955 ;
        RECT 2849.845 1427.405 2850.015 1427.575 ;
        RECT 2849.845 1369.945 2850.015 1370.115 ;
        RECT 2850.305 1369.265 2850.475 1369.435 ;
        RECT 2849.845 1336.285 2850.015 1336.455 ;
        RECT 2850.305 1134.325 2850.475 1134.495 ;
        RECT 2851.225 1027.225 2851.395 1027.395 ;
        RECT 2852.145 963.645 2852.315 963.815 ;
        RECT 2849.845 886.465 2850.015 886.635 ;
        RECT 2849.845 817.445 2850.015 817.615 ;
        RECT 2849.845 789.225 2850.015 789.395 ;
        RECT 2851.685 742.305 2851.855 742.475 ;
        RECT 2852.605 329.885 2852.775 330.055 ;
        RECT 2852.605 216.325 2852.775 216.495 ;
      LAYER met1 ;
        RECT 2849.770 2162.640 2850.090 2162.700 ;
        RECT 2849.575 2162.500 2850.090 2162.640 ;
        RECT 2849.770 2162.440 2850.090 2162.500 ;
        RECT 2849.770 2090.900 2850.090 2090.960 ;
        RECT 2849.575 2090.760 2850.090 2090.900 ;
        RECT 2849.770 2090.700 2850.090 2090.760 ;
        RECT 2849.770 2035.480 2850.090 2035.540 ;
        RECT 2850.230 2035.480 2850.550 2035.540 ;
        RECT 2849.770 2035.340 2850.550 2035.480 ;
        RECT 2849.770 2035.280 2850.090 2035.340 ;
        RECT 2850.230 2035.280 2850.550 2035.340 ;
        RECT 2849.785 1997.740 2850.075 1997.785 ;
        RECT 2850.230 1997.740 2850.550 1997.800 ;
        RECT 2849.785 1997.600 2850.550 1997.740 ;
        RECT 2849.785 1997.555 2850.075 1997.600 ;
        RECT 2850.230 1997.540 2850.550 1997.600 ;
        RECT 2849.325 1913.420 2849.615 1913.465 ;
        RECT 2849.770 1913.420 2850.090 1913.480 ;
        RECT 2849.325 1913.280 2850.090 1913.420 ;
        RECT 2849.325 1913.235 2849.615 1913.280 ;
        RECT 2849.770 1913.220 2850.090 1913.280 ;
        RECT 2849.770 1909.340 2850.090 1909.400 ;
        RECT 2850.245 1909.340 2850.535 1909.385 ;
        RECT 2849.770 1909.200 2850.535 1909.340 ;
        RECT 2849.770 1909.140 2850.090 1909.200 ;
        RECT 2850.245 1909.155 2850.535 1909.200 ;
        RECT 2849.770 1882.820 2850.090 1882.880 ;
        RECT 2850.245 1882.820 2850.535 1882.865 ;
        RECT 2849.770 1882.680 2850.535 1882.820 ;
        RECT 2849.770 1882.620 2850.090 1882.680 ;
        RECT 2850.245 1882.635 2850.535 1882.680 ;
        RECT 2849.770 1848.820 2850.090 1848.880 ;
        RECT 2850.705 1848.820 2850.995 1848.865 ;
        RECT 2849.770 1848.680 2850.995 1848.820 ;
        RECT 2849.770 1848.620 2850.090 1848.680 ;
        RECT 2850.705 1848.635 2850.995 1848.680 ;
        RECT 2849.770 1738.660 2850.090 1738.720 ;
        RECT 2850.705 1738.660 2850.995 1738.705 ;
        RECT 2849.770 1738.520 2850.995 1738.660 ;
        RECT 2849.770 1738.460 2850.090 1738.520 ;
        RECT 2850.705 1738.475 2850.995 1738.520 ;
        RECT 2851.150 1577.980 2851.470 1578.240 ;
        RECT 2850.230 1577.840 2850.550 1577.900 ;
        RECT 2851.240 1577.840 2851.380 1577.980 ;
        RECT 2850.230 1577.700 2851.380 1577.840 ;
        RECT 2850.230 1577.640 2850.550 1577.700 ;
        RECT 2849.785 1521.400 2850.075 1521.445 ;
        RECT 2850.230 1521.400 2850.550 1521.460 ;
        RECT 2849.785 1521.260 2850.550 1521.400 ;
        RECT 2849.785 1521.215 2850.075 1521.260 ;
        RECT 2850.230 1521.200 2850.550 1521.260 ;
        RECT 2849.785 1463.940 2850.075 1463.985 ;
        RECT 2851.150 1463.940 2851.470 1464.000 ;
        RECT 2849.785 1463.800 2851.470 1463.940 ;
        RECT 2849.785 1463.755 2850.075 1463.800 ;
        RECT 2851.150 1463.740 2851.470 1463.800 ;
        RECT 2849.785 1427.560 2850.075 1427.605 ;
        RECT 2851.150 1427.560 2851.470 1427.620 ;
        RECT 2849.785 1427.420 2851.470 1427.560 ;
        RECT 2849.785 1427.375 2850.075 1427.420 ;
        RECT 2851.150 1427.360 2851.470 1427.420 ;
        RECT 2849.785 1370.100 2850.075 1370.145 ;
        RECT 2849.785 1369.960 2850.460 1370.100 ;
        RECT 2849.785 1369.915 2850.075 1369.960 ;
        RECT 2850.320 1369.465 2850.460 1369.960 ;
        RECT 2850.245 1369.235 2850.535 1369.465 ;
        RECT 2849.770 1349.020 2850.090 1349.080 ;
        RECT 2850.245 1349.020 2850.535 1349.065 ;
        RECT 2849.770 1348.880 2850.535 1349.020 ;
        RECT 2849.770 1348.820 2850.090 1348.880 ;
        RECT 2850.245 1348.835 2850.535 1348.880 ;
        RECT 2849.770 1336.440 2850.090 1336.500 ;
        RECT 2849.575 1336.300 2850.090 1336.440 ;
        RECT 2849.770 1336.240 2850.090 1336.300 ;
        RECT 2849.770 1299.380 2850.090 1299.440 ;
        RECT 2849.575 1299.240 2850.090 1299.380 ;
        RECT 2849.770 1299.180 2850.090 1299.240 ;
        RECT 2849.770 1282.720 2850.090 1282.780 ;
        RECT 2851.150 1282.720 2851.470 1282.780 ;
        RECT 2849.770 1282.580 2851.470 1282.720 ;
        RECT 2849.770 1282.520 2850.090 1282.580 ;
        RECT 2851.150 1282.520 2851.470 1282.580 ;
        RECT 2850.245 1134.480 2850.535 1134.525 ;
        RECT 2851.150 1134.480 2851.470 1134.540 ;
        RECT 2850.245 1134.340 2851.470 1134.480 ;
        RECT 2850.245 1134.295 2850.535 1134.340 ;
        RECT 2851.150 1134.280 2851.470 1134.340 ;
        RECT 2850.245 1027.380 2850.535 1027.425 ;
        RECT 2851.165 1027.380 2851.455 1027.425 ;
        RECT 2850.245 1027.240 2851.455 1027.380 ;
        RECT 2850.245 1027.195 2850.535 1027.240 ;
        RECT 2851.165 1027.195 2851.455 1027.240 ;
        RECT 2850.230 1022.280 2850.550 1022.340 ;
        RECT 2851.165 1022.280 2851.455 1022.325 ;
        RECT 2850.230 1022.140 2851.455 1022.280 ;
        RECT 2850.230 1022.080 2850.550 1022.140 ;
        RECT 2851.165 1022.095 2851.455 1022.140 ;
        RECT 2849.770 963.800 2850.090 963.860 ;
        RECT 2852.085 963.800 2852.375 963.845 ;
        RECT 2849.770 963.660 2852.375 963.800 ;
        RECT 2849.770 963.600 2850.090 963.660 ;
        RECT 2852.085 963.615 2852.375 963.660 ;
        RECT 2850.690 957.680 2851.010 957.740 ;
        RECT 2852.085 957.680 2852.375 957.725 ;
        RECT 2850.690 957.540 2852.375 957.680 ;
        RECT 2850.690 957.480 2851.010 957.540 ;
        RECT 2852.085 957.495 2852.375 957.540 ;
        RECT 2849.785 886.620 2850.075 886.665 ;
        RECT 2850.690 886.620 2851.010 886.680 ;
        RECT 2849.785 886.480 2851.010 886.620 ;
        RECT 2849.785 886.435 2850.075 886.480 ;
        RECT 2850.690 886.420 2851.010 886.480 ;
        RECT 2849.770 817.600 2850.090 817.660 ;
        RECT 2849.575 817.460 2850.090 817.600 ;
        RECT 2849.770 817.400 2850.090 817.460 ;
        RECT 2849.770 789.380 2850.090 789.440 ;
        RECT 2849.770 789.240 2850.285 789.380 ;
        RECT 2849.770 789.180 2850.090 789.240 ;
        RECT 2849.770 746.540 2850.090 746.600 ;
        RECT 2849.770 746.400 2850.285 746.540 ;
        RECT 2849.770 746.340 2850.090 746.400 ;
        RECT 2849.770 742.460 2850.090 742.520 ;
        RECT 2851.625 742.460 2851.915 742.505 ;
        RECT 2849.770 742.320 2851.915 742.460 ;
        RECT 2849.770 742.260 2850.090 742.320 ;
        RECT 2851.625 742.275 2851.915 742.320 ;
        RECT 2849.770 665.620 2850.090 665.680 ;
        RECT 2851.625 665.620 2851.915 665.665 ;
        RECT 2849.770 665.480 2851.915 665.620 ;
        RECT 2849.770 665.420 2850.090 665.480 ;
        RECT 2851.625 665.435 2851.915 665.480 ;
        RECT 2850.230 330.040 2850.550 330.100 ;
        RECT 2852.545 330.040 2852.835 330.085 ;
        RECT 2850.230 329.900 2852.835 330.040 ;
        RECT 2850.230 329.840 2850.550 329.900 ;
        RECT 2852.545 329.855 2852.835 329.900 ;
        RECT 2852.545 282.935 2852.835 283.165 ;
        RECT 2849.770 282.780 2850.090 282.840 ;
        RECT 2852.620 282.780 2852.760 282.935 ;
        RECT 2849.770 282.640 2852.760 282.780 ;
        RECT 2849.770 282.580 2850.090 282.640 ;
        RECT 2849.770 216.480 2850.090 216.540 ;
        RECT 2852.545 216.480 2852.835 216.525 ;
        RECT 2849.770 216.340 2852.835 216.480 ;
        RECT 2849.770 216.280 2850.090 216.340 ;
        RECT 2852.545 216.295 2852.835 216.340 ;
        RECT 2851.150 195.400 2851.470 195.460 ;
        RECT 2852.545 195.400 2852.835 195.445 ;
        RECT 2851.150 195.260 2852.835 195.400 ;
        RECT 2851.150 195.200 2851.470 195.260 ;
        RECT 2852.545 195.215 2852.835 195.260 ;
      LAYER via ;
        RECT 2849.800 2162.440 2850.060 2162.700 ;
        RECT 2849.800 2090.700 2850.060 2090.960 ;
        RECT 2849.800 2035.280 2850.060 2035.540 ;
        RECT 2850.260 2035.280 2850.520 2035.540 ;
        RECT 2850.260 1997.540 2850.520 1997.800 ;
        RECT 2849.800 1913.220 2850.060 1913.480 ;
        RECT 2849.800 1909.140 2850.060 1909.400 ;
        RECT 2849.800 1882.620 2850.060 1882.880 ;
        RECT 2849.800 1848.620 2850.060 1848.880 ;
        RECT 2849.800 1738.460 2850.060 1738.720 ;
        RECT 2851.180 1577.980 2851.440 1578.240 ;
        RECT 2850.260 1577.640 2850.520 1577.900 ;
        RECT 2850.260 1521.200 2850.520 1521.460 ;
        RECT 2851.180 1463.740 2851.440 1464.000 ;
        RECT 2851.180 1427.360 2851.440 1427.620 ;
        RECT 2849.800 1348.820 2850.060 1349.080 ;
        RECT 2849.800 1336.240 2850.060 1336.500 ;
        RECT 2849.800 1299.180 2850.060 1299.440 ;
        RECT 2849.800 1282.520 2850.060 1282.780 ;
        RECT 2851.180 1282.520 2851.440 1282.780 ;
        RECT 2851.180 1134.280 2851.440 1134.540 ;
        RECT 2850.260 1022.080 2850.520 1022.340 ;
        RECT 2849.800 963.600 2850.060 963.860 ;
        RECT 2850.720 957.480 2850.980 957.740 ;
        RECT 2850.720 886.420 2850.980 886.680 ;
        RECT 2849.800 817.400 2850.060 817.660 ;
        RECT 2849.800 789.180 2850.060 789.440 ;
        RECT 2849.800 746.340 2850.060 746.600 ;
        RECT 2849.800 742.260 2850.060 742.520 ;
        RECT 2849.800 665.420 2850.060 665.680 ;
        RECT 2850.260 329.840 2850.520 330.100 ;
        RECT 2849.800 282.580 2850.060 282.840 ;
        RECT 2849.800 216.280 2850.060 216.540 ;
        RECT 2851.180 195.200 2851.440 195.460 ;
      LAYER met2 ;
        RECT 2851.630 2246.450 2851.910 2246.565 ;
        RECT 2848.940 2246.310 2851.910 2246.450 ;
        RECT 2848.940 2197.490 2849.080 2246.310 ;
        RECT 2851.630 2246.195 2851.910 2246.310 ;
        RECT 2848.940 2197.350 2849.540 2197.490 ;
        RECT 2849.400 2162.810 2849.540 2197.350 ;
        RECT 2849.400 2162.730 2850.000 2162.810 ;
        RECT 2849.400 2162.670 2850.060 2162.730 ;
        RECT 2849.800 2162.410 2850.060 2162.670 ;
        RECT 2849.800 2090.670 2850.060 2090.990 ;
        RECT 2849.860 2035.570 2850.000 2090.670 ;
        RECT 2849.800 2035.250 2850.060 2035.570 ;
        RECT 2850.260 2035.250 2850.520 2035.570 ;
        RECT 2850.320 1997.830 2850.460 2035.250 ;
        RECT 2850.260 1997.510 2850.520 1997.830 ;
        RECT 2849.800 1913.250 2850.060 1913.510 ;
        RECT 2848.940 1913.190 2850.060 1913.250 ;
        RECT 2848.940 1913.110 2850.000 1913.190 ;
        RECT 2848.940 1911.210 2849.080 1913.110 ;
        RECT 2848.940 1911.070 2850.000 1911.210 ;
        RECT 2849.860 1909.430 2850.000 1911.070 ;
        RECT 2849.800 1909.110 2850.060 1909.430 ;
        RECT 2849.800 1882.590 2850.060 1882.910 ;
        RECT 2849.860 1848.910 2850.000 1882.590 ;
        RECT 2849.800 1848.590 2850.060 1848.910 ;
        RECT 2849.800 1738.660 2850.060 1738.750 ;
        RECT 2849.400 1738.520 2850.060 1738.660 ;
        RECT 2849.400 1702.450 2849.540 1738.520 ;
        RECT 2849.800 1738.430 2850.060 1738.520 ;
        RECT 2849.400 1702.310 2850.000 1702.450 ;
        RECT 2849.860 1666.410 2850.000 1702.310 ;
        RECT 2848.940 1666.270 2850.000 1666.410 ;
        RECT 2848.940 1654.850 2849.080 1666.270 ;
        RECT 2848.940 1654.710 2851.380 1654.850 ;
        RECT 2851.240 1578.270 2851.380 1654.710 ;
        RECT 2851.180 1577.950 2851.440 1578.270 ;
        RECT 2850.260 1577.610 2850.520 1577.930 ;
        RECT 2850.320 1521.490 2850.460 1577.610 ;
        RECT 2850.260 1521.170 2850.520 1521.490 ;
        RECT 2851.180 1463.710 2851.440 1464.030 ;
        RECT 2851.240 1427.650 2851.380 1463.710 ;
        RECT 2851.180 1427.330 2851.440 1427.650 ;
        RECT 2849.800 1348.850 2850.060 1349.110 ;
        RECT 2848.940 1348.790 2850.060 1348.850 ;
        RECT 2848.940 1348.710 2850.000 1348.790 ;
        RECT 2848.940 1336.440 2849.080 1348.710 ;
        RECT 2849.800 1336.440 2850.060 1336.530 ;
        RECT 2848.940 1336.300 2850.060 1336.440 ;
        RECT 2849.800 1336.210 2850.060 1336.300 ;
        RECT 2849.800 1299.150 2850.060 1299.470 ;
        RECT 2849.860 1298.530 2850.000 1299.150 ;
        RECT 2849.400 1298.390 2850.000 1298.530 ;
        RECT 2849.400 1282.890 2849.540 1298.390 ;
        RECT 2849.400 1282.810 2850.000 1282.890 ;
        RECT 2849.400 1282.750 2850.060 1282.810 ;
        RECT 2849.800 1282.490 2850.060 1282.750 ;
        RECT 2851.180 1282.490 2851.440 1282.810 ;
        RECT 2851.240 1134.570 2851.380 1282.490 ;
        RECT 2851.180 1134.250 2851.440 1134.570 ;
        RECT 2850.260 1022.050 2850.520 1022.370 ;
        RECT 2850.320 994.570 2850.460 1022.050 ;
        RECT 2848.940 994.430 2850.460 994.570 ;
        RECT 2848.940 964.650 2849.080 994.430 ;
        RECT 2848.940 964.510 2850.000 964.650 ;
        RECT 2849.860 963.890 2850.000 964.510 ;
        RECT 2849.800 963.570 2850.060 963.890 ;
        RECT 2850.720 957.450 2850.980 957.770 ;
        RECT 2850.780 886.710 2850.920 957.450 ;
        RECT 2850.720 886.390 2850.980 886.710 ;
        RECT 2849.800 817.370 2850.060 817.690 ;
        RECT 2849.860 789.470 2850.000 817.370 ;
        RECT 2849.800 789.150 2850.060 789.470 ;
        RECT 2849.800 746.310 2850.060 746.630 ;
        RECT 2849.860 742.550 2850.000 746.310 ;
        RECT 2849.800 742.230 2850.060 742.550 ;
        RECT 2849.800 665.450 2850.060 665.710 ;
        RECT 2848.940 665.390 2850.060 665.450 ;
        RECT 2848.940 665.310 2850.000 665.390 ;
        RECT 2848.940 385.970 2849.080 665.310 ;
        RECT 2848.940 385.830 2850.460 385.970 ;
        RECT 2850.320 330.130 2850.460 385.830 ;
        RECT 2850.260 329.810 2850.520 330.130 ;
        RECT 2849.800 282.550 2850.060 282.870 ;
        RECT 2849.860 269.690 2850.000 282.550 ;
        RECT 2848.940 269.550 2850.000 269.690 ;
        RECT 2848.940 226.850 2849.080 269.550 ;
        RECT 2848.940 226.710 2850.000 226.850 ;
        RECT 2849.860 216.570 2850.000 226.710 ;
        RECT 2849.800 216.250 2850.060 216.570 ;
        RECT 2851.180 195.170 2851.440 195.490 ;
        RECT 2851.240 141.850 2851.380 195.170 ;
        RECT 2850.780 141.710 2851.380 141.850 ;
        RECT 2850.780 107.170 2850.920 141.710 ;
        RECT 2850.320 107.030 2850.920 107.170 ;
        RECT 2850.320 39.850 2850.460 107.030 ;
        RECT 2848.480 39.710 2850.460 39.850 ;
        RECT 597.240 2.820 598.300 2.960 ;
        RECT 597.240 2.400 597.380 2.820 ;
        RECT 597.030 -4.800 597.590 2.400 ;
        RECT 598.160 0.525 598.300 2.820 ;
        RECT 2848.480 0.525 2848.620 39.710 ;
        RECT 598.090 0.155 598.370 0.525 ;
        RECT 2848.410 0.155 2848.690 0.525 ;
      LAYER via2 ;
        RECT 2851.630 2246.240 2851.910 2246.520 ;
        RECT 598.090 0.200 598.370 0.480 ;
        RECT 2848.410 0.200 2848.690 0.480 ;
      LAYER met3 ;
        RECT 2851.000 2249.040 2855.000 2249.640 ;
        RECT 2851.390 2246.545 2851.690 2249.040 ;
        RECT 2851.390 2246.230 2851.935 2246.545 ;
        RECT 2851.605 2246.215 2851.935 2246.230 ;
        RECT 598.065 0.490 598.395 0.505 ;
        RECT 2848.385 0.490 2848.715 0.505 ;
        RECT 598.065 0.190 2848.715 0.490 ;
        RECT 598.065 0.175 598.395 0.190 ;
        RECT 2848.385 0.175 2848.715 0.190 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1972.625 3401.105 1972.795 3401.955 ;
        RECT 2063.245 3400.085 2063.415 3401.275 ;
        RECT 2256.445 3399.745 2256.615 3401.275 ;
        RECT 2307.965 3399.745 2308.135 3401.275 ;
        RECT 2347.985 3400.425 2348.155 3401.275 ;
        RECT 2452.405 3399.065 2452.575 3401.275 ;
        RECT 2501.165 3399.065 2501.335 3401.275 ;
        RECT 2549.005 3398.725 2549.175 3401.275 ;
        RECT 2581.665 3398.725 2581.835 3400.595 ;
        RECT 2645.145 3398.725 2645.315 3400.595 ;
        RECT 2669.985 3398.725 2670.155 3401.275 ;
        RECT 2694.365 3399.405 2694.535 3401.275 ;
        RECT 2734.385 3399.405 2734.555 3401.275 ;
        RECT 2767.045 3398.725 2767.215 3401.275 ;
        RECT 785.825 6.715 785.995 7.735 ;
        RECT 1326.325 7.565 1328.335 7.735 ;
        RECT 1326.325 7.225 1326.495 7.565 ;
        RECT 1328.165 7.395 1328.335 7.565 ;
        RECT 1328.165 7.225 1344.435 7.395 ;
        RECT 1410.965 7.225 1428.155 7.395 ;
        RECT 1428.445 7.225 1429.995 7.395 ;
        RECT 783.985 6.545 785.995 6.715 ;
        RECT 783.985 3.485 784.155 6.545 ;
        RECT 795.025 3.145 795.195 6.375 ;
        RECT 1410.045 5.695 1410.215 6.035 ;
        RECT 1410.965 5.695 1411.135 7.225 ;
        RECT 1410.045 5.525 1411.135 5.695 ;
        RECT 1446.385 4.335 1446.555 7.395 ;
        RECT 1790.465 6.885 1790.635 8.415 ;
        RECT 1836.465 6.205 1836.635 7.055 ;
        RECT 1873.725 5.865 1873.895 7.055 ;
        RECT 1942.265 6.885 1942.435 9.095 ;
        RECT 1957.905 6.885 1958.075 9.095 ;
        RECT 1446.385 4.165 1448.855 4.335 ;
      LAYER mcon ;
        RECT 1972.625 3401.785 1972.795 3401.955 ;
        RECT 2063.245 3401.105 2063.415 3401.275 ;
        RECT 2256.445 3401.105 2256.615 3401.275 ;
        RECT 2307.965 3401.105 2308.135 3401.275 ;
        RECT 2347.985 3401.105 2348.155 3401.275 ;
        RECT 2452.405 3401.105 2452.575 3401.275 ;
        RECT 2501.165 3401.105 2501.335 3401.275 ;
        RECT 2549.005 3401.105 2549.175 3401.275 ;
        RECT 2669.985 3401.105 2670.155 3401.275 ;
        RECT 2581.665 3400.425 2581.835 3400.595 ;
        RECT 2645.145 3400.425 2645.315 3400.595 ;
        RECT 2694.365 3401.105 2694.535 3401.275 ;
        RECT 2734.385 3401.105 2734.555 3401.275 ;
        RECT 2767.045 3401.105 2767.215 3401.275 ;
        RECT 1942.265 8.925 1942.435 9.095 ;
        RECT 1790.465 8.245 1790.635 8.415 ;
        RECT 785.825 7.565 785.995 7.735 ;
        RECT 1344.265 7.225 1344.435 7.395 ;
        RECT 1427.985 7.225 1428.155 7.395 ;
        RECT 1429.825 7.225 1429.995 7.395 ;
        RECT 1446.385 7.225 1446.555 7.395 ;
        RECT 795.025 6.205 795.195 6.375 ;
        RECT 1410.045 5.865 1410.215 6.035 ;
        RECT 1836.465 6.885 1836.635 7.055 ;
        RECT 1873.725 6.885 1873.895 7.055 ;
        RECT 1957.905 8.925 1958.075 9.095 ;
        RECT 1448.685 4.165 1448.855 4.335 ;
      LAYER met1 ;
        RECT 1921.030 3416.220 1921.350 3416.280 ;
        RECT 1955.990 3416.220 1956.310 3416.280 ;
        RECT 1921.030 3416.080 1956.310 3416.220 ;
        RECT 1921.030 3416.020 1921.350 3416.080 ;
        RECT 1955.990 3416.020 1956.310 3416.080 ;
        RECT 1955.990 3401.940 1956.310 3402.000 ;
        RECT 1972.565 3401.940 1972.855 3401.985 ;
        RECT 1955.990 3401.800 1972.855 3401.940 ;
        RECT 1955.990 3401.740 1956.310 3401.800 ;
        RECT 1972.565 3401.755 1972.855 3401.800 ;
        RECT 2831.830 3401.400 2832.150 3401.660 ;
        RECT 1972.565 3401.260 1972.855 3401.305 ;
        RECT 2063.185 3401.260 2063.475 3401.305 ;
        RECT 2256.385 3401.260 2256.675 3401.305 ;
        RECT 1972.565 3401.120 2039.020 3401.260 ;
        RECT 1972.565 3401.075 1972.855 3401.120 ;
        RECT 2038.880 3400.240 2039.020 3401.120 ;
        RECT 2063.185 3401.120 2256.675 3401.260 ;
        RECT 2063.185 3401.075 2063.475 3401.120 ;
        RECT 2256.385 3401.075 2256.675 3401.120 ;
        RECT 2307.905 3401.260 2308.195 3401.305 ;
        RECT 2347.925 3401.260 2348.215 3401.305 ;
        RECT 2452.345 3401.260 2452.635 3401.305 ;
        RECT 2307.905 3401.120 2348.215 3401.260 ;
        RECT 2307.905 3401.075 2308.195 3401.120 ;
        RECT 2347.925 3401.075 2348.215 3401.120 ;
        RECT 2390.320 3401.120 2452.635 3401.260 ;
        RECT 2347.925 3400.580 2348.215 3400.625 ;
        RECT 2390.320 3400.580 2390.460 3401.120 ;
        RECT 2452.345 3401.075 2452.635 3401.120 ;
        RECT 2501.105 3401.260 2501.395 3401.305 ;
        RECT 2548.945 3401.260 2549.235 3401.305 ;
        RECT 2501.105 3401.120 2549.235 3401.260 ;
        RECT 2501.105 3401.075 2501.395 3401.120 ;
        RECT 2548.945 3401.075 2549.235 3401.120 ;
        RECT 2669.925 3401.260 2670.215 3401.305 ;
        RECT 2694.305 3401.260 2694.595 3401.305 ;
        RECT 2669.925 3401.120 2694.595 3401.260 ;
        RECT 2669.925 3401.075 2670.215 3401.120 ;
        RECT 2694.305 3401.075 2694.595 3401.120 ;
        RECT 2734.325 3401.260 2734.615 3401.305 ;
        RECT 2766.985 3401.260 2767.275 3401.305 ;
        RECT 2734.325 3401.120 2767.275 3401.260 ;
        RECT 2734.325 3401.075 2734.615 3401.120 ;
        RECT 2766.985 3401.075 2767.275 3401.120 ;
        RECT 2347.925 3400.440 2390.460 3400.580 ;
        RECT 2581.605 3400.580 2581.895 3400.625 ;
        RECT 2645.085 3400.580 2645.375 3400.625 ;
        RECT 2581.605 3400.440 2645.375 3400.580 ;
        RECT 2347.925 3400.395 2348.215 3400.440 ;
        RECT 2581.605 3400.395 2581.895 3400.440 ;
        RECT 2645.085 3400.395 2645.375 3400.440 ;
        RECT 2063.185 3400.240 2063.475 3400.285 ;
        RECT 2038.880 3400.100 2063.475 3400.240 ;
        RECT 2063.185 3400.055 2063.475 3400.100 ;
        RECT 2256.385 3399.900 2256.675 3399.945 ;
        RECT 2307.905 3399.900 2308.195 3399.945 ;
        RECT 2256.385 3399.760 2308.195 3399.900 ;
        RECT 2256.385 3399.715 2256.675 3399.760 ;
        RECT 2307.905 3399.715 2308.195 3399.760 ;
        RECT 2694.305 3399.560 2694.595 3399.605 ;
        RECT 2734.325 3399.560 2734.615 3399.605 ;
        RECT 2694.305 3399.420 2734.615 3399.560 ;
        RECT 2694.305 3399.375 2694.595 3399.420 ;
        RECT 2734.325 3399.375 2734.615 3399.420 ;
        RECT 2452.345 3399.220 2452.635 3399.265 ;
        RECT 2501.105 3399.220 2501.395 3399.265 ;
        RECT 2452.345 3399.080 2501.395 3399.220 ;
        RECT 2452.345 3399.035 2452.635 3399.080 ;
        RECT 2501.105 3399.035 2501.395 3399.080 ;
        RECT 2548.945 3398.880 2549.235 3398.925 ;
        RECT 2581.605 3398.880 2581.895 3398.925 ;
        RECT 2548.945 3398.740 2581.895 3398.880 ;
        RECT 2548.945 3398.695 2549.235 3398.740 ;
        RECT 2581.605 3398.695 2581.895 3398.740 ;
        RECT 2645.085 3398.880 2645.375 3398.925 ;
        RECT 2669.925 3398.880 2670.215 3398.925 ;
        RECT 2645.085 3398.740 2670.215 3398.880 ;
        RECT 2645.085 3398.695 2645.375 3398.740 ;
        RECT 2669.925 3398.695 2670.215 3398.740 ;
        RECT 2766.985 3398.880 2767.275 3398.925 ;
        RECT 2831.920 3398.880 2832.060 3401.400 ;
        RECT 2766.985 3398.740 2832.060 3398.880 ;
        RECT 2766.985 3398.695 2767.275 3398.740 ;
        RECT 1942.205 9.080 1942.495 9.125 ;
        RECT 1957.845 9.080 1958.135 9.125 ;
        RECT 1942.205 8.940 1958.135 9.080 ;
        RECT 1942.205 8.895 1942.495 8.940 ;
        RECT 1957.845 8.895 1958.135 8.940 ;
        RECT 746.650 8.740 746.970 8.800 ;
        RECT 749.870 8.740 750.190 8.800 ;
        RECT 746.650 8.600 750.190 8.740 ;
        RECT 746.650 8.540 746.970 8.600 ;
        RECT 749.870 8.540 750.190 8.600 ;
        RECT 1743.470 8.400 1743.790 8.460 ;
        RECT 1790.405 8.400 1790.695 8.445 ;
        RECT 1743.470 8.260 1790.695 8.400 ;
        RECT 1743.470 8.200 1743.790 8.260 ;
        RECT 1790.405 8.215 1790.695 8.260 ;
        RECT 712.610 7.720 712.930 7.780 ;
        RECT 714.450 7.720 714.770 7.780 ;
        RECT 785.750 7.720 786.070 7.780 ;
        RECT 712.610 7.580 714.770 7.720 ;
        RECT 785.555 7.580 786.070 7.720 ;
        RECT 712.610 7.520 712.930 7.580 ;
        RECT 714.450 7.520 714.770 7.580 ;
        RECT 785.750 7.520 786.070 7.580 ;
        RECT 1325.790 7.380 1326.110 7.440 ;
        RECT 1326.265 7.380 1326.555 7.425 ;
        RECT 1344.190 7.380 1344.510 7.440 ;
        RECT 1325.790 7.240 1326.555 7.380 ;
        RECT 1343.995 7.240 1344.510 7.380 ;
        RECT 1325.790 7.180 1326.110 7.240 ;
        RECT 1326.265 7.195 1326.555 7.240 ;
        RECT 1344.190 7.180 1344.510 7.240 ;
        RECT 1427.925 7.380 1428.215 7.425 ;
        RECT 1428.385 7.380 1428.675 7.425 ;
        RECT 1427.925 7.240 1428.675 7.380 ;
        RECT 1427.925 7.195 1428.215 7.240 ;
        RECT 1428.385 7.195 1428.675 7.240 ;
        RECT 1429.765 7.380 1430.055 7.425 ;
        RECT 1446.325 7.380 1446.615 7.425 ;
        RECT 1429.765 7.240 1446.615 7.380 ;
        RECT 1429.765 7.195 1430.055 7.240 ;
        RECT 1446.325 7.195 1446.615 7.240 ;
        RECT 702.030 7.040 702.350 7.100 ;
        RECT 705.710 7.040 706.030 7.100 ;
        RECT 702.030 6.900 706.030 7.040 ;
        RECT 702.030 6.840 702.350 6.900 ;
        RECT 705.710 6.840 706.030 6.900 ;
        RECT 1790.405 7.040 1790.695 7.085 ;
        RECT 1836.405 7.040 1836.695 7.085 ;
        RECT 1790.405 6.900 1836.695 7.040 ;
        RECT 1790.405 6.855 1790.695 6.900 ;
        RECT 1836.405 6.855 1836.695 6.900 ;
        RECT 1873.665 7.040 1873.955 7.085 ;
        RECT 1942.205 7.040 1942.495 7.085 ;
        RECT 1873.665 6.900 1942.495 7.040 ;
        RECT 1873.665 6.855 1873.955 6.900 ;
        RECT 1942.205 6.855 1942.495 6.900 ;
        RECT 1957.845 7.040 1958.135 7.085 ;
        RECT 2829.070 7.040 2829.390 7.100 ;
        RECT 1957.845 6.900 2829.390 7.040 ;
        RECT 1957.845 6.855 1958.135 6.900 ;
        RECT 2829.070 6.840 2829.390 6.900 ;
        RECT 986.310 6.700 986.630 6.760 ;
        RECT 992.290 6.700 992.610 6.760 ;
        RECT 986.310 6.560 992.610 6.700 ;
        RECT 986.310 6.500 986.630 6.560 ;
        RECT 992.290 6.500 992.610 6.560 ;
        RECT 794.965 6.360 795.255 6.405 ;
        RECT 797.250 6.360 797.570 6.420 ;
        RECT 794.965 6.220 797.570 6.360 ;
        RECT 794.965 6.175 795.255 6.220 ;
        RECT 797.250 6.160 797.570 6.220 ;
        RECT 1836.405 6.360 1836.695 6.405 ;
        RECT 1836.405 6.220 1863.300 6.360 ;
        RECT 1836.405 6.175 1836.695 6.220 ;
        RECT 952.730 6.020 953.050 6.080 ;
        RECT 954.570 6.020 954.890 6.080 ;
        RECT 952.730 5.880 954.890 6.020 ;
        RECT 952.730 5.820 953.050 5.880 ;
        RECT 954.570 5.820 954.890 5.880 ;
        RECT 1409.510 6.020 1409.830 6.080 ;
        RECT 1409.985 6.020 1410.275 6.065 ;
        RECT 1409.510 5.880 1410.275 6.020 ;
        RECT 1863.160 6.020 1863.300 6.220 ;
        RECT 1873.665 6.020 1873.955 6.065 ;
        RECT 1863.160 5.880 1873.955 6.020 ;
        RECT 1409.510 5.820 1409.830 5.880 ;
        RECT 1409.985 5.835 1410.275 5.880 ;
        RECT 1873.665 5.835 1873.955 5.880 ;
        RECT 1448.625 4.320 1448.915 4.365 ;
        RECT 1468.850 4.320 1469.170 4.380 ;
        RECT 1448.625 4.180 1469.170 4.320 ;
        RECT 1448.625 4.135 1448.915 4.180 ;
        RECT 1468.850 4.120 1469.170 4.180 ;
        RECT 783.910 3.640 784.230 3.700 ;
        RECT 783.715 3.500 784.230 3.640 ;
        RECT 783.910 3.440 784.230 3.500 ;
        RECT 788.970 3.300 789.290 3.360 ;
        RECT 794.965 3.300 795.255 3.345 ;
        RECT 788.970 3.160 795.255 3.300 ;
        RECT 788.970 3.100 789.290 3.160 ;
        RECT 794.965 3.115 795.255 3.160 ;
      LAYER via ;
        RECT 1921.060 3416.020 1921.320 3416.280 ;
        RECT 1956.020 3416.020 1956.280 3416.280 ;
        RECT 1956.020 3401.740 1956.280 3402.000 ;
        RECT 2831.860 3401.400 2832.120 3401.660 ;
        RECT 746.680 8.540 746.940 8.800 ;
        RECT 749.900 8.540 750.160 8.800 ;
        RECT 1743.500 8.200 1743.760 8.460 ;
        RECT 712.640 7.520 712.900 7.780 ;
        RECT 714.480 7.520 714.740 7.780 ;
        RECT 785.780 7.520 786.040 7.780 ;
        RECT 1325.820 7.180 1326.080 7.440 ;
        RECT 1344.220 7.180 1344.480 7.440 ;
        RECT 702.060 6.840 702.320 7.100 ;
        RECT 705.740 6.840 706.000 7.100 ;
        RECT 2829.100 6.840 2829.360 7.100 ;
        RECT 986.340 6.500 986.600 6.760 ;
        RECT 992.320 6.500 992.580 6.760 ;
        RECT 797.280 6.160 797.540 6.420 ;
        RECT 952.760 5.820 953.020 6.080 ;
        RECT 954.600 5.820 954.860 6.080 ;
        RECT 1409.540 5.820 1409.800 6.080 ;
        RECT 1468.880 4.120 1469.140 4.380 ;
        RECT 783.940 3.440 784.200 3.700 ;
        RECT 789.000 3.100 789.260 3.360 ;
      LAYER met2 ;
        RECT 1921.060 3415.990 1921.320 3416.310 ;
        RECT 1956.020 3415.990 1956.280 3416.310 ;
        RECT 1921.120 3405.000 1921.260 3415.990 ;
        RECT 1920.990 3401.000 1921.270 3405.000 ;
        RECT 1956.080 3402.030 1956.220 3415.990 ;
        RECT 1956.020 3401.710 1956.280 3402.030 ;
        RECT 2831.850 3401.515 2832.130 3401.885 ;
        RECT 2831.860 3401.370 2832.120 3401.515 ;
        RECT 746.680 8.510 746.940 8.830 ;
        RECT 749.900 8.740 750.160 8.830 ;
        RECT 749.900 8.600 750.560 8.740 ;
        RECT 749.900 8.510 750.160 8.600 ;
        RECT 712.640 7.720 712.900 7.810 ;
        RECT 699.360 7.580 702.260 7.720 ;
        RECT 627.530 5.850 627.810 5.965 ;
        RECT 617.020 5.710 627.810 5.850 ;
        RECT 615.180 2.820 616.240 2.960 ;
        RECT 615.180 2.400 615.320 2.820 ;
        RECT 614.970 -4.800 615.530 2.400 ;
        RECT 616.100 1.090 616.240 2.820 ;
        RECT 617.020 1.090 617.160 5.710 ;
        RECT 627.530 5.595 627.810 5.710 ;
        RECT 633.510 5.850 633.790 5.965 ;
        RECT 642.250 5.850 642.530 5.965 ;
        RECT 633.510 5.710 642.530 5.850 ;
        RECT 633.510 5.595 633.790 5.710 ;
        RECT 642.250 5.595 642.530 5.710 ;
        RECT 677.670 5.595 677.950 5.965 ;
        RECT 677.740 5.170 677.880 5.595 ;
        RECT 699.360 5.340 699.500 7.580 ;
        RECT 702.120 7.130 702.260 7.580 ;
        RECT 705.800 7.580 712.900 7.720 ;
        RECT 705.800 7.130 705.940 7.580 ;
        RECT 712.640 7.490 712.900 7.580 ;
        RECT 714.480 7.490 714.740 7.810 ;
        RECT 702.060 6.810 702.320 7.130 ;
        RECT 705.740 6.810 706.000 7.130 ;
        RECT 679.050 5.170 679.330 5.285 ;
        RECT 677.740 5.030 679.330 5.170 ;
        RECT 679.050 4.915 679.330 5.030 ;
        RECT 695.150 5.170 695.430 5.285 ;
        RECT 697.060 5.200 699.500 5.340 ;
        RECT 697.060 5.170 697.200 5.200 ;
        RECT 695.150 5.030 697.200 5.170 ;
        RECT 695.150 4.915 695.430 5.030 ;
        RECT 714.540 5.000 714.680 7.490 ;
        RECT 726.960 6.220 728.940 6.360 ;
        RECT 726.960 5.000 727.100 6.220 ;
        RECT 714.540 4.860 727.100 5.000 ;
        RECT 728.800 3.925 728.940 6.220 ;
        RECT 728.730 3.555 729.010 3.925 ;
        RECT 734.710 3.640 734.990 3.925 ;
        RECT 746.740 3.640 746.880 8.510 ;
        RECT 750.420 7.890 750.560 8.600 ;
        RECT 993.690 8.570 993.970 8.685 ;
        RECT 784.460 8.430 785.980 8.570 ;
        RECT 753.640 8.260 771.260 8.400 ;
        RECT 753.640 7.890 753.780 8.260 ;
        RECT 771.120 8.060 771.260 8.260 ;
        RECT 784.460 8.060 784.600 8.430 ;
        RECT 771.120 7.920 784.600 8.060 ;
        RECT 750.420 7.750 753.780 7.890 ;
        RECT 785.840 7.810 785.980 8.430 ;
        RECT 992.380 8.430 993.970 8.570 ;
        RECT 785.780 7.490 786.040 7.810 ;
        RECT 923.310 7.635 923.590 8.005 ;
        RECT 797.280 6.130 797.540 6.450 ;
        RECT 797.340 5.965 797.480 6.130 ;
        RECT 797.270 5.595 797.550 5.965 ;
        RECT 923.380 4.490 923.520 7.635 ;
        RECT 992.380 6.790 992.520 8.430 ;
        RECT 993.690 8.315 993.970 8.430 ;
        RECT 1743.500 8.170 1743.760 8.490 ;
        RECT 1313.000 7.750 1325.560 7.890 ;
        RECT 1122.490 7.210 1122.770 7.325 ;
        RECT 1122.490 7.070 1123.160 7.210 ;
        RECT 1122.490 6.955 1122.770 7.070 ;
        RECT 986.340 6.470 986.600 6.790 ;
        RECT 992.320 6.470 992.580 6.790 ;
        RECT 952.760 6.020 953.020 6.110 ;
        RECT 952.360 5.880 953.020 6.020 ;
        RECT 952.360 4.490 952.500 5.880 ;
        RECT 952.760 5.790 953.020 5.880 ;
        RECT 954.600 5.790 954.860 6.110 ;
        RECT 954.660 5.170 954.800 5.790 ;
        RECT 956.890 5.170 957.170 5.285 ;
        RECT 954.660 5.030 957.170 5.170 ;
        RECT 956.890 4.915 957.170 5.030 ;
        RECT 985.870 5.170 986.150 5.285 ;
        RECT 986.400 5.170 986.540 6.470 ;
        RECT 985.870 5.030 986.540 5.170 ;
        RECT 985.870 4.915 986.150 5.030 ;
        RECT 923.380 4.350 952.500 4.490 ;
        RECT 1123.020 3.925 1123.160 7.070 ;
        RECT 784.000 3.730 789.200 3.810 ;
        RECT 734.710 3.555 746.880 3.640 ;
        RECT 734.780 3.500 746.880 3.555 ;
        RECT 783.940 3.670 789.200 3.730 ;
        RECT 783.940 3.410 784.200 3.670 ;
        RECT 789.060 3.390 789.200 3.670 ;
        RECT 1122.950 3.555 1123.230 3.925 ;
        RECT 789.000 3.070 789.260 3.390 ;
        RECT 1313.000 3.245 1313.140 7.750 ;
        RECT 1325.420 7.380 1325.560 7.750 ;
        RECT 1325.820 7.380 1326.080 7.470 ;
        RECT 1325.420 7.240 1326.080 7.380 ;
        RECT 1344.220 7.325 1344.480 7.470 ;
        RECT 1325.820 7.150 1326.080 7.240 ;
        RECT 1344.210 6.955 1344.490 7.325 ;
        RECT 1409.540 5.790 1409.800 6.110 ;
        RECT 1409.600 3.925 1409.740 5.790 ;
        RECT 1468.940 4.410 1473.680 4.490 ;
        RECT 1468.880 4.350 1473.680 4.410 ;
        RECT 1468.880 4.090 1469.140 4.350 ;
        RECT 1409.530 3.555 1409.810 3.925 ;
        RECT 1312.930 2.875 1313.210 3.245 ;
        RECT 1473.540 3.130 1473.680 4.350 ;
        RECT 1743.560 3.925 1743.700 8.170 ;
        RECT 2829.090 6.955 2829.370 7.325 ;
        RECT 2829.100 6.810 2829.360 6.955 ;
        RECT 1476.230 3.555 1476.510 3.925 ;
        RECT 1743.490 3.555 1743.770 3.925 ;
        RECT 1476.300 3.130 1476.440 3.555 ;
        RECT 1473.540 2.990 1476.440 3.130 ;
        RECT 616.100 0.950 617.160 1.090 ;
      LAYER via2 ;
        RECT 2831.850 3401.560 2832.130 3401.840 ;
        RECT 627.530 5.640 627.810 5.920 ;
        RECT 633.510 5.640 633.790 5.920 ;
        RECT 642.250 5.640 642.530 5.920 ;
        RECT 677.670 5.640 677.950 5.920 ;
        RECT 679.050 4.960 679.330 5.240 ;
        RECT 695.150 4.960 695.430 5.240 ;
        RECT 728.730 3.600 729.010 3.880 ;
        RECT 734.710 3.600 734.990 3.880 ;
        RECT 923.310 7.680 923.590 7.960 ;
        RECT 797.270 5.640 797.550 5.920 ;
        RECT 993.690 8.360 993.970 8.640 ;
        RECT 1122.490 7.000 1122.770 7.280 ;
        RECT 956.890 4.960 957.170 5.240 ;
        RECT 985.870 4.960 986.150 5.240 ;
        RECT 1122.950 3.600 1123.230 3.880 ;
        RECT 1344.210 7.000 1344.490 7.280 ;
        RECT 1409.530 3.600 1409.810 3.880 ;
        RECT 1312.930 2.920 1313.210 3.200 ;
        RECT 2829.090 7.000 2829.370 7.280 ;
        RECT 1476.230 3.600 1476.510 3.880 ;
        RECT 1743.490 3.600 1743.770 3.880 ;
      LAYER met3 ;
        RECT 2831.825 3401.860 2832.155 3401.865 ;
        RECT 2831.825 3401.850 2832.410 3401.860 ;
        RECT 2831.600 3401.550 2832.410 3401.850 ;
        RECT 2831.825 3401.540 2832.410 3401.550 ;
        RECT 2831.825 3401.535 2832.155 3401.540 ;
        RECT 993.665 8.650 993.995 8.665 ;
        RECT 993.665 8.350 999.730 8.650 ;
        RECT 993.665 8.335 993.995 8.350 ;
        RECT 890.830 7.970 891.210 7.980 ;
        RECT 889.030 7.670 891.210 7.970 ;
        RECT 885.310 7.290 885.690 7.300 ;
        RECT 889.030 7.290 889.330 7.670 ;
        RECT 890.830 7.660 891.210 7.670 ;
        RECT 920.270 7.970 920.650 7.980 ;
        RECT 923.285 7.970 923.615 7.985 ;
        RECT 920.270 7.670 923.615 7.970 ;
        RECT 999.430 7.970 999.730 8.350 ;
        RECT 1004.910 7.970 1005.290 7.980 ;
        RECT 999.430 7.670 1005.290 7.970 ;
        RECT 920.270 7.660 920.650 7.670 ;
        RECT 923.285 7.655 923.615 7.670 ;
        RECT 1004.910 7.660 1005.290 7.670 ;
        RECT 1195.350 7.970 1195.730 7.980 ;
        RECT 1209.150 7.970 1209.530 7.980 ;
        RECT 1195.350 7.670 1209.530 7.970 ;
        RECT 1195.350 7.660 1195.730 7.670 ;
        RECT 1209.150 7.660 1209.530 7.670 ;
        RECT 1122.465 7.300 1122.795 7.305 ;
        RECT 1344.185 7.300 1344.515 7.305 ;
        RECT 1122.465 7.290 1123.050 7.300 ;
        RECT 885.310 6.990 889.330 7.290 ;
        RECT 1122.240 6.990 1123.050 7.290 ;
        RECT 885.310 6.980 885.690 6.990 ;
        RECT 1122.465 6.980 1123.050 6.990 ;
        RECT 1215.590 7.290 1215.970 7.300 ;
        RECT 1225.710 7.290 1226.090 7.300 ;
        RECT 1344.185 7.290 1344.770 7.300 ;
        RECT 1215.590 6.990 1226.090 7.290 ;
        RECT 1343.960 6.990 1344.770 7.290 ;
        RECT 1215.590 6.980 1215.970 6.990 ;
        RECT 1225.710 6.980 1226.090 6.990 ;
        RECT 1344.185 6.980 1344.770 6.990 ;
        RECT 1359.110 7.290 1359.490 7.300 ;
        RECT 1366.470 7.290 1366.850 7.300 ;
        RECT 1359.110 6.990 1366.850 7.290 ;
        RECT 1359.110 6.980 1359.490 6.990 ;
        RECT 1366.470 6.980 1366.850 6.990 ;
        RECT 1368.310 7.290 1368.690 7.300 ;
        RECT 1396.830 7.290 1397.210 7.300 ;
        RECT 1368.310 6.990 1397.210 7.290 ;
        RECT 1368.310 6.980 1368.690 6.990 ;
        RECT 1396.830 6.980 1397.210 6.990 ;
        RECT 2829.065 7.290 2829.395 7.305 ;
        RECT 2832.030 7.290 2832.410 7.300 ;
        RECT 2829.065 6.990 2832.410 7.290 ;
        RECT 1122.465 6.975 1122.795 6.980 ;
        RECT 1344.185 6.975 1344.515 6.980 ;
        RECT 2829.065 6.975 2829.395 6.990 ;
        RECT 2832.030 6.980 2832.410 6.990 ;
        RECT 627.505 5.930 627.835 5.945 ;
        RECT 633.485 5.930 633.815 5.945 ;
        RECT 627.505 5.630 633.815 5.930 ;
        RECT 627.505 5.615 627.835 5.630 ;
        RECT 633.485 5.615 633.815 5.630 ;
        RECT 642.225 5.930 642.555 5.945 ;
        RECT 677.645 5.930 677.975 5.945 ;
        RECT 642.225 5.630 677.975 5.930 ;
        RECT 642.225 5.615 642.555 5.630 ;
        RECT 677.645 5.615 677.975 5.630 ;
        RECT 797.245 5.930 797.575 5.945 ;
        RECT 831.030 5.930 831.410 5.940 ;
        RECT 797.245 5.630 831.410 5.930 ;
        RECT 797.245 5.615 797.575 5.630 ;
        RECT 831.030 5.620 831.410 5.630 ;
        RECT 866.910 5.930 867.290 5.940 ;
        RECT 880.710 5.930 881.090 5.940 ;
        RECT 866.910 5.630 881.090 5.930 ;
        RECT 866.910 5.620 867.290 5.630 ;
        RECT 880.710 5.620 881.090 5.630 ;
        RECT 679.025 5.250 679.355 5.265 ;
        RECT 695.125 5.250 695.455 5.265 ;
        RECT 679.025 4.950 695.455 5.250 ;
        RECT 679.025 4.935 679.355 4.950 ;
        RECT 695.125 4.935 695.455 4.950 ;
        RECT 956.865 5.250 957.195 5.265 ;
        RECT 985.845 5.250 986.175 5.265 ;
        RECT 1263.430 5.250 1263.810 5.260 ;
        RECT 956.865 4.950 986.175 5.250 ;
        RECT 956.865 4.935 957.195 4.950 ;
        RECT 985.845 4.935 986.175 4.950 ;
        RECT 1258.870 4.950 1263.810 5.250 ;
        RECT 1251.470 4.570 1251.850 4.580 ;
        RECT 1258.870 4.570 1259.170 4.950 ;
        RECT 1263.430 4.940 1263.810 4.950 ;
        RECT 1251.470 4.270 1259.170 4.570 ;
        RECT 1268.950 4.570 1269.330 4.580 ;
        RECT 1278.150 4.570 1278.530 4.580 ;
        RECT 1268.950 4.270 1278.530 4.570 ;
        RECT 1251.470 4.260 1251.850 4.270 ;
        RECT 1268.950 4.260 1269.330 4.270 ;
        RECT 1278.150 4.260 1278.530 4.270 ;
        RECT 728.705 3.890 729.035 3.905 ;
        RECT 734.685 3.890 735.015 3.905 ;
        RECT 728.705 3.590 735.015 3.890 ;
        RECT 728.705 3.575 729.035 3.590 ;
        RECT 734.685 3.575 735.015 3.590 ;
        RECT 1122.925 3.890 1123.255 3.905 ;
        RECT 1155.790 3.890 1156.170 3.900 ;
        RECT 1122.925 3.590 1156.170 3.890 ;
        RECT 1122.925 3.575 1123.255 3.590 ;
        RECT 1155.790 3.580 1156.170 3.590 ;
        RECT 1305.750 3.890 1306.130 3.900 ;
        RECT 1403.270 3.890 1403.650 3.900 ;
        RECT 1409.505 3.890 1409.835 3.905 ;
        RECT 1305.750 3.590 1308.850 3.890 ;
        RECT 1305.750 3.580 1306.130 3.590 ;
        RECT 1308.550 3.210 1308.850 3.590 ;
        RECT 1403.270 3.590 1409.835 3.890 ;
        RECT 1403.270 3.580 1403.650 3.590 ;
        RECT 1409.505 3.575 1409.835 3.590 ;
        RECT 1476.205 3.890 1476.535 3.905 ;
        RECT 1743.465 3.890 1743.795 3.905 ;
        RECT 1476.205 3.590 1743.795 3.890 ;
        RECT 1476.205 3.575 1476.535 3.590 ;
        RECT 1743.465 3.575 1743.795 3.590 ;
        RECT 1312.905 3.210 1313.235 3.225 ;
        RECT 1308.550 2.910 1313.235 3.210 ;
        RECT 1312.905 2.895 1313.235 2.910 ;
      LAYER via3 ;
        RECT 2832.060 3401.540 2832.380 3401.860 ;
        RECT 885.340 6.980 885.660 7.300 ;
        RECT 890.860 7.660 891.180 7.980 ;
        RECT 920.300 7.660 920.620 7.980 ;
        RECT 1004.940 7.660 1005.260 7.980 ;
        RECT 1195.380 7.660 1195.700 7.980 ;
        RECT 1209.180 7.660 1209.500 7.980 ;
        RECT 1122.700 6.980 1123.020 7.300 ;
        RECT 1215.620 6.980 1215.940 7.300 ;
        RECT 1225.740 6.980 1226.060 7.300 ;
        RECT 1344.420 6.980 1344.740 7.300 ;
        RECT 1359.140 6.980 1359.460 7.300 ;
        RECT 1366.500 6.980 1366.820 7.300 ;
        RECT 1368.340 6.980 1368.660 7.300 ;
        RECT 1396.860 6.980 1397.180 7.300 ;
        RECT 2832.060 6.980 2832.380 7.300 ;
        RECT 831.060 5.620 831.380 5.940 ;
        RECT 866.940 5.620 867.260 5.940 ;
        RECT 880.740 5.620 881.060 5.940 ;
        RECT 1251.500 4.260 1251.820 4.580 ;
        RECT 1263.460 4.940 1263.780 5.260 ;
        RECT 1268.980 4.260 1269.300 4.580 ;
        RECT 1278.180 4.260 1278.500 4.580 ;
        RECT 1155.820 3.580 1156.140 3.900 ;
        RECT 1305.780 3.580 1306.100 3.900 ;
        RECT 1403.300 3.580 1403.620 3.900 ;
      LAYER met4 ;
        RECT 2832.055 3401.535 2832.385 3401.865 ;
        RECT 1004.510 14.710 1005.690 15.890 ;
        RECT 1120.430 14.710 1121.610 15.890 ;
        RECT 1004.950 7.985 1005.250 14.710 ;
        RECT 1120.870 12.050 1121.170 14.710 ;
        RECT 1120.870 11.750 1123.010 12.050 ;
        RECT 1122.710 9.330 1123.010 11.750 ;
        RECT 1225.750 11.750 1228.810 12.050 ;
        RECT 1122.710 9.030 1125.770 9.330 ;
        RECT 882.590 7.670 885.650 7.970 ;
        RECT 882.590 7.290 882.890 7.670 ;
        RECT 885.350 7.305 885.650 7.670 ;
        RECT 890.855 7.655 891.185 7.985 ;
        RECT 920.295 7.970 920.625 7.985 ;
        RECT 910.190 7.670 920.625 7.970 ;
        RECT 880.750 6.990 882.890 7.290 ;
        RECT 880.750 5.945 881.050 6.990 ;
        RECT 885.335 6.975 885.665 7.305 ;
        RECT 890.870 7.290 891.170 7.655 ;
        RECT 910.190 7.290 910.490 7.670 ;
        RECT 920.295 7.655 920.625 7.670 ;
        RECT 1004.935 7.655 1005.265 7.985 ;
        RECT 890.870 6.990 910.490 7.290 ;
        RECT 1122.695 7.290 1123.025 7.305 ;
        RECT 1125.470 7.290 1125.770 9.030 ;
        RECT 1122.695 6.990 1125.770 7.290 ;
        RECT 1155.830 8.350 1169.930 8.650 ;
        RECT 1122.695 6.975 1123.025 6.990 ;
        RECT 831.055 5.615 831.385 5.945 ;
        RECT 866.935 5.930 867.265 5.945 ;
        RECT 855.910 5.630 867.265 5.930 ;
        RECT 831.070 4.570 831.370 5.615 ;
        RECT 855.910 5.250 856.210 5.630 ;
        RECT 866.935 5.615 867.265 5.630 ;
        RECT 880.735 5.615 881.065 5.945 ;
        RECT 852.230 4.950 856.210 5.250 ;
        RECT 852.230 4.570 852.530 4.950 ;
        RECT 831.070 4.270 852.530 4.570 ;
        RECT 1155.830 3.905 1156.130 8.350 ;
        RECT 1169.630 7.970 1169.930 8.350 ;
        RECT 1169.630 7.670 1170.850 7.970 ;
        RECT 1170.550 7.290 1170.850 7.670 ;
        RECT 1195.375 7.655 1195.705 7.985 ;
        RECT 1209.175 7.655 1209.505 7.985 ;
        RECT 1195.390 7.290 1195.690 7.655 ;
        RECT 1170.550 6.990 1195.690 7.290 ;
        RECT 1209.190 7.290 1209.490 7.655 ;
        RECT 1225.750 7.305 1226.050 11.750 ;
        RECT 1228.510 9.330 1228.810 11.750 ;
        RECT 1228.510 9.030 1246.290 9.330 ;
        RECT 1215.615 7.290 1215.945 7.305 ;
        RECT 1209.190 6.990 1215.945 7.290 ;
        RECT 1215.615 6.975 1215.945 6.990 ;
        RECT 1225.735 6.975 1226.065 7.305 ;
        RECT 1245.990 4.570 1246.290 9.030 ;
        RECT 1398.710 9.030 1401.770 9.330 ;
        RECT 1344.430 7.670 1359.450 7.970 ;
        RECT 1344.430 7.305 1344.730 7.670 ;
        RECT 1359.150 7.305 1359.450 7.670 ;
        RECT 1344.415 6.975 1344.745 7.305 ;
        RECT 1359.135 6.975 1359.465 7.305 ;
        RECT 1366.495 6.975 1366.825 7.305 ;
        RECT 1368.335 6.975 1368.665 7.305 ;
        RECT 1396.855 7.290 1397.185 7.305 ;
        RECT 1398.710 7.290 1399.010 9.030 ;
        RECT 1401.470 8.650 1401.770 9.030 ;
        RECT 1401.470 8.350 1403.610 8.650 ;
        RECT 1396.855 6.990 1399.010 7.290 ;
        RECT 1396.855 6.975 1397.185 6.990 ;
        RECT 1291.070 6.310 1306.090 6.610 ;
        RECT 1263.455 4.935 1263.785 5.265 ;
        RECT 1291.070 5.250 1291.370 6.310 ;
        RECT 1290.150 4.950 1291.370 5.250 ;
        RECT 1251.495 4.570 1251.825 4.585 ;
        RECT 1245.990 4.270 1251.825 4.570 ;
        RECT 1263.470 4.570 1263.770 4.935 ;
        RECT 1268.975 4.570 1269.305 4.585 ;
        RECT 1263.470 4.270 1269.305 4.570 ;
        RECT 1251.495 4.255 1251.825 4.270 ;
        RECT 1268.975 4.255 1269.305 4.270 ;
        RECT 1278.175 4.255 1278.505 4.585 ;
        RECT 1155.815 3.575 1156.145 3.905 ;
        RECT 1278.190 3.210 1278.490 4.255 ;
        RECT 1290.150 3.210 1290.450 4.950 ;
        RECT 1305.790 3.905 1306.090 6.310 ;
        RECT 1366.510 5.250 1366.810 6.975 ;
        RECT 1368.350 5.250 1368.650 6.975 ;
        RECT 1366.510 4.950 1368.650 5.250 ;
        RECT 1403.310 3.905 1403.610 8.350 ;
        RECT 2832.070 7.305 2832.370 3401.535 ;
        RECT 2832.055 6.975 2832.385 7.305 ;
        RECT 1305.775 3.575 1306.105 3.905 ;
        RECT 1403.295 3.575 1403.625 3.905 ;
        RECT 1278.190 2.910 1290.450 3.210 ;
      LAYER met5 ;
        RECT 1004.300 14.500 1121.820 16.100 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 195.645 6.545 195.815 8.415 ;
        RECT 580.665 6.715 580.835 9.095 ;
        RECT 581.585 6.715 581.755 7.055 ;
        RECT 580.665 6.545 581.755 6.715 ;
        RECT 245.785 3.825 245.955 6.035 ;
        RECT 1598.185 4.165 1598.355 7.055 ;
        RECT 1880.165 5.185 1880.335 8.755 ;
      LAYER mcon ;
        RECT 580.665 8.925 580.835 9.095 ;
        RECT 195.645 8.245 195.815 8.415 ;
        RECT 1880.165 8.585 1880.335 8.755 ;
        RECT 581.585 6.885 581.755 7.055 ;
        RECT 1598.185 6.885 1598.355 7.055 ;
        RECT 245.785 5.865 245.955 6.035 ;
      LAYER met1 ;
        RECT 580.605 9.080 580.895 9.125 ;
        RECT 534.680 8.940 580.895 9.080 ;
        RECT 283.430 8.740 283.750 8.800 ;
        RECT 534.680 8.740 534.820 8.940 ;
        RECT 580.605 8.895 580.895 8.940 ;
        RECT 283.430 8.600 534.820 8.740 ;
        RECT 1880.105 8.740 1880.395 8.785 ;
        RECT 2022.230 8.740 2022.550 8.800 ;
        RECT 1880.105 8.600 2022.550 8.740 ;
        RECT 283.430 8.540 283.750 8.600 ;
        RECT 1880.105 8.555 1880.395 8.600 ;
        RECT 2022.230 8.540 2022.550 8.600 ;
        RECT 195.585 8.400 195.875 8.445 ;
        RECT 213.510 8.400 213.830 8.460 ;
        RECT 195.585 8.260 213.830 8.400 ;
        RECT 195.585 8.215 195.875 8.260 ;
        RECT 213.510 8.200 213.830 8.260 ;
        RECT 145.430 7.040 145.750 7.100 ;
        RECT 581.525 7.040 581.815 7.085 ;
        RECT 597.150 7.040 597.470 7.100 ;
        RECT 145.430 6.900 172.340 7.040 ;
        RECT 145.430 6.840 145.750 6.900 ;
        RECT 172.200 6.700 172.340 6.900 ;
        RECT 581.525 6.900 597.470 7.040 ;
        RECT 581.525 6.855 581.815 6.900 ;
        RECT 597.150 6.840 597.470 6.900 ;
        RECT 598.990 7.040 599.310 7.100 ;
        RECT 601.750 7.040 602.070 7.100 ;
        RECT 598.990 6.900 602.070 7.040 ;
        RECT 598.990 6.840 599.310 6.900 ;
        RECT 601.750 6.840 602.070 6.900 ;
        RECT 1548.890 7.040 1549.210 7.100 ;
        RECT 1598.125 7.040 1598.415 7.085 ;
        RECT 1548.890 6.900 1598.415 7.040 ;
        RECT 1548.890 6.840 1549.210 6.900 ;
        RECT 1598.125 6.855 1598.415 6.900 ;
        RECT 195.585 6.700 195.875 6.745 ;
        RECT 172.200 6.560 195.875 6.700 ;
        RECT 195.585 6.515 195.875 6.560 ;
        RECT 245.725 6.020 246.015 6.065 ;
        RECT 283.430 6.020 283.750 6.080 ;
        RECT 245.725 5.880 283.750 6.020 ;
        RECT 245.725 5.835 246.015 5.880 ;
        RECT 283.430 5.820 283.750 5.880 ;
        RECT 1880.105 5.340 1880.395 5.385 ;
        RECT 1864.540 5.200 1880.395 5.340 ;
        RECT 1864.540 5.000 1864.680 5.200 ;
        RECT 1880.105 5.155 1880.395 5.200 ;
        RECT 1864.080 4.860 1864.680 5.000 ;
        RECT 1864.080 4.660 1864.220 4.860 ;
        RECT 1863.620 4.520 1864.220 4.660 ;
        RECT 1598.125 4.320 1598.415 4.365 ;
        RECT 1863.620 4.320 1863.760 4.520 ;
        RECT 559.520 4.180 562.420 4.320 ;
        RECT 240.190 3.980 240.510 4.040 ;
        RECT 245.725 3.980 246.015 4.025 ;
        RECT 240.190 3.840 246.015 3.980 ;
        RECT 240.190 3.780 240.510 3.840 ;
        RECT 245.725 3.795 246.015 3.840 ;
        RECT 558.050 3.640 558.370 3.700 ;
        RECT 559.520 3.640 559.660 4.180 ;
        RECT 562.280 3.980 562.420 4.180 ;
        RECT 1598.125 4.180 1863.760 4.320 ;
        RECT 1598.125 4.135 1598.415 4.180 ;
        RECT 564.030 3.980 564.350 4.040 ;
        RECT 562.280 3.840 564.350 3.980 ;
        RECT 564.030 3.780 564.350 3.840 ;
        RECT 558.050 3.500 559.660 3.640 ;
        RECT 558.050 3.440 558.370 3.500 ;
        RECT 1235.170 2.620 1235.490 2.680 ;
        RECT 1237.470 2.620 1237.790 2.680 ;
        RECT 1235.170 2.480 1237.790 2.620 ;
        RECT 1235.170 2.420 1235.490 2.480 ;
        RECT 1237.470 2.420 1237.790 2.480 ;
      LAYER via ;
        RECT 283.460 8.540 283.720 8.800 ;
        RECT 2022.260 8.540 2022.520 8.800 ;
        RECT 213.540 8.200 213.800 8.460 ;
        RECT 145.460 6.840 145.720 7.100 ;
        RECT 597.180 6.840 597.440 7.100 ;
        RECT 599.020 6.840 599.280 7.100 ;
        RECT 601.780 6.840 602.040 7.100 ;
        RECT 1548.920 6.840 1549.180 7.100 ;
        RECT 283.460 5.820 283.720 6.080 ;
        RECT 240.220 3.780 240.480 4.040 ;
        RECT 558.080 3.440 558.340 3.700 ;
        RECT 564.060 3.780 564.320 4.040 ;
        RECT 1235.200 2.420 1235.460 2.680 ;
        RECT 1237.500 2.420 1237.760 2.680 ;
      LAYER met2 ;
        RECT 283.460 8.510 283.720 8.830 ;
        RECT 213.540 8.170 213.800 8.490 ;
        RECT 213.600 8.005 213.740 8.170 ;
        RECT 213.530 7.635 213.810 8.005 ;
        RECT 240.210 7.635 240.490 8.005 ;
        RECT 145.460 6.810 145.720 7.130 ;
        RECT 109.570 2.875 109.850 3.245 ;
        RECT 109.640 2.400 109.780 2.875 ;
        RECT 145.520 2.400 145.660 6.810 ;
        RECT 240.280 4.070 240.420 7.635 ;
        RECT 283.520 6.110 283.660 8.510 ;
        RECT 598.490 7.210 598.770 9.000 ;
        RECT 2022.260 8.570 2022.520 8.830 ;
        RECT 2023.570 8.570 2023.850 9.000 ;
        RECT 2022.260 8.510 2023.850 8.570 ;
        RECT 2022.320 8.430 2023.850 8.510 ;
        RECT 597.240 7.130 598.770 7.210 ;
        RECT 597.180 7.070 598.770 7.130 ;
        RECT 597.180 6.810 597.440 7.070 ;
        RECT 283.460 5.790 283.720 6.110 ;
        RECT 598.490 5.850 598.770 7.070 ;
        RECT 599.020 6.810 599.280 7.130 ;
        RECT 601.780 6.810 602.040 7.130 ;
        RECT 1548.920 6.810 1549.180 7.130 ;
        RECT 599.080 5.850 599.220 6.810 ;
        RECT 601.840 5.965 601.980 6.810 ;
        RECT 657.430 6.530 657.710 6.645 ;
        RECT 657.040 6.390 657.710 6.530 ;
        RECT 597.240 5.710 599.220 5.850 ;
        RECT 597.240 5.170 597.380 5.710 ;
        RECT 582.520 5.030 597.380 5.170 ;
        RECT 564.120 4.350 568.400 4.490 ;
        RECT 564.120 4.070 564.260 4.350 ;
        RECT 240.220 3.750 240.480 4.070 ;
        RECT 564.060 3.750 564.320 4.070 ;
        RECT 558.080 3.410 558.340 3.730 ;
        RECT 558.140 3.245 558.280 3.410 ;
        RECT 558.070 2.875 558.350 3.245 ;
        RECT 568.260 3.130 568.400 4.350 ;
        RECT 578.840 3.500 580.360 3.640 ;
        RECT 578.840 3.245 578.980 3.500 ;
        RECT 580.220 3.300 580.360 3.500 ;
        RECT 582.520 3.300 582.660 5.030 ;
        RECT 598.490 5.000 598.770 5.710 ;
        RECT 601.770 5.595 602.050 5.965 ;
        RECT 657.040 4.490 657.180 6.390 ;
        RECT 657.430 6.275 657.710 6.390 ;
        RECT 663.020 4.520 682.020 4.660 ;
        RECT 697.060 4.605 698.120 4.660 ;
        RECT 1548.980 4.605 1549.120 6.810 ;
        RECT 2023.570 5.000 2023.850 8.430 ;
        RECT 657.040 4.350 662.700 4.490 ;
        RECT 662.560 4.320 662.700 4.350 ;
        RECT 663.020 4.320 663.160 4.520 ;
        RECT 681.880 4.490 682.020 4.520 ;
        RECT 691.930 4.490 692.210 4.605 ;
        RECT 681.880 4.350 692.210 4.490 ;
        RECT 662.560 4.180 663.160 4.320 ;
        RECT 691.930 4.235 692.210 4.350 ;
        RECT 696.990 4.520 698.190 4.605 ;
        RECT 696.990 4.235 697.270 4.520 ;
        RECT 697.910 4.235 698.190 4.520 ;
        RECT 988.630 4.490 988.910 4.605 ;
        RECT 990.930 4.490 991.210 4.605 ;
        RECT 988.630 4.350 991.210 4.490 ;
        RECT 988.630 4.235 988.910 4.350 ;
        RECT 990.930 4.235 991.210 4.350 ;
        RECT 1233.810 4.235 1234.090 4.605 ;
        RECT 1548.910 4.235 1549.190 4.605 ;
        RECT 1233.880 3.980 1234.020 4.235 ;
        RECT 1233.880 3.840 1235.400 3.980 ;
        RECT 570.490 3.130 570.770 3.245 ;
        RECT 568.260 2.990 570.770 3.130 ;
        RECT 570.490 2.875 570.770 2.990 ;
        RECT 578.770 2.875 579.050 3.245 ;
        RECT 580.220 3.160 582.660 3.300 ;
        RECT 1235.260 2.710 1235.400 3.840 ;
        RECT 1239.330 3.810 1239.610 3.925 ;
        RECT 1237.560 3.670 1239.610 3.810 ;
        RECT 1237.560 2.710 1237.700 3.670 ;
        RECT 1239.330 3.555 1239.610 3.670 ;
        RECT 109.430 -4.800 109.990 2.400 ;
        RECT 145.310 -4.800 145.870 2.400 ;
        RECT 1235.200 2.390 1235.460 2.710 ;
        RECT 1237.500 2.390 1237.760 2.710 ;
      LAYER via2 ;
        RECT 213.530 7.680 213.810 7.960 ;
        RECT 240.210 7.680 240.490 7.960 ;
        RECT 109.570 2.920 109.850 3.200 ;
        RECT 558.070 2.920 558.350 3.200 ;
        RECT 601.770 5.640 602.050 5.920 ;
        RECT 657.430 6.320 657.710 6.600 ;
        RECT 691.930 4.280 692.210 4.560 ;
        RECT 696.990 4.280 697.270 4.560 ;
        RECT 697.910 4.280 698.190 4.560 ;
        RECT 988.630 4.280 988.910 4.560 ;
        RECT 990.930 4.280 991.210 4.560 ;
        RECT 1233.810 4.280 1234.090 4.560 ;
        RECT 1548.910 4.280 1549.190 4.560 ;
        RECT 570.490 2.920 570.770 3.200 ;
        RECT 578.770 2.920 579.050 3.200 ;
        RECT 1239.330 3.600 1239.610 3.880 ;
      LAYER met3 ;
        RECT 213.505 7.970 213.835 7.985 ;
        RECT 240.185 7.970 240.515 7.985 ;
        RECT 213.505 7.670 240.515 7.970 ;
        RECT 213.505 7.655 213.835 7.670 ;
        RECT 240.185 7.655 240.515 7.670 ;
        RECT 657.405 6.620 657.735 6.625 ;
        RECT 657.150 6.610 657.735 6.620 ;
        RECT 657.150 6.310 657.960 6.610 ;
        RECT 657.150 6.300 657.735 6.310 ;
        RECT 657.405 6.295 657.735 6.300 ;
        RECT 601.745 5.930 602.075 5.945 ;
        RECT 626.790 5.930 627.170 5.940 ;
        RECT 601.745 5.630 627.170 5.930 ;
        RECT 601.745 5.615 602.075 5.630 ;
        RECT 626.790 5.620 627.170 5.630 ;
        RECT 691.905 4.570 692.235 4.585 ;
        RECT 696.965 4.570 697.295 4.585 ;
        RECT 691.905 4.270 697.295 4.570 ;
        RECT 691.905 4.255 692.235 4.270 ;
        RECT 696.965 4.255 697.295 4.270 ;
        RECT 697.885 4.570 698.215 4.585 ;
        RECT 753.750 4.570 754.130 4.580 ;
        RECT 697.885 4.270 754.130 4.570 ;
        RECT 697.885 4.255 698.215 4.270 ;
        RECT 753.750 4.260 754.130 4.270 ;
        RECT 756.510 4.570 756.890 4.580 ;
        RECT 988.605 4.570 988.935 4.585 ;
        RECT 756.510 4.270 988.935 4.570 ;
        RECT 756.510 4.260 756.890 4.270 ;
        RECT 988.605 4.255 988.935 4.270 ;
        RECT 990.905 4.570 991.235 4.585 ;
        RECT 1156.710 4.570 1157.090 4.580 ;
        RECT 990.905 4.270 1157.090 4.570 ;
        RECT 990.905 4.255 991.235 4.270 ;
        RECT 1156.710 4.260 1157.090 4.270 ;
        RECT 1168.670 4.570 1169.050 4.580 ;
        RECT 1233.785 4.570 1234.115 4.585 ;
        RECT 1548.885 4.570 1549.215 4.585 ;
        RECT 1168.670 4.270 1234.115 4.570 ;
        RECT 1168.670 4.260 1169.050 4.270 ;
        RECT 1233.785 4.255 1234.115 4.270 ;
        RECT 1279.110 4.270 1549.215 4.570 ;
        RECT 1239.305 3.890 1239.635 3.905 ;
        RECT 1261.590 3.890 1261.970 3.900 ;
        RECT 1239.305 3.590 1261.970 3.890 ;
        RECT 1239.305 3.575 1239.635 3.590 ;
        RECT 1261.590 3.580 1261.970 3.590 ;
        RECT 1262.510 3.890 1262.890 3.900 ;
        RECT 1279.110 3.890 1279.410 4.270 ;
        RECT 1548.885 4.255 1549.215 4.270 ;
        RECT 1262.510 3.590 1279.410 3.890 ;
        RECT 1262.510 3.580 1262.890 3.590 ;
        RECT 109.545 3.210 109.875 3.225 ;
        RECT 558.045 3.210 558.375 3.225 ;
        RECT 109.545 2.910 513.970 3.210 ;
        RECT 109.545 2.895 109.875 2.910 ;
        RECT 513.670 2.530 513.970 2.910 ;
        RECT 515.510 2.910 558.375 3.210 ;
        RECT 515.510 2.530 515.810 2.910 ;
        RECT 558.045 2.895 558.375 2.910 ;
        RECT 570.465 3.210 570.795 3.225 ;
        RECT 578.745 3.210 579.075 3.225 ;
        RECT 570.465 2.910 579.075 3.210 ;
        RECT 570.465 2.895 570.795 2.910 ;
        RECT 578.745 2.895 579.075 2.910 ;
        RECT 513.670 2.230 515.810 2.530 ;
      LAYER via3 ;
        RECT 657.180 6.300 657.500 6.620 ;
        RECT 626.820 5.620 627.140 5.940 ;
        RECT 753.780 4.260 754.100 4.580 ;
        RECT 756.540 4.260 756.860 4.580 ;
        RECT 1156.740 4.260 1157.060 4.580 ;
        RECT 1168.700 4.260 1169.020 4.580 ;
        RECT 1261.620 3.580 1261.940 3.900 ;
        RECT 1262.540 3.580 1262.860 3.900 ;
      LAYER met4 ;
        RECT 1156.750 7.670 1169.010 7.970 ;
        RECT 657.175 6.610 657.505 6.625 ;
        RECT 636.030 6.310 657.505 6.610 ;
        RECT 626.815 5.615 627.145 5.945 ;
        RECT 626.830 4.570 627.130 5.615 ;
        RECT 636.030 4.570 636.330 6.310 ;
        RECT 657.175 6.295 657.505 6.310 ;
        RECT 753.790 4.950 755.930 5.250 ;
        RECT 753.790 4.585 754.090 4.950 ;
        RECT 626.830 4.270 636.330 4.570 ;
        RECT 753.775 4.255 754.105 4.585 ;
        RECT 755.630 4.570 755.930 4.950 ;
        RECT 1156.750 4.585 1157.050 7.670 ;
        RECT 1168.710 4.585 1169.010 7.670 ;
        RECT 756.535 4.570 756.865 4.585 ;
        RECT 755.630 4.270 756.865 4.570 ;
        RECT 756.535 4.255 756.865 4.270 ;
        RECT 1156.735 4.255 1157.065 4.585 ;
        RECT 1168.695 4.255 1169.025 4.585 ;
        RECT 1261.615 3.890 1261.945 3.905 ;
        RECT 1262.535 3.890 1262.865 3.905 ;
        RECT 1261.615 3.590 1262.865 3.890 ;
        RECT 1261.615 3.575 1261.945 3.590 ;
        RECT 1262.535 3.575 1262.865 3.590 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 812.505 4.335 812.675 4.675 ;
        RECT 807.445 4.165 812.675 4.335 ;
        RECT 789.965 3.315 790.135 3.995 ;
        RECT 802.845 3.825 803.935 3.995 ;
        RECT 788.125 3.145 790.135 3.315 ;
        RECT 803.765 2.975 803.935 3.825 ;
        RECT 803.765 2.805 804.395 2.975 ;
        RECT 804.225 2.635 804.395 2.805 ;
        RECT 807.445 2.635 807.615 4.165 ;
        RECT 804.225 2.465 807.615 2.635 ;
      LAYER mcon ;
        RECT 812.505 4.505 812.675 4.675 ;
        RECT 789.965 3.825 790.135 3.995 ;
      LAYER met1 ;
        RECT 1790.850 8.400 1791.170 8.460 ;
        RECT 2069.150 8.400 2069.470 8.460 ;
        RECT 1790.850 8.260 2069.470 8.400 ;
        RECT 1790.850 8.200 1791.170 8.260 ;
        RECT 2069.150 8.200 2069.470 8.260 ;
        RECT 771.950 4.660 772.270 4.720 ;
        RECT 775.630 4.660 775.950 4.720 ;
        RECT 771.950 4.520 775.950 4.660 ;
        RECT 771.950 4.460 772.270 4.520 ;
        RECT 775.630 4.460 775.950 4.520 ;
        RECT 812.445 4.660 812.735 4.705 ;
        RECT 812.890 4.660 813.210 4.720 ;
        RECT 812.445 4.520 813.210 4.660 ;
        RECT 812.445 4.475 812.735 4.520 ;
        RECT 812.890 4.460 813.210 4.520 ;
        RECT 789.905 3.980 790.195 4.025 ;
        RECT 802.785 3.980 803.075 4.025 ;
        RECT 789.905 3.840 803.075 3.980 ;
        RECT 789.905 3.795 790.195 3.840 ;
        RECT 802.785 3.795 803.075 3.840 ;
        RECT 788.050 3.300 788.370 3.360 ;
        RECT 787.855 3.160 788.370 3.300 ;
        RECT 788.050 3.100 788.370 3.160 ;
      LAYER via ;
        RECT 1790.880 8.200 1791.140 8.460 ;
        RECT 2069.180 8.200 2069.440 8.460 ;
        RECT 771.980 4.460 772.240 4.720 ;
        RECT 775.660 4.460 775.920 4.720 ;
        RECT 812.920 4.460 813.180 4.720 ;
        RECT 788.080 3.100 788.340 3.360 ;
      LAYER met2 ;
        RECT 2070.950 8.570 2071.230 9.000 ;
        RECT 2069.240 8.490 2071.230 8.570 ;
        RECT 1790.880 8.170 1791.140 8.490 ;
        RECT 2069.180 8.430 2071.230 8.490 ;
        RECT 2069.180 8.170 2069.440 8.430 ;
        RECT 771.980 4.430 772.240 4.750 ;
        RECT 775.660 4.430 775.920 4.750 ;
        RECT 812.920 4.660 813.180 4.750 ;
        RECT 812.920 4.520 816.800 4.660 ;
        RECT 812.920 4.430 813.180 4.520 ;
        RECT 614.260 3.670 616.700 3.810 ;
        RECT 151.500 2.990 152.560 3.130 ;
        RECT 151.500 2.400 151.640 2.990 ;
        RECT 151.290 -4.800 151.850 2.400 ;
        RECT 152.420 1.885 152.560 2.990 ;
        RECT 614.260 2.450 614.400 3.670 ;
        RECT 613.340 2.310 614.400 2.450 ;
        RECT 613.340 1.885 613.480 2.310 ;
        RECT 616.560 1.885 616.700 3.670 ;
        RECT 772.040 3.640 772.180 4.430 ;
        RECT 768.360 3.500 772.180 3.640 ;
        RECT 768.360 2.450 768.500 3.500 ;
        RECT 775.720 3.130 775.860 4.430 ;
        RECT 788.080 3.245 788.340 3.390 ;
        RECT 785.770 3.130 786.050 3.245 ;
        RECT 775.720 2.990 786.050 3.130 ;
        RECT 785.770 2.875 786.050 2.990 ;
        RECT 788.070 2.875 788.350 3.245 ;
        RECT 765.600 2.310 768.500 2.450 ;
        RECT 765.600 1.885 765.740 2.310 ;
        RECT 816.660 1.885 816.800 4.520 ;
        RECT 1790.940 1.885 1791.080 8.170 ;
        RECT 2070.950 5.000 2071.230 8.430 ;
        RECT 152.350 1.515 152.630 1.885 ;
        RECT 325.310 1.770 325.590 1.885 ;
        RECT 326.690 1.770 326.970 1.885 ;
        RECT 325.310 1.630 326.970 1.770 ;
        RECT 325.310 1.515 325.590 1.630 ;
        RECT 326.690 1.515 326.970 1.630 ;
        RECT 366.710 1.770 366.990 1.885 ;
        RECT 366.710 1.630 368.300 1.770 ;
        RECT 366.710 1.515 366.990 1.630 ;
        RECT 368.160 1.260 368.300 1.630 ;
        RECT 369.010 1.515 369.290 1.885 ;
        RECT 462.390 1.770 462.670 1.885 ;
        RECT 463.310 1.770 463.590 1.885 ;
        RECT 462.390 1.630 463.590 1.770 ;
        RECT 462.390 1.515 462.670 1.630 ;
        RECT 463.310 1.515 463.590 1.630 ;
        RECT 613.270 1.515 613.550 1.885 ;
        RECT 616.490 1.515 616.770 1.885 ;
        RECT 765.530 1.515 765.810 1.885 ;
        RECT 816.590 1.515 816.870 1.885 ;
        RECT 1121.570 1.515 1121.850 1.885 ;
        RECT 1123.410 1.770 1123.690 1.885 ;
        RECT 1123.020 1.630 1123.690 1.770 ;
        RECT 369.080 1.260 369.220 1.515 ;
        RECT 368.160 1.120 369.220 1.260 ;
        RECT 1121.640 1.090 1121.780 1.515 ;
        RECT 1123.020 1.090 1123.160 1.630 ;
        RECT 1123.410 1.515 1123.690 1.630 ;
        RECT 1241.630 1.770 1241.910 1.885 ;
        RECT 1243.930 1.770 1244.210 1.885 ;
        RECT 1241.630 1.630 1244.210 1.770 ;
        RECT 1241.630 1.515 1241.910 1.630 ;
        RECT 1243.930 1.515 1244.210 1.630 ;
        RECT 1790.870 1.515 1791.150 1.885 ;
        RECT 1121.640 0.950 1123.160 1.090 ;
      LAYER via2 ;
        RECT 785.770 2.920 786.050 3.200 ;
        RECT 788.070 2.920 788.350 3.200 ;
        RECT 152.350 1.560 152.630 1.840 ;
        RECT 325.310 1.560 325.590 1.840 ;
        RECT 326.690 1.560 326.970 1.840 ;
        RECT 366.710 1.560 366.990 1.840 ;
        RECT 369.010 1.560 369.290 1.840 ;
        RECT 462.390 1.560 462.670 1.840 ;
        RECT 463.310 1.560 463.590 1.840 ;
        RECT 613.270 1.560 613.550 1.840 ;
        RECT 616.490 1.560 616.770 1.840 ;
        RECT 765.530 1.560 765.810 1.840 ;
        RECT 816.590 1.560 816.870 1.840 ;
        RECT 1121.570 1.560 1121.850 1.840 ;
        RECT 1123.410 1.560 1123.690 1.840 ;
        RECT 1241.630 1.560 1241.910 1.840 ;
        RECT 1243.930 1.560 1244.210 1.840 ;
        RECT 1790.870 1.560 1791.150 1.840 ;
      LAYER met3 ;
        RECT 785.745 3.210 786.075 3.225 ;
        RECT 788.045 3.210 788.375 3.225 ;
        RECT 785.745 2.910 788.375 3.210 ;
        RECT 785.745 2.895 786.075 2.910 ;
        RECT 788.045 2.895 788.375 2.910 ;
        RECT 152.325 1.850 152.655 1.865 ;
        RECT 325.285 1.850 325.615 1.865 ;
        RECT 152.325 1.550 325.615 1.850 ;
        RECT 152.325 1.535 152.655 1.550 ;
        RECT 325.285 1.535 325.615 1.550 ;
        RECT 326.665 1.850 326.995 1.865 ;
        RECT 366.685 1.850 367.015 1.865 ;
        RECT 326.665 1.550 367.015 1.850 ;
        RECT 326.665 1.535 326.995 1.550 ;
        RECT 366.685 1.535 367.015 1.550 ;
        RECT 368.985 1.850 369.315 1.865 ;
        RECT 462.365 1.850 462.695 1.865 ;
        RECT 368.985 1.550 462.695 1.850 ;
        RECT 368.985 1.535 369.315 1.550 ;
        RECT 462.365 1.535 462.695 1.550 ;
        RECT 463.285 1.850 463.615 1.865 ;
        RECT 613.245 1.850 613.575 1.865 ;
        RECT 463.285 1.550 613.575 1.850 ;
        RECT 463.285 1.535 463.615 1.550 ;
        RECT 613.245 1.535 613.575 1.550 ;
        RECT 616.465 1.850 616.795 1.865 ;
        RECT 765.505 1.850 765.835 1.865 ;
        RECT 616.465 1.550 765.835 1.850 ;
        RECT 616.465 1.535 616.795 1.550 ;
        RECT 765.505 1.535 765.835 1.550 ;
        RECT 816.565 1.850 816.895 1.865 ;
        RECT 1121.545 1.850 1121.875 1.865 ;
        RECT 816.565 1.550 1121.875 1.850 ;
        RECT 816.565 1.535 816.895 1.550 ;
        RECT 1121.545 1.535 1121.875 1.550 ;
        RECT 1123.385 1.850 1123.715 1.865 ;
        RECT 1241.605 1.850 1241.935 1.865 ;
        RECT 1123.385 1.550 1241.935 1.850 ;
        RECT 1123.385 1.535 1123.715 1.550 ;
        RECT 1241.605 1.535 1241.935 1.550 ;
        RECT 1243.905 1.850 1244.235 1.865 ;
        RECT 1453.870 1.850 1454.250 1.860 ;
        RECT 1243.905 1.550 1454.250 1.850 ;
        RECT 1243.905 1.535 1244.235 1.550 ;
        RECT 1453.870 1.540 1454.250 1.550 ;
        RECT 1455.710 1.850 1456.090 1.860 ;
        RECT 1790.845 1.850 1791.175 1.865 ;
        RECT 1455.710 1.550 1791.175 1.850 ;
        RECT 1455.710 1.540 1456.090 1.550 ;
        RECT 1790.845 1.535 1791.175 1.550 ;
      LAYER via3 ;
        RECT 1453.900 1.540 1454.220 1.860 ;
        RECT 1455.740 1.540 1456.060 1.860 ;
      LAYER met4 ;
        RECT 1453.895 1.850 1454.225 1.865 ;
        RECT 1455.735 1.850 1456.065 1.865 ;
        RECT 1453.895 1.550 1456.065 1.850 ;
        RECT 1453.895 1.535 1454.225 1.550 ;
        RECT 1455.735 1.535 1456.065 1.550 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 8.885 1141.805 9.055 1210.995 ;
        RECT 8.885 881.025 9.055 892.075 ;
        RECT 8.885 623.645 9.055 667.335 ;
        RECT 7.965 91.885 8.135 148.495 ;
        RECT 5.205 8.245 5.375 51.935 ;
      LAYER mcon ;
        RECT 8.885 1210.825 9.055 1210.995 ;
        RECT 8.885 891.905 9.055 892.075 ;
        RECT 8.885 667.165 9.055 667.335 ;
        RECT 7.965 148.325 8.135 148.495 ;
        RECT 5.205 51.765 5.375 51.935 ;
      LAYER met1 ;
        RECT 6.970 1291.220 7.290 1291.280 ;
        RECT 8.810 1291.220 9.130 1291.280 ;
        RECT 6.970 1291.080 9.130 1291.220 ;
        RECT 6.970 1291.020 7.290 1291.080 ;
        RECT 8.810 1291.020 9.130 1291.080 ;
        RECT 8.810 1210.980 9.130 1211.040 ;
        RECT 8.615 1210.840 9.130 1210.980 ;
        RECT 8.810 1210.780 9.130 1210.840 ;
        RECT 8.810 1141.960 9.130 1142.020 ;
        RECT 8.615 1141.820 9.130 1141.960 ;
        RECT 8.810 1141.760 9.130 1141.820 ;
        RECT 8.810 892.060 9.130 892.120 ;
        RECT 8.615 891.920 9.130 892.060 ;
        RECT 8.810 891.860 9.130 891.920 ;
        RECT 8.810 881.180 9.130 881.240 ;
        RECT 8.615 881.040 9.130 881.180 ;
        RECT 8.810 880.980 9.130 881.040 ;
        RECT 8.810 667.320 9.130 667.380 ;
        RECT 8.615 667.180 9.130 667.320 ;
        RECT 8.810 667.120 9.130 667.180 ;
        RECT 8.810 623.800 9.130 623.860 ;
        RECT 8.810 623.660 9.325 623.800 ;
        RECT 8.810 623.600 9.130 623.660 ;
        RECT 7.905 148.480 8.195 148.525 ;
        RECT 8.810 148.480 9.130 148.540 ;
        RECT 7.905 148.340 9.130 148.480 ;
        RECT 7.905 148.295 8.195 148.340 ;
        RECT 8.810 148.280 9.130 148.340 ;
        RECT 5.130 92.040 5.450 92.100 ;
        RECT 7.905 92.040 8.195 92.085 ;
        RECT 5.130 91.900 8.195 92.040 ;
        RECT 5.130 91.840 5.450 91.900 ;
        RECT 7.905 91.855 8.195 91.900 ;
        RECT 5.130 51.920 5.450 51.980 ;
        RECT 4.935 51.780 5.450 51.920 ;
        RECT 5.130 51.720 5.450 51.780 ;
        RECT 5.145 8.400 5.435 8.445 ;
        RECT 7.430 8.400 7.750 8.460 ;
        RECT 5.145 8.260 7.750 8.400 ;
        RECT 5.145 8.215 5.435 8.260 ;
        RECT 7.430 8.200 7.750 8.260 ;
      LAYER via ;
        RECT 7.000 1291.020 7.260 1291.280 ;
        RECT 8.840 1291.020 9.100 1291.280 ;
        RECT 8.840 1210.780 9.100 1211.040 ;
        RECT 8.840 1141.760 9.100 1142.020 ;
        RECT 8.840 891.860 9.100 892.120 ;
        RECT 8.840 880.980 9.100 881.240 ;
        RECT 8.840 667.120 9.100 667.380 ;
        RECT 8.840 623.600 9.100 623.860 ;
        RECT 8.840 148.280 9.100 148.540 ;
        RECT 5.160 91.840 5.420 92.100 ;
        RECT 5.160 51.720 5.420 51.980 ;
        RECT 7.460 8.200 7.720 8.460 ;
      LAYER met2 ;
        RECT 6.990 1305.075 7.270 1305.445 ;
        RECT 7.060 1291.310 7.200 1305.075 ;
        RECT 7.000 1290.990 7.260 1291.310 ;
        RECT 8.840 1290.990 9.100 1291.310 ;
        RECT 8.900 1211.070 9.040 1290.990 ;
        RECT 8.840 1210.750 9.100 1211.070 ;
        RECT 8.840 1141.730 9.100 1142.050 ;
        RECT 8.900 892.150 9.040 1141.730 ;
        RECT 8.840 891.830 9.100 892.150 ;
        RECT 8.840 880.950 9.100 881.270 ;
        RECT 8.900 667.410 9.040 880.950 ;
        RECT 8.840 667.090 9.100 667.410 ;
        RECT 8.840 623.570 9.100 623.890 ;
        RECT 8.900 148.570 9.040 623.570 ;
        RECT 8.840 148.250 9.100 148.570 ;
        RECT 5.160 91.810 5.420 92.130 ;
        RECT 5.220 52.010 5.360 91.810 ;
        RECT 5.160 51.690 5.420 52.010 ;
        RECT 7.460 8.170 7.720 8.490 ;
        RECT 30.450 8.315 30.730 8.685 ;
        RECT 72.310 8.315 72.590 8.685 ;
        RECT 186.850 8.315 187.130 8.685 ;
        RECT 7.520 7.325 7.660 8.170 ;
        RECT 30.520 7.325 30.660 8.315 ;
        RECT 72.380 7.325 72.520 8.315 ;
        RECT 7.450 6.955 7.730 7.325 ;
        RECT 30.450 6.955 30.730 7.325 ;
        RECT 72.310 6.955 72.590 7.325 ;
        RECT 186.920 2.400 187.060 8.315 ;
        RECT 186.710 -4.800 187.270 2.400 ;
      LAYER via2 ;
        RECT 6.990 1305.120 7.270 1305.400 ;
        RECT 30.450 8.360 30.730 8.640 ;
        RECT 72.310 8.360 72.590 8.640 ;
        RECT 186.850 8.360 187.130 8.640 ;
        RECT 7.450 7.000 7.730 7.280 ;
        RECT 30.450 7.000 30.730 7.280 ;
        RECT 72.310 7.000 72.590 7.280 ;
      LAYER met3 ;
        RECT 5.000 1307.920 9.000 1308.520 ;
        RECT 6.750 1305.425 7.050 1307.920 ;
        RECT 6.750 1305.110 7.295 1305.425 ;
        RECT 6.965 1305.095 7.295 1305.110 ;
        RECT 14.990 8.650 15.370 8.660 ;
        RECT 30.425 8.650 30.755 8.665 ;
        RECT 14.990 8.350 30.755 8.650 ;
        RECT 14.990 8.340 15.370 8.350 ;
        RECT 30.425 8.335 30.755 8.350 ;
        RECT 72.285 8.650 72.615 8.665 ;
        RECT 186.825 8.650 187.155 8.665 ;
        RECT 72.285 8.350 187.155 8.650 ;
        RECT 72.285 8.335 72.615 8.350 ;
        RECT 186.825 8.335 187.155 8.350 ;
        RECT 7.425 7.290 7.755 7.305 ;
        RECT 14.990 7.290 15.370 7.300 ;
        RECT 7.425 6.990 15.370 7.290 ;
        RECT 7.425 6.975 7.755 6.990 ;
        RECT 14.990 6.980 15.370 6.990 ;
        RECT 30.425 7.290 30.755 7.305 ;
        RECT 72.285 7.290 72.615 7.305 ;
        RECT 30.425 6.990 72.615 7.290 ;
        RECT 30.425 6.975 30.755 6.990 ;
        RECT 72.285 6.975 72.615 6.990 ;
      LAYER via3 ;
        RECT 15.020 8.340 15.340 8.660 ;
        RECT 15.020 6.980 15.340 7.300 ;
      LAYER met4 ;
        RECT 15.015 8.335 15.345 8.665 ;
        RECT 15.030 7.305 15.330 8.335 ;
        RECT 15.015 6.975 15.345 7.305 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 4.285 1259.105 4.455 1307.895 ;
        RECT 6.585 989.995 6.755 1049.835 ;
        RECT 6.585 989.825 7.215 989.995 ;
        RECT 7.045 969.765 7.215 989.825 ;
        RECT 7.045 881.705 7.215 948.855 ;
        RECT 3.365 730.745 3.535 769.675 ;
        RECT 6.125 769.505 6.295 838.355 ;
        RECT 6.585 535.925 6.755 730.915 ;
        RECT 7.505 404.005 7.675 436.815 ;
        RECT 8.425 436.645 8.595 491.555 ;
        RECT 6.125 313.565 6.295 348.075 ;
        RECT 8.425 347.905 8.595 404.175 ;
        RECT 7.045 215.305 7.215 227.715 ;
        RECT 7.965 227.545 8.135 313.735 ;
        RECT 9.345 148.495 9.515 196.775 ;
        RECT 8.885 148.325 9.515 148.495 ;
        RECT 8.885 100.215 9.055 148.325 ;
        RECT 8.885 100.045 9.515 100.215 ;
        RECT 9.345 18.445 9.515 100.045 ;
        RECT 134.925 8.245 135.095 9.095 ;
      LAYER mcon ;
        RECT 4.285 1307.725 4.455 1307.895 ;
        RECT 6.585 1049.665 6.755 1049.835 ;
        RECT 7.045 948.685 7.215 948.855 ;
        RECT 6.125 838.185 6.295 838.355 ;
        RECT 3.365 769.505 3.535 769.675 ;
        RECT 6.585 730.745 6.755 730.915 ;
        RECT 8.425 491.385 8.595 491.555 ;
        RECT 7.505 436.645 7.675 436.815 ;
        RECT 8.425 404.005 8.595 404.175 ;
        RECT 6.125 347.905 6.295 348.075 ;
        RECT 7.965 313.565 8.135 313.735 ;
        RECT 7.045 227.545 7.215 227.715 ;
        RECT 9.345 196.605 9.515 196.775 ;
        RECT 134.925 8.925 135.095 9.095 ;
      LAYER met1 ;
        RECT 4.225 1307.880 4.515 1307.925 ;
        RECT 6.970 1307.880 7.290 1307.940 ;
        RECT 4.225 1307.740 7.290 1307.880 ;
        RECT 4.225 1307.695 4.515 1307.740 ;
        RECT 6.970 1307.680 7.290 1307.740 ;
        RECT 4.210 1259.260 4.530 1259.320 ;
        RECT 4.015 1259.120 4.530 1259.260 ;
        RECT 4.210 1259.060 4.530 1259.120 ;
        RECT 4.210 1049.820 4.530 1049.880 ;
        RECT 6.525 1049.820 6.815 1049.865 ;
        RECT 4.210 1049.680 6.815 1049.820 ;
        RECT 4.210 1049.620 4.530 1049.680 ;
        RECT 6.525 1049.635 6.815 1049.680 ;
        RECT 6.985 969.920 7.275 969.965 ;
        RECT 9.730 969.920 10.050 969.980 ;
        RECT 6.985 969.780 10.050 969.920 ;
        RECT 6.985 969.735 7.275 969.780 ;
        RECT 9.730 969.720 10.050 969.780 ;
        RECT 6.985 948.840 7.275 948.885 ;
        RECT 9.730 948.840 10.050 948.900 ;
        RECT 6.985 948.700 10.050 948.840 ;
        RECT 6.985 948.655 7.275 948.700 ;
        RECT 9.730 948.640 10.050 948.700 ;
        RECT 6.985 881.860 7.275 881.905 ;
        RECT 9.730 881.860 10.050 881.920 ;
        RECT 6.985 881.720 10.050 881.860 ;
        RECT 6.985 881.675 7.275 881.720 ;
        RECT 9.730 881.660 10.050 881.720 ;
        RECT 6.065 838.340 6.355 838.385 ;
        RECT 9.730 838.340 10.050 838.400 ;
        RECT 6.065 838.200 10.050 838.340 ;
        RECT 6.065 838.155 6.355 838.200 ;
        RECT 9.730 838.140 10.050 838.200 ;
        RECT 3.305 769.660 3.595 769.705 ;
        RECT 6.065 769.660 6.355 769.705 ;
        RECT 3.305 769.520 6.355 769.660 ;
        RECT 3.305 769.475 3.595 769.520 ;
        RECT 6.065 769.475 6.355 769.520 ;
        RECT 3.305 730.900 3.595 730.945 ;
        RECT 6.525 730.900 6.815 730.945 ;
        RECT 3.305 730.760 6.815 730.900 ;
        RECT 3.305 730.715 3.595 730.760 ;
        RECT 6.525 730.715 6.815 730.760 ;
        RECT 6.525 536.080 6.815 536.125 ;
        RECT 9.730 536.080 10.050 536.140 ;
        RECT 6.525 535.940 10.050 536.080 ;
        RECT 6.525 535.895 6.815 535.940 ;
        RECT 9.730 535.880 10.050 535.940 ;
        RECT 8.365 491.540 8.655 491.585 ;
        RECT 9.730 491.540 10.050 491.600 ;
        RECT 8.365 491.400 10.050 491.540 ;
        RECT 8.365 491.355 8.655 491.400 ;
        RECT 9.730 491.340 10.050 491.400 ;
        RECT 7.445 436.800 7.735 436.845 ;
        RECT 8.365 436.800 8.655 436.845 ;
        RECT 7.445 436.660 8.655 436.800 ;
        RECT 7.445 436.615 7.735 436.660 ;
        RECT 8.365 436.615 8.655 436.660 ;
        RECT 7.445 404.160 7.735 404.205 ;
        RECT 8.365 404.160 8.655 404.205 ;
        RECT 7.445 404.020 8.655 404.160 ;
        RECT 7.445 403.975 7.735 404.020 ;
        RECT 8.365 403.975 8.655 404.020 ;
        RECT 6.065 348.060 6.355 348.105 ;
        RECT 8.365 348.060 8.655 348.105 ;
        RECT 6.065 347.920 8.655 348.060 ;
        RECT 6.065 347.875 6.355 347.920 ;
        RECT 8.365 347.875 8.655 347.920 ;
        RECT 6.065 313.720 6.355 313.765 ;
        RECT 7.905 313.720 8.195 313.765 ;
        RECT 6.065 313.580 8.195 313.720 ;
        RECT 6.065 313.535 6.355 313.580 ;
        RECT 7.905 313.535 8.195 313.580 ;
        RECT 6.985 227.700 7.275 227.745 ;
        RECT 7.905 227.700 8.195 227.745 ;
        RECT 6.985 227.560 8.195 227.700 ;
        RECT 6.985 227.515 7.275 227.560 ;
        RECT 7.905 227.515 8.195 227.560 ;
        RECT 6.985 215.460 7.275 215.505 ;
        RECT 9.730 215.460 10.050 215.520 ;
        RECT 6.985 215.320 10.050 215.460 ;
        RECT 6.985 215.275 7.275 215.320 ;
        RECT 9.730 215.260 10.050 215.320 ;
        RECT 9.285 196.760 9.575 196.805 ;
        RECT 9.730 196.760 10.050 196.820 ;
        RECT 9.285 196.620 10.050 196.760 ;
        RECT 9.285 196.575 9.575 196.620 ;
        RECT 9.730 196.560 10.050 196.620 ;
        RECT 9.270 18.600 9.590 18.660 ;
        RECT 9.075 18.460 9.590 18.600 ;
        RECT 9.270 18.400 9.590 18.460 ;
        RECT 134.865 9.080 135.155 9.125 ;
        RECT 134.865 8.940 176.020 9.080 ;
        RECT 134.865 8.895 135.155 8.940 ;
        RECT 132.090 8.740 132.410 8.800 ;
        RECT 132.090 8.600 133.700 8.740 ;
        RECT 132.090 8.540 132.410 8.600 ;
        RECT 133.560 8.400 133.700 8.600 ;
        RECT 134.865 8.400 135.155 8.445 ;
        RECT 133.560 8.260 135.155 8.400 ;
        RECT 175.880 8.400 176.020 8.940 ;
        RECT 188.670 8.400 188.990 8.460 ;
        RECT 175.880 8.260 188.990 8.400 ;
        RECT 134.865 8.215 135.155 8.260 ;
        RECT 188.670 8.200 188.990 8.260 ;
      LAYER via ;
        RECT 7.000 1307.680 7.260 1307.940 ;
        RECT 4.240 1259.060 4.500 1259.320 ;
        RECT 4.240 1049.620 4.500 1049.880 ;
        RECT 9.760 969.720 10.020 969.980 ;
        RECT 9.760 948.640 10.020 948.900 ;
        RECT 9.760 881.660 10.020 881.920 ;
        RECT 9.760 838.140 10.020 838.400 ;
        RECT 9.760 535.880 10.020 536.140 ;
        RECT 9.760 491.340 10.020 491.600 ;
        RECT 9.760 215.260 10.020 215.520 ;
        RECT 9.760 196.560 10.020 196.820 ;
        RECT 9.300 18.400 9.560 18.660 ;
        RECT 132.120 8.540 132.380 8.800 ;
        RECT 188.700 8.200 188.960 8.460 ;
      LAYER met2 ;
        RECT 6.990 1418.635 7.270 1419.005 ;
        RECT 7.060 1307.970 7.200 1418.635 ;
        RECT 7.000 1307.650 7.260 1307.970 ;
        RECT 4.240 1259.030 4.500 1259.350 ;
        RECT 4.300 1049.910 4.440 1259.030 ;
        RECT 4.240 1049.590 4.500 1049.910 ;
        RECT 9.760 969.920 10.020 970.010 ;
        RECT 9.760 969.780 10.420 969.920 ;
        RECT 9.760 969.690 10.020 969.780 ;
        RECT 10.280 949.690 10.420 969.780 ;
        RECT 9.820 949.550 10.420 949.690 ;
        RECT 9.820 948.930 9.960 949.550 ;
        RECT 9.760 948.610 10.020 948.930 ;
        RECT 9.760 881.860 10.020 881.950 ;
        RECT 9.760 881.720 10.880 881.860 ;
        RECT 9.760 881.630 10.020 881.720 ;
        RECT 10.740 881.180 10.880 881.720 ;
        RECT 10.740 881.040 11.340 881.180 ;
        RECT 9.760 838.340 10.020 838.430 ;
        RECT 11.200 838.340 11.340 881.040 ;
        RECT 9.760 838.200 11.340 838.340 ;
        RECT 9.760 838.110 10.020 838.200 ;
        RECT 9.760 536.080 10.020 536.170 ;
        RECT 9.760 535.940 10.880 536.080 ;
        RECT 9.760 535.850 10.020 535.940 ;
        RECT 10.740 517.890 10.880 535.940 ;
        RECT 10.280 517.750 10.880 517.890 ;
        RECT 9.760 491.540 10.020 491.630 ;
        RECT 10.280 491.540 10.420 517.750 ;
        RECT 9.760 491.400 10.420 491.540 ;
        RECT 9.760 491.310 10.020 491.400 ;
        RECT 9.760 215.230 10.020 215.550 ;
        RECT 9.820 214.610 9.960 215.230 ;
        RECT 9.820 214.470 10.880 214.610 ;
        RECT 10.740 196.930 10.880 214.470 ;
        RECT 9.820 196.850 10.880 196.930 ;
        RECT 9.760 196.790 10.880 196.850 ;
        RECT 9.760 196.530 10.020 196.790 ;
        RECT 9.300 18.370 9.560 18.690 ;
        RECT 9.360 8.005 9.500 18.370 ;
        RECT 132.120 8.510 132.380 8.830 ;
        RECT 132.180 8.005 132.320 8.510 ;
        RECT 188.690 8.315 188.970 8.685 ;
        RECT 204.790 8.315 205.070 8.685 ;
        RECT 188.700 8.170 188.960 8.315 ;
        RECT 9.290 7.635 9.570 8.005 ;
        RECT 132.110 7.635 132.390 8.005 ;
        RECT 204.860 2.400 205.000 8.315 ;
        RECT 204.650 -4.800 205.210 2.400 ;
      LAYER via2 ;
        RECT 6.990 1418.680 7.270 1418.960 ;
        RECT 188.690 8.360 188.970 8.640 ;
        RECT 204.790 8.360 205.070 8.640 ;
        RECT 9.290 7.680 9.570 7.960 ;
        RECT 132.110 7.680 132.390 7.960 ;
      LAYER met3 ;
        RECT 5.000 1421.480 9.000 1422.080 ;
        RECT 6.750 1418.985 7.050 1421.480 ;
        RECT 6.750 1418.670 7.295 1418.985 ;
        RECT 6.965 1418.655 7.295 1418.670 ;
        RECT 188.665 8.650 188.995 8.665 ;
        RECT 204.765 8.650 205.095 8.665 ;
        RECT 188.665 8.350 205.095 8.650 ;
        RECT 188.665 8.335 188.995 8.350 ;
        RECT 204.765 8.335 205.095 8.350 ;
        RECT 9.265 7.970 9.595 7.985 ;
        RECT 132.085 7.970 132.415 7.985 ;
        RECT 9.265 7.670 132.415 7.970 ;
        RECT 9.265 7.655 9.595 7.670 ;
        RECT 132.085 7.655 132.415 7.670 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 58.565 3398.385 58.735 3399.235 ;
        RECT 82.945 3398.385 83.115 3399.235 ;
        RECT 155.165 3398.385 155.335 3399.235 ;
        RECT 179.545 3398.385 179.715 3399.235 ;
        RECT 251.765 3398.385 251.935 3399.235 ;
        RECT 276.145 3398.385 276.315 3399.235 ;
        RECT 348.365 3398.385 348.535 3399.235 ;
        RECT 372.745 3398.385 372.915 3399.235 ;
        RECT 444.965 3398.385 445.135 3399.235 ;
        RECT 469.345 3398.385 469.515 3399.235 ;
        RECT 541.565 3398.385 541.735 3399.235 ;
        RECT 565.945 3398.385 566.115 3399.235 ;
        RECT 638.165 3398.385 638.335 3399.235 ;
        RECT 662.545 3398.385 662.715 3399.235 ;
        RECT 734.765 3398.385 734.935 3399.235 ;
        RECT 759.145 3398.385 759.315 3399.235 ;
        RECT 831.365 3398.385 831.535 3399.235 ;
        RECT 855.745 3398.385 855.915 3399.235 ;
        RECT 927.965 3398.385 928.135 3399.235 ;
        RECT 952.345 3398.385 952.515 3399.235 ;
        RECT 1024.565 3398.385 1024.735 3399.235 ;
        RECT 1048.945 3398.385 1049.115 3399.235 ;
        RECT 1110.125 3399.065 1110.755 3399.235 ;
        RECT 1110.585 3398.725 1110.755 3399.065 ;
        RECT 1111.045 3397.705 1111.215 3398.555 ;
        RECT 1158.885 3397.705 1159.055 3398.895 ;
        RECT 1159.805 3398.725 1159.975 3401.955 ;
        RECT 9.805 3196.425 9.975 3240.455 ;
        RECT 9.345 2984.945 9.515 3011.975 ;
        RECT 9.805 2832.795 9.975 2901.135 ;
        RECT 9.345 2832.625 9.975 2832.795 ;
        RECT 9.345 2805.425 9.515 2832.625 ;
        RECT 9.345 2611.625 9.515 2638.655 ;
        RECT 9.345 2522.205 9.515 2549.575 ;
        RECT 9.345 2337.925 9.515 2370.395 ;
        RECT 7.965 2245.105 8.135 2253.775 ;
        RECT 8.885 2207.025 9.055 2211.615 ;
        RECT 7.965 1895.585 8.135 1907.315 ;
        RECT 9.805 1907.145 9.975 1935.535 ;
        RECT 8.885 1791.715 9.055 1851.215 ;
        RECT 8.425 1791.545 9.055 1791.715 ;
        RECT 8.425 1729.155 8.595 1791.545 ;
        RECT 7.965 1728.985 8.595 1729.155 ;
        RECT 7.965 1631.745 8.135 1728.985 ;
        RECT 8.425 1557.625 8.595 1569.695 ;
        RECT 9.345 1569.525 9.515 1631.915 ;
        RECT 8.885 1516.145 9.055 1527.535 ;
        RECT 8.425 1416.695 8.595 1479.255 ;
        RECT 8.425 1416.525 9.055 1416.695 ;
        RECT 8.885 1348.865 9.055 1416.525 ;
        RECT 7.965 1112.905 8.135 1210.655 ;
        RECT 9.345 1210.485 9.515 1332.375 ;
        RECT 9.345 1028.925 9.515 1113.075 ;
        RECT 8.885 976.395 9.055 1028.415 ;
        RECT 8.885 976.225 9.975 976.395 ;
        RECT 2.445 851.445 2.615 896.155 ;
        RECT 9.805 895.985 9.975 976.225 ;
        RECT 5.665 769.335 5.835 830.875 ;
        RECT 5.665 769.165 6.755 769.335 ;
        RECT 4.285 703.715 4.455 731.595 ;
        RECT 6.585 731.425 6.755 769.165 ;
        RECT 4.285 703.545 4.915 703.715 ;
        RECT 4.745 695.385 4.915 703.545 ;
        RECT 7.505 582.165 7.675 630.615 ;
        RECT 6.125 403.325 6.295 443.955 ;
        RECT 9.805 443.785 9.975 490.875 ;
        RECT 7.505 334.645 7.675 403.495 ;
        RECT 25.445 2.295 25.615 2.635 ;
        RECT 25.445 2.125 27.455 2.295 ;
        RECT 51.205 1.615 51.375 2.295 ;
        RECT 51.205 1.445 53.215 1.615 ;
        RECT 53.045 0.425 53.215 1.445 ;
      LAYER mcon ;
        RECT 1159.805 3401.785 1159.975 3401.955 ;
        RECT 58.565 3399.065 58.735 3399.235 ;
        RECT 82.945 3399.065 83.115 3399.235 ;
        RECT 155.165 3399.065 155.335 3399.235 ;
        RECT 179.545 3399.065 179.715 3399.235 ;
        RECT 251.765 3399.065 251.935 3399.235 ;
        RECT 276.145 3399.065 276.315 3399.235 ;
        RECT 348.365 3399.065 348.535 3399.235 ;
        RECT 372.745 3399.065 372.915 3399.235 ;
        RECT 444.965 3399.065 445.135 3399.235 ;
        RECT 469.345 3399.065 469.515 3399.235 ;
        RECT 541.565 3399.065 541.735 3399.235 ;
        RECT 565.945 3399.065 566.115 3399.235 ;
        RECT 638.165 3399.065 638.335 3399.235 ;
        RECT 662.545 3399.065 662.715 3399.235 ;
        RECT 734.765 3399.065 734.935 3399.235 ;
        RECT 759.145 3399.065 759.315 3399.235 ;
        RECT 831.365 3399.065 831.535 3399.235 ;
        RECT 855.745 3399.065 855.915 3399.235 ;
        RECT 927.965 3399.065 928.135 3399.235 ;
        RECT 952.345 3399.065 952.515 3399.235 ;
        RECT 1024.565 3399.065 1024.735 3399.235 ;
        RECT 1048.945 3399.065 1049.115 3399.235 ;
        RECT 1158.885 3398.725 1159.055 3398.895 ;
        RECT 1111.045 3398.385 1111.215 3398.555 ;
        RECT 9.805 3240.285 9.975 3240.455 ;
        RECT 9.345 3011.805 9.515 3011.975 ;
        RECT 9.805 2900.965 9.975 2901.135 ;
        RECT 9.345 2638.485 9.515 2638.655 ;
        RECT 9.345 2549.405 9.515 2549.575 ;
        RECT 9.345 2370.225 9.515 2370.395 ;
        RECT 7.965 2253.605 8.135 2253.775 ;
        RECT 8.885 2211.445 9.055 2211.615 ;
        RECT 9.805 1935.365 9.975 1935.535 ;
        RECT 7.965 1907.145 8.135 1907.315 ;
        RECT 8.885 1851.045 9.055 1851.215 ;
        RECT 9.345 1631.745 9.515 1631.915 ;
        RECT 8.425 1569.525 8.595 1569.695 ;
        RECT 8.885 1527.365 9.055 1527.535 ;
        RECT 8.425 1479.085 8.595 1479.255 ;
        RECT 9.345 1332.205 9.515 1332.375 ;
        RECT 7.965 1210.485 8.135 1210.655 ;
        RECT 9.345 1112.905 9.515 1113.075 ;
        RECT 8.885 1028.245 9.055 1028.415 ;
        RECT 2.445 895.985 2.615 896.155 ;
        RECT 5.665 830.705 5.835 830.875 ;
        RECT 4.285 731.425 4.455 731.595 ;
        RECT 7.505 630.445 7.675 630.615 ;
        RECT 9.805 490.705 9.975 490.875 ;
        RECT 6.125 443.785 6.295 443.955 ;
        RECT 7.505 403.325 7.675 403.495 ;
        RECT 25.445 2.465 25.615 2.635 ;
        RECT 27.285 2.125 27.455 2.295 ;
        RECT 51.205 2.125 51.375 2.295 ;
      LAYER met1 ;
        RECT 1159.745 3401.940 1160.035 3401.985 ;
        RECT 1231.030 3401.940 1231.350 3402.000 ;
        RECT 1159.745 3401.800 1231.350 3401.940 ;
        RECT 1159.745 3401.755 1160.035 3401.800 ;
        RECT 1231.030 3401.740 1231.350 3401.800 ;
        RECT 9.730 3399.220 10.050 3399.280 ;
        RECT 58.505 3399.220 58.795 3399.265 ;
        RECT 9.730 3399.080 58.795 3399.220 ;
        RECT 9.730 3399.020 10.050 3399.080 ;
        RECT 58.505 3399.035 58.795 3399.080 ;
        RECT 82.885 3399.220 83.175 3399.265 ;
        RECT 155.105 3399.220 155.395 3399.265 ;
        RECT 82.885 3399.080 155.395 3399.220 ;
        RECT 82.885 3399.035 83.175 3399.080 ;
        RECT 155.105 3399.035 155.395 3399.080 ;
        RECT 179.485 3399.220 179.775 3399.265 ;
        RECT 251.705 3399.220 251.995 3399.265 ;
        RECT 179.485 3399.080 251.995 3399.220 ;
        RECT 179.485 3399.035 179.775 3399.080 ;
        RECT 251.705 3399.035 251.995 3399.080 ;
        RECT 276.085 3399.220 276.375 3399.265 ;
        RECT 348.305 3399.220 348.595 3399.265 ;
        RECT 276.085 3399.080 348.595 3399.220 ;
        RECT 276.085 3399.035 276.375 3399.080 ;
        RECT 348.305 3399.035 348.595 3399.080 ;
        RECT 372.685 3399.220 372.975 3399.265 ;
        RECT 444.905 3399.220 445.195 3399.265 ;
        RECT 372.685 3399.080 445.195 3399.220 ;
        RECT 372.685 3399.035 372.975 3399.080 ;
        RECT 444.905 3399.035 445.195 3399.080 ;
        RECT 469.285 3399.220 469.575 3399.265 ;
        RECT 541.505 3399.220 541.795 3399.265 ;
        RECT 469.285 3399.080 541.795 3399.220 ;
        RECT 469.285 3399.035 469.575 3399.080 ;
        RECT 541.505 3399.035 541.795 3399.080 ;
        RECT 565.885 3399.220 566.175 3399.265 ;
        RECT 638.105 3399.220 638.395 3399.265 ;
        RECT 565.885 3399.080 638.395 3399.220 ;
        RECT 565.885 3399.035 566.175 3399.080 ;
        RECT 638.105 3399.035 638.395 3399.080 ;
        RECT 662.485 3399.220 662.775 3399.265 ;
        RECT 734.705 3399.220 734.995 3399.265 ;
        RECT 662.485 3399.080 734.995 3399.220 ;
        RECT 662.485 3399.035 662.775 3399.080 ;
        RECT 734.705 3399.035 734.995 3399.080 ;
        RECT 759.085 3399.220 759.375 3399.265 ;
        RECT 831.305 3399.220 831.595 3399.265 ;
        RECT 759.085 3399.080 831.595 3399.220 ;
        RECT 759.085 3399.035 759.375 3399.080 ;
        RECT 831.305 3399.035 831.595 3399.080 ;
        RECT 855.685 3399.220 855.975 3399.265 ;
        RECT 927.905 3399.220 928.195 3399.265 ;
        RECT 855.685 3399.080 928.195 3399.220 ;
        RECT 855.685 3399.035 855.975 3399.080 ;
        RECT 927.905 3399.035 928.195 3399.080 ;
        RECT 952.285 3399.220 952.575 3399.265 ;
        RECT 1024.505 3399.220 1024.795 3399.265 ;
        RECT 952.285 3399.080 1024.795 3399.220 ;
        RECT 952.285 3399.035 952.575 3399.080 ;
        RECT 1024.505 3399.035 1024.795 3399.080 ;
        RECT 1048.885 3399.220 1049.175 3399.265 ;
        RECT 1110.065 3399.220 1110.355 3399.265 ;
        RECT 1048.885 3399.080 1110.355 3399.220 ;
        RECT 1048.885 3399.035 1049.175 3399.080 ;
        RECT 1110.065 3399.035 1110.355 3399.080 ;
        RECT 1110.525 3398.695 1110.815 3398.925 ;
        RECT 1158.825 3398.880 1159.115 3398.925 ;
        RECT 1159.745 3398.880 1160.035 3398.925 ;
        RECT 1158.825 3398.740 1160.035 3398.880 ;
        RECT 1158.825 3398.695 1159.115 3398.740 ;
        RECT 1159.745 3398.695 1160.035 3398.740 ;
        RECT 58.505 3398.540 58.795 3398.585 ;
        RECT 82.885 3398.540 83.175 3398.585 ;
        RECT 58.505 3398.400 83.175 3398.540 ;
        RECT 58.505 3398.355 58.795 3398.400 ;
        RECT 82.885 3398.355 83.175 3398.400 ;
        RECT 155.105 3398.540 155.395 3398.585 ;
        RECT 179.485 3398.540 179.775 3398.585 ;
        RECT 155.105 3398.400 179.775 3398.540 ;
        RECT 155.105 3398.355 155.395 3398.400 ;
        RECT 179.485 3398.355 179.775 3398.400 ;
        RECT 251.705 3398.540 251.995 3398.585 ;
        RECT 276.085 3398.540 276.375 3398.585 ;
        RECT 251.705 3398.400 276.375 3398.540 ;
        RECT 251.705 3398.355 251.995 3398.400 ;
        RECT 276.085 3398.355 276.375 3398.400 ;
        RECT 348.305 3398.540 348.595 3398.585 ;
        RECT 372.685 3398.540 372.975 3398.585 ;
        RECT 348.305 3398.400 372.975 3398.540 ;
        RECT 348.305 3398.355 348.595 3398.400 ;
        RECT 372.685 3398.355 372.975 3398.400 ;
        RECT 444.905 3398.540 445.195 3398.585 ;
        RECT 469.285 3398.540 469.575 3398.585 ;
        RECT 444.905 3398.400 469.575 3398.540 ;
        RECT 444.905 3398.355 445.195 3398.400 ;
        RECT 469.285 3398.355 469.575 3398.400 ;
        RECT 541.505 3398.540 541.795 3398.585 ;
        RECT 565.885 3398.540 566.175 3398.585 ;
        RECT 541.505 3398.400 566.175 3398.540 ;
        RECT 541.505 3398.355 541.795 3398.400 ;
        RECT 565.885 3398.355 566.175 3398.400 ;
        RECT 638.105 3398.540 638.395 3398.585 ;
        RECT 662.485 3398.540 662.775 3398.585 ;
        RECT 638.105 3398.400 662.775 3398.540 ;
        RECT 638.105 3398.355 638.395 3398.400 ;
        RECT 662.485 3398.355 662.775 3398.400 ;
        RECT 734.705 3398.540 734.995 3398.585 ;
        RECT 759.085 3398.540 759.375 3398.585 ;
        RECT 734.705 3398.400 759.375 3398.540 ;
        RECT 734.705 3398.355 734.995 3398.400 ;
        RECT 759.085 3398.355 759.375 3398.400 ;
        RECT 831.305 3398.540 831.595 3398.585 ;
        RECT 855.685 3398.540 855.975 3398.585 ;
        RECT 831.305 3398.400 855.975 3398.540 ;
        RECT 831.305 3398.355 831.595 3398.400 ;
        RECT 855.685 3398.355 855.975 3398.400 ;
        RECT 927.905 3398.540 928.195 3398.585 ;
        RECT 952.285 3398.540 952.575 3398.585 ;
        RECT 927.905 3398.400 952.575 3398.540 ;
        RECT 927.905 3398.355 928.195 3398.400 ;
        RECT 952.285 3398.355 952.575 3398.400 ;
        RECT 1024.505 3398.540 1024.795 3398.585 ;
        RECT 1048.885 3398.540 1049.175 3398.585 ;
        RECT 1024.505 3398.400 1049.175 3398.540 ;
        RECT 1110.600 3398.540 1110.740 3398.695 ;
        RECT 1110.985 3398.540 1111.275 3398.585 ;
        RECT 1110.600 3398.400 1111.275 3398.540 ;
        RECT 1024.505 3398.355 1024.795 3398.400 ;
        RECT 1048.885 3398.355 1049.175 3398.400 ;
        RECT 1110.985 3398.355 1111.275 3398.400 ;
        RECT 1110.985 3397.860 1111.275 3397.905 ;
        RECT 1158.825 3397.860 1159.115 3397.905 ;
        RECT 1110.985 3397.720 1159.115 3397.860 ;
        RECT 1110.985 3397.675 1111.275 3397.720 ;
        RECT 1158.825 3397.675 1159.115 3397.720 ;
        RECT 9.730 3380.660 10.050 3380.920 ;
        RECT 9.820 3380.240 9.960 3380.660 ;
        RECT 9.730 3379.980 10.050 3380.240 ;
        RECT 9.730 3240.440 10.050 3240.500 ;
        RECT 9.535 3240.300 10.050 3240.440 ;
        RECT 9.730 3240.240 10.050 3240.300 ;
        RECT 9.730 3196.580 10.050 3196.640 ;
        RECT 9.535 3196.440 10.050 3196.580 ;
        RECT 9.730 3196.380 10.050 3196.440 ;
        RECT 9.285 3011.960 9.575 3012.005 ;
        RECT 9.730 3011.960 10.050 3012.020 ;
        RECT 9.285 3011.820 10.050 3011.960 ;
        RECT 9.285 3011.775 9.575 3011.820 ;
        RECT 9.730 3011.760 10.050 3011.820 ;
        RECT 9.285 2985.100 9.575 2985.145 ;
        RECT 9.730 2985.100 10.050 2985.160 ;
        RECT 9.285 2984.960 10.050 2985.100 ;
        RECT 9.285 2984.915 9.575 2984.960 ;
        RECT 9.730 2984.900 10.050 2984.960 ;
        RECT 9.730 2901.120 10.050 2901.180 ;
        RECT 9.535 2900.980 10.050 2901.120 ;
        RECT 9.730 2900.920 10.050 2900.980 ;
        RECT 9.285 2805.580 9.575 2805.625 ;
        RECT 9.730 2805.580 10.050 2805.640 ;
        RECT 9.285 2805.440 10.050 2805.580 ;
        RECT 9.285 2805.395 9.575 2805.440 ;
        RECT 9.730 2805.380 10.050 2805.440 ;
        RECT 9.285 2638.640 9.575 2638.685 ;
        RECT 9.730 2638.640 10.050 2638.700 ;
        RECT 9.285 2638.500 10.050 2638.640 ;
        RECT 9.285 2638.455 9.575 2638.500 ;
        RECT 9.730 2638.440 10.050 2638.500 ;
        RECT 9.285 2611.780 9.575 2611.825 ;
        RECT 9.730 2611.780 10.050 2611.840 ;
        RECT 9.285 2611.640 10.050 2611.780 ;
        RECT 9.285 2611.595 9.575 2611.640 ;
        RECT 9.730 2611.580 10.050 2611.640 ;
        RECT 9.285 2549.560 9.575 2549.605 ;
        RECT 9.730 2549.560 10.050 2549.620 ;
        RECT 9.285 2549.420 10.050 2549.560 ;
        RECT 9.285 2549.375 9.575 2549.420 ;
        RECT 9.730 2549.360 10.050 2549.420 ;
        RECT 9.270 2522.360 9.590 2522.420 ;
        RECT 9.075 2522.220 9.590 2522.360 ;
        RECT 9.270 2522.160 9.590 2522.220 ;
        RECT 9.270 2370.380 9.590 2370.440 ;
        RECT 9.075 2370.240 9.590 2370.380 ;
        RECT 9.270 2370.180 9.590 2370.240 ;
        RECT 9.285 2338.080 9.575 2338.125 ;
        RECT 9.730 2338.080 10.050 2338.140 ;
        RECT 9.285 2337.940 10.050 2338.080 ;
        RECT 9.285 2337.895 9.575 2337.940 ;
        RECT 9.730 2337.880 10.050 2337.940 ;
        RECT 7.905 2253.760 8.195 2253.805 ;
        RECT 9.730 2253.760 10.050 2253.820 ;
        RECT 7.905 2253.620 10.050 2253.760 ;
        RECT 7.905 2253.575 8.195 2253.620 ;
        RECT 9.730 2253.560 10.050 2253.620 ;
        RECT 7.905 2245.260 8.195 2245.305 ;
        RECT 9.270 2245.260 9.590 2245.320 ;
        RECT 7.905 2245.120 9.590 2245.260 ;
        RECT 7.905 2245.075 8.195 2245.120 ;
        RECT 9.270 2245.060 9.590 2245.120 ;
        RECT 8.825 2211.600 9.115 2211.645 ;
        RECT 9.270 2211.600 9.590 2211.660 ;
        RECT 8.825 2211.460 9.590 2211.600 ;
        RECT 8.825 2211.415 9.115 2211.460 ;
        RECT 9.270 2211.400 9.590 2211.460 ;
        RECT 8.825 2207.180 9.115 2207.225 ;
        RECT 9.730 2207.180 10.050 2207.240 ;
        RECT 8.825 2207.040 10.050 2207.180 ;
        RECT 8.825 2206.995 9.115 2207.040 ;
        RECT 9.730 2206.980 10.050 2207.040 ;
        RECT 9.730 1935.520 10.050 1935.580 ;
        RECT 9.535 1935.380 10.050 1935.520 ;
        RECT 9.730 1935.320 10.050 1935.380 ;
        RECT 7.905 1907.300 8.195 1907.345 ;
        RECT 9.745 1907.300 10.035 1907.345 ;
        RECT 7.905 1907.160 10.035 1907.300 ;
        RECT 7.905 1907.115 8.195 1907.160 ;
        RECT 9.745 1907.115 10.035 1907.160 ;
        RECT 7.905 1895.740 8.195 1895.785 ;
        RECT 9.730 1895.740 10.050 1895.800 ;
        RECT 7.905 1895.600 10.050 1895.740 ;
        RECT 7.905 1895.555 8.195 1895.600 ;
        RECT 9.730 1895.540 10.050 1895.600 ;
        RECT 8.825 1851.200 9.115 1851.245 ;
        RECT 9.730 1851.200 10.050 1851.260 ;
        RECT 8.825 1851.060 10.050 1851.200 ;
        RECT 8.825 1851.015 9.115 1851.060 ;
        RECT 9.730 1851.000 10.050 1851.060 ;
        RECT 7.905 1631.900 8.195 1631.945 ;
        RECT 9.285 1631.900 9.575 1631.945 ;
        RECT 7.905 1631.760 9.575 1631.900 ;
        RECT 7.905 1631.715 8.195 1631.760 ;
        RECT 9.285 1631.715 9.575 1631.760 ;
        RECT 8.365 1569.680 8.655 1569.725 ;
        RECT 9.285 1569.680 9.575 1569.725 ;
        RECT 8.365 1569.540 9.575 1569.680 ;
        RECT 8.365 1569.495 8.655 1569.540 ;
        RECT 9.285 1569.495 9.575 1569.540 ;
        RECT 8.365 1557.780 8.655 1557.825 ;
        RECT 9.730 1557.780 10.050 1557.840 ;
        RECT 8.365 1557.640 10.050 1557.780 ;
        RECT 8.365 1557.595 8.655 1557.640 ;
        RECT 9.730 1557.580 10.050 1557.640 ;
        RECT 8.825 1527.520 9.115 1527.565 ;
        RECT 9.730 1527.520 10.050 1527.580 ;
        RECT 8.825 1527.380 10.050 1527.520 ;
        RECT 8.825 1527.335 9.115 1527.380 ;
        RECT 9.730 1527.320 10.050 1527.380 ;
        RECT 8.825 1516.300 9.115 1516.345 ;
        RECT 9.730 1516.300 10.050 1516.360 ;
        RECT 8.825 1516.160 10.050 1516.300 ;
        RECT 8.825 1516.115 9.115 1516.160 ;
        RECT 9.730 1516.100 10.050 1516.160 ;
        RECT 8.365 1479.240 8.655 1479.285 ;
        RECT 9.730 1479.240 10.050 1479.300 ;
        RECT 8.365 1479.100 10.050 1479.240 ;
        RECT 8.365 1479.055 8.655 1479.100 ;
        RECT 9.730 1479.040 10.050 1479.100 ;
        RECT 8.825 1349.020 9.115 1349.065 ;
        RECT 9.730 1349.020 10.050 1349.080 ;
        RECT 8.825 1348.880 10.050 1349.020 ;
        RECT 8.825 1348.835 9.115 1348.880 ;
        RECT 9.730 1348.820 10.050 1348.880 ;
        RECT 9.285 1332.360 9.575 1332.405 ;
        RECT 9.730 1332.360 10.050 1332.420 ;
        RECT 9.285 1332.220 10.050 1332.360 ;
        RECT 9.285 1332.175 9.575 1332.220 ;
        RECT 9.730 1332.160 10.050 1332.220 ;
        RECT 7.905 1210.640 8.195 1210.685 ;
        RECT 9.285 1210.640 9.575 1210.685 ;
        RECT 7.905 1210.500 9.575 1210.640 ;
        RECT 7.905 1210.455 8.195 1210.500 ;
        RECT 9.285 1210.455 9.575 1210.500 ;
        RECT 7.905 1113.060 8.195 1113.105 ;
        RECT 9.285 1113.060 9.575 1113.105 ;
        RECT 7.905 1112.920 9.575 1113.060 ;
        RECT 7.905 1112.875 8.195 1112.920 ;
        RECT 9.285 1112.875 9.575 1112.920 ;
        RECT 9.285 1029.080 9.575 1029.125 ;
        RECT 8.900 1028.940 9.575 1029.080 ;
        RECT 8.900 1028.445 9.040 1028.940 ;
        RECT 9.285 1028.895 9.575 1028.940 ;
        RECT 8.825 1028.215 9.115 1028.445 ;
        RECT 2.385 896.140 2.675 896.185 ;
        RECT 9.745 896.140 10.035 896.185 ;
        RECT 2.385 896.000 10.035 896.140 ;
        RECT 2.385 895.955 2.675 896.000 ;
        RECT 9.745 895.955 10.035 896.000 ;
        RECT 2.370 851.600 2.690 851.660 ;
        RECT 2.175 851.460 2.690 851.600 ;
        RECT 2.370 851.400 2.690 851.460 ;
        RECT 2.370 830.860 2.690 830.920 ;
        RECT 5.605 830.860 5.895 830.905 ;
        RECT 2.370 830.720 5.895 830.860 ;
        RECT 2.370 830.660 2.690 830.720 ;
        RECT 5.605 830.675 5.895 830.720 ;
        RECT 4.225 731.580 4.515 731.625 ;
        RECT 6.525 731.580 6.815 731.625 ;
        RECT 4.225 731.440 6.815 731.580 ;
        RECT 4.225 731.395 4.515 731.440 ;
        RECT 6.525 731.395 6.815 731.440 ;
        RECT 4.685 695.540 4.975 695.585 ;
        RECT 9.730 695.540 10.050 695.600 ;
        RECT 4.685 695.400 10.050 695.540 ;
        RECT 4.685 695.355 4.975 695.400 ;
        RECT 9.730 695.340 10.050 695.400 ;
        RECT 7.445 630.600 7.735 630.645 ;
        RECT 9.730 630.600 10.050 630.660 ;
        RECT 7.445 630.460 10.050 630.600 ;
        RECT 7.445 630.415 7.735 630.460 ;
        RECT 9.730 630.400 10.050 630.460 ;
        RECT 6.510 582.320 6.830 582.380 ;
        RECT 7.445 582.320 7.735 582.365 ;
        RECT 6.510 582.180 7.735 582.320 ;
        RECT 6.510 582.120 6.830 582.180 ;
        RECT 7.445 582.135 7.735 582.180 ;
        RECT 6.510 536.760 6.830 536.820 ;
        RECT 9.730 536.760 10.050 536.820 ;
        RECT 6.510 536.620 10.050 536.760 ;
        RECT 6.510 536.560 6.830 536.620 ;
        RECT 9.730 536.560 10.050 536.620 ;
        RECT 9.730 490.860 10.050 490.920 ;
        RECT 9.535 490.720 10.050 490.860 ;
        RECT 9.730 490.660 10.050 490.720 ;
        RECT 6.065 443.940 6.355 443.985 ;
        RECT 9.745 443.940 10.035 443.985 ;
        RECT 6.065 443.800 10.035 443.940 ;
        RECT 6.065 443.755 6.355 443.800 ;
        RECT 9.745 443.755 10.035 443.800 ;
        RECT 6.065 403.480 6.355 403.525 ;
        RECT 7.445 403.480 7.735 403.525 ;
        RECT 6.065 403.340 7.735 403.480 ;
        RECT 6.065 403.295 6.355 403.340 ;
        RECT 7.445 403.295 7.735 403.340 ;
        RECT 0.990 334.800 1.310 334.860 ;
        RECT 7.445 334.800 7.735 334.845 ;
        RECT 0.990 334.660 7.735 334.800 ;
        RECT 0.990 334.600 1.310 334.660 ;
        RECT 7.445 334.615 7.735 334.660 ;
        RECT 24.910 2.620 25.230 2.680 ;
        RECT 25.385 2.620 25.675 2.665 ;
        RECT 24.910 2.480 25.675 2.620 ;
        RECT 24.910 2.420 25.230 2.480 ;
        RECT 25.385 2.435 25.675 2.480 ;
        RECT 27.225 2.280 27.515 2.325 ;
        RECT 51.145 2.280 51.435 2.325 ;
        RECT 27.225 2.140 51.435 2.280 ;
        RECT 27.225 2.095 27.515 2.140 ;
        RECT 51.145 2.095 51.435 2.140 ;
        RECT 52.985 0.580 53.275 0.625 ;
        RECT 221.790 0.580 222.110 0.640 ;
        RECT 52.985 0.440 222.110 0.580 ;
        RECT 52.985 0.395 53.275 0.440 ;
        RECT 221.790 0.380 222.110 0.440 ;
      LAYER via ;
        RECT 1231.060 3401.740 1231.320 3402.000 ;
        RECT 9.760 3399.020 10.020 3399.280 ;
        RECT 9.760 3380.660 10.020 3380.920 ;
        RECT 9.760 3379.980 10.020 3380.240 ;
        RECT 9.760 3240.240 10.020 3240.500 ;
        RECT 9.760 3196.380 10.020 3196.640 ;
        RECT 9.760 3011.760 10.020 3012.020 ;
        RECT 9.760 2984.900 10.020 2985.160 ;
        RECT 9.760 2900.920 10.020 2901.180 ;
        RECT 9.760 2805.380 10.020 2805.640 ;
        RECT 9.760 2638.440 10.020 2638.700 ;
        RECT 9.760 2611.580 10.020 2611.840 ;
        RECT 9.760 2549.360 10.020 2549.620 ;
        RECT 9.300 2522.160 9.560 2522.420 ;
        RECT 9.300 2370.180 9.560 2370.440 ;
        RECT 9.760 2337.880 10.020 2338.140 ;
        RECT 9.760 2253.560 10.020 2253.820 ;
        RECT 9.300 2245.060 9.560 2245.320 ;
        RECT 9.300 2211.400 9.560 2211.660 ;
        RECT 9.760 2206.980 10.020 2207.240 ;
        RECT 9.760 1935.320 10.020 1935.580 ;
        RECT 9.760 1895.540 10.020 1895.800 ;
        RECT 9.760 1851.000 10.020 1851.260 ;
        RECT 9.760 1557.580 10.020 1557.840 ;
        RECT 9.760 1527.320 10.020 1527.580 ;
        RECT 9.760 1516.100 10.020 1516.360 ;
        RECT 9.760 1479.040 10.020 1479.300 ;
        RECT 9.760 1348.820 10.020 1349.080 ;
        RECT 9.760 1332.160 10.020 1332.420 ;
        RECT 2.400 851.400 2.660 851.660 ;
        RECT 2.400 830.660 2.660 830.920 ;
        RECT 9.760 695.340 10.020 695.600 ;
        RECT 9.760 630.400 10.020 630.660 ;
        RECT 6.540 582.120 6.800 582.380 ;
        RECT 6.540 536.560 6.800 536.820 ;
        RECT 9.760 536.560 10.020 536.820 ;
        RECT 9.760 490.660 10.020 490.920 ;
        RECT 1.020 334.600 1.280 334.860 ;
        RECT 24.940 2.420 25.200 2.680 ;
        RECT 221.820 0.380 222.080 0.640 ;
      LAYER met2 ;
        RECT 1231.060 3401.770 1231.320 3402.030 ;
        RECT 1232.830 3401.770 1233.110 3405.000 ;
        RECT 1231.060 3401.710 1233.110 3401.770 ;
        RECT 1231.120 3401.630 1233.110 3401.710 ;
        RECT 1232.830 3401.000 1233.110 3401.630 ;
        RECT 9.760 3398.990 10.020 3399.310 ;
        RECT 9.820 3380.950 9.960 3398.990 ;
        RECT 9.760 3380.630 10.020 3380.950 ;
        RECT 9.760 3379.950 10.020 3380.270 ;
        RECT 9.820 3371.850 9.960 3379.950 ;
        RECT 9.820 3371.710 10.880 3371.850 ;
        RECT 9.760 3240.440 10.020 3240.530 ;
        RECT 10.740 3240.440 10.880 3371.710 ;
        RECT 9.760 3240.300 10.880 3240.440 ;
        RECT 9.760 3240.210 10.020 3240.300 ;
        RECT 9.760 3196.350 10.020 3196.670 ;
        RECT 9.820 3162.410 9.960 3196.350 ;
        RECT 9.820 3162.270 10.880 3162.410 ;
        RECT 10.740 3094.410 10.880 3162.270 ;
        RECT 10.740 3094.270 11.340 3094.410 ;
        RECT 11.200 3093.050 11.340 3094.270 ;
        RECT 10.740 3092.910 11.340 3093.050 ;
        RECT 10.740 3012.810 10.880 3092.910 ;
        RECT 9.820 3012.670 10.880 3012.810 ;
        RECT 9.820 3012.050 9.960 3012.670 ;
        RECT 9.760 3011.730 10.020 3012.050 ;
        RECT 9.760 2984.870 10.020 2985.190 ;
        RECT 9.820 2982.890 9.960 2984.870 ;
        RECT 9.820 2982.750 10.880 2982.890 ;
        RECT 10.740 2981.530 10.880 2982.750 ;
        RECT 10.740 2981.390 11.800 2981.530 ;
        RECT 11.660 2959.770 11.800 2981.390 ;
        RECT 10.740 2959.630 11.800 2959.770 ;
        RECT 10.740 2901.290 10.880 2959.630 ;
        RECT 9.820 2901.210 10.880 2901.290 ;
        RECT 9.760 2901.150 10.880 2901.210 ;
        RECT 9.760 2900.890 10.020 2901.150 ;
        RECT 9.760 2805.410 10.020 2805.670 ;
        RECT 9.760 2805.350 10.880 2805.410 ;
        RECT 9.820 2805.270 10.880 2805.350 ;
        RECT 10.740 2638.810 10.880 2805.270 ;
        RECT 9.820 2638.730 10.880 2638.810 ;
        RECT 9.760 2638.670 10.880 2638.730 ;
        RECT 9.760 2638.410 10.020 2638.670 ;
        RECT 9.760 2611.610 10.020 2611.870 ;
        RECT 9.760 2611.550 10.880 2611.610 ;
        RECT 9.820 2611.470 10.880 2611.550 ;
        RECT 9.760 2549.560 10.020 2549.650 ;
        RECT 10.740 2549.560 10.880 2611.470 ;
        RECT 9.760 2549.420 10.880 2549.560 ;
        RECT 9.760 2549.330 10.020 2549.420 ;
        RECT 9.300 2522.130 9.560 2522.450 ;
        RECT 9.360 2489.210 9.500 2522.130 ;
        RECT 9.360 2489.070 10.880 2489.210 ;
        RECT 10.740 2445.690 10.880 2489.070 ;
        RECT 10.280 2445.550 10.880 2445.690 ;
        RECT 10.280 2438.210 10.420 2445.550 ;
        RECT 10.280 2438.070 10.880 2438.210 ;
        RECT 10.740 2372.930 10.880 2438.070 ;
        RECT 9.360 2372.790 10.880 2372.930 ;
        RECT 9.360 2370.470 9.500 2372.790 ;
        RECT 9.300 2370.150 9.560 2370.470 ;
        RECT 9.760 2338.080 10.020 2338.170 ;
        RECT 9.760 2337.940 10.880 2338.080 ;
        RECT 9.760 2337.850 10.020 2337.940 ;
        RECT 10.740 2253.930 10.880 2337.940 ;
        RECT 9.820 2253.850 10.880 2253.930 ;
        RECT 9.760 2253.790 10.880 2253.850 ;
        RECT 9.760 2253.530 10.020 2253.790 ;
        RECT 9.300 2245.030 9.560 2245.350 ;
        RECT 9.360 2211.690 9.500 2245.030 ;
        RECT 9.300 2211.370 9.560 2211.690 ;
        RECT 9.760 2207.010 10.020 2207.270 ;
        RECT 9.760 2206.950 10.880 2207.010 ;
        RECT 9.820 2206.870 10.880 2206.950 ;
        RECT 10.740 1935.690 10.880 2206.870 ;
        RECT 9.820 1935.610 10.880 1935.690 ;
        RECT 9.760 1935.550 10.880 1935.610 ;
        RECT 9.760 1935.290 10.020 1935.550 ;
        RECT 9.760 1895.570 10.020 1895.830 ;
        RECT 9.760 1895.510 10.880 1895.570 ;
        RECT 9.820 1895.430 10.880 1895.510 ;
        RECT 10.740 1852.050 10.880 1895.430 ;
        RECT 10.280 1851.910 10.880 1852.050 ;
        RECT 10.280 1851.370 10.420 1851.910 ;
        RECT 9.820 1851.290 10.420 1851.370 ;
        RECT 9.760 1851.230 10.420 1851.290 ;
        RECT 9.760 1850.970 10.020 1851.230 ;
        RECT 9.760 1557.610 10.020 1557.870 ;
        RECT 9.760 1557.550 10.880 1557.610 ;
        RECT 9.820 1557.470 10.880 1557.550 ;
        RECT 9.760 1527.520 10.020 1527.610 ;
        RECT 10.740 1527.520 10.880 1557.470 ;
        RECT 9.760 1527.380 10.880 1527.520 ;
        RECT 9.760 1527.290 10.020 1527.380 ;
        RECT 9.760 1516.070 10.020 1516.390 ;
        RECT 9.820 1510.690 9.960 1516.070 ;
        RECT 9.820 1510.550 10.880 1510.690 ;
        RECT 10.740 1479.410 10.880 1510.550 ;
        RECT 9.820 1479.330 10.880 1479.410 ;
        RECT 9.760 1479.270 10.880 1479.330 ;
        RECT 9.760 1479.010 10.020 1479.270 ;
        RECT 9.760 1349.020 10.020 1349.110 ;
        RECT 9.760 1348.880 10.880 1349.020 ;
        RECT 9.760 1348.790 10.020 1348.880 ;
        RECT 10.740 1333.210 10.880 1348.880 ;
        RECT 10.280 1333.070 10.880 1333.210 ;
        RECT 10.280 1332.530 10.420 1333.070 ;
        RECT 9.820 1332.450 10.420 1332.530 ;
        RECT 9.760 1332.390 10.420 1332.450 ;
        RECT 9.760 1332.130 10.020 1332.390 ;
        RECT 2.400 851.370 2.660 851.690 ;
        RECT 2.460 830.950 2.600 851.370 ;
        RECT 2.400 830.630 2.660 830.950 ;
        RECT 9.760 695.370 10.020 695.630 ;
        RECT 9.760 695.310 12.260 695.370 ;
        RECT 9.820 695.230 12.260 695.310 ;
        RECT 12.120 658.650 12.260 695.230 ;
        RECT 8.900 658.510 12.260 658.650 ;
        RECT 8.900 642.330 9.040 658.510 ;
        RECT 8.900 642.190 9.960 642.330 ;
        RECT 9.820 630.690 9.960 642.190 ;
        RECT 9.760 630.370 10.020 630.690 ;
        RECT 6.540 582.090 6.800 582.410 ;
        RECT 6.600 536.850 6.740 582.090 ;
        RECT 6.540 536.530 6.800 536.850 ;
        RECT 9.760 536.760 10.020 536.850 ;
        RECT 9.760 536.620 11.340 536.760 ;
        RECT 9.760 536.530 10.020 536.620 ;
        RECT 11.200 517.210 11.340 536.620 ;
        RECT 10.740 517.070 11.340 517.210 ;
        RECT 9.760 490.860 10.020 490.950 ;
        RECT 10.740 490.860 10.880 517.070 ;
        RECT 9.760 490.720 10.880 490.860 ;
        RECT 9.760 490.630 10.020 490.720 ;
        RECT 1.020 334.570 1.280 334.890 ;
        RECT 1.080 3.245 1.220 334.570 ;
        RECT 1.010 2.875 1.290 3.245 ;
        RECT 24.930 2.875 25.210 3.245 ;
        RECT 221.880 2.990 222.940 3.130 ;
        RECT 25.000 2.710 25.140 2.875 ;
        RECT 24.940 2.390 25.200 2.710 ;
        RECT 221.880 0.670 222.020 2.990 ;
        RECT 222.800 2.400 222.940 2.990 ;
        RECT 221.820 0.350 222.080 0.670 ;
        RECT 222.590 -4.800 223.150 2.400 ;
      LAYER via2 ;
        RECT 1.010 2.920 1.290 3.200 ;
        RECT 24.930 2.920 25.210 3.200 ;
      LAYER met3 ;
        RECT 0.985 3.210 1.315 3.225 ;
        RECT 24.905 3.210 25.235 3.225 ;
        RECT 0.985 2.910 25.235 3.210 ;
        RECT 0.985 2.895 1.315 2.910 ;
        RECT 24.905 2.895 25.235 2.910 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 9.805 1214.565 9.975 1215.415 ;
        RECT 8.425 987.445 8.595 1107.635 ;
        RECT 9.805 1107.465 9.975 1212.695 ;
        RECT 8.425 540.345 8.595 623.815 ;
        RECT 5.665 458.065 5.835 470.135 ;
        RECT 5.665 351.985 5.835 423.215 ;
        RECT 6.585 263.585 6.755 351.475 ;
        RECT 5.205 147.645 5.375 177.055 ;
      LAYER mcon ;
        RECT 9.805 1215.245 9.975 1215.415 ;
        RECT 9.805 1212.525 9.975 1212.695 ;
        RECT 8.425 1107.465 8.595 1107.635 ;
        RECT 8.425 623.645 8.595 623.815 ;
        RECT 5.665 469.965 5.835 470.135 ;
        RECT 5.665 423.045 5.835 423.215 ;
        RECT 6.585 351.305 6.755 351.475 ;
        RECT 5.205 176.885 5.375 177.055 ;
      LAYER met1 ;
        RECT 3.750 1287.140 4.070 1287.200 ;
        RECT 6.970 1287.140 7.290 1287.200 ;
        RECT 3.750 1287.000 7.290 1287.140 ;
        RECT 3.750 1286.940 4.070 1287.000 ;
        RECT 6.970 1286.940 7.290 1287.000 ;
        RECT 6.510 1244.980 6.830 1245.040 ;
        RECT 9.730 1244.980 10.050 1245.040 ;
        RECT 6.510 1244.840 10.050 1244.980 ;
        RECT 6.510 1244.780 6.830 1244.840 ;
        RECT 9.730 1244.780 10.050 1244.840 ;
        RECT 9.730 1215.400 10.050 1215.460 ;
        RECT 9.535 1215.260 10.050 1215.400 ;
        RECT 9.730 1215.200 10.050 1215.260 ;
        RECT 9.730 1214.720 10.050 1214.780 ;
        RECT 9.730 1214.580 10.245 1214.720 ;
        RECT 9.730 1214.520 10.050 1214.580 ;
        RECT 9.730 1212.680 10.050 1212.740 ;
        RECT 9.535 1212.540 10.050 1212.680 ;
        RECT 9.730 1212.480 10.050 1212.540 ;
        RECT 8.365 1107.620 8.655 1107.665 ;
        RECT 9.745 1107.620 10.035 1107.665 ;
        RECT 8.365 1107.480 10.035 1107.620 ;
        RECT 8.365 1107.435 8.655 1107.480 ;
        RECT 9.745 1107.435 10.035 1107.480 ;
        RECT 4.670 987.600 4.990 987.660 ;
        RECT 8.365 987.600 8.655 987.645 ;
        RECT 4.670 987.460 8.655 987.600 ;
        RECT 4.670 987.400 4.990 987.460 ;
        RECT 8.365 987.415 8.655 987.460 ;
        RECT 4.670 673.440 4.990 673.500 ;
        RECT 6.970 673.440 7.290 673.500 ;
        RECT 4.670 673.300 7.290 673.440 ;
        RECT 4.670 673.240 4.990 673.300 ;
        RECT 6.970 673.240 7.290 673.300 ;
        RECT 6.970 623.800 7.290 623.860 ;
        RECT 8.365 623.800 8.655 623.845 ;
        RECT 6.970 623.660 8.655 623.800 ;
        RECT 6.970 623.600 7.290 623.660 ;
        RECT 8.365 623.615 8.655 623.660 ;
        RECT 8.365 540.500 8.655 540.545 ;
        RECT 9.730 540.500 10.050 540.560 ;
        RECT 8.365 540.360 10.050 540.500 ;
        RECT 8.365 540.315 8.655 540.360 ;
        RECT 9.730 540.300 10.050 540.360 ;
        RECT 5.605 470.120 5.895 470.165 ;
        RECT 9.730 470.120 10.050 470.180 ;
        RECT 5.605 469.980 10.050 470.120 ;
        RECT 5.605 469.935 5.895 469.980 ;
        RECT 9.730 469.920 10.050 469.980 ;
        RECT 5.605 458.220 5.895 458.265 ;
        RECT 9.730 458.220 10.050 458.280 ;
        RECT 5.605 458.080 10.050 458.220 ;
        RECT 5.605 458.035 5.895 458.080 ;
        RECT 9.730 458.020 10.050 458.080 ;
        RECT 5.605 423.200 5.895 423.245 ;
        RECT 9.730 423.200 10.050 423.260 ;
        RECT 5.605 423.060 10.050 423.200 ;
        RECT 5.605 423.015 5.895 423.060 ;
        RECT 9.730 423.000 10.050 423.060 ;
        RECT 5.605 351.955 5.895 352.185 ;
        RECT 5.680 351.460 5.820 351.955 ;
        RECT 6.525 351.460 6.815 351.505 ;
        RECT 5.680 351.320 6.815 351.460 ;
        RECT 6.525 351.275 6.815 351.320 ;
        RECT 6.525 263.740 6.815 263.785 ;
        RECT 9.730 263.740 10.050 263.800 ;
        RECT 6.525 263.600 10.050 263.740 ;
        RECT 6.525 263.555 6.815 263.600 ;
        RECT 9.730 263.540 10.050 263.600 ;
        RECT 5.145 177.040 5.435 177.085 ;
        RECT 9.730 177.040 10.050 177.100 ;
        RECT 5.145 176.900 10.050 177.040 ;
        RECT 5.145 176.855 5.435 176.900 ;
        RECT 9.730 176.840 10.050 176.900 ;
        RECT 5.145 147.800 5.435 147.845 ;
        RECT 8.810 147.800 9.130 147.860 ;
        RECT 5.145 147.660 9.130 147.800 ;
        RECT 5.145 147.615 5.435 147.660 ;
        RECT 8.810 147.600 9.130 147.660 ;
        RECT 7.430 75.040 7.750 75.100 ;
        RECT 8.810 75.040 9.130 75.100 ;
        RECT 7.430 74.900 9.130 75.040 ;
        RECT 7.430 74.840 7.750 74.900 ;
        RECT 8.810 74.840 9.130 74.900 ;
        RECT 7.430 62.460 7.750 62.520 ;
        RECT 9.730 62.460 10.050 62.520 ;
        RECT 7.430 62.320 10.050 62.460 ;
        RECT 7.430 62.260 7.750 62.320 ;
        RECT 9.730 62.260 10.050 62.320 ;
        RECT 14.790 8.400 15.110 8.460 ;
        RECT 20.310 8.400 20.630 8.460 ;
        RECT 14.790 8.260 20.630 8.400 ;
        RECT 14.790 8.200 15.110 8.260 ;
        RECT 20.310 8.200 20.630 8.260 ;
      LAYER via ;
        RECT 3.780 1286.940 4.040 1287.200 ;
        RECT 7.000 1286.940 7.260 1287.200 ;
        RECT 6.540 1244.780 6.800 1245.040 ;
        RECT 9.760 1244.780 10.020 1245.040 ;
        RECT 9.760 1215.200 10.020 1215.460 ;
        RECT 9.760 1214.520 10.020 1214.780 ;
        RECT 9.760 1212.480 10.020 1212.740 ;
        RECT 4.700 987.400 4.960 987.660 ;
        RECT 4.700 673.240 4.960 673.500 ;
        RECT 7.000 673.240 7.260 673.500 ;
        RECT 7.000 623.600 7.260 623.860 ;
        RECT 9.760 540.300 10.020 540.560 ;
        RECT 9.760 469.920 10.020 470.180 ;
        RECT 9.760 458.020 10.020 458.280 ;
        RECT 9.760 423.000 10.020 423.260 ;
        RECT 9.760 263.540 10.020 263.800 ;
        RECT 9.760 176.840 10.020 177.100 ;
        RECT 8.840 147.600 9.100 147.860 ;
        RECT 7.460 74.840 7.720 75.100 ;
        RECT 8.840 74.840 9.100 75.100 ;
        RECT 7.460 62.260 7.720 62.520 ;
        RECT 9.760 62.260 10.020 62.520 ;
        RECT 14.820 8.200 15.080 8.460 ;
        RECT 20.340 8.200 20.600 8.460 ;
      LAYER met2 ;
        RECT 3.770 2211.515 4.050 2211.885 ;
        RECT 3.840 1287.230 3.980 2211.515 ;
        RECT 3.780 1286.910 4.040 1287.230 ;
        RECT 7.000 1286.910 7.260 1287.230 ;
        RECT 7.060 1259.090 7.200 1286.910 ;
        RECT 6.600 1258.950 7.200 1259.090 ;
        RECT 6.600 1245.070 6.740 1258.950 ;
        RECT 6.540 1244.750 6.800 1245.070 ;
        RECT 9.760 1244.750 10.020 1245.070 ;
        RECT 9.820 1215.490 9.960 1244.750 ;
        RECT 9.760 1215.170 10.020 1215.490 ;
        RECT 9.760 1214.490 10.020 1214.810 ;
        RECT 9.820 1212.770 9.960 1214.490 ;
        RECT 9.760 1212.450 10.020 1212.770 ;
        RECT 4.700 987.370 4.960 987.690 ;
        RECT 4.760 673.530 4.900 987.370 ;
        RECT 4.700 673.210 4.960 673.530 ;
        RECT 7.000 673.210 7.260 673.530 ;
        RECT 7.060 623.890 7.200 673.210 ;
        RECT 7.000 623.570 7.260 623.890 ;
        RECT 9.760 540.330 10.020 540.590 ;
        RECT 9.760 540.270 13.180 540.330 ;
        RECT 9.820 540.190 13.180 540.270 ;
        RECT 9.760 470.120 10.020 470.210 ;
        RECT 13.040 470.120 13.180 540.190 ;
        RECT 9.760 469.980 13.180 470.120 ;
        RECT 9.760 469.890 10.020 469.980 ;
        RECT 9.760 458.220 10.020 458.310 ;
        RECT 9.760 458.080 13.180 458.220 ;
        RECT 9.760 457.990 10.020 458.080 ;
        RECT 13.040 423.370 13.180 458.080 ;
        RECT 9.820 423.290 13.180 423.370 ;
        RECT 9.760 423.230 13.180 423.290 ;
        RECT 9.760 422.970 10.020 423.230 ;
        RECT 9.760 263.740 10.020 263.830 ;
        RECT 9.760 263.600 10.420 263.740 ;
        RECT 9.760 263.510 10.020 263.600 ;
        RECT 10.280 257.450 10.420 263.600 ;
        RECT 10.280 257.310 10.880 257.450 ;
        RECT 10.740 217.330 10.880 257.310 ;
        RECT 10.740 217.190 11.800 217.330 ;
        RECT 11.660 215.970 11.800 217.190 ;
        RECT 11.660 215.830 13.180 215.970 ;
        RECT 13.040 177.210 13.180 215.830 ;
        RECT 9.820 177.130 13.180 177.210 ;
        RECT 9.760 177.070 13.180 177.130 ;
        RECT 9.760 176.810 10.020 177.070 ;
        RECT 8.840 147.570 9.100 147.890 ;
        RECT 8.900 75.130 9.040 147.570 ;
        RECT 7.460 74.810 7.720 75.130 ;
        RECT 8.840 74.810 9.100 75.130 ;
        RECT 7.520 62.550 7.660 74.810 ;
        RECT 7.460 62.230 7.720 62.550 ;
        RECT 9.760 62.460 10.020 62.550 ;
        RECT 9.760 62.320 15.020 62.460 ;
        RECT 9.760 62.230 10.020 62.320 ;
        RECT 14.880 8.490 15.020 62.320 ;
        RECT 14.820 8.170 15.080 8.490 ;
        RECT 20.340 8.170 20.600 8.490 ;
        RECT 20.400 2.400 20.540 8.170 ;
        RECT 20.190 -4.800 20.750 2.400 ;
      LAYER via2 ;
        RECT 3.770 2211.560 4.050 2211.840 ;
      LAYER met3 ;
        RECT 5.000 2214.360 9.000 2214.960 ;
        RECT 3.745 2211.850 4.075 2211.865 ;
        RECT 5.830 2211.850 6.130 2214.360 ;
        RECT 3.745 2211.550 6.130 2211.850 ;
        RECT 3.745 2211.535 4.075 2211.550 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2217.805 3395.665 2217.975 3401.955 ;
        RECT 2373.745 3400.085 2373.915 3401.955 ;
        RECT 2774.405 3395.665 2774.575 3401.615 ;
        RECT 5.205 92.905 5.375 135.575 ;
        RECT 7.505 73.185 7.675 79.815 ;
        RECT 28.205 6.885 28.375 9.095 ;
        RECT 243.485 8.925 245.035 9.095 ;
        RECT 129.405 4.165 129.575 5.015 ;
        RECT 140.905 0.765 141.075 4.335 ;
        RECT 174.945 1.615 175.115 8.755 ;
        RECT 243.485 8.585 243.655 8.925 ;
        RECT 174.945 1.445 176.495 1.615 ;
        RECT 190.125 0.765 190.295 8.415 ;
        RECT 196.105 0.595 196.275 1.955 ;
        RECT 199.325 0.595 199.495 1.615 ;
        RECT 196.105 0.425 199.495 0.595 ;
      LAYER mcon ;
        RECT 2217.805 3401.785 2217.975 3401.955 ;
        RECT 2373.745 3401.785 2373.915 3401.955 ;
        RECT 2774.405 3401.445 2774.575 3401.615 ;
        RECT 5.205 135.405 5.375 135.575 ;
        RECT 7.505 79.645 7.675 79.815 ;
        RECT 28.205 8.925 28.375 9.095 ;
        RECT 244.865 8.925 245.035 9.095 ;
        RECT 174.945 8.585 175.115 8.755 ;
        RECT 129.405 4.845 129.575 5.015 ;
        RECT 140.905 4.165 141.075 4.335 ;
        RECT 190.125 8.245 190.295 8.415 ;
        RECT 176.325 1.445 176.495 1.615 ;
        RECT 196.105 1.785 196.275 1.955 ;
        RECT 199.325 1.445 199.495 1.615 ;
      LAYER met1 ;
        RECT 2314.330 3416.220 2314.650 3416.280 ;
        RECT 2359.870 3416.220 2360.190 3416.280 ;
        RECT 2314.330 3416.080 2360.190 3416.220 ;
        RECT 2314.330 3416.020 2314.650 3416.080 ;
        RECT 2359.870 3416.020 2360.190 3416.080 ;
        RECT 2217.730 3401.940 2218.050 3402.000 ;
        RECT 2217.535 3401.800 2218.050 3401.940 ;
        RECT 2217.730 3401.740 2218.050 3401.800 ;
        RECT 2359.870 3401.940 2360.190 3402.000 ;
        RECT 2373.685 3401.940 2373.975 3401.985 ;
        RECT 2359.870 3401.800 2373.975 3401.940 ;
        RECT 2359.870 3401.740 2360.190 3401.800 ;
        RECT 2373.685 3401.755 2373.975 3401.800 ;
        RECT 2774.330 3401.600 2774.650 3401.660 ;
        RECT 2774.330 3401.460 2774.845 3401.600 ;
        RECT 2774.330 3401.400 2774.650 3401.460 ;
        RECT 2792.730 3401.400 2793.050 3401.660 ;
        RECT 2373.685 3400.240 2373.975 3400.285 ;
        RECT 2792.820 3400.240 2792.960 3401.400 ;
        RECT 2373.685 3400.100 2792.960 3400.240 ;
        RECT 2373.685 3400.055 2373.975 3400.100 ;
        RECT 2217.745 3395.820 2218.035 3395.865 ;
        RECT 2774.345 3395.820 2774.635 3395.865 ;
        RECT 2217.745 3395.680 2774.635 3395.820 ;
        RECT 2217.745 3395.635 2218.035 3395.680 ;
        RECT 2774.345 3395.635 2774.635 3395.680 ;
        RECT 5.145 135.560 5.435 135.605 ;
        RECT 6.050 135.560 6.370 135.620 ;
        RECT 5.145 135.420 6.370 135.560 ;
        RECT 5.145 135.375 5.435 135.420 ;
        RECT 6.050 135.360 6.370 135.420 ;
        RECT 0.530 100.880 0.850 100.940 ;
        RECT 6.970 100.880 7.290 100.940 ;
        RECT 0.530 100.740 7.290 100.880 ;
        RECT 0.530 100.680 0.850 100.740 ;
        RECT 6.970 100.680 7.290 100.740 ;
        RECT 5.145 93.060 5.435 93.105 ;
        RECT 6.970 93.060 7.290 93.120 ;
        RECT 5.145 92.920 7.290 93.060 ;
        RECT 5.145 92.875 5.435 92.920 ;
        RECT 6.970 92.860 7.290 92.920 ;
        RECT 6.970 79.800 7.290 79.860 ;
        RECT 7.445 79.800 7.735 79.845 ;
        RECT 6.970 79.660 7.735 79.800 ;
        RECT 6.970 79.600 7.290 79.660 ;
        RECT 7.445 79.615 7.735 79.660 ;
        RECT 5.590 73.340 5.910 73.400 ;
        RECT 7.445 73.340 7.735 73.385 ;
        RECT 5.590 73.200 7.735 73.340 ;
        RECT 5.590 73.140 5.910 73.200 ;
        RECT 7.445 73.155 7.735 73.200 ;
        RECT 5.590 65.180 5.910 65.240 ;
        RECT 9.730 65.180 10.050 65.240 ;
        RECT 5.590 65.040 10.050 65.180 ;
        RECT 5.590 64.980 5.910 65.040 ;
        RECT 9.730 64.980 10.050 65.040 ;
        RECT 28.145 9.080 28.435 9.125 ;
        RECT 244.805 9.080 245.095 9.125 ;
        RECT 28.145 8.940 134.620 9.080 ;
        RECT 28.145 8.895 28.435 8.940 ;
        RECT 134.480 8.740 134.620 8.940 ;
        RECT 244.805 8.940 282.280 9.080 ;
        RECT 244.805 8.895 245.095 8.940 ;
        RECT 282.140 8.800 282.280 8.940 ;
        RECT 174.885 8.740 175.175 8.785 ;
        RECT 134.480 8.600 175.175 8.740 ;
        RECT 174.885 8.555 175.175 8.600 ;
        RECT 243.410 8.740 243.730 8.800 ;
        RECT 243.410 8.600 243.925 8.740 ;
        RECT 243.410 8.540 243.730 8.600 ;
        RECT 282.050 8.540 282.370 8.800 ;
        RECT 190.065 8.400 190.355 8.445 ;
        RECT 195.110 8.400 195.430 8.460 ;
        RECT 190.065 8.260 195.430 8.400 ;
        RECT 190.065 8.215 190.355 8.260 ;
        RECT 195.110 8.200 195.430 8.260 ;
        RECT 197.870 7.720 198.190 7.780 ;
        RECT 205.690 7.720 206.010 7.780 ;
        RECT 197.870 7.580 206.010 7.720 ;
        RECT 197.870 7.520 198.190 7.580 ;
        RECT 205.690 7.520 206.010 7.580 ;
        RECT 26.290 7.040 26.610 7.100 ;
        RECT 28.145 7.040 28.435 7.085 ;
        RECT 26.290 6.900 28.435 7.040 ;
        RECT 26.290 6.840 26.610 6.900 ;
        RECT 28.145 6.855 28.435 6.900 ;
        RECT 16.170 5.000 16.490 5.060 ;
        RECT 129.345 5.000 129.635 5.045 ;
        RECT 16.170 4.860 129.635 5.000 ;
        RECT 16.170 4.800 16.490 4.860 ;
        RECT 129.345 4.815 129.635 4.860 ;
        RECT 129.345 4.320 129.635 4.365 ;
        RECT 140.845 4.320 141.135 4.365 ;
        RECT 129.345 4.180 141.135 4.320 ;
        RECT 129.345 4.135 129.635 4.180 ;
        RECT 140.845 4.135 141.135 4.180 ;
        RECT 0.530 2.960 0.850 3.020 ;
        RECT 24.450 2.960 24.770 3.020 ;
        RECT 0.530 2.820 24.770 2.960 ;
        RECT 0.530 2.760 0.850 2.820 ;
        RECT 24.450 2.760 24.770 2.820 ;
        RECT 196.045 1.940 196.335 1.985 ;
        RECT 193.820 1.800 196.335 1.940 ;
        RECT 176.265 1.600 176.555 1.645 ;
        RECT 193.820 1.600 193.960 1.800 ;
        RECT 196.045 1.755 196.335 1.800 ;
        RECT 176.265 1.460 193.960 1.600 ;
        RECT 199.265 1.600 199.555 1.645 ;
        RECT 245.710 1.600 246.030 1.660 ;
        RECT 199.265 1.460 246.030 1.600 ;
        RECT 176.265 1.415 176.555 1.460 ;
        RECT 199.265 1.415 199.555 1.460 ;
        RECT 245.710 1.400 246.030 1.460 ;
        RECT 140.845 0.920 141.135 0.965 ;
        RECT 190.065 0.920 190.355 0.965 ;
        RECT 140.845 0.780 190.355 0.920 ;
        RECT 140.845 0.735 141.135 0.780 ;
        RECT 190.065 0.735 190.355 0.780 ;
      LAYER via ;
        RECT 2314.360 3416.020 2314.620 3416.280 ;
        RECT 2359.900 3416.020 2360.160 3416.280 ;
        RECT 2217.760 3401.740 2218.020 3402.000 ;
        RECT 2359.900 3401.740 2360.160 3402.000 ;
        RECT 2774.360 3401.400 2774.620 3401.660 ;
        RECT 2792.760 3401.400 2793.020 3401.660 ;
        RECT 6.080 135.360 6.340 135.620 ;
        RECT 0.560 100.680 0.820 100.940 ;
        RECT 7.000 100.680 7.260 100.940 ;
        RECT 7.000 92.860 7.260 93.120 ;
        RECT 7.000 79.600 7.260 79.860 ;
        RECT 5.620 73.140 5.880 73.400 ;
        RECT 5.620 64.980 5.880 65.240 ;
        RECT 9.760 64.980 10.020 65.240 ;
        RECT 243.440 8.540 243.700 8.800 ;
        RECT 282.080 8.540 282.340 8.800 ;
        RECT 195.140 8.200 195.400 8.460 ;
        RECT 197.900 7.520 198.160 7.780 ;
        RECT 205.720 7.520 205.980 7.780 ;
        RECT 26.320 6.840 26.580 7.100 ;
        RECT 16.200 4.800 16.460 5.060 ;
        RECT 0.560 2.760 0.820 3.020 ;
        RECT 24.480 2.760 24.740 3.020 ;
        RECT 245.740 1.400 246.000 1.660 ;
      LAYER met2 ;
        RECT 2314.360 3415.990 2314.620 3416.310 ;
        RECT 2359.900 3415.990 2360.160 3416.310 ;
        RECT 2314.420 3405.000 2314.560 3415.990 ;
        RECT 2215.850 3401.770 2216.130 3405.000 ;
        RECT 2217.760 3401.770 2218.020 3402.030 ;
        RECT 2215.850 3401.710 2218.020 3401.770 ;
        RECT 2215.850 3401.630 2217.960 3401.710 ;
        RECT 2215.850 3401.000 2216.130 3401.630 ;
        RECT 2314.290 3401.000 2314.570 3405.000 ;
        RECT 2359.960 3402.030 2360.100 3415.990 ;
        RECT 2359.900 3401.710 2360.160 3402.030 ;
        RECT 2774.350 3401.515 2774.630 3401.885 ;
        RECT 2792.750 3401.515 2793.030 3401.885 ;
        RECT 2774.360 3401.370 2774.620 3401.515 ;
        RECT 2792.760 3401.370 2793.020 3401.515 ;
        RECT 6.070 166.075 6.350 166.445 ;
        RECT 6.140 135.650 6.280 166.075 ;
        RECT 6.990 148.395 7.270 148.765 ;
        RECT 6.080 135.330 6.340 135.650 ;
        RECT 7.060 100.970 7.200 148.395 ;
        RECT 0.560 100.650 0.820 100.970 ;
        RECT 7.000 100.650 7.260 100.970 ;
        RECT 0.620 3.050 0.760 100.650 ;
        RECT 7.000 92.830 7.260 93.150 ;
        RECT 7.060 79.890 7.200 92.830 ;
        RECT 7.000 79.570 7.260 79.890 ;
        RECT 5.620 73.110 5.880 73.430 ;
        RECT 5.680 65.270 5.820 73.110 ;
        RECT 5.620 64.950 5.880 65.270 ;
        RECT 9.760 65.180 10.020 65.270 ;
        RECT 9.760 65.040 16.400 65.180 ;
        RECT 9.760 64.950 10.020 65.040 ;
        RECT 16.260 5.090 16.400 65.040 ;
        RECT 243.440 8.685 243.700 8.830 ;
        RECT 195.200 8.490 198.100 8.570 ;
        RECT 195.140 8.430 198.100 8.490 ;
        RECT 195.140 8.170 195.400 8.430 ;
        RECT 197.960 7.810 198.100 8.430 ;
        RECT 205.710 8.315 205.990 8.685 ;
        RECT 243.430 8.315 243.710 8.685 ;
        RECT 282.080 8.510 282.340 8.830 ;
        RECT 205.780 7.810 205.920 8.315 ;
        RECT 197.900 7.490 198.160 7.810 ;
        RECT 205.720 7.490 205.980 7.810 ;
        RECT 24.540 7.130 26.520 7.210 ;
        RECT 24.540 7.070 26.580 7.130 ;
        RECT 16.200 4.770 16.460 5.090 ;
        RECT 24.540 3.050 24.680 7.070 ;
        RECT 26.320 6.810 26.580 7.070 ;
        RECT 0.560 2.730 0.820 3.050 ;
        RECT 24.480 2.730 24.740 3.050 ;
        RECT 245.800 2.990 246.860 3.130 ;
        RECT 245.800 1.690 245.940 2.990 ;
        RECT 246.720 2.400 246.860 2.990 ;
        RECT 282.140 2.400 282.280 8.510 ;
        RECT 245.740 1.370 246.000 1.690 ;
        RECT 246.510 -4.800 247.070 2.400 ;
        RECT 281.930 -4.800 282.490 2.400 ;
      LAYER via2 ;
        RECT 2774.350 3401.560 2774.630 3401.840 ;
        RECT 2792.750 3401.560 2793.030 3401.840 ;
        RECT 6.070 166.120 6.350 166.400 ;
        RECT 6.990 148.440 7.270 148.720 ;
        RECT 205.710 8.360 205.990 8.640 ;
        RECT 243.430 8.360 243.710 8.640 ;
      LAYER met3 ;
        RECT 2795.230 3402.530 2795.610 3402.540 ;
        RECT 2791.590 3402.230 2795.610 3402.530 ;
        RECT 2774.325 3401.850 2774.655 3401.865 ;
        RECT 2791.590 3401.850 2791.890 3402.230 ;
        RECT 2795.230 3402.220 2795.610 3402.230 ;
        RECT 2774.325 3401.550 2791.890 3401.850 ;
        RECT 2792.725 3401.850 2793.055 3401.865 ;
        RECT 2797.070 3401.850 2797.450 3401.860 ;
        RECT 2792.725 3401.550 2797.450 3401.850 ;
        RECT 2774.325 3401.535 2774.655 3401.550 ;
        RECT 2792.725 3401.535 2793.055 3401.550 ;
        RECT 2797.070 3401.540 2797.450 3401.550 ;
        RECT 6.045 166.410 6.375 166.425 ;
        RECT 7.630 166.410 8.010 166.420 ;
        RECT 6.045 166.110 8.010 166.410 ;
        RECT 6.045 166.095 6.375 166.110 ;
        RECT 7.630 166.100 8.010 166.110 ;
        RECT 6.965 148.740 7.295 148.745 ;
        RECT 6.710 148.730 7.295 148.740 ;
        RECT 6.510 148.430 7.295 148.730 ;
        RECT 6.710 148.420 7.295 148.430 ;
        RECT 6.965 148.415 7.295 148.420 ;
        RECT 205.685 8.650 206.015 8.665 ;
        RECT 243.405 8.650 243.735 8.665 ;
        RECT 205.685 8.350 243.735 8.650 ;
        RECT 205.685 8.335 206.015 8.350 ;
        RECT 243.405 8.335 243.735 8.350 ;
      LAYER via3 ;
        RECT 2795.260 3402.220 2795.580 3402.540 ;
        RECT 2797.100 3401.540 2797.420 3401.860 ;
        RECT 7.660 166.100 7.980 166.420 ;
        RECT 6.740 148.420 7.060 148.740 ;
      LAYER met4 ;
        RECT 2795.255 3402.530 2795.585 3402.545 ;
        RECT 2795.255 3402.230 2796.490 3402.530 ;
        RECT 2795.255 3402.215 2795.585 3402.230 ;
        RECT 2796.190 3330.890 2796.490 3402.230 ;
        RECT 2797.095 3401.535 2797.425 3401.865 ;
        RECT 2797.110 3371.250 2797.410 3401.535 ;
        RECT 2797.110 3370.950 2798.330 3371.250 ;
        RECT 2795.750 3329.710 2796.930 3330.890 ;
        RECT 2798.030 3235.250 2798.330 3370.950 ;
        RECT 2801.270 3330.450 2802.450 3330.890 ;
        RECT 2799.870 3330.150 2802.450 3330.450 ;
        RECT 2799.870 3265.850 2800.170 3330.150 ;
        RECT 2801.270 3329.710 2802.450 3330.150 ;
        RECT 2796.190 3234.950 2798.330 3235.250 ;
        RECT 2798.950 3265.550 2800.170 3265.850 ;
        RECT 2796.190 3191.050 2796.490 3234.950 ;
        RECT 2798.950 3231.850 2799.250 3265.550 ;
        RECT 2798.950 3231.550 2800.170 3231.850 ;
        RECT 2799.870 3211.450 2800.170 3231.550 ;
        RECT 2799.870 3211.150 2802.010 3211.450 ;
        RECT 2801.710 3191.050 2802.010 3211.150 ;
        RECT 2796.190 3190.750 2803.850 3191.050 ;
        RECT 2795.270 3163.550 2800.170 3163.850 ;
        RECT 2795.270 3136.650 2795.570 3163.550 ;
        RECT 2799.870 3153.650 2800.170 3163.550 ;
        RECT 2801.710 3153.650 2802.010 3190.750 ;
        RECT 2799.870 3153.350 2802.010 3153.650 ;
        RECT 2803.550 3146.850 2803.850 3190.750 ;
        RECT 2796.190 3146.550 2803.850 3146.850 ;
        RECT 2796.190 3143.450 2796.490 3146.550 ;
        RECT 2796.190 3143.150 2799.250 3143.450 ;
        RECT 2795.270 3136.350 2796.490 3136.650 ;
        RECT 2796.190 2704.850 2796.490 3136.350 ;
        RECT 2798.950 3092.450 2799.250 3143.150 ;
        RECT 2798.030 3092.150 2799.250 3092.450 ;
        RECT 2796.190 2704.550 2797.410 2704.850 ;
        RECT 2797.110 2660.650 2797.410 2704.550 ;
        RECT 2798.030 2674.250 2798.330 3092.150 ;
        RECT 2798.030 2673.950 2799.250 2674.250 ;
        RECT 2798.950 2660.650 2799.250 2673.950 ;
        RECT 2796.190 2660.350 2797.410 2660.650 ;
        RECT 2798.030 2660.350 2799.250 2660.650 ;
        RECT 2796.190 1062.650 2796.490 2660.350 ;
        RECT 2798.030 2497.450 2798.330 2660.350 ;
        RECT 2798.030 2497.150 2800.170 2497.450 ;
        RECT 2799.870 2449.850 2800.170 2497.150 ;
        RECT 2798.030 2449.550 2800.170 2449.850 ;
        RECT 2798.030 2256.050 2798.330 2449.550 ;
        RECT 2798.030 2255.750 2799.250 2256.050 ;
        RECT 2798.950 2208.450 2799.250 2255.750 ;
        RECT 2798.030 2208.150 2799.250 2208.450 ;
        RECT 2798.030 2014.650 2798.330 2208.150 ;
        RECT 2798.030 2014.350 2800.170 2014.650 ;
        RECT 2799.870 1967.050 2800.170 2014.350 ;
        RECT 2798.030 1966.750 2800.170 1967.050 ;
        RECT 2798.030 1773.250 2798.330 1966.750 ;
        RECT 2798.030 1772.950 2799.250 1773.250 ;
        RECT 2798.950 1718.850 2799.250 1772.950 ;
        RECT 2798.030 1718.550 2799.250 1718.850 ;
        RECT 2798.030 1433.250 2798.330 1718.550 ;
        RECT 2797.110 1432.950 2798.330 1433.250 ;
        RECT 2797.110 1392.450 2797.410 1432.950 ;
        RECT 2797.110 1392.150 2798.330 1392.450 ;
        RECT 2798.030 1385.650 2798.330 1392.150 ;
        RECT 2798.030 1385.350 2799.250 1385.650 ;
        RECT 2798.950 1341.450 2799.250 1385.350 ;
        RECT 2798.030 1341.150 2799.250 1341.450 ;
        RECT 2796.190 1062.350 2797.410 1062.650 ;
        RECT 2797.110 1038.850 2797.410 1062.350 ;
        RECT 2796.190 1038.550 2797.410 1038.850 ;
        RECT 2796.190 182.490 2796.490 1038.550 ;
        RECT 6.310 181.310 7.490 182.490 ;
        RECT 2795.750 181.310 2796.930 182.490 ;
        RECT 6.750 148.745 7.050 181.310 ;
        RECT 2798.030 179.090 2798.330 1341.150 ;
        RECT 8.150 177.910 9.330 179.090 ;
        RECT 2797.590 177.910 2798.770 179.090 ;
        RECT 8.590 168.450 8.890 177.910 ;
        RECT 7.670 168.150 8.890 168.450 ;
        RECT 7.670 166.425 7.970 168.150 ;
        RECT 7.655 166.095 7.985 166.425 ;
        RECT 6.735 148.415 7.065 148.745 ;
      LAYER met5 ;
        RECT 2795.540 3329.500 2802.660 3331.100 ;
        RECT 6.100 181.100 2797.140 182.700 ;
        RECT 7.940 177.700 2798.980 179.300 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 490.965 0.255 491.135 2.975 ;
        RECT 562.265 0.595 562.435 2.975 ;
        RECT 750.405 2.635 750.575 3.315 ;
        RECT 878.285 3.145 881.215 3.315 ;
        RECT 757.305 2.635 757.475 2.975 ;
        RECT 878.285 2.805 878.455 3.145 ;
        RECT 1677.305 2.805 1678.855 2.975 ;
        RECT 1736.645 2.805 1737.735 2.975 ;
        RECT 2367.305 2.805 2367.935 2.975 ;
        RECT 750.405 2.465 757.475 2.635 ;
        RECT 559.965 0.425 562.435 0.595 ;
        RECT 559.965 0.255 560.135 0.425 ;
        RECT 490.965 0.085 560.135 0.255 ;
      LAYER mcon ;
        RECT 750.405 3.145 750.575 3.315 ;
        RECT 490.965 2.805 491.135 2.975 ;
        RECT 562.265 2.805 562.435 2.975 ;
        RECT 881.045 3.145 881.215 3.315 ;
        RECT 757.305 2.805 757.475 2.975 ;
        RECT 1678.685 2.805 1678.855 2.975 ;
        RECT 1737.565 2.805 1737.735 2.975 ;
        RECT 2367.765 2.805 2367.935 2.975 ;
      LAYER met1 ;
        RECT 750.345 3.300 750.635 3.345 ;
        RECT 880.985 3.300 881.275 3.345 ;
        RECT 749.040 3.160 750.635 3.300 ;
        RECT 264.110 2.960 264.430 3.020 ;
        RECT 490.905 2.960 491.195 3.005 ;
        RECT 264.110 2.820 466.740 2.960 ;
        RECT 264.110 2.760 264.430 2.820 ;
        RECT 466.600 2.620 466.740 2.820 ;
        RECT 471.200 2.820 491.195 2.960 ;
        RECT 471.200 2.620 471.340 2.820 ;
        RECT 490.905 2.775 491.195 2.820 ;
        RECT 562.205 2.960 562.495 3.005 ;
        RECT 749.040 2.960 749.180 3.160 ;
        RECT 750.345 3.115 750.635 3.160 ;
        RECT 784.000 3.160 785.060 3.300 ;
        RECT 562.205 2.820 749.180 2.960 ;
        RECT 757.245 2.960 757.535 3.005 ;
        RECT 757.245 2.820 783.220 2.960 ;
        RECT 562.205 2.775 562.495 2.820 ;
        RECT 757.245 2.775 757.535 2.820 ;
        RECT 466.600 2.480 471.340 2.620 ;
        RECT 783.080 2.620 783.220 2.820 ;
        RECT 784.000 2.620 784.140 3.160 ;
        RECT 784.920 2.960 785.060 3.160 ;
        RECT 880.985 3.160 883.040 3.300 ;
        RECT 880.985 3.115 881.275 3.160 ;
        RECT 878.225 2.960 878.515 3.005 ;
        RECT 784.920 2.820 878.515 2.960 ;
        RECT 882.900 2.960 883.040 3.160 ;
        RECT 1677.245 2.960 1677.535 3.005 ;
        RECT 882.900 2.820 918.920 2.960 ;
        RECT 878.225 2.775 878.515 2.820 ;
        RECT 783.080 2.480 784.140 2.620 ;
        RECT 918.780 2.620 918.920 2.820 ;
        RECT 919.700 2.820 1677.535 2.960 ;
        RECT 919.700 2.620 919.840 2.820 ;
        RECT 1677.245 2.775 1677.535 2.820 ;
        RECT 1678.625 2.960 1678.915 3.005 ;
        RECT 1736.585 2.960 1736.875 3.005 ;
        RECT 1678.625 2.820 1736.875 2.960 ;
        RECT 1678.625 2.775 1678.915 2.820 ;
        RECT 1736.585 2.775 1736.875 2.820 ;
        RECT 1737.505 2.960 1737.795 3.005 ;
        RECT 2367.245 2.960 2367.535 3.005 ;
        RECT 1737.505 2.820 2367.535 2.960 ;
        RECT 1737.505 2.775 1737.795 2.820 ;
        RECT 2367.245 2.775 2367.535 2.820 ;
        RECT 2367.705 2.960 2367.995 3.005 ;
        RECT 2403.570 2.960 2403.890 3.020 ;
        RECT 2367.705 2.820 2403.890 2.960 ;
        RECT 2367.705 2.775 2367.995 2.820 ;
        RECT 2403.570 2.760 2403.890 2.820 ;
        RECT 918.780 2.480 919.840 2.620 ;
      LAYER via ;
        RECT 264.140 2.760 264.400 3.020 ;
        RECT 2403.600 2.760 2403.860 3.020 ;
      LAYER met2 ;
        RECT 2403.530 5.000 2403.810 9.000 ;
        RECT 2403.660 3.050 2403.800 5.000 ;
        RECT 264.140 2.730 264.400 3.050 ;
        RECT 2403.600 2.730 2403.860 3.050 ;
        RECT 264.200 2.400 264.340 2.730 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1648.325 7.225 1648.955 7.395 ;
        RECT 1648.785 6.205 1648.955 7.225 ;
        RECT 1679.145 6.205 1680.695 6.375 ;
        RECT 365.845 3.485 366.935 3.655 ;
        RECT 365.845 3.145 366.015 3.485 ;
        RECT 366.765 2.465 366.935 3.485 ;
        RECT 466.125 2.465 471.815 2.635 ;
        RECT 1680.525 2.465 1680.695 6.205 ;
        RECT 559.045 2.125 561.515 2.295 ;
        RECT 676.805 2.125 724.355 2.295 ;
        RECT 917.385 2.125 918.475 2.295 ;
        RECT 967.065 2.125 980.575 2.295 ;
        RECT 918.305 1.785 918.475 2.125 ;
        RECT 980.405 0.935 980.575 2.125 ;
        RECT 996.965 0.935 997.135 2.295 ;
        RECT 1015.365 2.125 1062.455 2.295 ;
        RECT 1208.105 2.125 1255.195 2.295 ;
        RECT 1256.865 2.125 1303.495 2.295 ;
        RECT 1304.705 2.125 1325.575 2.295 ;
        RECT 1344.725 2.125 1351.795 2.295 ;
        RECT 1353.005 2.125 1400.095 2.295 ;
        RECT 1401.305 2.125 1408.375 2.295 ;
        RECT 1427.525 2.125 1429.075 2.295 ;
        RECT 1449.605 2.125 1484.275 2.295 ;
        RECT 1484.105 1.275 1484.275 2.125 ;
        RECT 1485.025 1.275 1485.195 2.295 ;
        RECT 1546.205 2.125 1593.295 2.295 ;
        RECT 1687.425 1.955 1687.595 2.635 ;
        RECT 1689.725 1.955 1689.895 2.295 ;
        RECT 1863.145 2.125 1863.775 2.295 ;
        RECT 2297.845 2.125 2298.935 2.295 ;
        RECT 2367.305 2.125 2367.935 2.295 ;
        RECT 1687.425 1.785 1689.895 1.955 ;
        RECT 1863.605 1.955 1863.775 2.125 ;
        RECT 1863.605 1.785 1864.235 1.955 ;
        RECT 1484.105 1.105 1485.195 1.275 ;
        RECT 980.405 0.765 997.135 0.935 ;
      LAYER mcon ;
        RECT 471.645 2.465 471.815 2.635 ;
        RECT 1687.425 2.465 1687.595 2.635 ;
        RECT 561.345 2.125 561.515 2.295 ;
        RECT 724.185 2.125 724.355 2.295 ;
        RECT 996.965 2.125 997.135 2.295 ;
        RECT 1062.285 2.125 1062.455 2.295 ;
        RECT 1255.025 2.125 1255.195 2.295 ;
        RECT 1303.325 2.125 1303.495 2.295 ;
        RECT 1325.405 2.125 1325.575 2.295 ;
        RECT 1351.625 2.125 1351.795 2.295 ;
        RECT 1399.925 2.125 1400.095 2.295 ;
        RECT 1408.205 2.125 1408.375 2.295 ;
        RECT 1428.905 2.125 1429.075 2.295 ;
        RECT 1485.025 2.125 1485.195 2.295 ;
        RECT 1593.125 2.125 1593.295 2.295 ;
        RECT 1689.725 2.125 1689.895 2.295 ;
        RECT 2298.765 2.125 2298.935 2.295 ;
        RECT 2367.765 2.125 2367.935 2.295 ;
        RECT 1864.065 1.785 1864.235 1.955 ;
      LAYER met1 ;
        RECT 1601.330 7.380 1601.650 7.440 ;
        RECT 1648.265 7.380 1648.555 7.425 ;
        RECT 1601.330 7.240 1648.555 7.380 ;
        RECT 1601.330 7.180 1601.650 7.240 ;
        RECT 1648.265 7.195 1648.555 7.240 ;
        RECT 1648.725 6.360 1649.015 6.405 ;
        RECT 1679.085 6.360 1679.375 6.405 ;
        RECT 1648.725 6.220 1679.375 6.360 ;
        RECT 1648.725 6.175 1649.015 6.220 ;
        RECT 1679.085 6.175 1679.375 6.220 ;
        RECT 299.990 3.300 300.310 3.360 ;
        RECT 365.785 3.300 366.075 3.345 ;
        RECT 299.990 3.160 366.075 3.300 ;
        RECT 299.990 3.100 300.310 3.160 ;
        RECT 365.785 3.115 366.075 3.160 ;
        RECT 366.705 2.620 366.995 2.665 ;
        RECT 466.065 2.620 466.355 2.665 ;
        RECT 366.705 2.480 466.355 2.620 ;
        RECT 366.705 2.435 366.995 2.480 ;
        RECT 466.065 2.435 466.355 2.480 ;
        RECT 471.585 2.620 471.875 2.665 ;
        RECT 1680.465 2.620 1680.755 2.665 ;
        RECT 1687.365 2.620 1687.655 2.665 ;
        RECT 471.585 2.480 486.520 2.620 ;
        RECT 471.585 2.435 471.875 2.480 ;
        RECT 486.380 2.280 486.520 2.480 ;
        RECT 1680.465 2.480 1687.655 2.620 ;
        RECT 1680.465 2.435 1680.755 2.480 ;
        RECT 1687.365 2.435 1687.655 2.480 ;
        RECT 558.985 2.280 559.275 2.325 ;
        RECT 486.380 2.140 559.275 2.280 ;
        RECT 558.985 2.095 559.275 2.140 ;
        RECT 561.285 2.280 561.575 2.325 ;
        RECT 676.745 2.280 677.035 2.325 ;
        RECT 561.285 2.140 677.035 2.280 ;
        RECT 561.285 2.095 561.575 2.140 ;
        RECT 676.745 2.095 677.035 2.140 ;
        RECT 724.125 2.280 724.415 2.325 ;
        RECT 917.325 2.280 917.615 2.325 ;
        RECT 967.005 2.280 967.295 2.325 ;
        RECT 724.125 2.140 917.615 2.280 ;
        RECT 724.125 2.095 724.415 2.140 ;
        RECT 917.325 2.095 917.615 2.140 ;
        RECT 918.320 2.140 967.295 2.280 ;
        RECT 918.320 1.985 918.460 2.140 ;
        RECT 967.005 2.095 967.295 2.140 ;
        RECT 996.905 2.280 997.195 2.325 ;
        RECT 1015.305 2.280 1015.595 2.325 ;
        RECT 996.905 2.140 1015.595 2.280 ;
        RECT 996.905 2.095 997.195 2.140 ;
        RECT 1015.305 2.095 1015.595 2.140 ;
        RECT 1062.225 2.280 1062.515 2.325 ;
        RECT 1208.045 2.280 1208.335 2.325 ;
        RECT 1062.225 2.140 1208.335 2.280 ;
        RECT 1062.225 2.095 1062.515 2.140 ;
        RECT 1208.045 2.095 1208.335 2.140 ;
        RECT 1254.965 2.280 1255.255 2.325 ;
        RECT 1256.805 2.280 1257.095 2.325 ;
        RECT 1254.965 2.140 1257.095 2.280 ;
        RECT 1254.965 2.095 1255.255 2.140 ;
        RECT 1256.805 2.095 1257.095 2.140 ;
        RECT 1303.265 2.280 1303.555 2.325 ;
        RECT 1304.645 2.280 1304.935 2.325 ;
        RECT 1303.265 2.140 1304.935 2.280 ;
        RECT 1303.265 2.095 1303.555 2.140 ;
        RECT 1304.645 2.095 1304.935 2.140 ;
        RECT 1325.345 2.280 1325.635 2.325 ;
        RECT 1344.665 2.280 1344.955 2.325 ;
        RECT 1325.345 2.140 1344.955 2.280 ;
        RECT 1325.345 2.095 1325.635 2.140 ;
        RECT 1344.665 2.095 1344.955 2.140 ;
        RECT 1351.565 2.280 1351.855 2.325 ;
        RECT 1352.945 2.280 1353.235 2.325 ;
        RECT 1351.565 2.140 1353.235 2.280 ;
        RECT 1351.565 2.095 1351.855 2.140 ;
        RECT 1352.945 2.095 1353.235 2.140 ;
        RECT 1399.865 2.280 1400.155 2.325 ;
        RECT 1401.245 2.280 1401.535 2.325 ;
        RECT 1399.865 2.140 1401.535 2.280 ;
        RECT 1399.865 2.095 1400.155 2.140 ;
        RECT 1401.245 2.095 1401.535 2.140 ;
        RECT 1408.145 2.280 1408.435 2.325 ;
        RECT 1427.465 2.280 1427.755 2.325 ;
        RECT 1408.145 2.140 1427.755 2.280 ;
        RECT 1408.145 2.095 1408.435 2.140 ;
        RECT 1427.465 2.095 1427.755 2.140 ;
        RECT 1428.845 2.280 1429.135 2.325 ;
        RECT 1449.545 2.280 1449.835 2.325 ;
        RECT 1428.845 2.140 1449.835 2.280 ;
        RECT 1428.845 2.095 1429.135 2.140 ;
        RECT 1449.545 2.095 1449.835 2.140 ;
        RECT 1484.965 2.280 1485.255 2.325 ;
        RECT 1546.145 2.280 1546.435 2.325 ;
        RECT 1484.965 2.140 1546.435 2.280 ;
        RECT 1484.965 2.095 1485.255 2.140 ;
        RECT 1546.145 2.095 1546.435 2.140 ;
        RECT 1593.065 2.280 1593.355 2.325 ;
        RECT 1594.430 2.280 1594.750 2.340 ;
        RECT 1593.065 2.140 1594.750 2.280 ;
        RECT 1593.065 2.095 1593.355 2.140 ;
        RECT 1594.430 2.080 1594.750 2.140 ;
        RECT 1689.665 2.280 1689.955 2.325 ;
        RECT 1863.085 2.280 1863.375 2.325 ;
        RECT 2297.785 2.280 2298.075 2.325 ;
        RECT 1689.665 2.140 1863.375 2.280 ;
        RECT 1689.665 2.095 1689.955 2.140 ;
        RECT 1863.085 2.095 1863.375 2.140 ;
        RECT 1864.080 2.140 2298.075 2.280 ;
        RECT 1864.080 1.985 1864.220 2.140 ;
        RECT 2297.785 2.095 2298.075 2.140 ;
        RECT 2298.705 2.280 2298.995 2.325 ;
        RECT 2367.245 2.280 2367.535 2.325 ;
        RECT 2298.705 2.140 2367.535 2.280 ;
        RECT 2298.705 2.095 2298.995 2.140 ;
        RECT 2367.245 2.095 2367.535 2.140 ;
        RECT 2367.705 2.280 2367.995 2.325 ;
        RECT 2449.110 2.280 2449.430 2.340 ;
        RECT 2367.705 2.140 2449.430 2.280 ;
        RECT 2367.705 2.095 2367.995 2.140 ;
        RECT 2449.110 2.080 2449.430 2.140 ;
        RECT 918.245 1.755 918.535 1.985 ;
        RECT 1864.005 1.755 1864.295 1.985 ;
      LAYER via ;
        RECT 1601.360 7.180 1601.620 7.440 ;
        RECT 300.020 3.100 300.280 3.360 ;
        RECT 1594.460 2.080 1594.720 2.340 ;
        RECT 2449.140 2.080 2449.400 2.340 ;
      LAYER met2 ;
        RECT 1601.360 7.380 1601.620 7.470 ;
        RECT 1599.120 7.240 1601.620 7.380 ;
        RECT 300.020 3.070 300.280 3.390 ;
        RECT 1599.120 3.130 1599.260 7.240 ;
        RECT 1601.360 7.150 1601.620 7.240 ;
        RECT 2450.910 5.170 2451.190 9.000 ;
        RECT 300.080 2.400 300.220 3.070 ;
        RECT 1594.520 2.990 1599.260 3.130 ;
        RECT 2449.200 5.030 2451.190 5.170 ;
        RECT 299.870 -4.800 300.430 2.400 ;
        RECT 1594.520 2.370 1594.660 2.990 ;
        RECT 2449.200 2.370 2449.340 5.030 ;
        RECT 2450.910 5.000 2451.190 5.030 ;
        RECT 1594.460 2.050 1594.720 2.370 ;
        RECT 2449.140 2.050 2449.400 2.370 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 364.005 4.165 365.555 4.335 ;
        RECT 365.385 1.445 365.555 4.165 ;
        RECT 1770.685 1.615 1770.855 6.035 ;
        RECT 1428.905 1.275 1429.075 1.615 ;
        RECT 1429.825 1.445 1446.095 1.615 ;
        RECT 1759.645 1.445 1770.855 1.615 ;
        RECT 1779.885 1.445 1780.055 6.035 ;
        RECT 2367.305 1.445 2368.855 1.615 ;
        RECT 1429.825 1.275 1429.995 1.445 ;
        RECT 1428.905 1.105 1429.995 1.275 ;
      LAYER mcon ;
        RECT 1770.685 5.865 1770.855 6.035 ;
        RECT 1428.905 1.445 1429.075 1.615 ;
        RECT 1445.925 1.445 1446.095 1.615 ;
        RECT 1779.885 5.865 1780.055 6.035 ;
        RECT 2368.685 1.445 2368.855 1.615 ;
      LAYER met1 ;
        RECT 1770.625 6.020 1770.915 6.065 ;
        RECT 1779.825 6.020 1780.115 6.065 ;
        RECT 1770.625 5.880 1780.115 6.020 ;
        RECT 1770.625 5.835 1770.915 5.880 ;
        RECT 1779.825 5.835 1780.115 5.880 ;
        RECT 319.310 4.320 319.630 4.380 ;
        RECT 363.945 4.320 364.235 4.365 ;
        RECT 319.310 4.180 364.235 4.320 ;
        RECT 319.310 4.120 319.630 4.180 ;
        RECT 363.945 4.135 364.235 4.180 ;
        RECT 1842.460 1.800 1862.380 1.940 ;
        RECT 365.325 1.600 365.615 1.645 ;
        RECT 1428.845 1.600 1429.135 1.645 ;
        RECT 365.325 1.460 534.820 1.600 ;
        RECT 365.325 1.415 365.615 1.460 ;
        RECT 534.680 1.260 534.820 1.460 ;
        RECT 560.900 1.460 918.460 1.600 ;
        RECT 560.900 1.260 561.040 1.460 ;
        RECT 534.680 1.120 561.040 1.260 ;
        RECT 918.320 1.260 918.460 1.460 ;
        RECT 920.620 1.460 1429.135 1.600 ;
        RECT 920.620 1.260 920.760 1.460 ;
        RECT 1428.845 1.415 1429.135 1.460 ;
        RECT 1445.865 1.600 1446.155 1.645 ;
        RECT 1759.585 1.600 1759.875 1.645 ;
        RECT 1445.865 1.460 1759.875 1.600 ;
        RECT 1445.865 1.415 1446.155 1.460 ;
        RECT 1759.585 1.415 1759.875 1.460 ;
        RECT 1779.825 1.600 1780.115 1.645 ;
        RECT 1842.460 1.600 1842.600 1.800 ;
        RECT 1779.825 1.460 1842.600 1.600 ;
        RECT 1862.240 1.600 1862.380 1.800 ;
        RECT 2367.245 1.600 2367.535 1.645 ;
        RECT 1862.240 1.460 2367.535 1.600 ;
        RECT 1779.825 1.415 1780.115 1.460 ;
        RECT 2367.245 1.415 2367.535 1.460 ;
        RECT 2368.625 1.600 2368.915 1.645 ;
        RECT 2498.330 1.600 2498.650 1.660 ;
        RECT 2368.625 1.460 2498.650 1.600 ;
        RECT 2368.625 1.415 2368.915 1.460 ;
        RECT 2498.330 1.400 2498.650 1.460 ;
        RECT 918.320 1.120 920.760 1.260 ;
      LAYER via ;
        RECT 319.340 4.120 319.600 4.380 ;
        RECT 2498.360 1.400 2498.620 1.660 ;
      LAYER met2 ;
        RECT 2498.290 5.000 2498.570 9.000 ;
        RECT 319.340 4.090 319.600 4.410 ;
        RECT 319.400 3.810 319.540 4.090 ;
        RECT 318.020 3.670 319.540 3.810 ;
        RECT 318.020 2.400 318.160 3.670 ;
        RECT 317.810 -4.800 318.370 2.400 ;
        RECT 2498.420 1.690 2498.560 5.000 ;
        RECT 2498.360 1.370 2498.620 1.690 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 534.205 1.445 535.295 1.615 ;
        RECT 559.965 1.445 561.515 1.615 ;
        RECT 367.225 0.935 367.395 1.275 ;
        RECT 368.605 0.935 368.775 1.275 ;
        RECT 534.205 1.105 534.375 1.445 ;
        RECT 561.345 1.105 561.515 1.445 ;
        RECT 756.385 1.105 759.315 1.275 ;
        RECT 917.845 1.105 921.235 1.275 ;
        RECT 1862.685 1.105 1865.155 1.275 ;
        RECT 367.225 0.765 368.775 0.935 ;
      LAYER mcon ;
        RECT 535.125 1.445 535.295 1.615 ;
        RECT 367.225 1.105 367.395 1.275 ;
        RECT 368.605 1.105 368.775 1.275 ;
        RECT 759.145 1.105 759.315 1.275 ;
        RECT 921.065 1.105 921.235 1.275 ;
        RECT 1864.985 1.105 1865.155 1.275 ;
      LAYER met1 ;
        RECT 535.065 1.600 535.355 1.645 ;
        RECT 559.905 1.600 560.195 1.645 ;
        RECT 535.065 1.460 560.195 1.600 ;
        RECT 535.065 1.415 535.355 1.460 ;
        RECT 559.905 1.415 560.195 1.460 ;
        RECT 336.790 1.260 337.110 1.320 ;
        RECT 367.165 1.260 367.455 1.305 ;
        RECT 336.790 1.120 367.455 1.260 ;
        RECT 336.790 1.060 337.110 1.120 ;
        RECT 367.165 1.075 367.455 1.120 ;
        RECT 368.545 1.260 368.835 1.305 ;
        RECT 534.145 1.260 534.435 1.305 ;
        RECT 368.545 1.120 534.435 1.260 ;
        RECT 368.545 1.075 368.835 1.120 ;
        RECT 534.145 1.075 534.435 1.120 ;
        RECT 561.285 1.260 561.575 1.305 ;
        RECT 756.325 1.260 756.615 1.305 ;
        RECT 561.285 1.120 756.615 1.260 ;
        RECT 561.285 1.075 561.575 1.120 ;
        RECT 756.325 1.075 756.615 1.120 ;
        RECT 759.085 1.260 759.375 1.305 ;
        RECT 917.785 1.260 918.075 1.305 ;
        RECT 759.085 1.120 918.075 1.260 ;
        RECT 759.085 1.075 759.375 1.120 ;
        RECT 917.785 1.075 918.075 1.120 ;
        RECT 921.005 1.260 921.295 1.305 ;
        RECT 1862.625 1.260 1862.915 1.305 ;
        RECT 921.005 1.120 1862.915 1.260 ;
        RECT 921.005 1.075 921.295 1.120 ;
        RECT 1862.625 1.075 1862.915 1.120 ;
        RECT 1864.925 1.260 1865.215 1.305 ;
        RECT 2546.170 1.260 2546.490 1.320 ;
        RECT 1864.925 1.120 2546.490 1.260 ;
        RECT 1864.925 1.075 1865.215 1.120 ;
        RECT 2546.170 1.060 2546.490 1.120 ;
      LAYER via ;
        RECT 336.820 1.060 337.080 1.320 ;
        RECT 2546.200 1.060 2546.460 1.320 ;
      LAYER met2 ;
        RECT 2546.130 5.000 2546.410 9.000 ;
        RECT 335.960 2.990 337.020 3.130 ;
        RECT 335.960 2.400 336.100 2.990 ;
        RECT 335.750 -4.800 336.310 2.400 ;
        RECT 336.880 1.350 337.020 2.990 ;
        RECT 2546.260 1.350 2546.400 5.000 ;
        RECT 336.820 1.030 337.080 1.350 ;
        RECT 2546.200 1.030 2546.460 1.350 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2850.305 2317.865 2850.475 2326.195 ;
        RECT 2849.845 1949.305 2850.015 1968.515 ;
        RECT 2849.845 1744.625 2850.015 1763.155 ;
        RECT 2850.305 1624.945 2850.475 1648.575 ;
        RECT 2850.765 1524.985 2850.935 1603.695 ;
        RECT 2852.605 1480.445 2852.775 1524.815 ;
        RECT 2851.225 1351.585 2851.395 1417.375 ;
        RECT 2851.225 1297.865 2851.395 1320.135 ;
        RECT 2849.845 1229.865 2850.015 1273.895 ;
        RECT 2851.225 1218.305 2851.395 1230.035 ;
        RECT 2852.605 1146.225 2852.775 1168.495 ;
        RECT 2850.765 809.795 2850.935 890.375 ;
        RECT 2851.685 890.205 2851.855 960.415 ;
        RECT 2850.765 809.625 2851.395 809.795 ;
        RECT 2851.225 767.125 2851.395 809.625 ;
        RECT 2849.385 381.565 2850.015 381.735 ;
        RECT 2849.385 294.185 2849.555 381.565 ;
        RECT 2850.765 116.025 2850.935 198.815 ;
        RECT 2851.685 198.645 2851.855 209.015 ;
        RECT 809.285 10.285 850.855 10.455 ;
        RECT 797.785 5.015 797.955 6.375 ;
        RECT 807.445 5.695 807.615 6.375 ;
        RECT 809.285 5.695 809.455 10.285 ;
        RECT 850.685 10.115 850.855 10.285 ;
        RECT 850.685 9.945 852.695 10.115 ;
        RECT 852.525 8.755 852.695 9.945 ;
        RECT 869.545 9.605 891.795 9.775 ;
        RECT 869.545 8.755 869.715 9.605 ;
        RECT 891.625 9.095 891.795 9.605 ;
        RECT 891.625 8.925 895.475 9.095 ;
        RECT 852.525 8.585 869.715 8.755 ;
        RECT 807.445 5.525 809.455 5.695 ;
        RECT 797.785 4.845 799.335 5.015 ;
        RECT 379.645 3.145 379.815 4.335 ;
        RECT 411.385 2.975 411.555 3.315 ;
        RECT 413.685 2.975 413.855 3.315 ;
        RECT 460.605 3.145 462.615 3.315 ;
        RECT 411.385 2.805 413.855 2.975 ;
        RECT 607.345 2.295 607.515 3.315 ;
        RECT 623.445 2.295 623.615 3.315 ;
        RECT 607.345 2.125 623.615 2.295 ;
        RECT 748.565 0.935 748.735 3.315 ;
        RECT 767.425 1.785 769.435 1.955 ;
        RECT 767.425 1.275 767.595 1.785 ;
        RECT 760.065 1.105 767.595 1.275 ;
        RECT 760.065 0.935 760.235 1.105 ;
        RECT 748.565 0.765 760.235 0.935 ;
        RECT 772.945 0.935 773.115 1.955 ;
        RECT 799.165 0.935 799.335 4.845 ;
        RECT 895.305 4.335 895.475 8.925 ;
        RECT 902.205 8.925 903.295 9.095 ;
        RECT 898.525 4.335 898.695 8.755 ;
        RECT 902.205 8.585 902.375 8.925 ;
        RECT 903.125 5.865 903.295 8.925 ;
        RECT 920.145 7.565 920.775 7.735 ;
        RECT 919.225 5.695 919.395 6.035 ;
        RECT 920.145 5.695 920.315 7.565 ;
        RECT 919.225 5.525 920.315 5.695 ;
        RECT 947.285 5.355 947.455 7.735 ;
        RECT 1121.625 6.545 1123.175 6.715 ;
        RECT 1127.145 6.545 1129.155 6.715 ;
        RECT 954.645 5.865 955.275 6.035 ;
        RECT 954.645 5.355 954.815 5.865 ;
        RECT 1120.705 5.695 1120.875 6.035 ;
        RECT 1121.625 5.695 1121.795 6.545 ;
        RECT 1120.705 5.525 1121.795 5.695 ;
        RECT 1128.985 5.695 1129.155 6.545 ;
        RECT 1141.865 5.695 1142.035 6.035 ;
        RECT 1183.265 5.865 1183.435 7.395 ;
        RECT 1409.125 6.205 1410.675 6.375 ;
        RECT 1128.985 5.525 1142.035 5.695 ;
        RECT 947.285 5.185 954.815 5.355 ;
        RECT 895.305 4.165 898.695 4.335 ;
        RECT 1255.945 2.635 1256.115 6.035 ;
        RECT 1298.265 5.865 1303.955 6.035 ;
        RECT 1255.945 2.465 1258.415 2.635 ;
        RECT 1298.265 2.465 1298.435 5.865 ;
        RECT 1400.385 3.995 1400.555 6.035 ;
        RECT 1407.745 5.695 1407.915 6.035 ;
        RECT 1409.125 5.695 1409.295 6.205 ;
        RECT 1410.505 5.865 1410.675 6.205 ;
        RECT 1635.445 6.035 1635.615 6.375 ;
        RECT 1503.425 5.865 1504.055 6.035 ;
        RECT 1634.525 5.865 1635.615 6.035 ;
        RECT 1407.745 5.525 1409.295 5.695 ;
        RECT 1399.465 3.825 1400.555 3.995 ;
        RECT 1399.465 2.635 1399.635 3.825 ;
        RECT 1399.005 2.465 1399.635 2.635 ;
        RECT 1487.325 2.805 1488.415 2.975 ;
        RECT 1487.325 2.465 1487.495 2.805 ;
        RECT 1488.245 1.785 1488.415 2.805 ;
        RECT 1503.425 1.785 1503.595 5.865 ;
        RECT 1637.285 2.635 1637.455 6.375 ;
        RECT 1637.285 2.465 1640.215 2.635 ;
        RECT 1677.765 2.465 1678.855 2.635 ;
        RECT 1742.625 2.465 1742.795 6.035 ;
        RECT 1763.325 2.465 1763.495 5.355 ;
        RECT 1785.405 5.185 1785.575 6.035 ;
        RECT 1835.085 5.865 1835.715 6.035 ;
        RECT 1841.985 5.865 1842.155 9.095 ;
        RECT 1874.185 5.865 1874.355 9.095 ;
        RECT 1932.605 5.865 1932.775 7.395 ;
        RECT 1956.065 5.865 1956.235 7.395 ;
        RECT 1678.685 2.125 1678.855 2.465 ;
        RECT 772.945 0.765 799.335 0.935 ;
      LAYER mcon ;
        RECT 2850.305 2326.025 2850.475 2326.195 ;
        RECT 2849.845 1968.345 2850.015 1968.515 ;
        RECT 2849.845 1762.985 2850.015 1763.155 ;
        RECT 2850.305 1648.405 2850.475 1648.575 ;
        RECT 2850.765 1603.525 2850.935 1603.695 ;
        RECT 2852.605 1524.645 2852.775 1524.815 ;
        RECT 2851.225 1417.205 2851.395 1417.375 ;
        RECT 2851.225 1319.965 2851.395 1320.135 ;
        RECT 2849.845 1273.725 2850.015 1273.895 ;
        RECT 2851.225 1229.865 2851.395 1230.035 ;
        RECT 2852.605 1168.325 2852.775 1168.495 ;
        RECT 2851.685 960.245 2851.855 960.415 ;
        RECT 2850.765 890.205 2850.935 890.375 ;
        RECT 2849.845 381.565 2850.015 381.735 ;
        RECT 2851.685 208.845 2851.855 209.015 ;
        RECT 2850.765 198.645 2850.935 198.815 ;
        RECT 797.785 6.205 797.955 6.375 ;
        RECT 807.445 6.205 807.615 6.375 ;
        RECT 379.645 4.165 379.815 4.335 ;
        RECT 411.385 3.145 411.555 3.315 ;
        RECT 413.685 3.145 413.855 3.315 ;
        RECT 462.445 3.145 462.615 3.315 ;
        RECT 607.345 3.145 607.515 3.315 ;
        RECT 623.445 3.145 623.615 3.315 ;
        RECT 748.565 3.145 748.735 3.315 ;
        RECT 769.265 1.785 769.435 1.955 ;
        RECT 772.945 1.785 773.115 1.955 ;
        RECT 898.525 8.585 898.695 8.755 ;
        RECT 1841.985 8.925 1842.155 9.095 ;
        RECT 920.605 7.565 920.775 7.735 ;
        RECT 947.285 7.565 947.455 7.735 ;
        RECT 919.225 5.865 919.395 6.035 ;
        RECT 1183.265 7.225 1183.435 7.395 ;
        RECT 1123.005 6.545 1123.175 6.715 ;
        RECT 955.105 5.865 955.275 6.035 ;
        RECT 1120.705 5.865 1120.875 6.035 ;
        RECT 1141.865 5.865 1142.035 6.035 ;
        RECT 1255.945 5.865 1256.115 6.035 ;
        RECT 1303.785 5.865 1303.955 6.035 ;
        RECT 1400.385 5.865 1400.555 6.035 ;
        RECT 1407.745 5.865 1407.915 6.035 ;
        RECT 1635.445 6.205 1635.615 6.375 ;
        RECT 1503.885 5.865 1504.055 6.035 ;
        RECT 1637.285 6.205 1637.455 6.375 ;
        RECT 1258.245 2.465 1258.415 2.635 ;
        RECT 1742.625 5.865 1742.795 6.035 ;
        RECT 1785.405 5.865 1785.575 6.035 ;
        RECT 1835.545 5.865 1835.715 6.035 ;
        RECT 1874.185 8.925 1874.355 9.095 ;
        RECT 1932.605 7.225 1932.775 7.395 ;
        RECT 1956.065 7.225 1956.235 7.395 ;
        RECT 1640.045 2.465 1640.215 2.635 ;
        RECT 1763.325 5.185 1763.495 5.355 ;
      LAYER met1 ;
        RECT 2849.770 2759.340 2850.090 2759.400 ;
        RECT 2863.570 2759.340 2863.890 2759.400 ;
        RECT 2849.770 2759.200 2863.890 2759.340 ;
        RECT 2849.770 2759.140 2850.090 2759.200 ;
        RECT 2863.570 2759.140 2863.890 2759.200 ;
        RECT 2849.770 2326.180 2850.090 2326.240 ;
        RECT 2850.245 2326.180 2850.535 2326.225 ;
        RECT 2849.770 2326.040 2850.535 2326.180 ;
        RECT 2849.770 2325.980 2850.090 2326.040 ;
        RECT 2850.245 2325.995 2850.535 2326.040 ;
        RECT 2849.770 2318.020 2850.090 2318.080 ;
        RECT 2850.245 2318.020 2850.535 2318.065 ;
        RECT 2849.770 2317.880 2850.535 2318.020 ;
        RECT 2849.770 2317.820 2850.090 2317.880 ;
        RECT 2850.245 2317.835 2850.535 2317.880 ;
        RECT 2849.770 1968.500 2850.090 1968.560 ;
        RECT 2849.575 1968.360 2850.090 1968.500 ;
        RECT 2849.770 1968.300 2850.090 1968.360 ;
        RECT 2849.770 1949.460 2850.090 1949.520 ;
        RECT 2849.575 1949.320 2850.090 1949.460 ;
        RECT 2849.770 1949.260 2850.090 1949.320 ;
        RECT 2849.770 1840.320 2850.090 1840.380 ;
        RECT 2850.690 1840.320 2851.010 1840.380 ;
        RECT 2849.770 1840.180 2851.010 1840.320 ;
        RECT 2849.770 1840.120 2850.090 1840.180 ;
        RECT 2850.690 1840.120 2851.010 1840.180 ;
        RECT 2850.230 1790.480 2850.550 1790.740 ;
        RECT 2850.320 1789.720 2850.460 1790.480 ;
        RECT 2850.230 1789.460 2850.550 1789.720 ;
        RECT 2849.785 1763.140 2850.075 1763.185 ;
        RECT 2850.230 1763.140 2850.550 1763.200 ;
        RECT 2849.785 1763.000 2850.550 1763.140 ;
        RECT 2849.785 1762.955 2850.075 1763.000 ;
        RECT 2850.230 1762.940 2850.550 1763.000 ;
        RECT 2849.770 1744.780 2850.090 1744.840 ;
        RECT 2849.575 1744.640 2850.090 1744.780 ;
        RECT 2849.770 1744.580 2850.090 1744.640 ;
        RECT 2849.770 1648.560 2850.090 1648.620 ;
        RECT 2850.245 1648.560 2850.535 1648.605 ;
        RECT 2849.770 1648.420 2850.535 1648.560 ;
        RECT 2849.770 1648.360 2850.090 1648.420 ;
        RECT 2850.245 1648.375 2850.535 1648.420 ;
        RECT 2850.230 1625.100 2850.550 1625.160 ;
        RECT 2850.035 1624.960 2850.550 1625.100 ;
        RECT 2850.230 1624.900 2850.550 1624.960 ;
        RECT 2850.230 1603.680 2850.550 1603.740 ;
        RECT 2850.705 1603.680 2850.995 1603.725 ;
        RECT 2850.230 1603.540 2850.995 1603.680 ;
        RECT 2850.230 1603.480 2850.550 1603.540 ;
        RECT 2850.705 1603.495 2850.995 1603.540 ;
        RECT 2850.705 1525.140 2850.995 1525.185 ;
        RECT 2849.400 1525.000 2850.995 1525.140 ;
        RECT 2849.400 1524.800 2849.540 1525.000 ;
        RECT 2850.705 1524.955 2850.995 1525.000 ;
        RECT 2852.545 1524.800 2852.835 1524.845 ;
        RECT 2849.400 1524.660 2852.835 1524.800 ;
        RECT 2852.545 1524.615 2852.835 1524.660 ;
        RECT 2849.770 1480.600 2850.090 1480.660 ;
        RECT 2852.545 1480.600 2852.835 1480.645 ;
        RECT 2849.770 1480.460 2852.835 1480.600 ;
        RECT 2849.770 1480.400 2850.090 1480.460 ;
        RECT 2852.545 1480.415 2852.835 1480.460 ;
        RECT 2850.230 1417.360 2850.550 1417.420 ;
        RECT 2851.165 1417.360 2851.455 1417.405 ;
        RECT 2850.230 1417.220 2851.455 1417.360 ;
        RECT 2850.230 1417.160 2850.550 1417.220 ;
        RECT 2851.165 1417.175 2851.455 1417.220 ;
        RECT 2849.770 1351.740 2850.090 1351.800 ;
        RECT 2851.165 1351.740 2851.455 1351.785 ;
        RECT 2849.770 1351.600 2851.455 1351.740 ;
        RECT 2849.770 1351.540 2850.090 1351.600 ;
        RECT 2851.165 1351.555 2851.455 1351.600 ;
        RECT 2849.770 1320.120 2850.090 1320.180 ;
        RECT 2851.165 1320.120 2851.455 1320.165 ;
        RECT 2849.770 1319.980 2851.455 1320.120 ;
        RECT 2849.770 1319.920 2850.090 1319.980 ;
        RECT 2851.165 1319.935 2851.455 1319.980 ;
        RECT 2849.770 1298.020 2850.090 1298.080 ;
        RECT 2851.165 1298.020 2851.455 1298.065 ;
        RECT 2849.770 1297.880 2851.455 1298.020 ;
        RECT 2849.770 1297.820 2850.090 1297.880 ;
        RECT 2851.165 1297.835 2851.455 1297.880 ;
        RECT 2849.785 1273.880 2850.075 1273.925 ;
        RECT 2850.230 1273.880 2850.550 1273.940 ;
        RECT 2849.785 1273.740 2850.550 1273.880 ;
        RECT 2849.785 1273.695 2850.075 1273.740 ;
        RECT 2850.230 1273.680 2850.550 1273.740 ;
        RECT 2849.785 1230.020 2850.075 1230.065 ;
        RECT 2851.165 1230.020 2851.455 1230.065 ;
        RECT 2849.785 1229.880 2851.455 1230.020 ;
        RECT 2849.785 1229.835 2850.075 1229.880 ;
        RECT 2851.165 1229.835 2851.455 1229.880 ;
        RECT 2849.770 1218.460 2850.090 1218.520 ;
        RECT 2851.165 1218.460 2851.455 1218.505 ;
        RECT 2849.770 1218.320 2851.455 1218.460 ;
        RECT 2849.770 1218.260 2850.090 1218.320 ;
        RECT 2851.165 1218.275 2851.455 1218.320 ;
        RECT 2849.770 1168.480 2850.090 1168.540 ;
        RECT 2852.545 1168.480 2852.835 1168.525 ;
        RECT 2849.770 1168.340 2852.835 1168.480 ;
        RECT 2849.770 1168.280 2850.090 1168.340 ;
        RECT 2852.545 1168.295 2852.835 1168.340 ;
        RECT 2849.770 1146.380 2850.090 1146.440 ;
        RECT 2852.545 1146.380 2852.835 1146.425 ;
        RECT 2849.770 1146.240 2852.835 1146.380 ;
        RECT 2849.770 1146.180 2850.090 1146.240 ;
        RECT 2852.545 1146.195 2852.835 1146.240 ;
        RECT 2849.770 1130.060 2850.090 1130.120 ;
        RECT 2851.150 1130.060 2851.470 1130.120 ;
        RECT 2849.770 1129.920 2851.470 1130.060 ;
        RECT 2849.770 1129.860 2850.090 1129.920 ;
        RECT 2851.150 1129.860 2851.470 1129.920 ;
        RECT 2849.770 1070.220 2850.090 1070.280 ;
        RECT 2851.150 1070.220 2851.470 1070.280 ;
        RECT 2849.770 1070.080 2851.470 1070.220 ;
        RECT 2849.770 1070.020 2850.090 1070.080 ;
        RECT 2851.150 1070.020 2851.470 1070.080 ;
        RECT 2849.770 1025.340 2850.090 1025.400 ;
        RECT 2851.150 1025.340 2851.470 1025.400 ;
        RECT 2849.770 1025.200 2851.470 1025.340 ;
        RECT 2849.770 1025.140 2850.090 1025.200 ;
        RECT 2851.150 1025.140 2851.470 1025.200 ;
        RECT 2849.770 1017.180 2850.090 1017.240 ;
        RECT 2851.150 1017.180 2851.470 1017.240 ;
        RECT 2849.770 1017.040 2851.470 1017.180 ;
        RECT 2849.770 1016.980 2850.090 1017.040 ;
        RECT 2851.150 1016.980 2851.470 1017.040 ;
        RECT 2849.770 960.400 2850.090 960.460 ;
        RECT 2851.625 960.400 2851.915 960.445 ;
        RECT 2849.770 960.260 2851.915 960.400 ;
        RECT 2849.770 960.200 2850.090 960.260 ;
        RECT 2851.625 960.215 2851.915 960.260 ;
        RECT 2850.705 890.360 2850.995 890.405 ;
        RECT 2851.625 890.360 2851.915 890.405 ;
        RECT 2850.705 890.220 2851.915 890.360 ;
        RECT 2850.705 890.175 2850.995 890.220 ;
        RECT 2851.625 890.175 2851.915 890.220 ;
        RECT 2851.150 767.280 2851.470 767.340 ;
        RECT 2850.955 767.140 2851.470 767.280 ;
        RECT 2851.150 767.080 2851.470 767.140 ;
        RECT 2849.770 721.380 2850.090 721.440 ;
        RECT 2851.610 721.380 2851.930 721.440 ;
        RECT 2849.770 721.240 2851.930 721.380 ;
        RECT 2849.770 721.180 2850.090 721.240 ;
        RECT 2851.610 721.180 2851.930 721.240 ;
        RECT 2849.770 381.720 2850.090 381.780 ;
        RECT 2849.575 381.580 2850.090 381.720 ;
        RECT 2849.770 381.520 2850.090 381.580 ;
        RECT 2849.325 294.340 2849.615 294.385 ;
        RECT 2849.770 294.340 2850.090 294.400 ;
        RECT 2849.325 294.200 2850.090 294.340 ;
        RECT 2849.325 294.155 2849.615 294.200 ;
        RECT 2849.770 294.140 2850.090 294.200 ;
        RECT 2849.770 209.000 2850.090 209.060 ;
        RECT 2851.625 209.000 2851.915 209.045 ;
        RECT 2849.770 208.860 2851.915 209.000 ;
        RECT 2849.770 208.800 2850.090 208.860 ;
        RECT 2851.625 208.815 2851.915 208.860 ;
        RECT 2850.705 198.800 2850.995 198.845 ;
        RECT 2851.625 198.800 2851.915 198.845 ;
        RECT 2850.705 198.660 2851.915 198.800 ;
        RECT 2850.705 198.615 2850.995 198.660 ;
        RECT 2851.625 198.615 2851.915 198.660 ;
        RECT 2849.770 116.180 2850.090 116.240 ;
        RECT 2850.705 116.180 2850.995 116.225 ;
        RECT 2849.770 116.040 2850.995 116.180 ;
        RECT 2849.770 115.980 2850.090 116.040 ;
        RECT 2850.705 115.995 2850.995 116.040 ;
        RECT 1841.925 9.080 1842.215 9.125 ;
        RECT 1874.125 9.080 1874.415 9.125 ;
        RECT 1841.925 8.940 1874.415 9.080 ;
        RECT 1841.925 8.895 1842.215 8.940 ;
        RECT 1874.125 8.895 1874.415 8.940 ;
        RECT 898.465 8.740 898.755 8.785 ;
        RECT 902.145 8.740 902.435 8.785 ;
        RECT 898.465 8.600 902.435 8.740 ;
        RECT 898.465 8.555 898.755 8.600 ;
        RECT 902.145 8.555 902.435 8.600 ;
        RECT 920.545 7.720 920.835 7.765 ;
        RECT 947.225 7.720 947.515 7.765 ;
        RECT 920.545 7.580 947.515 7.720 ;
        RECT 920.545 7.535 920.835 7.580 ;
        RECT 947.225 7.535 947.515 7.580 ;
        RECT 1183.205 7.380 1183.495 7.425 ;
        RECT 1194.690 7.380 1195.010 7.440 ;
        RECT 1183.205 7.240 1195.010 7.380 ;
        RECT 1183.205 7.195 1183.495 7.240 ;
        RECT 1194.690 7.180 1195.010 7.240 ;
        RECT 1932.545 7.380 1932.835 7.425 ;
        RECT 1956.005 7.380 1956.295 7.425 ;
        RECT 1932.545 7.240 1956.295 7.380 ;
        RECT 1932.545 7.195 1932.835 7.240 ;
        RECT 1956.005 7.195 1956.295 7.240 ;
        RECT 1122.945 6.700 1123.235 6.745 ;
        RECT 1127.085 6.700 1127.375 6.745 ;
        RECT 1122.945 6.560 1127.375 6.700 ;
        RECT 1122.945 6.515 1123.235 6.560 ;
        RECT 1127.085 6.515 1127.375 6.560 ;
        RECT 797.725 6.360 798.015 6.405 ;
        RECT 807.385 6.360 807.675 6.405 ;
        RECT 1635.385 6.360 1635.675 6.405 ;
        RECT 1637.225 6.360 1637.515 6.405 ;
        RECT 797.725 6.220 807.675 6.360 ;
        RECT 797.725 6.175 798.015 6.220 ;
        RECT 807.385 6.175 807.675 6.220 ;
        RECT 1546.680 6.220 1592.820 6.360 ;
        RECT 903.065 6.020 903.355 6.065 ;
        RECT 919.165 6.020 919.455 6.065 ;
        RECT 903.065 5.880 919.455 6.020 ;
        RECT 903.065 5.835 903.355 5.880 ;
        RECT 919.165 5.835 919.455 5.880 ;
        RECT 955.045 6.020 955.335 6.065 ;
        RECT 1120.645 6.020 1120.935 6.065 ;
        RECT 955.045 5.880 1120.935 6.020 ;
        RECT 955.045 5.835 955.335 5.880 ;
        RECT 1120.645 5.835 1120.935 5.880 ;
        RECT 1141.805 6.020 1142.095 6.065 ;
        RECT 1183.205 6.020 1183.495 6.065 ;
        RECT 1141.805 5.880 1183.495 6.020 ;
        RECT 1141.805 5.835 1142.095 5.880 ;
        RECT 1183.205 5.835 1183.495 5.880 ;
        RECT 1194.690 6.020 1195.010 6.080 ;
        RECT 1255.885 6.020 1256.175 6.065 ;
        RECT 1194.690 5.880 1256.175 6.020 ;
        RECT 1194.690 5.820 1195.010 5.880 ;
        RECT 1255.885 5.835 1256.175 5.880 ;
        RECT 1303.725 6.020 1304.015 6.065 ;
        RECT 1352.930 6.020 1353.250 6.080 ;
        RECT 1303.725 5.880 1353.250 6.020 ;
        RECT 1303.725 5.835 1304.015 5.880 ;
        RECT 1352.930 5.820 1353.250 5.880 ;
        RECT 1400.325 6.020 1400.615 6.065 ;
        RECT 1407.685 6.020 1407.975 6.065 ;
        RECT 1400.325 5.880 1407.975 6.020 ;
        RECT 1400.325 5.835 1400.615 5.880 ;
        RECT 1407.685 5.835 1407.975 5.880 ;
        RECT 1410.445 6.020 1410.735 6.065 ;
        RECT 1450.910 6.020 1451.230 6.080 ;
        RECT 1410.445 5.880 1451.230 6.020 ;
        RECT 1410.445 5.835 1410.735 5.880 ;
        RECT 1450.910 5.820 1451.230 5.880 ;
        RECT 1503.825 6.020 1504.115 6.065 ;
        RECT 1546.680 6.020 1546.820 6.220 ;
        RECT 1503.825 5.880 1546.820 6.020 ;
        RECT 1592.680 6.020 1592.820 6.220 ;
        RECT 1635.385 6.220 1637.515 6.360 ;
        RECT 1635.385 6.175 1635.675 6.220 ;
        RECT 1637.225 6.175 1637.515 6.220 ;
        RECT 1634.465 6.020 1634.755 6.065 ;
        RECT 1592.680 5.880 1634.755 6.020 ;
        RECT 1503.825 5.835 1504.115 5.880 ;
        RECT 1634.465 5.835 1634.755 5.880 ;
        RECT 1691.490 6.020 1691.810 6.080 ;
        RECT 1742.565 6.020 1742.855 6.065 ;
        RECT 1691.490 5.880 1742.855 6.020 ;
        RECT 1691.490 5.820 1691.810 5.880 ;
        RECT 1742.565 5.835 1742.855 5.880 ;
        RECT 1785.345 6.020 1785.635 6.065 ;
        RECT 1835.025 6.020 1835.315 6.065 ;
        RECT 1785.345 5.880 1835.315 6.020 ;
        RECT 1785.345 5.835 1785.635 5.880 ;
        RECT 1835.025 5.835 1835.315 5.880 ;
        RECT 1835.485 6.020 1835.775 6.065 ;
        RECT 1841.925 6.020 1842.215 6.065 ;
        RECT 1835.485 5.880 1842.215 6.020 ;
        RECT 1835.485 5.835 1835.775 5.880 ;
        RECT 1841.925 5.835 1842.215 5.880 ;
        RECT 1874.125 6.020 1874.415 6.065 ;
        RECT 1932.545 6.020 1932.835 6.065 ;
        RECT 1874.125 5.880 1932.835 6.020 ;
        RECT 1874.125 5.835 1874.415 5.880 ;
        RECT 1932.545 5.835 1932.835 5.880 ;
        RECT 1956.005 6.020 1956.295 6.065 ;
        RECT 2469.810 6.020 2470.130 6.080 ;
        RECT 1956.005 5.880 2470.130 6.020 ;
        RECT 1956.005 5.835 1956.295 5.880 ;
        RECT 2469.810 5.820 2470.130 5.880 ;
        RECT 2471.190 6.020 2471.510 6.080 ;
        RECT 2847.470 6.020 2847.790 6.080 ;
        RECT 2471.190 5.880 2847.790 6.020 ;
        RECT 2471.190 5.820 2471.510 5.880 ;
        RECT 2847.470 5.820 2847.790 5.880 ;
        RECT 1763.265 5.340 1763.555 5.385 ;
        RECT 1785.345 5.340 1785.635 5.385 ;
        RECT 1763.265 5.200 1785.635 5.340 ;
        RECT 1763.265 5.155 1763.555 5.200 ;
        RECT 1785.345 5.155 1785.635 5.200 ;
        RECT 353.350 4.660 353.670 4.720 ;
        RECT 353.350 4.520 364.620 4.660 ;
        RECT 353.350 4.460 353.670 4.520 ;
        RECT 364.480 4.320 364.620 4.520 ;
        RECT 379.585 4.320 379.875 4.365 ;
        RECT 364.480 4.180 379.875 4.320 ;
        RECT 379.585 4.135 379.875 4.180 ;
        RECT 379.585 3.300 379.875 3.345 ;
        RECT 411.325 3.300 411.615 3.345 ;
        RECT 379.585 3.160 411.615 3.300 ;
        RECT 379.585 3.115 379.875 3.160 ;
        RECT 411.325 3.115 411.615 3.160 ;
        RECT 413.625 3.300 413.915 3.345 ;
        RECT 460.545 3.300 460.835 3.345 ;
        RECT 413.625 3.160 460.835 3.300 ;
        RECT 413.625 3.115 413.915 3.160 ;
        RECT 460.545 3.115 460.835 3.160 ;
        RECT 462.385 3.300 462.675 3.345 ;
        RECT 607.285 3.300 607.575 3.345 ;
        RECT 462.385 3.160 557.820 3.300 ;
        RECT 462.385 3.115 462.675 3.160 ;
        RECT 557.680 2.960 557.820 3.160 ;
        RECT 561.360 3.160 607.575 3.300 ;
        RECT 561.360 2.960 561.500 3.160 ;
        RECT 607.285 3.115 607.575 3.160 ;
        RECT 623.385 3.300 623.675 3.345 ;
        RECT 748.505 3.300 748.795 3.345 ;
        RECT 623.385 3.160 748.795 3.300 ;
        RECT 623.385 3.115 623.675 3.160 ;
        RECT 748.505 3.115 748.795 3.160 ;
        RECT 557.680 2.820 561.500 2.960 ;
        RECT 1258.185 2.620 1258.475 2.665 ;
        RECT 1298.205 2.620 1298.495 2.665 ;
        RECT 1258.185 2.480 1298.495 2.620 ;
        RECT 1258.185 2.435 1258.475 2.480 ;
        RECT 1298.205 2.435 1298.495 2.480 ;
        RECT 1398.945 2.435 1399.235 2.665 ;
        RECT 1487.265 2.620 1487.555 2.665 ;
        RECT 1484.120 2.480 1487.555 2.620 ;
        RECT 1353.390 2.280 1353.710 2.340 ;
        RECT 1399.020 2.280 1399.160 2.435 ;
        RECT 1353.390 2.140 1399.160 2.280 ;
        RECT 1450.910 2.280 1451.230 2.340 ;
        RECT 1484.120 2.280 1484.260 2.480 ;
        RECT 1487.265 2.435 1487.555 2.480 ;
        RECT 1639.985 2.620 1640.275 2.665 ;
        RECT 1677.705 2.620 1677.995 2.665 ;
        RECT 1639.985 2.480 1677.995 2.620 ;
        RECT 1639.985 2.435 1640.275 2.480 ;
        RECT 1677.705 2.435 1677.995 2.480 ;
        RECT 1742.565 2.620 1742.855 2.665 ;
        RECT 1763.265 2.620 1763.555 2.665 ;
        RECT 1742.565 2.480 1763.555 2.620 ;
        RECT 1742.565 2.435 1742.855 2.480 ;
        RECT 1763.265 2.435 1763.555 2.480 ;
        RECT 1450.910 2.140 1484.260 2.280 ;
        RECT 1678.625 2.280 1678.915 2.325 ;
        RECT 1689.190 2.280 1689.510 2.340 ;
        RECT 1678.625 2.140 1689.510 2.280 ;
        RECT 1353.390 2.080 1353.710 2.140 ;
        RECT 1450.910 2.080 1451.230 2.140 ;
        RECT 1678.625 2.095 1678.915 2.140 ;
        RECT 1689.190 2.080 1689.510 2.140 ;
        RECT 769.205 1.940 769.495 1.985 ;
        RECT 772.885 1.940 773.175 1.985 ;
        RECT 769.205 1.800 773.175 1.940 ;
        RECT 769.205 1.755 769.495 1.800 ;
        RECT 772.885 1.755 773.175 1.800 ;
        RECT 1488.185 1.940 1488.475 1.985 ;
        RECT 1503.365 1.940 1503.655 1.985 ;
        RECT 1488.185 1.800 1503.655 1.940 ;
        RECT 1488.185 1.755 1488.475 1.800 ;
        RECT 1503.365 1.755 1503.655 1.800 ;
      LAYER via ;
        RECT 2849.800 2759.140 2850.060 2759.400 ;
        RECT 2863.600 2759.140 2863.860 2759.400 ;
        RECT 2849.800 2325.980 2850.060 2326.240 ;
        RECT 2849.800 2317.820 2850.060 2318.080 ;
        RECT 2849.800 1968.300 2850.060 1968.560 ;
        RECT 2849.800 1949.260 2850.060 1949.520 ;
        RECT 2849.800 1840.120 2850.060 1840.380 ;
        RECT 2850.720 1840.120 2850.980 1840.380 ;
        RECT 2850.260 1790.480 2850.520 1790.740 ;
        RECT 2850.260 1789.460 2850.520 1789.720 ;
        RECT 2850.260 1762.940 2850.520 1763.200 ;
        RECT 2849.800 1744.580 2850.060 1744.840 ;
        RECT 2849.800 1648.360 2850.060 1648.620 ;
        RECT 2850.260 1624.900 2850.520 1625.160 ;
        RECT 2850.260 1603.480 2850.520 1603.740 ;
        RECT 2849.800 1480.400 2850.060 1480.660 ;
        RECT 2850.260 1417.160 2850.520 1417.420 ;
        RECT 2849.800 1351.540 2850.060 1351.800 ;
        RECT 2849.800 1319.920 2850.060 1320.180 ;
        RECT 2849.800 1297.820 2850.060 1298.080 ;
        RECT 2850.260 1273.680 2850.520 1273.940 ;
        RECT 2849.800 1218.260 2850.060 1218.520 ;
        RECT 2849.800 1168.280 2850.060 1168.540 ;
        RECT 2849.800 1146.180 2850.060 1146.440 ;
        RECT 2849.800 1129.860 2850.060 1130.120 ;
        RECT 2851.180 1129.860 2851.440 1130.120 ;
        RECT 2849.800 1070.020 2850.060 1070.280 ;
        RECT 2851.180 1070.020 2851.440 1070.280 ;
        RECT 2849.800 1025.140 2850.060 1025.400 ;
        RECT 2851.180 1025.140 2851.440 1025.400 ;
        RECT 2849.800 1016.980 2850.060 1017.240 ;
        RECT 2851.180 1016.980 2851.440 1017.240 ;
        RECT 2849.800 960.200 2850.060 960.460 ;
        RECT 2851.180 767.080 2851.440 767.340 ;
        RECT 2849.800 721.180 2850.060 721.440 ;
        RECT 2851.640 721.180 2851.900 721.440 ;
        RECT 2849.800 381.520 2850.060 381.780 ;
        RECT 2849.800 294.140 2850.060 294.400 ;
        RECT 2849.800 208.800 2850.060 209.060 ;
        RECT 2849.800 115.980 2850.060 116.240 ;
        RECT 1194.720 7.180 1194.980 7.440 ;
        RECT 1194.720 5.820 1194.980 6.080 ;
        RECT 1352.960 5.820 1353.220 6.080 ;
        RECT 1450.940 5.820 1451.200 6.080 ;
        RECT 1691.520 5.820 1691.780 6.080 ;
        RECT 2469.840 5.820 2470.100 6.080 ;
        RECT 2471.220 5.820 2471.480 6.080 ;
        RECT 2847.500 5.820 2847.760 6.080 ;
        RECT 353.380 4.460 353.640 4.720 ;
        RECT 1353.420 2.080 1353.680 2.340 ;
        RECT 1450.940 2.080 1451.200 2.340 ;
        RECT 1689.220 2.080 1689.480 2.340 ;
      LAYER met2 ;
        RECT 2863.590 2792.915 2863.870 2793.285 ;
        RECT 2863.660 2759.430 2863.800 2792.915 ;
        RECT 2849.800 2759.340 2850.060 2759.430 ;
        RECT 2849.400 2759.200 2850.060 2759.340 ;
        RECT 2849.400 2758.490 2849.540 2759.200 ;
        RECT 2849.800 2759.110 2850.060 2759.200 ;
        RECT 2863.600 2759.110 2863.860 2759.430 ;
        RECT 2847.100 2758.350 2849.540 2758.490 ;
        RECT 2847.100 2326.180 2847.240 2758.350 ;
        RECT 2849.800 2326.180 2850.060 2326.270 ;
        RECT 2847.100 2326.040 2850.060 2326.180 ;
        RECT 2849.800 2325.950 2850.060 2326.040 ;
        RECT 2849.800 2317.790 2850.060 2318.110 ;
        RECT 2849.860 2315.130 2850.000 2317.790 ;
        RECT 2847.100 2314.990 2850.000 2315.130 ;
        RECT 2847.100 1969.180 2847.240 2314.990 ;
        RECT 2847.100 1969.040 2849.540 1969.180 ;
        RECT 2849.400 1968.500 2849.540 1969.040 ;
        RECT 2849.800 1968.500 2850.060 1968.590 ;
        RECT 2849.400 1968.360 2850.060 1968.500 ;
        RECT 2849.800 1968.270 2850.060 1968.360 ;
        RECT 2849.800 1949.230 2850.060 1949.550 ;
        RECT 2849.860 1945.890 2850.000 1949.230 ;
        RECT 2847.100 1945.750 2850.000 1945.890 ;
        RECT 2847.100 1890.130 2847.240 1945.750 ;
        RECT 2847.100 1889.990 2847.700 1890.130 ;
        RECT 2847.560 1886.730 2847.700 1889.990 ;
        RECT 2847.100 1886.590 2847.700 1886.730 ;
        RECT 2847.100 1840.320 2847.240 1886.590 ;
        RECT 2849.800 1840.320 2850.060 1840.410 ;
        RECT 2847.100 1840.180 2850.060 1840.320 ;
        RECT 2849.800 1840.090 2850.060 1840.180 ;
        RECT 2850.720 1840.090 2850.980 1840.410 ;
        RECT 2850.780 1811.250 2850.920 1840.090 ;
        RECT 2850.320 1811.110 2850.920 1811.250 ;
        RECT 2850.320 1790.770 2850.460 1811.110 ;
        RECT 2850.260 1790.450 2850.520 1790.770 ;
        RECT 2850.260 1789.430 2850.520 1789.750 ;
        RECT 2850.320 1763.230 2850.460 1789.430 ;
        RECT 2850.260 1762.910 2850.520 1763.230 ;
        RECT 2849.800 1744.780 2850.060 1744.870 ;
        RECT 2848.020 1744.640 2850.060 1744.780 ;
        RECT 2848.020 1741.210 2848.160 1744.640 ;
        RECT 2849.800 1744.550 2850.060 1744.640 ;
        RECT 2847.100 1741.070 2848.160 1741.210 ;
        RECT 2847.100 1699.730 2847.240 1741.070 ;
        RECT 2847.100 1699.590 2848.160 1699.730 ;
        RECT 2848.020 1686.130 2848.160 1699.590 ;
        RECT 2847.100 1685.990 2848.160 1686.130 ;
        RECT 2847.100 1650.090 2847.240 1685.990 ;
        RECT 2847.100 1649.950 2850.000 1650.090 ;
        RECT 2849.860 1648.650 2850.000 1649.950 ;
        RECT 2849.800 1648.330 2850.060 1648.650 ;
        RECT 2850.260 1624.870 2850.520 1625.190 ;
        RECT 2850.320 1603.770 2850.460 1624.870 ;
        RECT 2850.260 1603.450 2850.520 1603.770 ;
        RECT 2849.800 1480.370 2850.060 1480.690 ;
        RECT 2849.860 1480.090 2850.000 1480.370 ;
        RECT 2848.480 1479.950 2850.000 1480.090 ;
        RECT 2848.480 1464.450 2848.620 1479.950 ;
        RECT 2848.020 1464.310 2848.620 1464.450 ;
        RECT 2848.020 1426.370 2848.160 1464.310 ;
        RECT 2848.020 1426.230 2850.460 1426.370 ;
        RECT 2850.320 1417.450 2850.460 1426.230 ;
        RECT 2850.260 1417.130 2850.520 1417.450 ;
        RECT 2849.800 1351.570 2850.060 1351.830 ;
        RECT 2847.100 1351.510 2850.060 1351.570 ;
        RECT 2847.100 1351.430 2850.000 1351.510 ;
        RECT 2847.100 1320.120 2847.240 1351.430 ;
        RECT 2849.800 1320.120 2850.060 1320.210 ;
        RECT 2847.100 1319.980 2850.060 1320.120 ;
        RECT 2849.800 1319.890 2850.060 1319.980 ;
        RECT 2849.800 1297.790 2850.060 1298.110 ;
        RECT 2849.860 1286.290 2850.000 1297.790 ;
        RECT 2849.860 1286.150 2850.460 1286.290 ;
        RECT 2850.320 1273.970 2850.460 1286.150 ;
        RECT 2850.260 1273.650 2850.520 1273.970 ;
        RECT 2849.800 1218.460 2850.060 1218.550 ;
        RECT 2848.940 1218.320 2850.060 1218.460 ;
        RECT 2848.940 1214.210 2849.080 1218.320 ;
        RECT 2849.800 1218.230 2850.060 1218.320 ;
        RECT 2848.480 1214.070 2849.080 1214.210 ;
        RECT 2848.480 1168.650 2848.620 1214.070 ;
        RECT 2848.480 1168.570 2850.000 1168.650 ;
        RECT 2848.480 1168.510 2850.060 1168.570 ;
        RECT 2849.800 1168.250 2850.060 1168.510 ;
        RECT 2849.800 1146.150 2850.060 1146.470 ;
        RECT 2849.860 1142.130 2850.000 1146.150 ;
        RECT 2849.400 1141.990 2850.000 1142.130 ;
        RECT 2849.400 1135.330 2849.540 1141.990 ;
        RECT 2849.400 1135.190 2850.000 1135.330 ;
        RECT 2849.860 1130.150 2850.000 1135.190 ;
        RECT 2849.800 1129.830 2850.060 1130.150 ;
        RECT 2851.180 1129.830 2851.440 1130.150 ;
        RECT 2851.240 1070.310 2851.380 1129.830 ;
        RECT 2849.800 1070.050 2850.060 1070.310 ;
        RECT 2848.940 1069.990 2850.060 1070.050 ;
        RECT 2851.180 1069.990 2851.440 1070.310 ;
        RECT 2848.940 1069.910 2850.000 1069.990 ;
        RECT 2848.940 1064.610 2849.080 1069.910 ;
        RECT 2848.940 1064.470 2849.540 1064.610 ;
        RECT 2849.400 1055.770 2849.540 1064.470 ;
        RECT 2849.400 1055.630 2850.000 1055.770 ;
        RECT 2849.860 1048.970 2850.000 1055.630 ;
        RECT 2848.480 1048.830 2850.000 1048.970 ;
        RECT 2848.480 1025.340 2848.620 1048.830 ;
        RECT 2849.800 1025.340 2850.060 1025.430 ;
        RECT 2848.480 1025.200 2850.060 1025.340 ;
        RECT 2849.800 1025.110 2850.060 1025.200 ;
        RECT 2851.180 1025.110 2851.440 1025.430 ;
        RECT 2851.240 1017.270 2851.380 1025.110 ;
        RECT 2849.800 1017.010 2850.060 1017.270 ;
        RECT 2847.100 1016.950 2850.060 1017.010 ;
        RECT 2851.180 1016.950 2851.440 1017.270 ;
        RECT 2847.100 1016.870 2850.000 1016.950 ;
        RECT 2847.100 961.250 2847.240 1016.870 ;
        RECT 2847.100 961.110 2847.700 961.250 ;
        RECT 2847.560 960.570 2847.700 961.110 ;
        RECT 2847.560 960.490 2850.000 960.570 ;
        RECT 2847.560 960.430 2850.060 960.490 ;
        RECT 2849.800 960.170 2850.060 960.430 ;
        RECT 2851.180 767.050 2851.440 767.370 ;
        RECT 2851.240 746.540 2851.380 767.050 ;
        RECT 2851.240 746.400 2851.840 746.540 ;
        RECT 2851.700 721.470 2851.840 746.400 ;
        RECT 2849.800 721.210 2850.060 721.470 ;
        RECT 2849.400 721.150 2850.060 721.210 ;
        RECT 2851.640 721.150 2851.900 721.470 ;
        RECT 2849.400 721.070 2850.000 721.150 ;
        RECT 2849.400 679.050 2849.540 721.070 ;
        RECT 2849.400 678.910 2850.460 679.050 ;
        RECT 2850.320 674.290 2850.460 678.910 ;
        RECT 2848.940 674.150 2850.460 674.290 ;
        RECT 2848.940 673.610 2849.080 674.150 ;
        RECT 2847.100 673.470 2849.080 673.610 ;
        RECT 2847.100 382.400 2847.240 673.470 ;
        RECT 2847.100 382.260 2847.700 382.400 ;
        RECT 2847.560 381.720 2847.700 382.260 ;
        RECT 2848.940 381.810 2850.000 381.890 ;
        RECT 2848.940 381.750 2850.060 381.810 ;
        RECT 2848.940 381.720 2849.080 381.750 ;
        RECT 2847.560 381.580 2849.080 381.720 ;
        RECT 2849.800 381.490 2850.060 381.750 ;
        RECT 2849.800 294.170 2850.060 294.430 ;
        RECT 2847.100 294.110 2850.060 294.170 ;
        RECT 2847.100 294.030 2850.000 294.110 ;
        RECT 2847.100 209.000 2847.240 294.030 ;
        RECT 2849.800 209.000 2850.060 209.090 ;
        RECT 2847.100 208.860 2850.060 209.000 ;
        RECT 2849.800 208.770 2850.060 208.860 ;
        RECT 2849.800 115.950 2850.060 116.270 ;
        RECT 2849.860 88.810 2850.000 115.950 ;
        RECT 2848.020 88.670 2850.000 88.810 ;
        RECT 2848.020 75.890 2848.160 88.670 ;
        RECT 2847.560 75.750 2848.160 75.890 ;
        RECT 2847.560 42.570 2847.700 75.750 ;
        RECT 2847.560 42.430 2848.160 42.570 ;
        RECT 2848.020 41.210 2848.160 42.430 ;
        RECT 2847.560 41.070 2848.160 41.210 ;
        RECT 1194.720 7.150 1194.980 7.470 ;
        RECT 1194.780 6.110 1194.920 7.150 ;
        RECT 2847.560 6.110 2847.700 41.070 ;
        RECT 1194.720 5.790 1194.980 6.110 ;
        RECT 1352.960 5.850 1353.220 6.110 ;
        RECT 1352.960 5.790 1353.620 5.850 ;
        RECT 1450.940 5.790 1451.200 6.110 ;
        RECT 1353.020 5.710 1353.620 5.790 ;
        RECT 353.380 4.430 353.640 4.750 ;
        RECT 353.440 2.400 353.580 4.430 ;
        RECT 353.230 -4.800 353.790 2.400 ;
        RECT 1353.480 2.370 1353.620 5.710 ;
        RECT 1451.000 2.370 1451.140 5.790 ;
        RECT 1689.280 5.710 1690.800 5.850 ;
        RECT 1691.520 5.790 1691.780 6.110 ;
        RECT 2469.840 5.850 2470.100 6.110 ;
        RECT 2471.220 5.850 2471.480 6.110 ;
        RECT 2469.840 5.790 2471.480 5.850 ;
        RECT 2847.500 5.790 2847.760 6.110 ;
        RECT 1689.280 2.370 1689.420 5.710 ;
        RECT 1690.660 4.660 1690.800 5.710 ;
        RECT 1691.580 4.660 1691.720 5.790 ;
        RECT 2469.900 5.710 2471.420 5.790 ;
        RECT 1690.660 4.520 1691.720 4.660 ;
        RECT 1353.420 2.050 1353.680 2.370 ;
        RECT 1450.940 2.050 1451.200 2.370 ;
        RECT 1689.220 2.050 1689.480 2.370 ;
      LAYER via2 ;
        RECT 2863.590 2792.960 2863.870 2793.240 ;
      LAYER met3 ;
        RECT 2851.000 2793.250 2855.000 2793.640 ;
        RECT 2863.565 2793.250 2863.895 2793.265 ;
        RECT 2851.000 2793.040 2863.895 2793.250 ;
        RECT 2854.300 2792.950 2863.895 2793.040 ;
        RECT 2863.565 2792.935 2863.895 2792.950 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2470.345 3399.745 2470.515 3401.955 ;
        RECT 2796.025 3399.745 2796.195 3401.615 ;
        RECT 2.445 1.445 2.615 43.435 ;
        RECT 26.365 0.255 26.535 1.615 ;
        RECT 30.045 0.255 30.215 0.595 ;
        RECT 48.905 0.425 49.075 1.615 ;
        RECT 134.005 1.445 134.175 7.055 ;
        RECT 135.385 6.885 135.555 8.415 ;
        RECT 175.405 6.885 175.575 8.415 ;
        RECT 195.185 1.445 195.355 7.055 ;
        RECT 198.865 0.765 199.035 1.615 ;
        RECT 249.005 0.765 249.175 3.315 ;
        RECT 26.365 0.085 30.215 0.255 ;
      LAYER mcon ;
        RECT 2470.345 3401.785 2470.515 3401.955 ;
        RECT 2796.025 3401.445 2796.195 3401.615 ;
        RECT 2.445 43.265 2.615 43.435 ;
        RECT 135.385 8.245 135.555 8.415 ;
        RECT 134.005 6.885 134.175 7.055 ;
        RECT 175.405 8.245 175.575 8.415 ;
        RECT 195.185 6.885 195.355 7.055 ;
        RECT 26.365 1.445 26.535 1.615 ;
        RECT 48.905 1.445 49.075 1.615 ;
        RECT 249.005 3.145 249.175 3.315 ;
        RECT 198.865 1.445 199.035 1.615 ;
        RECT 30.045 0.425 30.215 0.595 ;
      LAYER met1 ;
        RECT 2412.310 3416.220 2412.630 3416.280 ;
        RECT 2470.270 3416.220 2470.590 3416.280 ;
        RECT 2412.310 3416.080 2470.590 3416.220 ;
        RECT 2412.310 3416.020 2412.630 3416.080 ;
        RECT 2470.270 3416.020 2470.590 3416.080 ;
        RECT 2470.270 3401.940 2470.590 3402.000 ;
        RECT 2470.075 3401.800 2470.590 3401.940 ;
        RECT 2470.270 3401.740 2470.590 3401.800 ;
        RECT 2795.950 3401.600 2796.270 3401.660 ;
        RECT 2795.755 3401.460 2796.270 3401.600 ;
        RECT 2795.950 3401.400 2796.270 3401.460 ;
        RECT 2470.285 3399.900 2470.575 3399.945 ;
        RECT 2795.965 3399.900 2796.255 3399.945 ;
        RECT 2470.285 3399.760 2796.255 3399.900 ;
        RECT 2470.285 3399.715 2470.575 3399.760 ;
        RECT 2795.965 3399.715 2796.255 3399.760 ;
        RECT 3.290 51.720 3.610 51.980 ;
        RECT 2.370 50.900 2.690 50.960 ;
        RECT 3.380 50.900 3.520 51.720 ;
        RECT 2.370 50.760 3.520 50.900 ;
        RECT 2.370 50.700 2.690 50.760 ;
        RECT 2.370 43.420 2.690 43.480 ;
        RECT 2.175 43.280 2.690 43.420 ;
        RECT 2.370 43.220 2.690 43.280 ;
        RECT 135.325 8.400 135.615 8.445 ;
        RECT 175.345 8.400 175.635 8.445 ;
        RECT 135.325 8.260 175.635 8.400 ;
        RECT 135.325 8.215 135.615 8.260 ;
        RECT 175.345 8.215 175.635 8.260 ;
        RECT 296.770 7.720 297.090 7.780 ;
        RECT 334.490 7.720 334.810 7.780 ;
        RECT 296.770 7.580 334.810 7.720 ;
        RECT 296.770 7.520 297.090 7.580 ;
        RECT 334.490 7.520 334.810 7.580 ;
        RECT 133.945 7.040 134.235 7.085 ;
        RECT 135.325 7.040 135.615 7.085 ;
        RECT 133.945 6.900 135.615 7.040 ;
        RECT 133.945 6.855 134.235 6.900 ;
        RECT 135.325 6.855 135.615 6.900 ;
        RECT 175.345 7.040 175.635 7.085 ;
        RECT 195.125 7.040 195.415 7.085 ;
        RECT 175.345 6.900 195.415 7.040 ;
        RECT 175.345 6.855 175.635 6.900 ;
        RECT 195.125 6.855 195.415 6.900 ;
        RECT 248.945 3.300 249.235 3.345 ;
        RECT 296.770 3.300 297.090 3.360 ;
        RECT 248.945 3.160 297.090 3.300 ;
        RECT 248.945 3.115 249.235 3.160 ;
        RECT 296.770 3.100 297.090 3.160 ;
        RECT 2.385 1.600 2.675 1.645 ;
        RECT 26.305 1.600 26.595 1.645 ;
        RECT 2.385 1.460 26.595 1.600 ;
        RECT 2.385 1.415 2.675 1.460 ;
        RECT 26.305 1.415 26.595 1.460 ;
        RECT 48.845 1.600 49.135 1.645 ;
        RECT 133.945 1.600 134.235 1.645 ;
        RECT 48.845 1.460 134.235 1.600 ;
        RECT 48.845 1.415 49.135 1.460 ;
        RECT 133.945 1.415 134.235 1.460 ;
        RECT 195.125 1.600 195.415 1.645 ;
        RECT 198.805 1.600 199.095 1.645 ;
        RECT 195.125 1.460 199.095 1.600 ;
        RECT 195.125 1.415 195.415 1.460 ;
        RECT 198.805 1.415 199.095 1.460 ;
        RECT 198.805 0.920 199.095 0.965 ;
        RECT 248.945 0.920 249.235 0.965 ;
        RECT 198.805 0.780 249.235 0.920 ;
        RECT 198.805 0.735 199.095 0.780 ;
        RECT 248.945 0.735 249.235 0.780 ;
        RECT 29.985 0.580 30.275 0.625 ;
        RECT 48.845 0.580 49.135 0.625 ;
        RECT 29.985 0.440 49.135 0.580 ;
        RECT 29.985 0.395 30.275 0.440 ;
        RECT 48.845 0.395 49.135 0.440 ;
      LAYER via ;
        RECT 2412.340 3416.020 2412.600 3416.280 ;
        RECT 2470.300 3416.020 2470.560 3416.280 ;
        RECT 2470.300 3401.740 2470.560 3402.000 ;
        RECT 2795.980 3401.400 2796.240 3401.660 ;
        RECT 3.320 51.720 3.580 51.980 ;
        RECT 2.400 50.700 2.660 50.960 ;
        RECT 2.400 43.220 2.660 43.480 ;
        RECT 296.800 7.520 297.060 7.780 ;
        RECT 334.520 7.520 334.780 7.780 ;
        RECT 296.800 3.100 297.060 3.360 ;
      LAYER met2 ;
        RECT 2412.340 3415.990 2412.600 3416.310 ;
        RECT 2470.300 3415.990 2470.560 3416.310 ;
        RECT 2412.400 3405.000 2412.540 3415.990 ;
        RECT 2412.270 3401.000 2412.550 3405.000 ;
        RECT 2470.360 3402.030 2470.500 3415.990 ;
        RECT 2795.970 3402.195 2796.250 3402.565 ;
        RECT 2470.300 3401.710 2470.560 3402.030 ;
        RECT 2796.040 3401.690 2796.180 3402.195 ;
        RECT 2795.980 3401.370 2796.240 3401.690 ;
        RECT 3.310 161.315 3.590 161.685 ;
        RECT 3.380 52.010 3.520 161.315 ;
        RECT 3.320 51.690 3.580 52.010 ;
        RECT 2.400 50.670 2.660 50.990 ;
        RECT 2.460 43.510 2.600 50.670 ;
        RECT 2.400 43.190 2.660 43.510 ;
        RECT 296.800 7.490 297.060 7.810 ;
        RECT 334.510 7.635 334.790 8.005 ;
        RECT 334.520 7.490 334.780 7.635 ;
        RECT 296.860 3.390 297.000 7.490 ;
        RECT 366.710 4.915 366.990 5.285 ;
        RECT 296.800 3.070 297.060 3.390 ;
        RECT 366.780 3.130 366.920 4.915 ;
        RECT 366.780 2.990 371.520 3.130 ;
        RECT 371.380 2.400 371.520 2.990 ;
        RECT 371.170 -4.800 371.730 2.400 ;
      LAYER via2 ;
        RECT 2795.970 3402.240 2796.250 3402.520 ;
        RECT 3.310 161.360 3.590 161.640 ;
        RECT 334.510 7.680 334.790 7.960 ;
        RECT 366.710 4.960 366.990 5.240 ;
      LAYER met3 ;
        RECT 2795.945 3402.530 2796.275 3402.545 ;
        RECT 2806.270 3402.530 2806.650 3402.540 ;
        RECT 2795.945 3402.230 2806.650 3402.530 ;
        RECT 2795.945 3402.215 2796.275 3402.230 ;
        RECT 2806.270 3402.220 2806.650 3402.230 ;
        RECT 3.285 161.660 3.615 161.665 ;
        RECT 3.030 161.650 3.615 161.660 ;
        RECT 3.030 161.350 3.840 161.650 ;
        RECT 3.030 161.340 3.615 161.350 ;
        RECT 3.285 161.335 3.615 161.340 ;
        RECT 334.485 7.970 334.815 7.985 ;
        RECT 365.510 7.970 365.890 7.980 ;
        RECT 334.485 7.670 365.890 7.970 ;
        RECT 334.485 7.655 334.815 7.670 ;
        RECT 365.510 7.660 365.890 7.670 ;
        RECT 365.510 5.250 365.890 5.260 ;
        RECT 366.685 5.250 367.015 5.265 ;
        RECT 365.510 4.950 367.015 5.250 ;
        RECT 365.510 4.940 365.890 4.950 ;
        RECT 366.685 4.935 367.015 4.950 ;
      LAYER via3 ;
        RECT 2806.300 3402.220 2806.620 3402.540 ;
        RECT 3.060 161.340 3.380 161.660 ;
        RECT 365.540 7.660 365.860 7.980 ;
        RECT 365.540 4.940 365.860 5.260 ;
      LAYER met4 ;
        RECT 2806.295 3402.215 2806.625 3402.545 ;
        RECT 2806.310 981.050 2806.610 3402.215 ;
        RECT 2805.390 980.750 2806.610 981.050 ;
        RECT 2805.390 974.250 2805.690 980.750 ;
        RECT 2805.390 973.950 2806.610 974.250 ;
        RECT 2806.310 168.450 2806.610 973.950 ;
        RECT 2806.310 168.150 2807.530 168.450 ;
        RECT 2807.230 162.090 2807.530 168.150 ;
        RECT 2.630 160.910 3.810 162.090 ;
        RECT 2806.790 160.910 2807.970 162.090 ;
        RECT 365.535 7.655 365.865 7.985 ;
        RECT 365.550 5.265 365.850 7.655 ;
        RECT 365.535 4.935 365.865 5.265 ;
      LAYER met5 ;
        RECT 2.420 160.700 2808.180 162.300 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 9.805 2553.145 9.975 2646.135 ;
        RECT 9.805 2487.525 9.975 2550.255 ;
        RECT 9.805 2311.745 9.975 2373.455 ;
        RECT 9.805 2195.805 9.975 2273.155 ;
        RECT 9.805 2128.485 9.975 2171.155 ;
        RECT 9.805 2036.345 9.975 2074.935 ;
        RECT 9.805 1967.325 9.975 2028.355 ;
        RECT 8.885 1883.685 9.055 1936.895 ;
        RECT 9.805 1701.105 9.975 1853.255 ;
        RECT 9.805 1645.685 9.975 1690.395 ;
        RECT 9.805 1574.965 9.975 1595.875 ;
        RECT 9.345 1548.105 9.515 1562.895 ;
        RECT 9.805 1346.825 9.975 1533.315 ;
        RECT 2.905 1259.105 3.075 1333.055 ;
        RECT 5.205 994.245 5.375 1004.275 ;
        RECT 7.505 1004.105 7.675 1023.655 ;
        RECT 7.965 990.845 8.135 993.735 ;
        RECT 9.345 980.305 9.515 991.015 ;
        RECT 5.665 694.365 5.835 728.535 ;
        RECT 3.365 587.095 3.535 630.275 ;
        RECT 3.365 586.925 4.455 587.095 ;
        RECT 4.285 538.305 4.455 586.925 ;
        RECT 5.205 451.945 5.375 473.535 ;
        RECT 7.045 347.225 7.215 452.115 ;
        RECT 8.425 331.585 8.595 347.395 ;
        RECT 9.805 238.595 9.975 331.755 ;
        RECT 9.345 238.425 9.975 238.595 ;
        RECT 9.345 217.175 9.515 238.425 ;
        RECT 9.345 217.005 9.975 217.175 ;
        RECT 9.805 149.345 9.975 217.005 ;
        RECT 0.605 84.745 0.775 121.295 ;
        RECT 7.045 5.185 7.215 51.935 ;
        RECT 8.425 51.765 8.595 84.915 ;
      LAYER mcon ;
        RECT 9.805 2645.965 9.975 2646.135 ;
        RECT 9.805 2550.085 9.975 2550.255 ;
        RECT 9.805 2373.285 9.975 2373.455 ;
        RECT 9.805 2272.985 9.975 2273.155 ;
        RECT 9.805 2170.985 9.975 2171.155 ;
        RECT 9.805 2074.765 9.975 2074.935 ;
        RECT 9.805 2028.185 9.975 2028.355 ;
        RECT 8.885 1936.725 9.055 1936.895 ;
        RECT 9.805 1853.085 9.975 1853.255 ;
        RECT 9.805 1690.225 9.975 1690.395 ;
        RECT 9.805 1595.705 9.975 1595.875 ;
        RECT 9.345 1562.725 9.515 1562.895 ;
        RECT 9.805 1533.145 9.975 1533.315 ;
        RECT 2.905 1332.885 3.075 1333.055 ;
        RECT 7.505 1023.485 7.675 1023.655 ;
        RECT 5.205 1004.105 5.375 1004.275 ;
        RECT 7.965 993.565 8.135 993.735 ;
        RECT 9.345 990.845 9.515 991.015 ;
        RECT 5.665 728.365 5.835 728.535 ;
        RECT 3.365 630.105 3.535 630.275 ;
        RECT 5.205 473.365 5.375 473.535 ;
        RECT 7.045 451.945 7.215 452.115 ;
        RECT 8.425 347.225 8.595 347.395 ;
        RECT 9.805 331.585 9.975 331.755 ;
        RECT 0.605 121.125 0.775 121.295 ;
        RECT 8.425 84.745 8.595 84.915 ;
        RECT 7.045 51.765 7.215 51.935 ;
      LAYER met1 ;
        RECT 7.890 2781.100 8.210 2781.160 ;
        RECT 9.730 2781.100 10.050 2781.160 ;
        RECT 7.890 2780.960 10.050 2781.100 ;
        RECT 7.890 2780.900 8.210 2780.960 ;
        RECT 9.730 2780.900 10.050 2780.960 ;
        RECT 9.730 2646.120 10.050 2646.180 ;
        RECT 9.535 2645.980 10.050 2646.120 ;
        RECT 9.730 2645.920 10.050 2645.980 ;
        RECT 9.730 2553.300 10.050 2553.360 ;
        RECT 9.535 2553.160 10.050 2553.300 ;
        RECT 9.730 2553.100 10.050 2553.160 ;
        RECT 9.730 2550.240 10.050 2550.300 ;
        RECT 9.535 2550.100 10.050 2550.240 ;
        RECT 9.730 2550.040 10.050 2550.100 ;
        RECT 9.730 2487.680 10.050 2487.740 ;
        RECT 9.535 2487.540 10.050 2487.680 ;
        RECT 9.730 2487.480 10.050 2487.540 ;
        RECT 9.730 2397.720 10.050 2397.980 ;
        RECT 9.820 2396.960 9.960 2397.720 ;
        RECT 9.730 2396.700 10.050 2396.960 ;
        RECT 9.730 2373.440 10.050 2373.500 ;
        RECT 9.535 2373.300 10.050 2373.440 ;
        RECT 9.730 2373.240 10.050 2373.300 ;
        RECT 9.730 2311.900 10.050 2311.960 ;
        RECT 9.535 2311.760 10.050 2311.900 ;
        RECT 9.730 2311.700 10.050 2311.760 ;
        RECT 9.730 2273.140 10.050 2273.200 ;
        RECT 9.535 2273.000 10.050 2273.140 ;
        RECT 9.730 2272.940 10.050 2273.000 ;
        RECT 9.730 2195.960 10.050 2196.020 ;
        RECT 9.535 2195.820 10.050 2195.960 ;
        RECT 9.730 2195.760 10.050 2195.820 ;
        RECT 9.730 2171.140 10.050 2171.200 ;
        RECT 9.535 2171.000 10.050 2171.140 ;
        RECT 9.730 2170.940 10.050 2171.000 ;
        RECT 9.730 2128.640 10.050 2128.700 ;
        RECT 9.535 2128.500 10.050 2128.640 ;
        RECT 9.730 2128.440 10.050 2128.500 ;
        RECT 9.730 2074.920 10.050 2074.980 ;
        RECT 9.730 2074.780 10.245 2074.920 ;
        RECT 9.730 2074.720 10.050 2074.780 ;
        RECT 9.730 2036.500 10.050 2036.560 ;
        RECT 9.535 2036.360 10.050 2036.500 ;
        RECT 9.730 2036.300 10.050 2036.360 ;
        RECT 9.730 2028.340 10.050 2028.400 ;
        RECT 9.535 2028.200 10.050 2028.340 ;
        RECT 9.730 2028.140 10.050 2028.200 ;
        RECT 9.730 1967.480 10.050 1967.540 ;
        RECT 9.535 1967.340 10.050 1967.480 ;
        RECT 9.730 1967.280 10.050 1967.340 ;
        RECT 8.825 1936.880 9.115 1936.925 ;
        RECT 9.730 1936.880 10.050 1936.940 ;
        RECT 8.825 1936.740 10.050 1936.880 ;
        RECT 8.825 1936.695 9.115 1936.740 ;
        RECT 9.730 1936.680 10.050 1936.740 ;
        RECT 8.825 1883.840 9.115 1883.885 ;
        RECT 9.730 1883.840 10.050 1883.900 ;
        RECT 8.825 1883.700 10.050 1883.840 ;
        RECT 8.825 1883.655 9.115 1883.700 ;
        RECT 9.730 1883.640 10.050 1883.700 ;
        RECT 9.730 1853.240 10.050 1853.300 ;
        RECT 9.535 1853.100 10.050 1853.240 ;
        RECT 9.730 1853.040 10.050 1853.100 ;
        RECT 9.730 1701.260 10.050 1701.320 ;
        RECT 9.535 1701.120 10.050 1701.260 ;
        RECT 9.730 1701.060 10.050 1701.120 ;
        RECT 9.730 1690.380 10.050 1690.440 ;
        RECT 9.535 1690.240 10.050 1690.380 ;
        RECT 9.730 1690.180 10.050 1690.240 ;
        RECT 9.730 1645.840 10.050 1645.900 ;
        RECT 9.535 1645.700 10.050 1645.840 ;
        RECT 9.730 1645.640 10.050 1645.700 ;
        RECT 9.730 1595.860 10.050 1595.920 ;
        RECT 9.535 1595.720 10.050 1595.860 ;
        RECT 9.730 1595.660 10.050 1595.720 ;
        RECT 9.730 1575.120 10.050 1575.180 ;
        RECT 9.535 1574.980 10.050 1575.120 ;
        RECT 9.730 1574.920 10.050 1574.980 ;
        RECT 9.285 1562.880 9.575 1562.925 ;
        RECT 9.730 1562.880 10.050 1562.940 ;
        RECT 9.285 1562.740 10.050 1562.880 ;
        RECT 9.285 1562.695 9.575 1562.740 ;
        RECT 9.730 1562.680 10.050 1562.740 ;
        RECT 9.285 1548.260 9.575 1548.305 ;
        RECT 9.730 1548.260 10.050 1548.320 ;
        RECT 9.285 1548.120 10.050 1548.260 ;
        RECT 9.285 1548.075 9.575 1548.120 ;
        RECT 9.730 1548.060 10.050 1548.120 ;
        RECT 9.730 1533.300 10.050 1533.360 ;
        RECT 9.535 1533.160 10.050 1533.300 ;
        RECT 9.730 1533.100 10.050 1533.160 ;
        RECT 9.730 1346.980 10.050 1347.040 ;
        RECT 9.535 1346.840 10.050 1346.980 ;
        RECT 9.730 1346.780 10.050 1346.840 ;
        RECT 2.845 1333.040 3.135 1333.085 ;
        RECT 9.730 1333.040 10.050 1333.100 ;
        RECT 2.845 1332.900 10.050 1333.040 ;
        RECT 2.845 1332.855 3.135 1332.900 ;
        RECT 9.730 1332.840 10.050 1332.900 ;
        RECT 2.830 1259.260 3.150 1259.320 ;
        RECT 2.635 1259.120 3.150 1259.260 ;
        RECT 2.830 1259.060 3.150 1259.120 ;
        RECT 2.830 1070.900 3.150 1070.960 ;
        RECT 9.730 1070.900 10.050 1070.960 ;
        RECT 2.830 1070.760 10.050 1070.900 ;
        RECT 2.830 1070.700 3.150 1070.760 ;
        RECT 9.730 1070.700 10.050 1070.760 ;
        RECT 7.445 1023.640 7.735 1023.685 ;
        RECT 9.730 1023.640 10.050 1023.700 ;
        RECT 7.445 1023.500 10.050 1023.640 ;
        RECT 7.445 1023.455 7.735 1023.500 ;
        RECT 9.730 1023.440 10.050 1023.500 ;
        RECT 5.145 1004.260 5.435 1004.305 ;
        RECT 7.445 1004.260 7.735 1004.305 ;
        RECT 5.145 1004.120 7.735 1004.260 ;
        RECT 5.145 1004.075 5.435 1004.120 ;
        RECT 7.445 1004.075 7.735 1004.120 ;
        RECT 5.145 994.400 5.435 994.445 ;
        RECT 5.145 994.260 5.820 994.400 ;
        RECT 5.145 994.215 5.435 994.260 ;
        RECT 5.680 993.720 5.820 994.260 ;
        RECT 7.905 993.720 8.195 993.765 ;
        RECT 5.680 993.580 8.195 993.720 ;
        RECT 7.905 993.535 8.195 993.580 ;
        RECT 7.905 991.000 8.195 991.045 ;
        RECT 9.285 991.000 9.575 991.045 ;
        RECT 7.905 990.860 9.575 991.000 ;
        RECT 7.905 990.815 8.195 990.860 ;
        RECT 9.285 990.815 9.575 990.860 ;
        RECT 9.285 980.460 9.575 980.505 ;
        RECT 9.730 980.460 10.050 980.520 ;
        RECT 9.285 980.320 10.050 980.460 ;
        RECT 9.285 980.275 9.575 980.320 ;
        RECT 9.730 980.260 10.050 980.320 ;
        RECT 5.130 833.920 5.450 833.980 ;
        RECT 9.730 833.920 10.050 833.980 ;
        RECT 5.130 833.780 10.050 833.920 ;
        RECT 5.130 833.720 5.450 833.780 ;
        RECT 9.730 833.720 10.050 833.780 ;
        RECT 5.130 818.960 5.450 819.020 ;
        RECT 7.430 818.960 7.750 819.020 ;
        RECT 5.130 818.820 7.750 818.960 ;
        RECT 5.130 818.760 5.450 818.820 ;
        RECT 7.430 818.760 7.750 818.820 ;
        RECT 7.430 800.600 7.750 800.660 ;
        RECT 7.060 800.460 7.750 800.600 ;
        RECT 7.060 799.580 7.200 800.460 ;
        RECT 7.430 800.400 7.750 800.460 ;
        RECT 7.060 799.440 9.960 799.580 ;
        RECT 9.820 799.300 9.960 799.440 ;
        RECT 9.730 799.040 10.050 799.300 ;
        RECT 5.605 728.520 5.895 728.565 ;
        RECT 9.270 728.520 9.590 728.580 ;
        RECT 5.605 728.380 9.590 728.520 ;
        RECT 5.605 728.335 5.895 728.380 ;
        RECT 9.270 728.320 9.590 728.380 ;
        RECT 5.605 694.520 5.895 694.565 ;
        RECT 9.730 694.520 10.050 694.580 ;
        RECT 5.605 694.380 10.050 694.520 ;
        RECT 5.605 694.335 5.895 694.380 ;
        RECT 9.730 694.320 10.050 694.380 ;
        RECT 3.305 630.260 3.595 630.305 ;
        RECT 8.350 630.260 8.670 630.320 ;
        RECT 3.305 630.120 8.670 630.260 ;
        RECT 3.305 630.075 3.595 630.120 ;
        RECT 8.350 630.060 8.670 630.120 ;
        RECT 4.225 538.460 4.515 538.505 ;
        RECT 9.730 538.460 10.050 538.520 ;
        RECT 4.225 538.320 10.050 538.460 ;
        RECT 4.225 538.275 4.515 538.320 ;
        RECT 9.730 538.260 10.050 538.320 ;
        RECT 5.145 473.520 5.435 473.565 ;
        RECT 9.730 473.520 10.050 473.580 ;
        RECT 5.145 473.380 10.050 473.520 ;
        RECT 5.145 473.335 5.435 473.380 ;
        RECT 9.730 473.320 10.050 473.380 ;
        RECT 5.145 452.100 5.435 452.145 ;
        RECT 6.985 452.100 7.275 452.145 ;
        RECT 5.145 451.960 7.275 452.100 ;
        RECT 5.145 451.915 5.435 451.960 ;
        RECT 6.985 451.915 7.275 451.960 ;
        RECT 6.985 347.380 7.275 347.425 ;
        RECT 8.365 347.380 8.655 347.425 ;
        RECT 6.985 347.240 8.655 347.380 ;
        RECT 6.985 347.195 7.275 347.240 ;
        RECT 8.365 347.195 8.655 347.240 ;
        RECT 8.365 331.740 8.655 331.785 ;
        RECT 9.745 331.740 10.035 331.785 ;
        RECT 8.365 331.600 10.035 331.740 ;
        RECT 8.365 331.555 8.655 331.600 ;
        RECT 9.745 331.555 10.035 331.600 ;
        RECT 0.530 149.500 0.850 149.560 ;
        RECT 9.745 149.500 10.035 149.545 ;
        RECT 0.530 149.360 10.035 149.500 ;
        RECT 0.530 149.300 0.850 149.360 ;
        RECT 9.745 149.315 10.035 149.360 ;
        RECT 0.530 121.280 0.850 121.340 ;
        RECT 0.335 121.140 0.850 121.280 ;
        RECT 0.530 121.080 0.850 121.140 ;
        RECT 0.545 84.900 0.835 84.945 ;
        RECT 8.365 84.900 8.655 84.945 ;
        RECT 0.545 84.760 8.655 84.900 ;
        RECT 0.545 84.715 0.835 84.760 ;
        RECT 8.365 84.715 8.655 84.760 ;
        RECT 6.985 51.920 7.275 51.965 ;
        RECT 8.365 51.920 8.655 51.965 ;
        RECT 6.985 51.780 8.655 51.920 ;
        RECT 6.985 51.735 7.275 51.780 ;
        RECT 8.365 51.735 8.655 51.780 ;
        RECT 311.490 7.040 311.810 7.100 ;
        RECT 344.150 7.040 344.470 7.100 ;
        RECT 311.490 6.900 344.470 7.040 ;
        RECT 311.490 6.840 311.810 6.900 ;
        RECT 344.150 6.840 344.470 6.900 ;
        RECT 6.985 5.340 7.275 5.385 ;
        RECT 25.370 5.340 25.690 5.400 ;
        RECT 6.985 5.200 25.690 5.340 ;
        RECT 6.985 5.155 7.275 5.200 ;
        RECT 25.370 5.140 25.690 5.200 ;
        RECT 27.670 5.340 27.990 5.400 ;
        RECT 311.490 5.340 311.810 5.400 ;
        RECT 27.670 5.200 311.810 5.340 ;
        RECT 27.670 5.140 27.990 5.200 ;
        RECT 311.490 5.140 311.810 5.200 ;
      LAYER via ;
        RECT 7.920 2780.900 8.180 2781.160 ;
        RECT 9.760 2780.900 10.020 2781.160 ;
        RECT 9.760 2645.920 10.020 2646.180 ;
        RECT 9.760 2553.100 10.020 2553.360 ;
        RECT 9.760 2550.040 10.020 2550.300 ;
        RECT 9.760 2487.480 10.020 2487.740 ;
        RECT 9.760 2397.720 10.020 2397.980 ;
        RECT 9.760 2396.700 10.020 2396.960 ;
        RECT 9.760 2373.240 10.020 2373.500 ;
        RECT 9.760 2311.700 10.020 2311.960 ;
        RECT 9.760 2272.940 10.020 2273.200 ;
        RECT 9.760 2195.760 10.020 2196.020 ;
        RECT 9.760 2170.940 10.020 2171.200 ;
        RECT 9.760 2128.440 10.020 2128.700 ;
        RECT 9.760 2074.720 10.020 2074.980 ;
        RECT 9.760 2036.300 10.020 2036.560 ;
        RECT 9.760 2028.140 10.020 2028.400 ;
        RECT 9.760 1967.280 10.020 1967.540 ;
        RECT 9.760 1936.680 10.020 1936.940 ;
        RECT 9.760 1883.640 10.020 1883.900 ;
        RECT 9.760 1853.040 10.020 1853.300 ;
        RECT 9.760 1701.060 10.020 1701.320 ;
        RECT 9.760 1690.180 10.020 1690.440 ;
        RECT 9.760 1645.640 10.020 1645.900 ;
        RECT 9.760 1595.660 10.020 1595.920 ;
        RECT 9.760 1574.920 10.020 1575.180 ;
        RECT 9.760 1562.680 10.020 1562.940 ;
        RECT 9.760 1548.060 10.020 1548.320 ;
        RECT 9.760 1533.100 10.020 1533.360 ;
        RECT 9.760 1346.780 10.020 1347.040 ;
        RECT 9.760 1332.840 10.020 1333.100 ;
        RECT 2.860 1259.060 3.120 1259.320 ;
        RECT 2.860 1070.700 3.120 1070.960 ;
        RECT 9.760 1070.700 10.020 1070.960 ;
        RECT 9.760 1023.440 10.020 1023.700 ;
        RECT 9.760 980.260 10.020 980.520 ;
        RECT 5.160 833.720 5.420 833.980 ;
        RECT 9.760 833.720 10.020 833.980 ;
        RECT 5.160 818.760 5.420 819.020 ;
        RECT 7.460 818.760 7.720 819.020 ;
        RECT 7.460 800.400 7.720 800.660 ;
        RECT 9.760 799.040 10.020 799.300 ;
        RECT 9.300 728.320 9.560 728.580 ;
        RECT 9.760 694.320 10.020 694.580 ;
        RECT 8.380 630.060 8.640 630.320 ;
        RECT 9.760 538.260 10.020 538.520 ;
        RECT 9.760 473.320 10.020 473.580 ;
        RECT 0.560 149.300 0.820 149.560 ;
        RECT 0.560 121.080 0.820 121.340 ;
        RECT 311.520 6.840 311.780 7.100 ;
        RECT 344.180 6.840 344.440 7.100 ;
        RECT 25.400 5.140 25.660 5.400 ;
        RECT 27.700 5.140 27.960 5.400 ;
        RECT 311.520 5.140 311.780 5.400 ;
      LAYER met2 ;
        RECT 7.920 2781.045 8.180 2781.190 ;
        RECT 7.910 2780.675 8.190 2781.045 ;
        RECT 9.760 2780.870 10.020 2781.190 ;
        RECT 9.820 2646.210 9.960 2780.870 ;
        RECT 9.760 2645.890 10.020 2646.210 ;
        RECT 9.760 2553.130 10.020 2553.390 ;
        RECT 9.760 2553.070 10.420 2553.130 ;
        RECT 9.820 2552.990 10.420 2553.070 ;
        RECT 10.280 2550.410 10.420 2552.990 ;
        RECT 9.820 2550.330 10.420 2550.410 ;
        RECT 9.760 2550.270 10.420 2550.330 ;
        RECT 9.760 2550.010 10.020 2550.270 ;
        RECT 9.760 2487.450 10.020 2487.770 ;
        RECT 9.820 2398.010 9.960 2487.450 ;
        RECT 9.760 2397.690 10.020 2398.010 ;
        RECT 9.760 2396.670 10.020 2396.990 ;
        RECT 9.820 2373.530 9.960 2396.670 ;
        RECT 9.760 2373.210 10.020 2373.530 ;
        RECT 9.760 2311.670 10.020 2311.990 ;
        RECT 9.820 2273.230 9.960 2311.670 ;
        RECT 9.760 2272.910 10.020 2273.230 ;
        RECT 9.760 2195.730 10.020 2196.050 ;
        RECT 9.820 2171.230 9.960 2195.730 ;
        RECT 9.760 2170.910 10.020 2171.230 ;
        RECT 9.760 2128.410 10.020 2128.730 ;
        RECT 9.820 2075.010 9.960 2128.410 ;
        RECT 9.760 2074.690 10.020 2075.010 ;
        RECT 9.760 2036.270 10.020 2036.590 ;
        RECT 9.820 2028.430 9.960 2036.270 ;
        RECT 9.760 2028.110 10.020 2028.430 ;
        RECT 9.760 1967.250 10.020 1967.570 ;
        RECT 9.820 1936.970 9.960 1967.250 ;
        RECT 9.760 1936.650 10.020 1936.970 ;
        RECT 9.760 1883.610 10.020 1883.930 ;
        RECT 9.820 1853.330 9.960 1883.610 ;
        RECT 9.760 1853.010 10.020 1853.330 ;
        RECT 9.760 1701.030 10.020 1701.350 ;
        RECT 9.820 1690.470 9.960 1701.030 ;
        RECT 9.760 1690.150 10.020 1690.470 ;
        RECT 9.760 1645.610 10.020 1645.930 ;
        RECT 9.820 1595.950 9.960 1645.610 ;
        RECT 9.760 1595.630 10.020 1595.950 ;
        RECT 9.760 1574.890 10.020 1575.210 ;
        RECT 9.820 1562.970 9.960 1574.890 ;
        RECT 9.760 1562.650 10.020 1562.970 ;
        RECT 9.760 1548.030 10.020 1548.350 ;
        RECT 9.820 1533.390 9.960 1548.030 ;
        RECT 9.760 1533.070 10.020 1533.390 ;
        RECT 9.760 1346.750 10.020 1347.070 ;
        RECT 9.820 1333.130 9.960 1346.750 ;
        RECT 9.760 1332.810 10.020 1333.130 ;
        RECT 2.860 1259.030 3.120 1259.350 ;
        RECT 2.920 1070.990 3.060 1259.030 ;
        RECT 2.860 1070.670 3.120 1070.990 ;
        RECT 9.760 1070.730 10.020 1070.990 ;
        RECT 9.760 1070.670 10.420 1070.730 ;
        RECT 9.820 1070.590 10.420 1070.670 ;
        RECT 10.280 1023.810 10.420 1070.590 ;
        RECT 9.820 1023.730 10.420 1023.810 ;
        RECT 9.760 1023.670 10.420 1023.730 ;
        RECT 9.760 1023.410 10.020 1023.670 ;
        RECT 9.760 980.290 10.020 980.550 ;
        RECT 9.760 980.230 13.640 980.290 ;
        RECT 9.820 980.150 13.640 980.230 ;
        RECT 13.500 931.330 13.640 980.150 ;
        RECT 13.040 931.190 13.640 931.330 ;
        RECT 13.040 930.650 13.180 931.190 ;
        RECT 11.660 930.510 13.180 930.650 ;
        RECT 11.660 886.450 11.800 930.510 ;
        RECT 11.660 886.310 13.640 886.450 ;
        RECT 13.500 834.090 13.640 886.310 ;
        RECT 9.820 834.010 13.640 834.090 ;
        RECT 5.160 833.690 5.420 834.010 ;
        RECT 9.760 833.950 13.640 834.010 ;
        RECT 9.760 833.690 10.020 833.950 ;
        RECT 5.220 819.050 5.360 833.690 ;
        RECT 5.160 818.730 5.420 819.050 ;
        RECT 7.460 818.730 7.720 819.050 ;
        RECT 7.520 800.690 7.660 818.730 ;
        RECT 7.460 800.370 7.720 800.690 ;
        RECT 9.760 799.240 10.020 799.330 ;
        RECT 9.760 799.100 10.420 799.240 ;
        RECT 9.760 799.010 10.020 799.100 ;
        RECT 10.280 797.880 10.420 799.100 ;
        RECT 10.280 797.740 11.340 797.880 ;
        RECT 11.200 754.530 11.340 797.740 ;
        RECT 10.280 754.390 11.340 754.530 ;
        RECT 10.280 728.690 10.420 754.390 ;
        RECT 9.360 728.610 10.420 728.690 ;
        RECT 9.300 728.550 10.420 728.610 ;
        RECT 9.300 728.290 9.560 728.550 ;
        RECT 9.760 694.520 10.020 694.610 ;
        RECT 9.760 694.380 11.800 694.520 ;
        RECT 9.760 694.290 10.020 694.380 ;
        RECT 11.660 659.330 11.800 694.380 ;
        RECT 8.440 659.190 11.800 659.330 ;
        RECT 8.440 630.350 8.580 659.190 ;
        RECT 8.380 630.030 8.640 630.350 ;
        RECT 9.760 538.460 10.020 538.550 ;
        RECT 9.760 538.320 11.800 538.460 ;
        RECT 9.760 538.230 10.020 538.320 ;
        RECT 9.760 473.520 10.020 473.610 ;
        RECT 11.660 473.520 11.800 538.320 ;
        RECT 9.760 473.380 11.800 473.520 ;
        RECT 9.760 473.290 10.020 473.380 ;
        RECT 0.560 149.270 0.820 149.590 ;
        RECT 0.620 121.370 0.760 149.270 ;
        RECT 0.560 121.050 0.820 121.370 ;
        RECT 344.240 7.580 360.480 7.720 ;
        RECT 344.240 7.130 344.380 7.580 ;
        RECT 311.520 6.810 311.780 7.130 ;
        RECT 344.180 6.810 344.440 7.130 ;
        RECT 311.580 5.430 311.720 6.810 ;
        RECT 25.400 5.170 25.660 5.430 ;
        RECT 27.700 5.170 27.960 5.430 ;
        RECT 25.400 5.110 27.960 5.170 ;
        RECT 311.520 5.110 311.780 5.430 ;
        RECT 25.460 5.030 27.900 5.110 ;
        RECT 360.340 1.770 360.480 7.580 ;
        RECT 388.400 2.990 389.460 3.130 ;
        RECT 363.950 2.450 364.230 2.565 ;
        RECT 363.560 2.310 364.230 2.450 ;
        RECT 363.560 1.770 363.700 2.310 ;
        RECT 363.950 2.195 364.230 2.310 ;
        RECT 370.390 2.195 370.670 2.565 ;
        RECT 360.340 1.630 363.700 1.770 ;
        RECT 370.460 1.205 370.600 2.195 ;
        RECT 388.400 1.205 388.540 2.990 ;
        RECT 389.320 2.400 389.460 2.990 ;
        RECT 370.390 0.835 370.670 1.205 ;
        RECT 388.330 0.835 388.610 1.205 ;
        RECT 389.110 -4.800 389.670 2.400 ;
      LAYER via2 ;
        RECT 7.910 2780.720 8.190 2781.000 ;
        RECT 363.950 2.240 364.230 2.520 ;
        RECT 370.390 2.240 370.670 2.520 ;
        RECT 370.390 0.880 370.670 1.160 ;
        RECT 388.330 0.880 388.610 1.160 ;
      LAYER met3 ;
        RECT 5.000 2781.480 9.000 2782.080 ;
        RECT 7.670 2781.025 7.970 2781.480 ;
        RECT 7.670 2780.710 8.215 2781.025 ;
        RECT 7.885 2780.695 8.215 2780.710 ;
        RECT 363.925 2.530 364.255 2.545 ;
        RECT 370.365 2.530 370.695 2.545 ;
        RECT 363.925 2.230 370.695 2.530 ;
        RECT 363.925 2.215 364.255 2.230 ;
        RECT 370.365 2.215 370.695 2.230 ;
        RECT 370.365 1.170 370.695 1.185 ;
        RECT 388.305 1.170 388.635 1.185 ;
        RECT 370.365 0.870 388.635 1.170 ;
        RECT 370.365 0.855 370.695 0.870 ;
        RECT 388.305 0.855 388.635 0.870 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.170 4.235 68.450 4.605 ;
        RECT 68.240 2.400 68.380 4.235 ;
        RECT 68.030 -4.800 68.590 2.400 ;
      LAYER via2 ;
        RECT 68.170 4.280 68.450 4.560 ;
      LAYER met3 ;
        RECT 99.980 39.640 100.190 39.920 ;
        RECT 52.710 4.570 53.090 4.580 ;
        RECT 68.145 4.570 68.475 4.585 ;
        RECT 52.710 4.270 68.475 4.570 ;
        RECT 52.710 4.260 53.090 4.270 ;
        RECT 68.145 4.255 68.475 4.270 ;
      LAYER via3 ;
        RECT 52.740 4.260 53.060 4.580 ;
      LAYER met4 ;
        RECT 99.655 39.690 99.985 39.945 ;
        RECT 99.230 38.510 100.410 39.690 ;
        RECT 23.790 35.110 24.970 36.290 ;
        RECT 24.230 5.690 24.530 35.110 ;
        RECT 23.790 4.510 24.970 5.690 ;
        RECT 52.310 4.510 53.490 5.690 ;
        RECT 52.735 4.255 53.065 4.510 ;
      LAYER via4 ;
        RECT 52.310 4.510 53.490 5.690 ;
      LAYER met5 ;
        RECT 99.020 36.500 100.620 39.900 ;
        RECT 23.580 34.900 100.620 36.500 ;
        RECT 23.580 4.300 53.700 5.900 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 458.305 3.485 458.475 6.035 ;
        RECT 486.825 2.465 486.995 3.655 ;
        RECT 502.465 2.975 502.635 3.655 ;
        RECT 501.545 2.805 502.635 2.975 ;
        RECT 501.545 2.465 501.715 2.805 ;
        RECT 503.385 2.465 503.555 3.655 ;
        RECT 1207.645 2.805 1235.415 2.975 ;
        RECT 559.965 2.465 561.055 2.635 ;
        RECT 782.605 2.295 782.775 2.635 ;
        RECT 784.905 2.295 785.075 2.635 ;
        RECT 881.045 2.465 882.595 2.635 ;
        RECT 918.305 2.465 919.395 2.635 ;
        RECT 1207.645 2.465 1207.815 2.805 ;
        RECT 1235.245 2.635 1235.415 2.805 ;
        RECT 1235.245 2.465 1238.175 2.635 ;
        RECT 1304.245 2.465 1327.875 2.635 ;
        RECT 1344.265 2.465 1352.255 2.635 ;
        RECT 1352.545 2.465 1354.095 2.635 ;
        RECT 782.605 2.125 785.075 2.295 ;
        RECT 919.225 1.445 919.395 2.465 ;
        RECT 1487.785 1.785 1487.955 2.635 ;
        RECT 1594.045 2.295 1594.215 2.635 ;
        RECT 1680.065 2.465 1680.235 6.035 ;
        RECT 1694.325 2.465 1694.495 6.375 ;
        RECT 1594.045 2.125 1616.295 2.295 ;
        RECT 1741.705 1.785 1741.875 2.635 ;
        RECT 1783.105 1.785 1783.275 2.635 ;
        RECT 1932.145 2.465 1932.315 3.995 ;
        RECT 1979.985 2.465 1980.155 3.995 ;
        RECT 2125.345 2.465 2125.515 4.335 ;
        RECT 2154.325 2.465 2154.495 4.335 ;
        RECT 2318.545 2.465 2318.715 3.995 ;
        RECT 2365.925 2.465 2366.095 3.995 ;
        RECT 2366.845 2.465 2368.395 2.635 ;
        RECT 2405.485 2.465 2405.655 4.335 ;
        RECT 2544.405 2.465 2544.575 4.335 ;
        RECT 2573.845 2.465 2574.015 3.995 ;
      LAYER mcon ;
        RECT 1694.325 6.205 1694.495 6.375 ;
        RECT 458.305 5.865 458.475 6.035 ;
        RECT 1680.065 5.865 1680.235 6.035 ;
        RECT 486.825 3.485 486.995 3.655 ;
        RECT 502.465 3.485 502.635 3.655 ;
        RECT 503.385 3.485 503.555 3.655 ;
        RECT 560.885 2.465 561.055 2.635 ;
        RECT 782.605 2.465 782.775 2.635 ;
        RECT 784.905 2.465 785.075 2.635 ;
        RECT 882.425 2.465 882.595 2.635 ;
        RECT 1238.005 2.465 1238.175 2.635 ;
        RECT 1327.705 2.465 1327.875 2.635 ;
        RECT 1352.085 2.465 1352.255 2.635 ;
        RECT 1353.925 2.465 1354.095 2.635 ;
        RECT 1487.785 2.465 1487.955 2.635 ;
        RECT 1594.045 2.465 1594.215 2.635 ;
        RECT 2125.345 4.165 2125.515 4.335 ;
        RECT 1932.145 3.825 1932.315 3.995 ;
        RECT 1741.705 2.465 1741.875 2.635 ;
        RECT 1616.125 2.125 1616.295 2.295 ;
        RECT 1783.105 2.465 1783.275 2.635 ;
        RECT 1979.985 3.825 1980.155 3.995 ;
        RECT 2154.325 4.165 2154.495 4.335 ;
        RECT 2405.485 4.165 2405.655 4.335 ;
        RECT 2318.545 3.825 2318.715 3.995 ;
        RECT 2365.925 3.825 2366.095 3.995 ;
        RECT 2368.225 2.465 2368.395 2.635 ;
        RECT 2544.405 4.165 2544.575 4.335 ;
        RECT 2573.845 3.825 2574.015 3.995 ;
      LAYER met1 ;
        RECT 1694.265 6.360 1694.555 6.405 ;
        RECT 1688.360 6.220 1694.555 6.360 ;
        RECT 443.050 6.020 443.370 6.080 ;
        RECT 458.245 6.020 458.535 6.065 ;
        RECT 443.050 5.880 458.535 6.020 ;
        RECT 443.050 5.820 443.370 5.880 ;
        RECT 458.245 5.835 458.535 5.880 ;
        RECT 1680.005 6.020 1680.295 6.065 ;
        RECT 1688.360 6.020 1688.500 6.220 ;
        RECT 1694.265 6.175 1694.555 6.220 ;
        RECT 1680.005 5.880 1688.500 6.020 ;
        RECT 1680.005 5.835 1680.295 5.880 ;
        RECT 2125.285 4.320 2125.575 4.365 ;
        RECT 2154.265 4.320 2154.555 4.365 ;
        RECT 2125.285 4.180 2154.555 4.320 ;
        RECT 2125.285 4.135 2125.575 4.180 ;
        RECT 2154.265 4.135 2154.555 4.180 ;
        RECT 2405.425 4.320 2405.715 4.365 ;
        RECT 2544.345 4.320 2544.635 4.365 ;
        RECT 2405.425 4.180 2544.635 4.320 ;
        RECT 2405.425 4.135 2405.715 4.180 ;
        RECT 2544.345 4.135 2544.635 4.180 ;
        RECT 1932.085 3.980 1932.375 4.025 ;
        RECT 1979.925 3.980 1980.215 4.025 ;
        RECT 1932.085 3.840 1980.215 3.980 ;
        RECT 1932.085 3.795 1932.375 3.840 ;
        RECT 1979.925 3.795 1980.215 3.840 ;
        RECT 2318.485 3.980 2318.775 4.025 ;
        RECT 2365.865 3.980 2366.155 4.025 ;
        RECT 2318.485 3.840 2366.155 3.980 ;
        RECT 2318.485 3.795 2318.775 3.840 ;
        RECT 2365.865 3.795 2366.155 3.840 ;
        RECT 2573.785 3.980 2574.075 4.025 ;
        RECT 2593.550 3.980 2593.870 4.040 ;
        RECT 2573.785 3.840 2593.870 3.980 ;
        RECT 2573.785 3.795 2574.075 3.840 ;
        RECT 2593.550 3.780 2593.870 3.840 ;
        RECT 458.245 3.640 458.535 3.685 ;
        RECT 486.765 3.640 487.055 3.685 ;
        RECT 458.245 3.500 487.055 3.640 ;
        RECT 458.245 3.455 458.535 3.500 ;
        RECT 486.765 3.455 487.055 3.500 ;
        RECT 502.405 3.640 502.695 3.685 ;
        RECT 503.325 3.640 503.615 3.685 ;
        RECT 502.405 3.500 503.615 3.640 ;
        RECT 502.405 3.455 502.695 3.500 ;
        RECT 503.325 3.455 503.615 3.500 ;
        RECT 486.765 2.620 487.055 2.665 ;
        RECT 501.485 2.620 501.775 2.665 ;
        RECT 486.765 2.480 501.775 2.620 ;
        RECT 486.765 2.435 487.055 2.480 ;
        RECT 501.485 2.435 501.775 2.480 ;
        RECT 503.325 2.620 503.615 2.665 ;
        RECT 559.905 2.620 560.195 2.665 ;
        RECT 503.325 2.480 560.195 2.620 ;
        RECT 503.325 2.435 503.615 2.480 ;
        RECT 559.905 2.435 560.195 2.480 ;
        RECT 560.825 2.620 561.115 2.665 ;
        RECT 782.545 2.620 782.835 2.665 ;
        RECT 560.825 2.480 782.835 2.620 ;
        RECT 560.825 2.435 561.115 2.480 ;
        RECT 782.545 2.435 782.835 2.480 ;
        RECT 784.845 2.620 785.135 2.665 ;
        RECT 878.670 2.620 878.990 2.680 ;
        RECT 784.845 2.480 878.990 2.620 ;
        RECT 784.845 2.435 785.135 2.480 ;
        RECT 878.670 2.420 878.990 2.480 ;
        RECT 880.970 2.620 881.290 2.680 ;
        RECT 882.365 2.620 882.655 2.665 ;
        RECT 918.245 2.620 918.535 2.665 ;
        RECT 880.970 2.480 881.485 2.620 ;
        RECT 882.365 2.480 918.535 2.620 ;
        RECT 880.970 2.420 881.290 2.480 ;
        RECT 882.365 2.435 882.655 2.480 ;
        RECT 918.245 2.435 918.535 2.480 ;
        RECT 920.070 2.620 920.390 2.680 ;
        RECT 1087.510 2.620 1087.830 2.680 ;
        RECT 920.070 2.480 1087.830 2.620 ;
        RECT 920.070 2.420 920.390 2.480 ;
        RECT 1087.510 2.420 1087.830 2.480 ;
        RECT 1089.810 2.620 1090.130 2.680 ;
        RECT 1207.585 2.620 1207.875 2.665 ;
        RECT 1089.810 2.480 1207.875 2.620 ;
        RECT 1089.810 2.420 1090.130 2.480 ;
        RECT 1207.585 2.435 1207.875 2.480 ;
        RECT 1237.945 2.620 1238.235 2.665 ;
        RECT 1304.185 2.620 1304.475 2.665 ;
        RECT 1237.945 2.480 1257.940 2.620 ;
        RECT 1237.945 2.435 1238.235 2.480 ;
        RECT 1257.800 2.280 1257.940 2.480 ;
        RECT 1298.740 2.480 1304.475 2.620 ;
        RECT 1257.800 2.140 1258.400 2.280 ;
        RECT 1258.260 1.940 1258.400 2.140 ;
        RECT 1298.740 1.940 1298.880 2.480 ;
        RECT 1304.185 2.435 1304.475 2.480 ;
        RECT 1327.645 2.620 1327.935 2.665 ;
        RECT 1344.205 2.620 1344.495 2.665 ;
        RECT 1327.645 2.480 1344.495 2.620 ;
        RECT 1327.645 2.435 1327.935 2.480 ;
        RECT 1344.205 2.435 1344.495 2.480 ;
        RECT 1352.025 2.620 1352.315 2.665 ;
        RECT 1352.485 2.620 1352.775 2.665 ;
        RECT 1352.025 2.480 1352.775 2.620 ;
        RECT 1352.025 2.435 1352.315 2.480 ;
        RECT 1352.485 2.435 1352.775 2.480 ;
        RECT 1353.850 2.620 1354.170 2.680 ;
        RECT 1487.725 2.620 1488.015 2.665 ;
        RECT 1593.985 2.620 1594.275 2.665 ;
        RECT 1680.005 2.620 1680.295 2.665 ;
        RECT 1353.850 2.480 1354.365 2.620 ;
        RECT 1399.480 2.480 1450.220 2.620 ;
        RECT 1353.850 2.420 1354.170 2.480 ;
        RECT 1258.260 1.800 1298.880 1.940 ;
        RECT 1353.850 1.940 1354.170 2.000 ;
        RECT 1399.480 1.940 1399.620 2.480 ;
        RECT 1353.850 1.800 1399.620 1.940 ;
        RECT 1450.080 1.940 1450.220 2.480 ;
        RECT 1487.725 2.480 1594.275 2.620 ;
        RECT 1487.725 2.435 1488.015 2.480 ;
        RECT 1593.985 2.435 1594.275 2.480 ;
        RECT 1678.240 2.480 1680.295 2.620 ;
        RECT 1616.065 2.280 1616.355 2.325 ;
        RECT 1678.240 2.280 1678.380 2.480 ;
        RECT 1680.005 2.435 1680.295 2.480 ;
        RECT 1694.265 2.620 1694.555 2.665 ;
        RECT 1741.645 2.620 1741.935 2.665 ;
        RECT 1694.265 2.480 1741.935 2.620 ;
        RECT 1694.265 2.435 1694.555 2.480 ;
        RECT 1741.645 2.435 1741.935 2.480 ;
        RECT 1783.045 2.620 1783.335 2.665 ;
        RECT 1883.310 2.620 1883.630 2.680 ;
        RECT 1783.045 2.480 1883.630 2.620 ;
        RECT 1783.045 2.435 1783.335 2.480 ;
        RECT 1883.310 2.420 1883.630 2.480 ;
        RECT 1907.690 2.620 1908.010 2.680 ;
        RECT 1932.085 2.620 1932.375 2.665 ;
        RECT 1907.690 2.480 1932.375 2.620 ;
        RECT 1907.690 2.420 1908.010 2.480 ;
        RECT 1932.085 2.435 1932.375 2.480 ;
        RECT 1979.925 2.620 1980.215 2.665 ;
        RECT 2125.285 2.620 2125.575 2.665 ;
        RECT 1979.925 2.480 2125.575 2.620 ;
        RECT 1979.925 2.435 1980.215 2.480 ;
        RECT 2125.285 2.435 2125.575 2.480 ;
        RECT 2154.265 2.620 2154.555 2.665 ;
        RECT 2318.485 2.620 2318.775 2.665 ;
        RECT 2154.265 2.480 2318.775 2.620 ;
        RECT 2154.265 2.435 2154.555 2.480 ;
        RECT 2318.485 2.435 2318.775 2.480 ;
        RECT 2365.865 2.620 2366.155 2.665 ;
        RECT 2366.785 2.620 2367.075 2.665 ;
        RECT 2365.865 2.480 2367.075 2.620 ;
        RECT 2365.865 2.435 2366.155 2.480 ;
        RECT 2366.785 2.435 2367.075 2.480 ;
        RECT 2368.165 2.620 2368.455 2.665 ;
        RECT 2405.425 2.620 2405.715 2.665 ;
        RECT 2368.165 2.480 2405.715 2.620 ;
        RECT 2368.165 2.435 2368.455 2.480 ;
        RECT 2405.425 2.435 2405.715 2.480 ;
        RECT 2544.345 2.620 2544.635 2.665 ;
        RECT 2573.785 2.620 2574.075 2.665 ;
        RECT 2544.345 2.480 2574.075 2.620 ;
        RECT 2544.345 2.435 2544.635 2.480 ;
        RECT 2573.785 2.435 2574.075 2.480 ;
        RECT 1616.065 2.140 1678.380 2.280 ;
        RECT 1616.065 2.095 1616.355 2.140 ;
        RECT 1487.725 1.940 1488.015 1.985 ;
        RECT 1450.080 1.800 1488.015 1.940 ;
        RECT 1353.850 1.740 1354.170 1.800 ;
        RECT 1487.725 1.755 1488.015 1.800 ;
        RECT 1741.645 1.940 1741.935 1.985 ;
        RECT 1783.045 1.940 1783.335 1.985 ;
        RECT 1741.645 1.800 1783.335 1.940 ;
        RECT 1741.645 1.755 1741.935 1.800 ;
        RECT 1783.045 1.755 1783.335 1.800 ;
        RECT 919.165 1.600 919.455 1.645 ;
        RECT 920.070 1.600 920.390 1.660 ;
        RECT 919.165 1.460 920.390 1.600 ;
        RECT 919.165 1.415 919.455 1.460 ;
        RECT 920.070 1.400 920.390 1.460 ;
      LAYER via ;
        RECT 443.080 5.820 443.340 6.080 ;
        RECT 2593.580 3.780 2593.840 4.040 ;
        RECT 878.700 2.420 878.960 2.680 ;
        RECT 881.000 2.420 881.260 2.680 ;
        RECT 920.100 2.420 920.360 2.680 ;
        RECT 1087.540 2.420 1087.800 2.680 ;
        RECT 1089.840 2.420 1090.100 2.680 ;
        RECT 1353.880 2.420 1354.140 2.680 ;
        RECT 1353.880 1.740 1354.140 2.000 ;
        RECT 1883.340 2.420 1883.600 2.680 ;
        RECT 1907.720 2.420 1907.980 2.680 ;
        RECT 920.100 1.400 920.360 1.660 ;
      LAYER met2 ;
        RECT 443.080 5.790 443.340 6.110 ;
        RECT 443.140 2.960 443.280 5.790 ;
        RECT 2593.510 5.000 2593.790 9.000 ;
        RECT 2593.640 4.070 2593.780 5.000 ;
        RECT 1883.790 3.555 1884.070 3.925 ;
        RECT 1907.710 3.555 1907.990 3.925 ;
        RECT 2593.580 3.750 2593.840 4.070 ;
        RECT 442.680 2.820 443.280 2.960 ;
        RECT 442.680 2.400 442.820 2.820 ;
        RECT 878.700 2.450 878.960 2.710 ;
        RECT 881.000 2.620 881.260 2.710 ;
        RECT 880.140 2.480 881.260 2.620 ;
        RECT 880.140 2.450 880.280 2.480 ;
        RECT 442.470 -4.800 443.030 2.400 ;
        RECT 878.700 2.390 880.280 2.450 ;
        RECT 881.000 2.390 881.260 2.480 ;
        RECT 920.100 2.390 920.360 2.710 ;
        RECT 1087.540 2.390 1087.800 2.710 ;
        RECT 1089.840 2.620 1090.100 2.710 ;
        RECT 1089.440 2.480 1090.100 2.620 ;
        RECT 878.760 2.310 880.280 2.390 ;
        RECT 920.160 1.690 920.300 2.390 ;
        RECT 1087.600 1.770 1087.740 2.390 ;
        RECT 1089.440 1.770 1089.580 2.480 ;
        RECT 1089.840 2.390 1090.100 2.480 ;
        RECT 1353.880 2.390 1354.140 2.710 ;
        RECT 1883.340 2.450 1883.600 2.710 ;
        RECT 1883.860 2.450 1884.000 3.555 ;
        RECT 1907.780 2.710 1907.920 3.555 ;
        RECT 1883.340 2.390 1884.000 2.450 ;
        RECT 1907.720 2.390 1907.980 2.710 ;
        RECT 1353.940 2.030 1354.080 2.390 ;
        RECT 1883.400 2.310 1884.000 2.390 ;
        RECT 920.100 1.370 920.360 1.690 ;
        RECT 1087.600 1.630 1089.580 1.770 ;
        RECT 1353.880 1.710 1354.140 2.030 ;
      LAYER via2 ;
        RECT 1883.790 3.600 1884.070 3.880 ;
        RECT 1907.710 3.600 1907.990 3.880 ;
      LAYER met3 ;
        RECT 1883.765 3.890 1884.095 3.905 ;
        RECT 1907.685 3.890 1908.015 3.905 ;
        RECT 1883.765 3.590 1908.015 3.890 ;
        RECT 1883.765 3.575 1884.095 3.590 ;
        RECT 1907.685 3.575 1908.015 3.590 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1493.305 7.565 1500.835 7.735 ;
        RECT 1455.585 4.335 1455.755 6.375 ;
        RECT 1454.205 4.165 1455.755 4.335 ;
        RECT 1454.205 2.635 1454.375 4.165 ;
        RECT 1449.145 2.465 1454.375 2.635 ;
        RECT 880.125 2.125 882.135 2.295 ;
        RECT 880.125 1.955 880.295 2.125 ;
        RECT 879.665 1.785 880.295 1.955 ;
        RECT 881.965 1.785 882.135 2.125 ;
        RECT 917.845 1.615 918.015 1.955 ;
        RECT 966.605 1.785 980.115 1.955 ;
        RECT 917.845 1.445 918.935 1.615 ;
        RECT 979.945 0.595 980.115 1.785 ;
        RECT 997.425 0.595 997.595 1.955 ;
        RECT 1257.785 1.785 1299.355 1.955 ;
        RECT 1352.545 1.785 1400.555 1.955 ;
        RECT 1449.145 1.785 1449.315 2.465 ;
        RECT 1500.665 1.615 1500.835 7.565 ;
        RECT 1503.885 1.615 1504.055 1.955 ;
        RECT 1500.665 1.445 1504.055 1.615 ;
        RECT 1614.745 1.615 1614.915 1.955 ;
        RECT 1617.045 1.615 1617.215 1.955 ;
        RECT 1741.245 1.785 1741.415 4.675 ;
        RECT 1747.225 4.505 1747.395 8.755 ;
        RECT 1764.245 2.465 1764.415 8.755 ;
        RECT 1782.645 2.805 1783.735 2.975 ;
        RECT 1782.645 2.465 1782.815 2.805 ;
        RECT 1783.565 1.785 1783.735 2.805 ;
        RECT 1835.545 1.785 1843.075 1.955 ;
        RECT 1614.745 1.445 1617.215 1.615 ;
        RECT 1842.905 1.445 1843.075 1.785 ;
        RECT 1861.765 1.785 1863.315 1.955 ;
        RECT 1861.765 1.445 1861.935 1.785 ;
        RECT 1863.145 1.615 1863.315 1.785 ;
        RECT 1864.985 1.785 1866.075 1.955 ;
        RECT 2366.845 1.785 2368.395 1.955 ;
        RECT 2538.885 1.785 2539.515 1.955 ;
        RECT 1864.985 1.615 1865.155 1.785 ;
        RECT 1863.145 1.445 1865.155 1.615 ;
        RECT 979.945 0.425 997.595 0.595 ;
      LAYER mcon ;
        RECT 1747.225 8.585 1747.395 8.755 ;
        RECT 1455.585 6.205 1455.755 6.375 ;
        RECT 917.845 1.785 918.015 1.955 ;
        RECT 918.765 1.445 918.935 1.615 ;
        RECT 997.425 1.785 997.595 1.955 ;
        RECT 1299.185 1.785 1299.355 1.955 ;
        RECT 1400.385 1.785 1400.555 1.955 ;
        RECT 1741.245 4.505 1741.415 4.675 ;
        RECT 1764.245 8.585 1764.415 8.755 ;
        RECT 1503.885 1.785 1504.055 1.955 ;
        RECT 1614.745 1.785 1614.915 1.955 ;
        RECT 1617.045 1.785 1617.215 1.955 ;
        RECT 1865.905 1.785 1866.075 1.955 ;
        RECT 2368.225 1.785 2368.395 1.955 ;
        RECT 2539.345 1.785 2539.515 1.955 ;
      LAYER met1 ;
        RECT 1747.165 8.740 1747.455 8.785 ;
        RECT 1764.185 8.740 1764.475 8.785 ;
        RECT 1747.165 8.600 1764.475 8.740 ;
        RECT 1747.165 8.555 1747.455 8.600 ;
        RECT 1764.185 8.555 1764.475 8.600 ;
        RECT 1492.770 7.720 1493.090 7.780 ;
        RECT 1493.245 7.720 1493.535 7.765 ;
        RECT 1492.770 7.580 1493.535 7.720 ;
        RECT 1492.770 7.520 1493.090 7.580 ;
        RECT 1493.245 7.535 1493.535 7.580 ;
        RECT 1455.525 6.360 1455.815 6.405 ;
        RECT 1483.570 6.360 1483.890 6.420 ;
        RECT 1455.525 6.220 1483.890 6.360 ;
        RECT 1455.525 6.175 1455.815 6.220 ;
        RECT 1483.570 6.160 1483.890 6.220 ;
        RECT 1741.185 4.660 1741.475 4.705 ;
        RECT 1747.165 4.660 1747.455 4.705 ;
        RECT 1741.185 4.520 1747.455 4.660 ;
        RECT 1741.185 4.475 1741.475 4.520 ;
        RECT 1747.165 4.475 1747.455 4.520 ;
        RECT 1764.185 2.620 1764.475 2.665 ;
        RECT 1782.585 2.620 1782.875 2.665 ;
        RECT 1764.185 2.480 1782.875 2.620 ;
        RECT 1764.185 2.435 1764.475 2.480 ;
        RECT 1782.585 2.435 1782.875 2.480 ;
        RECT 479.390 1.940 479.710 2.000 ;
        RECT 559.430 1.940 559.750 2.000 ;
        RECT 479.390 1.800 559.750 1.940 ;
        RECT 479.390 1.740 479.710 1.800 ;
        RECT 559.430 1.740 559.750 1.800 ;
        RECT 560.350 1.940 560.670 2.000 ;
        RECT 765.970 1.940 766.290 2.000 ;
        RECT 560.350 1.800 766.290 1.940 ;
        RECT 560.350 1.740 560.670 1.800 ;
        RECT 765.970 1.740 766.290 1.800 ;
        RECT 786.210 1.940 786.530 2.000 ;
        RECT 879.605 1.940 879.895 1.985 ;
        RECT 786.210 1.800 879.895 1.940 ;
        RECT 786.210 1.740 786.530 1.800 ;
        RECT 879.605 1.755 879.895 1.800 ;
        RECT 881.905 1.940 882.195 1.985 ;
        RECT 917.785 1.940 918.075 1.985 ;
        RECT 966.545 1.940 966.835 1.985 ;
        RECT 881.905 1.800 918.075 1.940 ;
        RECT 881.905 1.755 882.195 1.800 ;
        RECT 917.785 1.755 918.075 1.800 ;
        RECT 918.780 1.800 966.835 1.940 ;
        RECT 918.780 1.645 918.920 1.800 ;
        RECT 966.545 1.755 966.835 1.800 ;
        RECT 997.365 1.940 997.655 1.985 ;
        RECT 1257.725 1.940 1258.015 1.985 ;
        RECT 997.365 1.800 1258.015 1.940 ;
        RECT 997.365 1.755 997.655 1.800 ;
        RECT 1257.725 1.755 1258.015 1.800 ;
        RECT 1299.125 1.940 1299.415 1.985 ;
        RECT 1352.485 1.940 1352.775 1.985 ;
        RECT 1299.125 1.800 1352.775 1.940 ;
        RECT 1299.125 1.755 1299.415 1.800 ;
        RECT 1352.485 1.755 1352.775 1.800 ;
        RECT 1400.325 1.940 1400.615 1.985 ;
        RECT 1449.085 1.940 1449.375 1.985 ;
        RECT 1400.325 1.800 1449.375 1.940 ;
        RECT 1400.325 1.755 1400.615 1.800 ;
        RECT 1449.085 1.755 1449.375 1.800 ;
        RECT 1503.825 1.940 1504.115 1.985 ;
        RECT 1614.685 1.940 1614.975 1.985 ;
        RECT 1503.825 1.800 1614.975 1.940 ;
        RECT 1503.825 1.755 1504.115 1.800 ;
        RECT 1614.685 1.755 1614.975 1.800 ;
        RECT 1616.985 1.940 1617.275 1.985 ;
        RECT 1741.185 1.940 1741.475 1.985 ;
        RECT 1616.985 1.800 1741.475 1.940 ;
        RECT 1616.985 1.755 1617.275 1.800 ;
        RECT 1741.185 1.755 1741.475 1.800 ;
        RECT 1783.505 1.940 1783.795 1.985 ;
        RECT 1835.485 1.940 1835.775 1.985 ;
        RECT 1783.505 1.800 1835.775 1.940 ;
        RECT 1783.505 1.755 1783.795 1.800 ;
        RECT 1835.485 1.755 1835.775 1.800 ;
        RECT 1865.845 1.940 1866.135 1.985 ;
        RECT 1883.310 1.940 1883.630 2.000 ;
        RECT 1865.845 1.800 1883.630 1.940 ;
        RECT 1865.845 1.755 1866.135 1.800 ;
        RECT 1883.310 1.740 1883.630 1.800 ;
        RECT 1885.150 1.940 1885.470 2.000 ;
        RECT 2366.785 1.940 2367.075 1.985 ;
        RECT 1885.150 1.800 2367.075 1.940 ;
        RECT 1885.150 1.740 1885.470 1.800 ;
        RECT 2366.785 1.755 2367.075 1.800 ;
        RECT 2368.165 1.940 2368.455 1.985 ;
        RECT 2538.825 1.940 2539.115 1.985 ;
        RECT 2368.165 1.800 2539.115 1.940 ;
        RECT 2368.165 1.755 2368.455 1.800 ;
        RECT 2538.825 1.755 2539.115 1.800 ;
        RECT 2539.285 1.940 2539.575 1.985 ;
        RECT 2640.930 1.940 2641.250 2.000 ;
        RECT 2539.285 1.800 2641.250 1.940 ;
        RECT 2539.285 1.755 2539.575 1.800 ;
        RECT 2640.930 1.740 2641.250 1.800 ;
        RECT 918.705 1.415 918.995 1.645 ;
        RECT 1842.845 1.600 1843.135 1.645 ;
        RECT 1861.705 1.600 1861.995 1.645 ;
        RECT 1842.845 1.460 1861.995 1.600 ;
        RECT 1842.845 1.415 1843.135 1.460 ;
        RECT 1861.705 1.415 1861.995 1.460 ;
      LAYER via ;
        RECT 1492.800 7.520 1493.060 7.780 ;
        RECT 1483.600 6.160 1483.860 6.420 ;
        RECT 479.420 1.740 479.680 2.000 ;
        RECT 559.460 1.740 559.720 2.000 ;
        RECT 560.380 1.740 560.640 2.000 ;
        RECT 766.000 1.740 766.260 2.000 ;
        RECT 786.240 1.740 786.500 2.000 ;
        RECT 1883.340 1.740 1883.600 2.000 ;
        RECT 1885.180 1.740 1885.440 2.000 ;
        RECT 2640.960 1.740 2641.220 2.000 ;
      LAYER met2 ;
        RECT 1483.660 7.810 1493.000 7.890 ;
        RECT 1483.660 7.750 1493.060 7.810 ;
        RECT 1483.660 6.450 1483.800 7.750 ;
        RECT 1492.800 7.490 1493.060 7.750 ;
        RECT 1483.600 6.130 1483.860 6.450 ;
        RECT 2640.890 5.000 2641.170 9.000 ;
        RECT 478.560 2.820 479.620 2.960 ;
        RECT 478.560 2.400 478.700 2.820 ;
        RECT 478.350 -4.800 478.910 2.400 ;
        RECT 479.480 2.030 479.620 2.820 ;
        RECT 559.450 2.195 559.730 2.565 ;
        RECT 560.370 2.195 560.650 2.565 ;
        RECT 559.520 2.030 559.660 2.195 ;
        RECT 560.440 2.030 560.580 2.195 ;
        RECT 2641.020 2.030 2641.160 5.000 ;
        RECT 479.420 1.710 479.680 2.030 ;
        RECT 559.460 1.710 559.720 2.030 ;
        RECT 560.380 1.710 560.640 2.030 ;
        RECT 766.000 1.770 766.260 2.030 ;
        RECT 766.450 1.770 766.730 1.885 ;
        RECT 766.000 1.710 766.730 1.770 ;
        RECT 766.060 1.630 766.730 1.710 ;
        RECT 766.450 1.515 766.730 1.630 ;
        RECT 784.390 1.770 784.670 1.885 ;
        RECT 786.240 1.770 786.500 2.030 ;
        RECT 784.390 1.710 786.500 1.770 ;
        RECT 1883.340 1.770 1883.600 2.030 ;
        RECT 1885.180 1.770 1885.440 2.030 ;
        RECT 1883.340 1.710 1885.440 1.770 ;
        RECT 2640.960 1.710 2641.220 2.030 ;
        RECT 784.390 1.630 786.440 1.710 ;
        RECT 1883.400 1.630 1885.380 1.710 ;
        RECT 784.390 1.515 784.670 1.630 ;
      LAYER via2 ;
        RECT 559.450 2.240 559.730 2.520 ;
        RECT 560.370 2.240 560.650 2.520 ;
        RECT 766.450 1.560 766.730 1.840 ;
        RECT 784.390 1.560 784.670 1.840 ;
      LAYER met3 ;
        RECT 559.425 2.530 559.755 2.545 ;
        RECT 560.345 2.530 560.675 2.545 ;
        RECT 559.425 2.230 560.675 2.530 ;
        RECT 559.425 2.215 559.755 2.230 ;
        RECT 560.345 2.215 560.675 2.230 ;
        RECT 766.425 1.850 766.755 1.865 ;
        RECT 784.365 1.850 784.695 1.865 ;
        RECT 766.425 1.550 784.695 1.850 ;
        RECT 766.425 1.535 766.755 1.550 ;
        RECT 784.365 1.535 784.695 1.550 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1400.845 9.265 1410.675 9.435 ;
        RECT 1400.845 8.585 1401.015 9.265 ;
        RECT 1311.145 8.245 1312.695 8.415 ;
        RECT 1301.485 7.905 1304.415 8.075 ;
        RECT 1311.145 7.905 1311.315 8.245 ;
        RECT 1312.525 8.075 1312.695 8.245 ;
        RECT 1312.525 7.905 1314.075 8.075 ;
        RECT 899.445 7.395 899.615 7.735 ;
        RECT 1352.545 7.395 1352.715 8.075 ;
        RECT 1410.505 7.735 1410.675 9.265 ;
        RECT 1452.825 9.265 1470.475 9.435 ;
        RECT 1452.825 7.735 1452.995 9.265 ;
        RECT 1410.505 7.565 1429.535 7.735 ;
        RECT 1448.225 7.565 1452.995 7.735 ;
        RECT 851.605 7.225 858.215 7.395 ;
        RECT 851.605 3.995 851.775 7.225 ;
        RECT 867.245 7.055 867.415 7.395 ;
        RECT 868.625 7.055 868.795 7.395 ;
        RECT 899.445 7.225 902.375 7.395 ;
        RECT 867.245 6.885 868.795 7.055 ;
        RECT 850.225 3.825 851.775 3.995 ;
        RECT 850.225 3.485 850.395 3.825 ;
        RECT 903.585 3.655 903.755 7.395 ;
        RECT 1352.545 7.225 1357.315 7.395 ;
        RECT 1470.305 5.865 1470.475 9.265 ;
        RECT 917.845 4.165 951.595 4.335 ;
        RECT 917.845 3.655 918.015 4.165 ;
        RECT 951.425 3.825 951.595 4.165 ;
        RECT 903.585 3.485 918.015 3.655 ;
        RECT 1040.205 2.975 1040.375 3.995 ;
        RECT 1044.805 3.825 1050.035 3.995 ;
        RECT 1044.805 2.975 1044.975 3.825 ;
        RECT 1049.865 3.655 1050.035 3.825 ;
        RECT 1049.865 3.485 1063.375 3.655 ;
        RECT 1476.285 3.485 1476.455 6.035 ;
        RECT 1040.205 2.805 1044.975 2.975 ;
        RECT 1063.205 2.635 1063.375 3.485 ;
        RECT 2366.845 3.145 2367.015 3.995 ;
        RECT 1063.205 2.465 1088.215 2.635 ;
      LAYER mcon ;
        RECT 1304.245 7.905 1304.415 8.075 ;
        RECT 1313.905 7.905 1314.075 8.075 ;
        RECT 1352.545 7.905 1352.715 8.075 ;
        RECT 899.445 7.565 899.615 7.735 ;
        RECT 1429.365 7.565 1429.535 7.735 ;
        RECT 858.045 7.225 858.215 7.395 ;
        RECT 867.245 7.225 867.415 7.395 ;
        RECT 868.625 7.225 868.795 7.395 ;
        RECT 902.205 7.225 902.375 7.395 ;
        RECT 903.585 7.225 903.755 7.395 ;
        RECT 1357.145 7.225 1357.315 7.395 ;
        RECT 1476.285 5.865 1476.455 6.035 ;
        RECT 1040.205 3.825 1040.375 3.995 ;
        RECT 2366.845 3.825 2367.015 3.995 ;
        RECT 1088.045 2.465 1088.215 2.635 ;
      LAYER met1 ;
        RECT 1400.310 8.740 1400.630 8.800 ;
        RECT 1400.785 8.740 1401.075 8.785 ;
        RECT 1400.310 8.600 1401.075 8.740 ;
        RECT 1400.310 8.540 1400.630 8.600 ;
        RECT 1400.785 8.555 1401.075 8.600 ;
        RECT 1190.550 8.060 1190.870 8.120 ;
        RECT 1193.310 8.060 1193.630 8.120 ;
        RECT 1190.550 7.920 1193.630 8.060 ;
        RECT 1190.550 7.860 1190.870 7.920 ;
        RECT 1193.310 7.860 1193.630 7.920 ;
        RECT 1193.770 8.060 1194.090 8.120 ;
        RECT 1301.425 8.060 1301.715 8.105 ;
        RECT 1193.770 7.920 1301.715 8.060 ;
        RECT 1193.770 7.860 1194.090 7.920 ;
        RECT 1301.425 7.875 1301.715 7.920 ;
        RECT 1304.185 8.060 1304.475 8.105 ;
        RECT 1311.085 8.060 1311.375 8.105 ;
        RECT 1304.185 7.920 1311.375 8.060 ;
        RECT 1304.185 7.875 1304.475 7.920 ;
        RECT 1311.085 7.875 1311.375 7.920 ;
        RECT 1313.845 8.060 1314.135 8.105 ;
        RECT 1352.485 8.060 1352.775 8.105 ;
        RECT 1313.845 7.920 1352.775 8.060 ;
        RECT 1313.845 7.875 1314.135 7.920 ;
        RECT 1352.485 7.875 1352.775 7.920 ;
        RECT 899.385 7.720 899.675 7.765 ;
        RECT 883.360 7.580 899.675 7.720 ;
        RECT 857.985 7.380 858.275 7.425 ;
        RECT 867.185 7.380 867.475 7.425 ;
        RECT 857.985 7.240 867.475 7.380 ;
        RECT 857.985 7.195 858.275 7.240 ;
        RECT 867.185 7.195 867.475 7.240 ;
        RECT 868.565 7.380 868.855 7.425 ;
        RECT 883.360 7.380 883.500 7.580 ;
        RECT 899.385 7.535 899.675 7.580 ;
        RECT 1429.305 7.720 1429.595 7.765 ;
        RECT 1448.165 7.720 1448.455 7.765 ;
        RECT 1429.305 7.580 1448.455 7.720 ;
        RECT 1429.305 7.535 1429.595 7.580 ;
        RECT 1448.165 7.535 1448.455 7.580 ;
        RECT 868.565 7.240 883.500 7.380 ;
        RECT 902.145 7.380 902.435 7.425 ;
        RECT 903.525 7.380 903.815 7.425 ;
        RECT 902.145 7.240 903.815 7.380 ;
        RECT 868.565 7.195 868.855 7.240 ;
        RECT 902.145 7.195 902.435 7.240 ;
        RECT 903.525 7.195 903.815 7.240 ;
        RECT 1357.085 7.380 1357.375 7.425 ;
        RECT 1361.210 7.380 1361.530 7.440 ;
        RECT 1357.085 7.240 1361.530 7.380 ;
        RECT 1357.085 7.195 1357.375 7.240 ;
        RECT 1361.210 7.180 1361.530 7.240 ;
        RECT 1165.710 6.360 1166.030 6.420 ;
        RECT 1190.550 6.360 1190.870 6.420 ;
        RECT 1165.710 6.220 1190.870 6.360 ;
        RECT 1165.710 6.160 1166.030 6.220 ;
        RECT 1190.550 6.160 1190.870 6.220 ;
        RECT 1470.245 6.020 1470.535 6.065 ;
        RECT 1476.225 6.020 1476.515 6.065 ;
        RECT 1470.245 5.880 1476.515 6.020 ;
        RECT 1470.245 5.835 1470.535 5.880 ;
        RECT 1476.225 5.835 1476.515 5.880 ;
        RECT 535.050 3.980 535.370 4.040 ;
        RECT 951.365 3.980 951.655 4.025 ;
        RECT 1040.145 3.980 1040.435 4.025 ;
        RECT 535.050 3.840 539.880 3.980 ;
        RECT 535.050 3.780 535.370 3.840 ;
        RECT 539.740 3.640 539.880 3.840 ;
        RECT 951.365 3.840 1040.435 3.980 ;
        RECT 951.365 3.795 951.655 3.840 ;
        RECT 1040.145 3.795 1040.435 3.840 ;
        RECT 2366.785 3.980 2367.075 4.025 ;
        RECT 2366.785 3.840 2368.380 3.980 ;
        RECT 2366.785 3.795 2367.075 3.840 ;
        RECT 557.590 3.640 557.910 3.700 ;
        RECT 539.740 3.500 557.910 3.640 ;
        RECT 557.590 3.440 557.910 3.500 ;
        RECT 560.350 3.640 560.670 3.700 ;
        RECT 760.910 3.640 761.230 3.700 ;
        RECT 560.350 3.500 761.230 3.640 ;
        RECT 560.350 3.440 560.670 3.500 ;
        RECT 760.910 3.440 761.230 3.500 ;
        RECT 819.790 3.640 820.110 3.700 ;
        RECT 819.790 3.500 845.320 3.640 ;
        RECT 819.790 3.440 820.110 3.500 ;
        RECT 845.180 3.300 845.320 3.500 ;
        RECT 850.165 3.455 850.455 3.685 ;
        RECT 1476.225 3.640 1476.515 3.685 ;
        RECT 1476.225 3.500 1597.420 3.640 ;
        RECT 1476.225 3.455 1476.515 3.500 ;
        RECT 850.240 3.300 850.380 3.455 ;
        RECT 845.180 3.160 850.380 3.300 ;
        RECT 1597.280 3.300 1597.420 3.500 ;
        RECT 1676.770 3.300 1677.090 3.360 ;
        RECT 1597.280 3.160 1677.090 3.300 ;
        RECT 1676.770 3.100 1677.090 3.160 ;
        RECT 1677.690 3.300 1678.010 3.360 ;
        RECT 2366.785 3.300 2367.075 3.345 ;
        RECT 1677.690 3.160 2367.075 3.300 ;
        RECT 2368.240 3.300 2368.380 3.840 ;
        RECT 2736.150 3.300 2736.470 3.360 ;
        RECT 2368.240 3.160 2736.470 3.300 ;
        RECT 1677.690 3.100 1678.010 3.160 ;
        RECT 2366.785 3.115 2367.075 3.160 ;
        RECT 2736.150 3.100 2736.470 3.160 ;
        RECT 1087.985 2.620 1088.275 2.665 ;
        RECT 1088.430 2.620 1088.750 2.680 ;
        RECT 1087.985 2.480 1088.750 2.620 ;
        RECT 1087.985 2.435 1088.275 2.480 ;
        RECT 1088.430 2.420 1088.750 2.480 ;
      LAYER via ;
        RECT 1400.340 8.540 1400.600 8.800 ;
        RECT 1190.580 7.860 1190.840 8.120 ;
        RECT 1193.340 7.860 1193.600 8.120 ;
        RECT 1193.800 7.860 1194.060 8.120 ;
        RECT 1361.240 7.180 1361.500 7.440 ;
        RECT 1165.740 6.160 1166.000 6.420 ;
        RECT 1190.580 6.160 1190.840 6.420 ;
        RECT 535.080 3.780 535.340 4.040 ;
        RECT 557.620 3.440 557.880 3.700 ;
        RECT 560.380 3.440 560.640 3.700 ;
        RECT 760.940 3.440 761.200 3.700 ;
        RECT 819.820 3.440 820.080 3.700 ;
        RECT 1676.800 3.100 1677.060 3.360 ;
        RECT 1677.720 3.100 1677.980 3.360 ;
        RECT 2736.180 3.100 2736.440 3.360 ;
        RECT 1088.460 2.420 1088.720 2.680 ;
      LAYER met2 ;
        RECT 1400.340 8.570 1400.600 8.830 ;
        RECT 1361.300 8.430 1367.420 8.570 ;
        RECT 1190.580 7.830 1190.840 8.150 ;
        RECT 1193.340 8.060 1193.600 8.150 ;
        RECT 1193.800 8.060 1194.060 8.150 ;
        RECT 1193.340 7.920 1194.060 8.060 ;
        RECT 1193.340 7.830 1193.600 7.920 ;
        RECT 1193.800 7.830 1194.060 7.920 ;
        RECT 517.590 6.275 517.870 6.645 ;
        RECT 533.690 6.275 533.970 6.645 ;
        RECT 1190.640 6.450 1190.780 7.830 ;
        RECT 1361.300 7.470 1361.440 8.430 ;
        RECT 1361.240 7.150 1361.500 7.470 ;
        RECT 517.660 5.000 517.800 6.275 ;
        RECT 533.760 5.340 533.900 6.275 ;
        RECT 1165.740 6.130 1166.000 6.450 ;
        RECT 1190.580 6.130 1190.840 6.450 ;
        RECT 765.140 5.540 768.040 5.680 ;
        RECT 533.760 5.200 535.280 5.340 ;
        RECT 515.820 4.860 517.800 5.000 ;
        RECT 513.980 2.820 515.040 2.960 ;
        RECT 513.980 2.400 514.120 2.820 ;
        RECT 514.900 2.450 515.040 2.820 ;
        RECT 515.820 2.450 515.960 4.860 ;
        RECT 535.140 4.070 535.280 5.200 ;
        RECT 557.680 4.180 559.200 4.320 ;
        RECT 535.080 3.750 535.340 4.070 ;
        RECT 557.680 3.730 557.820 4.180 ;
        RECT 557.620 3.410 557.880 3.730 ;
        RECT 559.060 3.245 559.200 4.180 ;
        RECT 560.380 3.410 560.640 3.730 ;
        RECT 760.940 3.640 761.200 3.730 ;
        RECT 765.140 3.640 765.280 5.540 ;
        RECT 767.900 5.285 768.040 5.540 ;
        RECT 785.380 5.540 786.900 5.680 ;
        RECT 785.380 5.285 785.520 5.540 ;
        RECT 767.830 4.915 768.110 5.285 ;
        RECT 785.310 4.915 785.590 5.285 ;
        RECT 786.760 4.660 786.900 5.540 ;
        RECT 786.760 4.520 789.660 4.660 ;
        RECT 1165.800 4.605 1165.940 6.130 ;
        RECT 1367.280 5.965 1367.420 8.430 ;
        RECT 1397.180 8.510 1400.600 8.570 ;
        RECT 1397.180 8.430 1400.540 8.510 ;
        RECT 1397.180 5.965 1397.320 8.430 ;
        RECT 1367.210 5.595 1367.490 5.965 ;
        RECT 1397.110 5.595 1397.390 5.965 ;
        RECT 2736.110 5.000 2736.390 9.000 ;
        RECT 760.940 3.500 765.280 3.640 ;
        RECT 760.940 3.410 761.200 3.500 ;
        RECT 560.440 3.245 560.580 3.410 ;
        RECT 789.520 3.245 789.660 4.520 ;
        RECT 818.500 4.180 820.020 4.320 ;
        RECT 1165.730 4.235 1166.010 4.605 ;
        RECT 818.500 3.925 818.640 4.180 ;
        RECT 818.430 3.555 818.710 3.925 ;
        RECT 819.880 3.730 820.020 4.180 ;
        RECT 819.820 3.410 820.080 3.730 ;
        RECT 1676.860 3.670 1677.920 3.810 ;
        RECT 1088.520 3.500 1089.580 3.640 ;
        RECT 558.990 2.875 559.270 3.245 ;
        RECT 560.370 2.875 560.650 3.245 ;
        RECT 789.450 2.875 789.730 3.245 ;
        RECT 1088.520 2.710 1088.660 3.500 ;
        RECT 1089.440 3.130 1089.580 3.500 ;
        RECT 1676.860 3.390 1677.000 3.670 ;
        RECT 1677.780 3.390 1677.920 3.670 ;
        RECT 2736.240 3.390 2736.380 5.000 ;
        RECT 1089.830 3.130 1090.110 3.245 ;
        RECT 1089.440 2.990 1090.110 3.130 ;
        RECT 1676.800 3.070 1677.060 3.390 ;
        RECT 1677.720 3.070 1677.980 3.390 ;
        RECT 2736.180 3.070 2736.440 3.390 ;
        RECT 1089.830 2.875 1090.110 2.990 ;
        RECT 513.770 -4.800 514.330 2.400 ;
        RECT 514.900 2.310 515.960 2.450 ;
        RECT 1088.460 2.390 1088.720 2.710 ;
      LAYER via2 ;
        RECT 517.590 6.320 517.870 6.600 ;
        RECT 533.690 6.320 533.970 6.600 ;
        RECT 767.830 4.960 768.110 5.240 ;
        RECT 785.310 4.960 785.590 5.240 ;
        RECT 1367.210 5.640 1367.490 5.920 ;
        RECT 1397.110 5.640 1397.390 5.920 ;
        RECT 1165.730 4.280 1166.010 4.560 ;
        RECT 818.430 3.600 818.710 3.880 ;
        RECT 558.990 2.920 559.270 3.200 ;
        RECT 560.370 2.920 560.650 3.200 ;
        RECT 789.450 2.920 789.730 3.200 ;
        RECT 1089.830 2.920 1090.110 3.200 ;
      LAYER met3 ;
        RECT 517.565 6.610 517.895 6.625 ;
        RECT 533.665 6.610 533.995 6.625 ;
        RECT 517.565 6.310 533.995 6.610 ;
        RECT 517.565 6.295 517.895 6.310 ;
        RECT 533.665 6.295 533.995 6.310 ;
        RECT 1367.185 5.930 1367.515 5.945 ;
        RECT 1397.085 5.930 1397.415 5.945 ;
        RECT 1367.185 5.630 1397.415 5.930 ;
        RECT 1367.185 5.615 1367.515 5.630 ;
        RECT 1397.085 5.615 1397.415 5.630 ;
        RECT 767.805 5.250 768.135 5.265 ;
        RECT 785.285 5.250 785.615 5.265 ;
        RECT 767.805 4.950 785.615 5.250 ;
        RECT 767.805 4.935 768.135 4.950 ;
        RECT 785.285 4.935 785.615 4.950 ;
        RECT 1164.070 4.570 1164.450 4.580 ;
        RECT 1165.705 4.570 1166.035 4.585 ;
        RECT 1164.070 4.270 1166.035 4.570 ;
        RECT 1164.070 4.260 1164.450 4.270 ;
        RECT 1165.705 4.255 1166.035 4.270 ;
        RECT 816.310 3.890 816.690 3.900 ;
        RECT 818.405 3.890 818.735 3.905 ;
        RECT 816.310 3.590 818.735 3.890 ;
        RECT 816.310 3.580 816.690 3.590 ;
        RECT 818.405 3.575 818.735 3.590 ;
        RECT 558.965 3.210 559.295 3.225 ;
        RECT 560.345 3.210 560.675 3.225 ;
        RECT 789.425 3.220 789.755 3.225 ;
        RECT 789.425 3.210 790.010 3.220 ;
        RECT 558.965 2.910 560.675 3.210 ;
        RECT 789.200 2.910 790.010 3.210 ;
        RECT 558.965 2.895 559.295 2.910 ;
        RECT 560.345 2.895 560.675 2.910 ;
        RECT 789.425 2.900 790.010 2.910 ;
        RECT 1089.805 3.210 1090.135 3.225 ;
        RECT 1095.990 3.210 1096.370 3.220 ;
        RECT 1089.805 2.910 1096.370 3.210 ;
        RECT 789.425 2.895 789.755 2.900 ;
        RECT 1089.805 2.895 1090.135 2.910 ;
        RECT 1095.990 2.900 1096.370 2.910 ;
      LAYER via3 ;
        RECT 1164.100 4.260 1164.420 4.580 ;
        RECT 816.340 3.580 816.660 3.900 ;
        RECT 789.660 2.900 789.980 3.220 ;
        RECT 1096.020 2.900 1096.340 3.220 ;
      LAYER met4 ;
        RECT 1162.270 4.950 1164.410 5.250 ;
        RECT 816.335 3.890 816.665 3.905 ;
        RECT 808.990 3.590 816.665 3.890 ;
        RECT 789.655 3.210 789.985 3.225 ;
        RECT 808.990 3.210 809.290 3.590 ;
        RECT 816.335 3.575 816.665 3.590 ;
        RECT 789.655 2.910 809.290 3.210 ;
        RECT 1096.015 3.210 1096.345 3.225 ;
        RECT 1096.015 2.910 1106.450 3.210 ;
        RECT 789.655 2.895 789.985 2.910 ;
        RECT 1096.015 2.895 1096.345 2.910 ;
        RECT 1106.150 1.850 1106.450 2.910 ;
        RECT 1162.270 2.290 1162.570 4.950 ;
        RECT 1164.110 4.585 1164.410 4.950 ;
        RECT 1164.095 4.255 1164.425 4.585 ;
        RECT 1123.190 1.850 1124.370 2.290 ;
        RECT 1106.150 1.550 1124.370 1.850 ;
        RECT 1123.190 1.110 1124.370 1.550 ;
        RECT 1161.830 1.110 1163.010 2.290 ;
      LAYER met5 ;
        RECT 1122.980 0.900 1163.220 2.500 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 8.425 2634.745 8.595 2635.595 ;
        RECT 8.425 2466.785 8.595 2511.495 ;
        RECT 8.885 2321.775 9.055 2360.535 ;
        RECT 8.425 2321.605 9.055 2321.775 ;
        RECT 8.425 2243.405 8.595 2321.605 ;
        RECT 176.325 7.565 176.495 9.095 ;
        RECT 96.745 3.825 97.375 3.995 ;
        RECT 197.945 3.145 198.115 9.095 ;
        RECT 512.585 7.565 517.355 7.735 ;
        RECT 459.225 5.015 459.395 5.355 ;
        RECT 460.145 5.185 461.235 5.355 ;
        RECT 460.145 5.015 460.315 5.185 ;
        RECT 459.225 4.845 460.315 5.015 ;
        RECT 461.065 5.015 461.235 5.185 ;
        RECT 512.585 5.015 512.755 7.565 ;
        RECT 461.065 4.845 462.615 5.015 ;
        RECT 462.445 4.675 462.615 4.845 ;
        RECT 509.365 4.845 512.755 5.015 ;
        RECT 462.445 4.505 464.915 4.675 ;
        RECT 509.365 4.505 509.535 4.845 ;
        RECT 464.745 3.825 464.915 4.505 ;
      LAYER mcon ;
        RECT 8.425 2635.425 8.595 2635.595 ;
        RECT 8.425 2511.325 8.595 2511.495 ;
        RECT 8.885 2360.365 9.055 2360.535 ;
        RECT 176.325 8.925 176.495 9.095 ;
        RECT 197.945 8.925 198.115 9.095 ;
        RECT 97.205 3.825 97.375 3.995 ;
        RECT 517.185 7.565 517.355 7.735 ;
        RECT 459.225 5.185 459.395 5.355 ;
      LAYER met1 ;
        RECT 7.890 3091.520 8.210 3091.580 ;
        RECT 8.350 3091.520 8.670 3091.580 ;
        RECT 7.890 3091.380 8.670 3091.520 ;
        RECT 7.890 3091.320 8.210 3091.380 ;
        RECT 8.350 3091.320 8.670 3091.380 ;
        RECT 8.350 2959.940 8.670 2960.000 ;
        RECT 9.270 2959.940 9.590 2960.000 ;
        RECT 8.350 2959.800 9.590 2959.940 ;
        RECT 8.350 2959.740 8.670 2959.800 ;
        RECT 9.270 2959.740 9.590 2959.800 ;
        RECT 8.350 2635.580 8.670 2635.640 ;
        RECT 8.155 2635.440 8.670 2635.580 ;
        RECT 8.350 2635.380 8.670 2635.440 ;
        RECT 8.365 2634.900 8.655 2634.945 ;
        RECT 8.810 2634.900 9.130 2634.960 ;
        RECT 8.365 2634.760 9.130 2634.900 ;
        RECT 8.365 2634.715 8.655 2634.760 ;
        RECT 8.810 2634.700 9.130 2634.760 ;
        RECT 8.810 2549.560 9.130 2549.620 ;
        RECT 8.440 2549.420 9.130 2549.560 ;
        RECT 8.440 2547.920 8.580 2549.420 ;
        RECT 8.810 2549.360 9.130 2549.420 ;
        RECT 8.350 2547.660 8.670 2547.920 ;
        RECT 8.350 2511.480 8.670 2511.540 ;
        RECT 8.155 2511.340 8.670 2511.480 ;
        RECT 8.350 2511.280 8.670 2511.340 ;
        RECT 8.365 2466.940 8.655 2466.985 ;
        RECT 9.270 2466.940 9.590 2467.000 ;
        RECT 8.365 2466.800 9.590 2466.940 ;
        RECT 8.365 2466.755 8.655 2466.800 ;
        RECT 9.270 2466.740 9.590 2466.800 ;
        RECT 8.810 2360.520 9.130 2360.580 ;
        RECT 8.615 2360.380 9.130 2360.520 ;
        RECT 8.810 2360.320 9.130 2360.380 ;
        RECT 8.350 2243.560 8.670 2243.620 ;
        RECT 8.155 2243.420 8.670 2243.560 ;
        RECT 8.350 2243.360 8.670 2243.420 ;
        RECT 6.970 2127.960 7.290 2128.020 ;
        RECT 8.810 2127.960 9.130 2128.020 ;
        RECT 6.970 2127.820 9.130 2127.960 ;
        RECT 6.970 2127.760 7.290 2127.820 ;
        RECT 8.810 2127.760 9.130 2127.820 ;
        RECT 6.970 2099.400 7.290 2099.460 ;
        RECT 8.350 2099.400 8.670 2099.460 ;
        RECT 6.970 2099.260 8.670 2099.400 ;
        RECT 6.970 2099.200 7.290 2099.260 ;
        RECT 8.350 2099.200 8.670 2099.260 ;
        RECT 6.970 2027.320 7.290 2027.380 ;
        RECT 8.810 2027.320 9.130 2027.380 ;
        RECT 6.970 2027.180 9.130 2027.320 ;
        RECT 6.970 2027.120 7.290 2027.180 ;
        RECT 8.810 2027.120 9.130 2027.180 ;
        RECT 6.970 1992.300 7.290 1992.360 ;
        RECT 8.810 1992.300 9.130 1992.360 ;
        RECT 6.970 1992.160 9.130 1992.300 ;
        RECT 6.970 1992.100 7.290 1992.160 ;
        RECT 8.810 1992.100 9.130 1992.160 ;
        RECT 8.810 1935.320 9.130 1935.580 ;
        RECT 8.900 1935.180 9.040 1935.320 ;
        RECT 7.060 1935.040 9.040 1935.180 ;
        RECT 7.060 1934.900 7.200 1935.040 ;
        RECT 6.970 1934.640 7.290 1934.900 ;
        RECT 6.970 1902.880 7.290 1902.940 ;
        RECT 8.810 1902.880 9.130 1902.940 ;
        RECT 6.970 1902.740 9.130 1902.880 ;
        RECT 6.970 1902.680 7.290 1902.740 ;
        RECT 8.810 1902.680 9.130 1902.740 ;
        RECT 6.970 1792.040 7.290 1792.100 ;
        RECT 8.810 1792.040 9.130 1792.100 ;
        RECT 6.970 1791.900 9.130 1792.040 ;
        RECT 6.970 1791.840 7.290 1791.900 ;
        RECT 8.810 1791.840 9.130 1791.900 ;
        RECT 6.970 1764.840 7.290 1764.900 ;
        RECT 8.810 1764.840 9.130 1764.900 ;
        RECT 6.970 1764.700 9.130 1764.840 ;
        RECT 6.970 1764.640 7.290 1764.700 ;
        RECT 8.810 1764.640 9.130 1764.700 ;
        RECT 6.970 1700.920 7.290 1700.980 ;
        RECT 8.810 1700.920 9.130 1700.980 ;
        RECT 6.970 1700.780 9.130 1700.920 ;
        RECT 6.970 1700.720 7.290 1700.780 ;
        RECT 8.810 1700.720 9.130 1700.780 ;
        RECT 6.970 1657.740 7.290 1657.800 ;
        RECT 8.810 1657.740 9.130 1657.800 ;
        RECT 6.970 1657.600 9.130 1657.740 ;
        RECT 6.970 1657.540 7.290 1657.600 ;
        RECT 8.810 1657.540 9.130 1657.600 ;
        RECT 5.590 1303.800 5.910 1303.860 ;
        RECT 8.810 1303.800 9.130 1303.860 ;
        RECT 5.590 1303.660 9.130 1303.800 ;
        RECT 5.590 1303.600 5.910 1303.660 ;
        RECT 8.810 1303.600 9.130 1303.660 ;
        RECT 5.590 83.540 5.910 83.600 ;
        RECT 5.590 83.400 9.960 83.540 ;
        RECT 5.590 83.340 5.910 83.400 ;
        RECT 9.820 81.560 9.960 83.400 ;
        RECT 9.730 81.300 10.050 81.560 ;
        RECT 7.430 78.780 7.750 78.840 ;
        RECT 9.730 78.780 10.050 78.840 ;
        RECT 7.430 78.640 10.050 78.780 ;
        RECT 7.430 78.580 7.750 78.640 ;
        RECT 9.730 78.580 10.050 78.640 ;
        RECT 7.430 75.720 7.750 75.780 ;
        RECT 7.430 75.580 9.500 75.720 ;
        RECT 7.430 75.520 7.750 75.580 ;
        RECT 9.360 74.080 9.500 75.580 ;
        RECT 9.270 73.820 9.590 74.080 ;
        RECT 176.265 9.080 176.555 9.125 ;
        RECT 197.885 9.080 198.175 9.125 ;
        RECT 176.265 8.940 198.175 9.080 ;
        RECT 176.265 8.895 176.555 8.940 ;
        RECT 197.885 8.895 198.175 8.940 ;
        RECT 141.750 7.720 142.070 7.780 ;
        RECT 176.265 7.720 176.555 7.765 ;
        RECT 141.750 7.580 176.555 7.720 ;
        RECT 141.750 7.520 142.070 7.580 ;
        RECT 176.265 7.535 176.555 7.580 ;
        RECT 517.125 7.720 517.415 7.765 ;
        RECT 518.490 7.720 518.810 7.780 ;
        RECT 517.125 7.580 518.810 7.720 ;
        RECT 517.125 7.535 517.415 7.580 ;
        RECT 518.490 7.520 518.810 7.580 ;
        RECT 414.990 5.340 415.310 5.400 ;
        RECT 459.165 5.340 459.455 5.385 ;
        RECT 414.990 5.200 459.455 5.340 ;
        RECT 414.990 5.140 415.310 5.200 ;
        RECT 459.165 5.155 459.455 5.200 ;
        RECT 508.370 4.660 508.690 4.720 ;
        RECT 509.305 4.660 509.595 4.705 ;
        RECT 508.370 4.520 509.595 4.660 ;
        RECT 508.370 4.460 508.690 4.520 ;
        RECT 509.305 4.475 509.595 4.520 ;
        RECT 547.010 4.320 547.330 4.380 ;
        RECT 549.770 4.320 550.090 4.380 ;
        RECT 547.010 4.180 550.090 4.320 ;
        RECT 547.010 4.120 547.330 4.180 ;
        RECT 549.770 4.120 550.090 4.180 ;
        RECT 15.250 3.980 15.570 4.040 ;
        RECT 96.685 3.980 96.975 4.025 ;
        RECT 15.250 3.840 96.975 3.980 ;
        RECT 15.250 3.780 15.570 3.840 ;
        RECT 96.685 3.795 96.975 3.840 ;
        RECT 97.130 3.980 97.450 4.040 ;
        RECT 464.685 3.980 464.975 4.025 ;
        RECT 465.130 3.980 465.450 4.040 ;
        RECT 97.130 3.840 97.645 3.980 ;
        RECT 464.685 3.840 465.450 3.980 ;
        RECT 97.130 3.780 97.450 3.840 ;
        RECT 464.685 3.795 464.975 3.840 ;
        RECT 465.130 3.780 465.450 3.840 ;
        RECT 197.885 3.300 198.175 3.345 ;
        RECT 233.750 3.300 234.070 3.360 ;
        RECT 197.885 3.160 234.070 3.300 ;
        RECT 197.885 3.115 198.175 3.160 ;
        RECT 233.750 3.100 234.070 3.160 ;
      LAYER via ;
        RECT 7.920 3091.320 8.180 3091.580 ;
        RECT 8.380 3091.320 8.640 3091.580 ;
        RECT 8.380 2959.740 8.640 2960.000 ;
        RECT 9.300 2959.740 9.560 2960.000 ;
        RECT 8.380 2635.380 8.640 2635.640 ;
        RECT 8.840 2634.700 9.100 2634.960 ;
        RECT 8.840 2549.360 9.100 2549.620 ;
        RECT 8.380 2547.660 8.640 2547.920 ;
        RECT 8.380 2511.280 8.640 2511.540 ;
        RECT 9.300 2466.740 9.560 2467.000 ;
        RECT 8.840 2360.320 9.100 2360.580 ;
        RECT 8.380 2243.360 8.640 2243.620 ;
        RECT 7.000 2127.760 7.260 2128.020 ;
        RECT 8.840 2127.760 9.100 2128.020 ;
        RECT 7.000 2099.200 7.260 2099.460 ;
        RECT 8.380 2099.200 8.640 2099.460 ;
        RECT 7.000 2027.120 7.260 2027.380 ;
        RECT 8.840 2027.120 9.100 2027.380 ;
        RECT 7.000 1992.100 7.260 1992.360 ;
        RECT 8.840 1992.100 9.100 1992.360 ;
        RECT 8.840 1935.320 9.100 1935.580 ;
        RECT 7.000 1934.640 7.260 1934.900 ;
        RECT 7.000 1902.680 7.260 1902.940 ;
        RECT 8.840 1902.680 9.100 1902.940 ;
        RECT 7.000 1791.840 7.260 1792.100 ;
        RECT 8.840 1791.840 9.100 1792.100 ;
        RECT 7.000 1764.640 7.260 1764.900 ;
        RECT 8.840 1764.640 9.100 1764.900 ;
        RECT 7.000 1700.720 7.260 1700.980 ;
        RECT 8.840 1700.720 9.100 1700.980 ;
        RECT 7.000 1657.540 7.260 1657.800 ;
        RECT 8.840 1657.540 9.100 1657.800 ;
        RECT 5.620 1303.600 5.880 1303.860 ;
        RECT 8.840 1303.600 9.100 1303.860 ;
        RECT 5.620 83.340 5.880 83.600 ;
        RECT 9.760 81.300 10.020 81.560 ;
        RECT 7.460 78.580 7.720 78.840 ;
        RECT 9.760 78.580 10.020 78.840 ;
        RECT 7.460 75.520 7.720 75.780 ;
        RECT 9.300 73.820 9.560 74.080 ;
        RECT 141.780 7.520 142.040 7.780 ;
        RECT 518.520 7.520 518.780 7.780 ;
        RECT 415.020 5.140 415.280 5.400 ;
        RECT 508.400 4.460 508.660 4.720 ;
        RECT 547.040 4.120 547.300 4.380 ;
        RECT 549.800 4.120 550.060 4.380 ;
        RECT 15.280 3.780 15.540 4.040 ;
        RECT 97.160 3.780 97.420 4.040 ;
        RECT 465.160 3.780 465.420 4.040 ;
        RECT 233.780 3.100 234.040 3.360 ;
      LAYER met2 ;
        RECT 7.910 3118.635 8.190 3119.005 ;
        RECT 7.980 3091.610 8.120 3118.635 ;
        RECT 7.920 3091.290 8.180 3091.610 ;
        RECT 8.380 3091.290 8.640 3091.610 ;
        RECT 8.440 2960.030 8.580 3091.290 ;
        RECT 8.380 2959.710 8.640 2960.030 ;
        RECT 9.300 2959.710 9.560 2960.030 ;
        RECT 9.360 2901.290 9.500 2959.710 ;
        RECT 8.900 2901.150 9.500 2901.290 ;
        RECT 8.900 2846.210 9.040 2901.150 ;
        RECT 8.440 2846.070 9.040 2846.210 ;
        RECT 8.440 2635.670 8.580 2846.070 ;
        RECT 8.380 2635.350 8.640 2635.670 ;
        RECT 8.840 2634.670 9.100 2634.990 ;
        RECT 8.900 2549.650 9.040 2634.670 ;
        RECT 8.840 2549.330 9.100 2549.650 ;
        RECT 8.380 2547.630 8.640 2547.950 ;
        RECT 8.440 2511.570 8.580 2547.630 ;
        RECT 8.380 2511.250 8.640 2511.570 ;
        RECT 9.300 2466.710 9.560 2467.030 ;
        RECT 9.360 2417.810 9.500 2466.710 ;
        RECT 8.900 2417.670 9.500 2417.810 ;
        RECT 8.900 2360.610 9.040 2417.670 ;
        RECT 8.840 2360.290 9.100 2360.610 ;
        RECT 8.380 2243.330 8.640 2243.650 ;
        RECT 8.440 2210.410 8.580 2243.330 ;
        RECT 8.440 2210.270 9.040 2210.410 ;
        RECT 8.900 2128.050 9.040 2210.270 ;
        RECT 7.000 2127.730 7.260 2128.050 ;
        RECT 8.840 2127.730 9.100 2128.050 ;
        RECT 7.060 2099.490 7.200 2127.730 ;
        RECT 7.000 2099.170 7.260 2099.490 ;
        RECT 8.380 2099.170 8.640 2099.490 ;
        RECT 8.440 2073.730 8.580 2099.170 ;
        RECT 8.440 2073.590 9.040 2073.730 ;
        RECT 8.900 2027.410 9.040 2073.590 ;
        RECT 7.000 2027.090 7.260 2027.410 ;
        RECT 8.840 2027.090 9.100 2027.410 ;
        RECT 7.060 1992.390 7.200 2027.090 ;
        RECT 7.000 1992.070 7.260 1992.390 ;
        RECT 8.840 1992.070 9.100 1992.390 ;
        RECT 8.900 1935.610 9.040 1992.070 ;
        RECT 8.840 1935.290 9.100 1935.610 ;
        RECT 7.000 1934.610 7.260 1934.930 ;
        RECT 7.060 1902.970 7.200 1934.610 ;
        RECT 7.000 1902.650 7.260 1902.970 ;
        RECT 8.840 1902.650 9.100 1902.970 ;
        RECT 8.900 1792.130 9.040 1902.650 ;
        RECT 7.000 1791.810 7.260 1792.130 ;
        RECT 8.840 1791.810 9.100 1792.130 ;
        RECT 7.060 1764.930 7.200 1791.810 ;
        RECT 7.000 1764.610 7.260 1764.930 ;
        RECT 8.840 1764.610 9.100 1764.930 ;
        RECT 8.900 1701.010 9.040 1764.610 ;
        RECT 7.000 1700.690 7.260 1701.010 ;
        RECT 8.840 1700.690 9.100 1701.010 ;
        RECT 7.060 1657.830 7.200 1700.690 ;
        RECT 7.000 1657.510 7.260 1657.830 ;
        RECT 8.840 1657.510 9.100 1657.830 ;
        RECT 8.900 1303.890 9.040 1657.510 ;
        RECT 5.620 1303.570 5.880 1303.890 ;
        RECT 8.840 1303.570 9.100 1303.890 ;
        RECT 5.680 83.630 5.820 1303.570 ;
        RECT 5.620 83.310 5.880 83.630 ;
        RECT 9.760 81.270 10.020 81.590 ;
        RECT 9.820 78.870 9.960 81.270 ;
        RECT 7.460 78.550 7.720 78.870 ;
        RECT 9.760 78.550 10.020 78.870 ;
        RECT 7.520 75.810 7.660 78.550 ;
        RECT 7.460 75.490 7.720 75.810 ;
        RECT 9.300 73.790 9.560 74.110 ;
        RECT 9.360 62.970 9.500 73.790 ;
        RECT 9.360 62.830 15.480 62.970 ;
        RECT 15.340 4.070 15.480 62.830 ;
        RECT 518.580 8.260 535.740 8.400 ;
        RECT 518.580 7.810 518.720 8.260 ;
        RECT 141.780 7.490 142.040 7.810 ;
        RECT 518.520 7.490 518.780 7.810 ;
        RECT 15.280 3.750 15.540 4.070 ;
        RECT 97.160 3.980 97.420 4.070 ;
        RECT 97.160 3.840 99.200 3.980 ;
        RECT 97.160 3.750 97.420 3.840 ;
        RECT 99.060 1.885 99.200 3.840 ;
        RECT 141.840 1.885 141.980 7.490 ;
        RECT 410.870 5.595 411.150 5.965 ;
        RECT 412.780 5.710 415.220 5.850 ;
        RECT 410.940 5.340 411.080 5.595 ;
        RECT 412.780 5.340 412.920 5.710 ;
        RECT 415.080 5.430 415.220 5.710 ;
        RECT 233.770 4.915 234.050 5.285 ;
        RECT 410.940 5.200 412.920 5.340 ;
        RECT 415.020 5.110 415.280 5.430 ;
        RECT 535.600 5.285 535.740 8.260 ;
        RECT 465.220 5.030 470.880 5.170 ;
        RECT 233.840 3.390 233.980 4.915 ;
        RECT 465.220 4.070 465.360 5.030 ;
        RECT 465.160 3.750 465.420 4.070 ;
        RECT 233.780 3.070 234.040 3.390 ;
        RECT 98.990 1.515 99.270 1.885 ;
        RECT 141.770 1.515 142.050 1.885 ;
        RECT 470.740 0.525 470.880 5.030 ;
        RECT 535.530 4.915 535.810 5.285 ;
        RECT 545.190 4.915 545.470 5.285 ;
        RECT 508.400 4.660 508.660 4.750 ;
        RECT 505.700 4.520 508.660 4.660 ;
        RECT 505.700 1.770 505.840 4.520 ;
        RECT 508.400 4.430 508.660 4.520 ;
        RECT 545.260 4.320 545.400 4.915 ;
        RECT 547.040 4.320 547.300 4.410 ;
        RECT 545.260 4.180 547.300 4.320 ;
        RECT 547.040 4.090 547.300 4.180 ;
        RECT 549.800 4.090 550.060 4.410 ;
        RECT 549.860 2.400 550.000 4.090 ;
        RECT 505.240 1.630 505.840 1.770 ;
        RECT 505.240 0.525 505.380 1.630 ;
        RECT 470.670 0.155 470.950 0.525 ;
        RECT 505.170 0.155 505.450 0.525 ;
        RECT 549.650 -4.800 550.210 2.400 ;
      LAYER via2 ;
        RECT 7.910 3118.680 8.190 3118.960 ;
        RECT 410.870 5.640 411.150 5.920 ;
        RECT 233.770 4.960 234.050 5.240 ;
        RECT 98.990 1.560 99.270 1.840 ;
        RECT 141.770 1.560 142.050 1.840 ;
        RECT 535.530 4.960 535.810 5.240 ;
        RECT 545.190 4.960 545.470 5.240 ;
        RECT 470.670 0.200 470.950 0.480 ;
        RECT 505.170 0.200 505.450 0.480 ;
      LAYER met3 ;
        RECT 5.000 3121.480 9.000 3122.080 ;
        RECT 7.670 3118.985 7.970 3121.480 ;
        RECT 7.670 3118.670 8.215 3118.985 ;
        RECT 7.885 3118.655 8.215 3118.670 ;
        RECT 334.230 5.930 334.610 5.940 ;
        RECT 410.845 5.930 411.175 5.945 ;
        RECT 334.230 5.630 411.175 5.930 ;
        RECT 334.230 5.620 334.610 5.630 ;
        RECT 410.845 5.615 411.175 5.630 ;
        RECT 233.745 5.260 234.075 5.265 ;
        RECT 233.745 5.250 234.330 5.260 ;
        RECT 233.520 4.950 234.330 5.250 ;
        RECT 233.745 4.940 234.330 4.950 ;
        RECT 535.505 5.250 535.835 5.265 ;
        RECT 545.165 5.250 545.495 5.265 ;
        RECT 535.505 4.950 545.495 5.250 ;
        RECT 233.745 4.935 234.075 4.940 ;
        RECT 535.505 4.935 535.835 4.950 ;
        RECT 545.165 4.935 545.495 4.950 ;
        RECT 98.965 1.850 99.295 1.865 ;
        RECT 141.745 1.850 142.075 1.865 ;
        RECT 98.965 1.550 142.075 1.850 ;
        RECT 98.965 1.535 99.295 1.550 ;
        RECT 141.745 1.535 142.075 1.550 ;
        RECT 470.645 0.490 470.975 0.505 ;
        RECT 505.145 0.490 505.475 0.505 ;
        RECT 470.645 0.190 505.475 0.490 ;
        RECT 470.645 0.175 470.975 0.190 ;
        RECT 505.145 0.175 505.475 0.190 ;
      LAYER via3 ;
        RECT 334.260 5.620 334.580 5.940 ;
        RECT 233.980 4.940 234.300 5.260 ;
      LAYER met4 ;
        RECT 334.255 5.690 334.585 5.945 ;
        RECT 233.550 4.510 234.730 5.690 ;
        RECT 333.830 4.510 335.010 5.690 ;
      LAYER met5 ;
        RECT 233.340 4.300 335.220 5.900 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 6.125 975.205 6.295 1038.615 ;
        RECT 6.125 883.065 6.295 944.775 ;
        RECT 3.825 734.825 3.995 798.235 ;
        RECT 8.425 798.065 8.595 836.315 ;
        RECT 7.045 456.705 7.215 693.175 ;
        RECT 8.885 362.015 9.055 431.035 ;
        RECT 8.885 361.845 9.515 362.015 ;
        RECT 7.965 321.215 8.135 327.335 ;
        RECT 9.345 327.165 9.515 361.845 ;
        RECT 7.965 321.045 8.595 321.215 ;
        RECT 8.425 217.855 8.595 321.045 ;
        RECT 7.965 217.685 8.595 217.855 ;
        RECT 7.965 213.945 8.135 217.685 ;
        RECT 5.665 147.985 5.835 197.455 ;
        RECT 9.345 100.385 9.515 148.155 ;
        RECT 542.025 9.605 560.135 9.775 ;
        RECT 542.025 9.435 542.195 9.605 ;
        RECT 531.905 9.265 542.195 9.435 ;
        RECT 559.965 9.435 560.135 9.605 ;
        RECT 559.965 9.265 562.435 9.435 ;
        RECT 437.145 7.905 466.295 8.075 ;
        RECT 407.705 7.225 409.715 7.395 ;
        RECT 407.705 6.715 407.875 7.225 ;
        RECT 393.445 6.545 407.875 6.715 ;
        RECT 393.445 6.205 393.615 6.545 ;
        RECT 409.545 0.595 409.715 7.225 ;
        RECT 420.125 7.225 429.035 7.395 ;
        RECT 420.125 0.595 420.295 7.225 ;
        RECT 428.865 6.715 429.035 7.225 ;
        RECT 428.865 6.545 429.955 6.715 ;
        RECT 429.785 6.375 429.955 6.545 ;
        RECT 430.245 6.375 430.415 7.055 ;
        RECT 437.145 6.885 437.315 7.905 ;
        RECT 429.785 6.205 430.415 6.375 ;
        RECT 466.125 5.525 466.295 7.905 ;
        RECT 517.645 4.165 517.815 5.695 ;
        RECT 531.905 4.165 532.075 9.265 ;
        RECT 562.265 9.095 562.435 9.265 ;
        RECT 562.265 8.925 563.355 9.095 ;
        RECT 563.185 3.995 563.355 8.925 ;
        RECT 563.185 3.825 564.735 3.995 ;
        RECT 409.545 0.425 420.295 0.595 ;
      LAYER mcon ;
        RECT 6.125 1038.445 6.295 1038.615 ;
        RECT 6.125 944.605 6.295 944.775 ;
        RECT 8.425 836.145 8.595 836.315 ;
        RECT 3.825 798.065 3.995 798.235 ;
        RECT 7.045 693.005 7.215 693.175 ;
        RECT 8.885 430.865 9.055 431.035 ;
        RECT 7.965 327.165 8.135 327.335 ;
        RECT 5.665 197.285 5.835 197.455 ;
        RECT 9.345 147.985 9.515 148.155 ;
        RECT 430.245 6.885 430.415 7.055 ;
        RECT 517.645 5.525 517.815 5.695 ;
        RECT 564.565 3.825 564.735 3.995 ;
      LAYER met1 ;
        RECT 6.050 1038.600 6.370 1038.660 ;
        RECT 5.855 1038.460 6.370 1038.600 ;
        RECT 6.050 1038.400 6.370 1038.460 ;
        RECT 6.065 975.360 6.355 975.405 ;
        RECT 9.730 975.360 10.050 975.420 ;
        RECT 6.065 975.220 10.050 975.360 ;
        RECT 6.065 975.175 6.355 975.220 ;
        RECT 9.730 975.160 10.050 975.220 ;
        RECT 6.065 944.760 6.355 944.805 ;
        RECT 9.730 944.760 10.050 944.820 ;
        RECT 6.065 944.620 10.050 944.760 ;
        RECT 6.065 944.575 6.355 944.620 ;
        RECT 9.730 944.560 10.050 944.620 ;
        RECT 6.065 883.220 6.355 883.265 ;
        RECT 9.730 883.220 10.050 883.280 ;
        RECT 6.065 883.080 10.050 883.220 ;
        RECT 6.065 883.035 6.355 883.080 ;
        RECT 9.730 883.020 10.050 883.080 ;
        RECT 8.365 836.300 8.655 836.345 ;
        RECT 9.730 836.300 10.050 836.360 ;
        RECT 8.365 836.160 10.050 836.300 ;
        RECT 8.365 836.115 8.655 836.160 ;
        RECT 9.730 836.100 10.050 836.160 ;
        RECT 3.765 798.220 4.055 798.265 ;
        RECT 8.365 798.220 8.655 798.265 ;
        RECT 3.765 798.080 8.655 798.220 ;
        RECT 3.765 798.035 4.055 798.080 ;
        RECT 8.365 798.035 8.655 798.080 ;
        RECT 3.750 734.980 4.070 735.040 ;
        RECT 3.555 734.840 4.070 734.980 ;
        RECT 3.750 734.780 4.070 734.840 ;
        RECT 3.750 693.640 4.070 693.900 ;
        RECT 3.840 693.160 3.980 693.640 ;
        RECT 6.985 693.160 7.275 693.205 ;
        RECT 3.840 693.020 7.275 693.160 ;
        RECT 6.985 692.975 7.275 693.020 ;
        RECT 6.985 456.860 7.275 456.905 ;
        RECT 9.730 456.860 10.050 456.920 ;
        RECT 6.985 456.720 10.050 456.860 ;
        RECT 6.985 456.675 7.275 456.720 ;
        RECT 9.730 456.660 10.050 456.720 ;
        RECT 8.825 431.020 9.115 431.065 ;
        RECT 9.730 431.020 10.050 431.080 ;
        RECT 8.825 430.880 10.050 431.020 ;
        RECT 8.825 430.835 9.115 430.880 ;
        RECT 9.730 430.820 10.050 430.880 ;
        RECT 7.905 327.320 8.195 327.365 ;
        RECT 9.285 327.320 9.575 327.365 ;
        RECT 7.905 327.180 9.575 327.320 ;
        RECT 7.905 327.135 8.195 327.180 ;
        RECT 9.285 327.135 9.575 327.180 ;
        RECT 7.905 214.100 8.195 214.145 ;
        RECT 9.730 214.100 10.050 214.160 ;
        RECT 7.905 213.960 10.050 214.100 ;
        RECT 7.905 213.915 8.195 213.960 ;
        RECT 9.730 213.900 10.050 213.960 ;
        RECT 5.605 197.440 5.895 197.485 ;
        RECT 9.730 197.440 10.050 197.500 ;
        RECT 5.605 197.300 10.050 197.440 ;
        RECT 5.605 197.255 5.895 197.300 ;
        RECT 9.730 197.240 10.050 197.300 ;
        RECT 5.605 148.140 5.895 148.185 ;
        RECT 9.285 148.140 9.575 148.185 ;
        RECT 5.605 148.000 9.575 148.140 ;
        RECT 5.605 147.955 5.895 148.000 ;
        RECT 9.285 147.955 9.575 148.000 ;
        RECT 9.285 100.540 9.575 100.585 ;
        RECT 3.840 100.400 9.575 100.540 ;
        RECT 3.840 99.240 3.980 100.400 ;
        RECT 9.285 100.355 9.575 100.400 ;
        RECT 3.750 98.980 4.070 99.240 ;
        RECT 3.750 23.700 4.070 23.760 ;
        RECT 9.730 23.700 10.050 23.760 ;
        RECT 3.750 23.560 10.050 23.700 ;
        RECT 3.750 23.500 4.070 23.560 ;
        RECT 9.730 23.500 10.050 23.560 ;
        RECT 65.020 7.240 196.720 7.380 ;
        RECT 53.430 7.040 53.750 7.100 ;
        RECT 65.020 7.040 65.160 7.240 ;
        RECT 53.430 6.900 65.160 7.040 ;
        RECT 53.430 6.840 53.750 6.900 ;
        RECT 196.580 6.700 196.720 7.240 ;
        RECT 430.185 7.040 430.475 7.085 ;
        RECT 437.085 7.040 437.375 7.085 ;
        RECT 430.185 6.900 437.375 7.040 ;
        RECT 430.185 6.855 430.475 6.900 ;
        RECT 437.085 6.855 437.375 6.900 ;
        RECT 235.130 6.700 235.450 6.760 ;
        RECT 196.580 6.560 235.450 6.700 ;
        RECT 235.130 6.500 235.450 6.560 ;
        RECT 318.390 6.360 318.710 6.420 ;
        RECT 393.385 6.360 393.675 6.405 ;
        RECT 318.390 6.220 393.675 6.360 ;
        RECT 318.390 6.160 318.710 6.220 ;
        RECT 393.385 6.175 393.675 6.220 ;
        RECT 466.065 5.680 466.355 5.725 ;
        RECT 517.585 5.680 517.875 5.725 ;
        RECT 466.065 5.540 517.875 5.680 ;
        RECT 466.065 5.495 466.355 5.540 ;
        RECT 517.585 5.495 517.875 5.540 ;
        RECT 517.585 4.320 517.875 4.365 ;
        RECT 531.845 4.320 532.135 4.365 ;
        RECT 517.585 4.180 532.135 4.320 ;
        RECT 517.585 4.135 517.875 4.180 ;
        RECT 531.845 4.135 532.135 4.180 ;
        RECT 564.505 3.980 564.795 4.025 ;
        RECT 567.710 3.980 568.030 4.040 ;
        RECT 564.505 3.840 568.030 3.980 ;
        RECT 564.505 3.795 564.795 3.840 ;
        RECT 567.710 3.780 568.030 3.840 ;
      LAYER via ;
        RECT 6.080 1038.400 6.340 1038.660 ;
        RECT 9.760 975.160 10.020 975.420 ;
        RECT 9.760 944.560 10.020 944.820 ;
        RECT 9.760 883.020 10.020 883.280 ;
        RECT 9.760 836.100 10.020 836.360 ;
        RECT 3.780 734.780 4.040 735.040 ;
        RECT 3.780 693.640 4.040 693.900 ;
        RECT 9.760 456.660 10.020 456.920 ;
        RECT 9.760 430.820 10.020 431.080 ;
        RECT 9.760 213.900 10.020 214.160 ;
        RECT 9.760 197.240 10.020 197.500 ;
        RECT 3.780 98.980 4.040 99.240 ;
        RECT 3.780 23.500 4.040 23.760 ;
        RECT 9.760 23.500 10.020 23.760 ;
        RECT 53.460 6.840 53.720 7.100 ;
        RECT 235.160 6.500 235.420 6.760 ;
        RECT 318.420 6.160 318.680 6.420 ;
        RECT 567.740 3.780 568.000 4.040 ;
      LAYER met2 ;
        RECT 6.070 3233.555 6.350 3233.925 ;
        RECT 6.140 1038.690 6.280 3233.555 ;
        RECT 6.080 1038.370 6.340 1038.690 ;
        RECT 9.820 975.450 12.260 975.530 ;
        RECT 9.760 975.390 12.260 975.450 ;
        RECT 9.760 975.130 10.020 975.390 ;
        RECT 12.120 946.970 12.260 975.390 ;
        RECT 11.660 946.830 12.260 946.970 ;
        RECT 9.760 944.760 10.020 944.850 ;
        RECT 11.660 944.760 11.800 946.830 ;
        RECT 9.760 944.620 11.800 944.760 ;
        RECT 9.760 944.530 10.020 944.620 ;
        RECT 9.760 883.050 10.020 883.310 ;
        RECT 9.760 882.990 11.800 883.050 ;
        RECT 9.820 882.910 11.800 882.990 ;
        RECT 11.660 882.540 11.800 882.910 ;
        RECT 11.660 882.400 12.260 882.540 ;
        RECT 9.760 836.300 10.020 836.390 ;
        RECT 12.120 836.300 12.260 882.400 ;
        RECT 9.760 836.160 12.260 836.300 ;
        RECT 9.760 836.070 10.020 836.160 ;
        RECT 3.780 734.750 4.040 735.070 ;
        RECT 3.840 693.930 3.980 734.750 ;
        RECT 3.780 693.610 4.040 693.930 ;
        RECT 9.760 456.690 10.020 456.950 ;
        RECT 9.760 456.630 10.420 456.690 ;
        RECT 9.820 456.550 10.420 456.630 ;
        RECT 10.280 431.530 10.420 456.550 ;
        RECT 9.820 431.390 10.420 431.530 ;
        RECT 9.820 431.110 9.960 431.390 ;
        RECT 9.760 430.790 10.020 431.110 ;
        RECT 9.760 213.930 10.020 214.190 ;
        RECT 9.760 213.870 10.420 213.930 ;
        RECT 9.820 213.790 10.420 213.870 ;
        RECT 10.280 197.610 10.420 213.790 ;
        RECT 9.820 197.530 10.420 197.610 ;
        RECT 9.760 197.470 10.420 197.530 ;
        RECT 9.760 197.210 10.020 197.470 ;
        RECT 3.780 98.950 4.040 99.270 ;
        RECT 3.840 23.790 3.980 98.950 ;
        RECT 3.780 23.470 4.040 23.790 ;
        RECT 9.760 23.470 10.020 23.790 ;
        RECT 9.820 1.885 9.960 23.470 ;
        RECT 53.460 6.810 53.720 7.130 ;
        RECT 53.520 1.885 53.660 6.810 ;
        RECT 235.160 6.470 235.420 6.790 ;
        RECT 235.220 5.285 235.360 6.470 ;
        RECT 317.560 6.450 318.620 6.530 ;
        RECT 317.560 6.390 318.680 6.450 ;
        RECT 317.560 5.285 317.700 6.390 ;
        RECT 318.420 6.130 318.680 6.390 ;
        RECT 235.150 4.915 235.430 5.285 ;
        RECT 317.490 4.915 317.770 5.285 ;
        RECT 567.740 3.750 568.000 4.070 ;
        RECT 567.800 2.400 567.940 3.750 ;
        RECT 9.750 1.515 10.030 1.885 ;
        RECT 53.450 1.515 53.730 1.885 ;
        RECT 567.590 -4.800 568.150 2.400 ;
      LAYER via2 ;
        RECT 6.070 3233.600 6.350 3233.880 ;
        RECT 235.150 4.960 235.430 5.240 ;
        RECT 317.490 4.960 317.770 5.240 ;
        RECT 9.750 1.560 10.030 1.840 ;
        RECT 53.450 1.560 53.730 1.840 ;
      LAYER met3 ;
        RECT 5.000 3234.360 9.000 3234.960 ;
        RECT 5.830 3233.905 6.130 3234.360 ;
        RECT 5.830 3233.590 6.375 3233.905 ;
        RECT 6.045 3233.575 6.375 3233.590 ;
        RECT 235.125 5.250 235.455 5.265 ;
        RECT 317.465 5.250 317.795 5.265 ;
        RECT 235.125 4.950 317.795 5.250 ;
        RECT 235.125 4.935 235.455 4.950 ;
        RECT 317.465 4.935 317.795 4.950 ;
        RECT 9.725 1.850 10.055 1.865 ;
        RECT 53.425 1.850 53.755 1.865 ;
        RECT 9.725 1.550 53.755 1.850 ;
        RECT 9.725 1.535 10.055 1.550 ;
        RECT 53.425 1.535 53.755 1.550 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2511.285 3396.005 2511.455 3401.955 ;
        RECT 2812.585 3396.005 2812.755 3401.615 ;
        RECT 1157.965 10.965 1162.275 11.135 ;
        RECT 1101.385 9.265 1103.855 9.435 ;
        RECT 1101.385 8.925 1101.555 9.265 ;
        RECT 1103.685 8.925 1103.855 9.265 ;
        RECT 1157.965 8.925 1158.135 10.965 ;
        RECT 760.065 3.825 761.615 3.995 ;
        RECT 761.445 3.485 761.615 3.825 ;
        RECT 785.825 3.315 785.995 3.655 ;
        RECT 772.485 3.145 773.115 3.315 ;
        RECT 783.525 3.145 785.995 3.315 ;
        RECT 799.625 0.935 799.795 3.655 ;
        RECT 830.905 3.485 831.995 3.655 ;
        RECT 811.585 0.935 811.755 3.315 ;
        RECT 815.265 2.975 815.435 3.315 ;
        RECT 830.905 2.975 831.075 3.485 ;
        RECT 815.265 2.805 831.075 2.975 ;
        RECT 831.825 2.635 831.995 3.485 ;
        RECT 851.605 2.635 851.775 3.315 ;
        RECT 831.825 2.465 851.775 2.635 ;
        RECT 881.505 1.615 881.675 1.955 ;
        RECT 900.825 1.615 900.995 6.035 ;
        RECT 902.665 5.865 902.835 8.755 ;
        RECT 1162.105 8.585 1162.275 10.965 ;
        RECT 1195.685 7.055 1195.855 8.755 ;
        RECT 1195.685 6.885 1197.235 7.055 ;
        RECT 1197.065 5.695 1197.235 6.885 ;
        RECT 1196.145 5.525 1197.235 5.695 ;
        RECT 1196.145 5.185 1196.315 5.525 ;
        RECT 881.505 1.445 900.995 1.615 ;
        RECT 799.625 0.765 811.755 0.935 ;
      LAYER mcon ;
        RECT 2511.285 3401.785 2511.455 3401.955 ;
        RECT 2812.585 3401.445 2812.755 3401.615 ;
        RECT 902.665 8.585 902.835 8.755 ;
        RECT 1195.685 8.585 1195.855 8.755 ;
        RECT 900.825 5.865 900.995 6.035 ;
        RECT 785.825 3.485 785.995 3.655 ;
        RECT 772.945 3.145 773.115 3.315 ;
        RECT 799.625 3.485 799.795 3.655 ;
        RECT 811.585 3.145 811.755 3.315 ;
        RECT 815.265 3.145 815.435 3.315 ;
        RECT 851.605 3.145 851.775 3.315 ;
        RECT 881.505 1.785 881.675 1.955 ;
      LAYER met1 ;
        RECT 2511.210 3401.940 2511.530 3402.000 ;
        RECT 2511.015 3401.800 2511.530 3401.940 ;
        RECT 2511.210 3401.740 2511.530 3401.800 ;
        RECT 2812.510 3401.600 2812.830 3401.660 ;
        RECT 2812.315 3401.460 2812.830 3401.600 ;
        RECT 2812.510 3401.400 2812.830 3401.460 ;
        RECT 2511.225 3396.160 2511.515 3396.205 ;
        RECT 2812.525 3396.160 2812.815 3396.205 ;
        RECT 2511.225 3396.020 2812.815 3396.160 ;
        RECT 2511.225 3395.975 2511.515 3396.020 ;
        RECT 2812.525 3395.975 2812.815 3396.020 ;
        RECT 1101.325 9.080 1101.615 9.125 ;
        RECT 918.320 8.940 1101.615 9.080 ;
        RECT 902.605 8.740 902.895 8.785 ;
        RECT 918.320 8.740 918.460 8.940 ;
        RECT 1101.325 8.895 1101.615 8.940 ;
        RECT 1103.625 9.080 1103.915 9.125 ;
        RECT 1157.905 9.080 1158.195 9.125 ;
        RECT 1103.625 8.940 1158.195 9.080 ;
        RECT 1103.625 8.895 1103.915 8.940 ;
        RECT 1157.905 8.895 1158.195 8.940 ;
        RECT 1163.500 8.940 1183.420 9.080 ;
        RECT 902.605 8.600 918.460 8.740 ;
        RECT 1162.045 8.740 1162.335 8.785 ;
        RECT 1163.500 8.740 1163.640 8.940 ;
        RECT 1162.045 8.600 1163.640 8.740 ;
        RECT 1183.280 8.740 1183.420 8.940 ;
        RECT 1195.625 8.740 1195.915 8.785 ;
        RECT 1183.280 8.600 1195.915 8.740 ;
        RECT 902.605 8.555 902.895 8.600 ;
        RECT 1162.045 8.555 1162.335 8.600 ;
        RECT 1195.625 8.555 1195.915 8.600 ;
        RECT 1648.710 7.380 1649.030 7.440 ;
        RECT 1781.650 7.380 1781.970 7.440 ;
        RECT 1648.710 7.240 1781.970 7.380 ;
        RECT 1648.710 7.180 1649.030 7.240 ;
        RECT 1781.650 7.180 1781.970 7.240 ;
        RECT 1266.450 6.360 1266.770 6.420 ;
        RECT 1270.130 6.360 1270.450 6.420 ;
        RECT 1266.450 6.220 1270.450 6.360 ;
        RECT 1266.450 6.160 1266.770 6.220 ;
        RECT 1270.130 6.160 1270.450 6.220 ;
        RECT 900.765 6.020 901.055 6.065 ;
        RECT 902.605 6.020 902.895 6.065 ;
        RECT 900.765 5.880 902.895 6.020 ;
        RECT 900.765 5.835 901.055 5.880 ;
        RECT 902.605 5.835 902.895 5.880 ;
        RECT 1196.070 5.340 1196.390 5.400 ;
        RECT 1195.875 5.200 1196.390 5.340 ;
        RECT 1196.070 5.140 1196.390 5.200 ;
        RECT 1209.870 4.800 1210.190 5.060 ;
        RECT 1639.050 5.000 1639.370 5.060 ;
        RECT 1647.790 5.000 1648.110 5.060 ;
        RECT 1639.050 4.860 1648.110 5.000 ;
        RECT 1639.050 4.800 1639.370 4.860 ;
        RECT 1647.790 4.800 1648.110 4.860 ;
        RECT 585.650 4.660 585.970 4.720 ;
        RECT 612.790 4.660 613.110 4.720 ;
        RECT 585.650 4.520 613.110 4.660 ;
        RECT 585.650 4.460 585.970 4.520 ;
        RECT 612.790 4.460 613.110 4.520 ;
        RECT 1209.960 4.320 1210.100 4.800 ;
        RECT 1209.040 4.180 1210.100 4.320 ;
        RECT 612.790 3.980 613.110 4.040 ;
        RECT 760.005 3.980 760.295 4.025 ;
        RECT 612.790 3.840 760.295 3.980 ;
        RECT 612.790 3.780 613.110 3.840 ;
        RECT 760.005 3.795 760.295 3.840 ;
        RECT 1196.070 3.980 1196.390 4.040 ;
        RECT 1209.040 3.980 1209.180 4.180 ;
        RECT 1196.070 3.840 1209.180 3.980 ;
        RECT 1196.070 3.780 1196.390 3.840 ;
        RECT 761.385 3.640 761.675 3.685 ;
        RECT 785.765 3.640 786.055 3.685 ;
        RECT 799.565 3.640 799.855 3.685 ;
        RECT 761.385 3.500 767.580 3.640 ;
        RECT 761.385 3.455 761.675 3.500 ;
        RECT 767.440 3.300 767.580 3.500 ;
        RECT 785.765 3.500 799.855 3.640 ;
        RECT 785.765 3.455 786.055 3.500 ;
        RECT 799.565 3.455 799.855 3.500 ;
        RECT 772.425 3.300 772.715 3.345 ;
        RECT 767.440 3.160 772.715 3.300 ;
        RECT 772.425 3.115 772.715 3.160 ;
        RECT 772.885 3.300 773.175 3.345 ;
        RECT 783.465 3.300 783.755 3.345 ;
        RECT 772.885 3.160 783.755 3.300 ;
        RECT 772.885 3.115 773.175 3.160 ;
        RECT 783.465 3.115 783.755 3.160 ;
        RECT 811.525 3.300 811.815 3.345 ;
        RECT 815.205 3.300 815.495 3.345 ;
        RECT 811.525 3.160 815.495 3.300 ;
        RECT 811.525 3.115 811.815 3.160 ;
        RECT 815.205 3.115 815.495 3.160 ;
        RECT 851.545 3.300 851.835 3.345 ;
        RECT 880.510 3.300 880.830 3.360 ;
        RECT 851.545 3.160 880.830 3.300 ;
        RECT 851.545 3.115 851.835 3.160 ;
        RECT 880.510 3.100 880.830 3.160 ;
        RECT 881.430 1.940 881.750 2.000 ;
        RECT 881.235 1.800 881.750 1.940 ;
        RECT 881.430 1.740 881.750 1.800 ;
      LAYER via ;
        RECT 2511.240 3401.740 2511.500 3402.000 ;
        RECT 2812.540 3401.400 2812.800 3401.660 ;
        RECT 1648.740 7.180 1649.000 7.440 ;
        RECT 1781.680 7.180 1781.940 7.440 ;
        RECT 1266.480 6.160 1266.740 6.420 ;
        RECT 1270.160 6.160 1270.420 6.420 ;
        RECT 1196.100 5.140 1196.360 5.400 ;
        RECT 1209.900 4.800 1210.160 5.060 ;
        RECT 1639.080 4.800 1639.340 5.060 ;
        RECT 1647.820 4.800 1648.080 5.060 ;
        RECT 585.680 4.460 585.940 4.720 ;
        RECT 612.820 4.460 613.080 4.720 ;
        RECT 612.820 3.780 613.080 4.040 ;
        RECT 1196.100 3.780 1196.360 4.040 ;
        RECT 880.540 3.100 880.800 3.360 ;
        RECT 881.460 1.740 881.720 2.000 ;
      LAYER met2 ;
        RECT 2510.710 3401.770 2510.990 3405.000 ;
        RECT 2511.240 3401.770 2511.500 3402.030 ;
        RECT 2510.710 3401.710 2511.500 3401.770 ;
        RECT 2510.710 3401.630 2511.440 3401.710 ;
        RECT 2510.710 3401.000 2510.990 3401.630 ;
        RECT 2812.530 3401.515 2812.810 3401.885 ;
        RECT 2812.540 3401.370 2812.800 3401.515 ;
        RECT 1210.350 7.635 1210.630 8.005 ;
        RECT 1210.420 5.680 1210.560 7.635 ;
        RECT 1648.740 7.210 1649.000 7.470 ;
        RECT 1263.780 7.070 1266.680 7.210 ;
        RECT 1263.780 6.645 1263.920 7.070 ;
        RECT 1263.710 6.275 1263.990 6.645 ;
        RECT 1266.540 6.450 1266.680 7.070 ;
        RECT 1647.880 7.150 1649.000 7.210 ;
        RECT 1781.680 7.150 1781.940 7.470 ;
        RECT 1647.880 7.070 1648.940 7.150 ;
        RECT 1266.480 6.130 1266.740 6.450 ;
        RECT 1270.150 6.275 1270.430 6.645 ;
        RECT 1270.160 6.130 1270.420 6.275 ;
        RECT 1209.960 5.540 1210.560 5.680 ;
        RECT 1196.100 5.110 1196.360 5.430 ;
        RECT 585.680 4.430 585.940 4.750 ;
        RECT 612.820 4.430 613.080 4.750 ;
        RECT 585.740 2.400 585.880 4.430 ;
        RECT 612.880 4.070 613.020 4.430 ;
        RECT 1196.160 4.070 1196.300 5.110 ;
        RECT 1209.960 5.090 1210.100 5.540 ;
        RECT 1209.900 4.770 1210.160 5.090 ;
        RECT 1635.390 4.915 1635.670 5.285 ;
        RECT 1647.880 5.090 1648.020 7.070 ;
        RECT 1635.460 4.490 1635.600 4.915 ;
        RECT 1639.080 4.770 1639.340 5.090 ;
        RECT 1647.820 4.770 1648.080 5.090 ;
        RECT 1639.140 4.490 1639.280 4.770 ;
        RECT 1635.460 4.350 1639.280 4.490 ;
        RECT 1781.740 4.490 1781.880 7.150 ;
        RECT 1782.130 4.490 1782.410 4.605 ;
        RECT 1781.740 4.350 1782.410 4.490 ;
        RECT 1782.130 4.235 1782.410 4.350 ;
        RECT 612.820 3.750 613.080 4.070 ;
        RECT 1196.100 3.750 1196.360 4.070 ;
        RECT 880.540 3.300 880.800 3.390 ;
        RECT 880.540 3.160 881.660 3.300 ;
        RECT 880.540 3.070 880.800 3.160 ;
        RECT 585.530 -4.800 586.090 2.400 ;
        RECT 881.520 2.030 881.660 3.160 ;
        RECT 881.460 1.710 881.720 2.030 ;
      LAYER via2 ;
        RECT 2812.530 3401.560 2812.810 3401.840 ;
        RECT 1210.350 7.680 1210.630 7.960 ;
        RECT 1263.710 6.320 1263.990 6.600 ;
        RECT 1270.150 6.320 1270.430 6.600 ;
        RECT 1635.390 4.960 1635.670 5.240 ;
        RECT 1782.130 4.280 1782.410 4.560 ;
      LAYER met3 ;
        RECT 2812.505 3401.850 2812.835 3401.865 ;
        RECT 2818.230 3401.850 2818.610 3401.860 ;
        RECT 2812.505 3401.550 2818.610 3401.850 ;
        RECT 2812.505 3401.535 2812.835 3401.550 ;
        RECT 2818.230 3401.540 2818.610 3401.550 ;
        RECT 1210.325 7.970 1210.655 7.985 ;
        RECT 1248.710 7.970 1249.090 7.980 ;
        RECT 1210.325 7.670 1249.090 7.970 ;
        RECT 1210.325 7.655 1210.655 7.670 ;
        RECT 1248.710 7.660 1249.090 7.670 ;
        RECT 1250.550 7.290 1250.930 7.300 ;
        RECT 1250.550 6.990 1257.330 7.290 ;
        RECT 1250.550 6.980 1250.930 6.990 ;
        RECT 1257.030 6.610 1257.330 6.990 ;
        RECT 1263.685 6.610 1264.015 6.625 ;
        RECT 1257.030 6.310 1264.015 6.610 ;
        RECT 1263.685 6.295 1264.015 6.310 ;
        RECT 1270.125 6.610 1270.455 6.625 ;
        RECT 1281.830 6.610 1282.210 6.620 ;
        RECT 1270.125 6.310 1282.210 6.610 ;
        RECT 1270.125 6.295 1270.455 6.310 ;
        RECT 1281.830 6.300 1282.210 6.310 ;
        RECT 1635.365 5.260 1635.695 5.265 ;
        RECT 1635.110 5.250 1635.695 5.260 ;
        RECT 1635.110 4.950 1635.920 5.250 ;
        RECT 1635.110 4.940 1635.695 4.950 ;
        RECT 1635.365 4.935 1635.695 4.940 ;
        RECT 1782.105 4.570 1782.435 4.585 ;
        RECT 1782.105 4.270 1789.090 4.570 ;
        RECT 1782.105 4.255 1782.435 4.270 ;
        RECT 1788.790 3.890 1789.090 4.270 ;
        RECT 1813.590 3.890 1813.970 3.900 ;
        RECT 1788.790 3.590 1813.970 3.890 ;
        RECT 1813.590 3.580 1813.970 3.590 ;
        RECT 2200.910 3.890 2201.290 3.900 ;
        RECT 2248.750 3.890 2249.130 3.900 ;
        RECT 2200.910 3.590 2249.130 3.890 ;
        RECT 2200.910 3.580 2201.290 3.590 ;
        RECT 2248.750 3.580 2249.130 3.590 ;
        RECT 2153.070 3.210 2153.450 3.220 ;
        RECT 2172.390 3.210 2172.770 3.220 ;
        RECT 2153.070 2.910 2172.770 3.210 ;
        RECT 2153.070 2.900 2153.450 2.910 ;
        RECT 2172.390 2.900 2172.770 2.910 ;
        RECT 2314.990 2.530 2315.370 2.540 ;
        RECT 2345.350 2.530 2345.730 2.540 ;
        RECT 2611.230 2.530 2611.610 2.540 ;
        RECT 2314.990 2.230 2345.730 2.530 ;
        RECT 2314.990 2.220 2315.370 2.230 ;
        RECT 2345.350 2.220 2345.730 2.230 ;
        RECT 2564.350 2.230 2611.610 2.530 ;
        RECT 2094.190 1.850 2094.570 1.860 ;
        RECT 2110.750 1.850 2111.130 1.860 ;
        RECT 2094.190 1.550 2111.130 1.850 ;
        RECT 2094.190 1.540 2094.570 1.550 ;
        RECT 2110.750 1.540 2111.130 1.550 ;
        RECT 2383.990 1.850 2384.370 1.860 ;
        RECT 2452.990 1.850 2453.370 1.860 ;
        RECT 2383.990 1.550 2453.370 1.850 ;
        RECT 2383.990 1.540 2384.370 1.550 ;
        RECT 2452.990 1.540 2453.370 1.550 ;
        RECT 2521.990 1.170 2522.370 1.180 ;
        RECT 2564.350 1.170 2564.650 2.230 ;
        RECT 2611.230 2.220 2611.610 2.230 ;
        RECT 2521.990 0.870 2564.650 1.170 ;
        RECT 2521.990 0.860 2522.370 0.870 ;
      LAYER via3 ;
        RECT 2818.260 3401.540 2818.580 3401.860 ;
        RECT 1248.740 7.660 1249.060 7.980 ;
        RECT 1250.580 6.980 1250.900 7.300 ;
        RECT 1281.860 6.300 1282.180 6.620 ;
        RECT 1635.140 4.940 1635.460 5.260 ;
        RECT 1813.620 3.580 1813.940 3.900 ;
        RECT 2200.940 3.580 2201.260 3.900 ;
        RECT 2248.780 3.580 2249.100 3.900 ;
        RECT 2153.100 2.900 2153.420 3.220 ;
        RECT 2172.420 2.900 2172.740 3.220 ;
        RECT 2315.020 2.220 2315.340 2.540 ;
        RECT 2345.380 2.220 2345.700 2.540 ;
        RECT 2094.220 1.540 2094.540 1.860 ;
        RECT 2110.780 1.540 2111.100 1.860 ;
        RECT 2384.020 1.540 2384.340 1.860 ;
        RECT 2453.020 1.540 2453.340 1.860 ;
        RECT 2522.020 0.860 2522.340 1.180 ;
        RECT 2611.260 2.220 2611.580 2.540 ;
      LAYER met4 ;
        RECT 2818.255 3401.535 2818.585 3401.865 ;
        RECT 1248.735 7.970 1249.065 7.985 ;
        RECT 1248.735 7.670 1250.890 7.970 ;
        RECT 1248.735 7.655 1249.065 7.670 ;
        RECT 1250.590 7.305 1250.890 7.670 ;
        RECT 1250.575 6.975 1250.905 7.305 ;
        RECT 1281.855 6.295 1282.185 6.625 ;
        RECT 1281.870 5.690 1282.170 6.295 ;
        RECT 2818.270 5.690 2818.570 3401.535 ;
        RECT 1281.430 4.510 1282.610 5.690 ;
        RECT 1325.590 5.250 1326.770 5.690 ;
        RECT 1334.790 5.250 1335.970 5.690 ;
        RECT 1325.590 4.950 1335.970 5.250 ;
        RECT 1325.590 4.510 1326.770 4.950 ;
        RECT 1334.790 4.510 1335.970 4.950 ;
        RECT 1634.710 4.510 1635.890 5.690 ;
        RECT 1813.630 4.950 1815.770 5.250 ;
        RECT 1813.630 3.905 1813.930 4.950 ;
        RECT 1813.615 3.575 1813.945 3.905 ;
        RECT 1815.470 2.290 1815.770 4.950 ;
        RECT 2072.630 4.510 2073.810 5.690 ;
        RECT 2093.790 4.510 2094.970 5.690 ;
        RECT 2200.510 4.510 2201.690 5.690 ;
        RECT 2314.590 4.510 2315.770 5.690 ;
        RECT 2610.830 4.510 2612.010 5.690 ;
        RECT 2817.830 4.510 2819.010 5.690 ;
        RECT 1815.030 1.110 1816.210 2.290 ;
        RECT 2069.870 1.850 2071.050 2.290 ;
        RECT 2073.070 1.850 2073.370 4.510 ;
        RECT 2094.230 1.865 2094.530 4.510 ;
        RECT 2200.950 3.905 2201.250 4.510 ;
        RECT 2200.935 3.575 2201.265 3.905 ;
        RECT 2248.775 3.575 2249.105 3.905 ;
        RECT 2153.095 2.895 2153.425 3.225 ;
        RECT 2172.415 2.895 2172.745 3.225 ;
        RECT 2153.110 2.290 2153.410 2.895 ;
        RECT 2172.430 2.290 2172.730 2.895 ;
        RECT 2248.790 2.290 2249.090 3.575 ;
        RECT 2315.030 2.545 2315.330 4.510 ;
        RECT 2611.270 2.545 2611.570 4.510 ;
        RECT 2069.870 1.550 2073.370 1.850 ;
        RECT 2069.870 1.110 2071.050 1.550 ;
        RECT 2094.215 1.535 2094.545 1.865 ;
        RECT 2110.350 1.110 2111.530 2.290 ;
        RECT 2152.670 1.110 2153.850 2.290 ;
        RECT 2171.990 1.110 2173.170 2.290 ;
        RECT 2248.350 1.110 2249.530 2.290 ;
        RECT 2315.015 2.215 2315.345 2.545 ;
        RECT 2345.375 2.290 2345.705 2.545 ;
        RECT 2344.950 1.110 2346.130 2.290 ;
        RECT 2383.590 1.110 2384.770 2.290 ;
        RECT 2452.590 1.110 2453.770 2.290 ;
        RECT 2521.590 1.110 2522.770 2.290 ;
        RECT 2611.255 2.215 2611.585 2.545 ;
        RECT 2522.015 0.855 2522.345 1.110 ;
      LAYER via4 ;
        RECT 2521.590 1.110 2522.770 2.290 ;
      LAYER met5 ;
        RECT 1281.220 4.300 1326.980 5.900 ;
        RECT 1334.580 4.300 1636.100 5.900 ;
        RECT 1920.620 4.300 1947.060 5.900 ;
        RECT 1920.620 2.500 1922.220 4.300 ;
        RECT 1814.820 0.900 1922.220 2.500 ;
        RECT 1945.460 2.500 1947.060 4.300 ;
        RECT 1994.220 4.300 2056.540 5.900 ;
        RECT 2072.420 4.300 2095.180 5.900 ;
        RECT 2171.780 4.300 2201.900 5.900 ;
        RECT 2251.820 4.300 2315.980 5.900 ;
        RECT 2610.620 4.300 2819.220 5.900 ;
        RECT 1994.220 2.500 1995.820 4.300 ;
        RECT 1945.460 0.900 1995.820 2.500 ;
        RECT 2054.940 2.500 2056.540 4.300 ;
        RECT 2054.940 0.900 2071.260 2.500 ;
        RECT 2110.140 0.900 2154.060 2.500 ;
        RECT 2171.780 0.900 2173.380 4.300 ;
        RECT 2251.820 3.180 2253.420 4.300 ;
        RECT 2249.060 2.500 2253.420 3.180 ;
        RECT 2248.140 1.580 2253.420 2.500 ;
        RECT 2248.140 0.900 2250.660 1.580 ;
        RECT 2344.740 0.900 2384.980 2.500 ;
        RECT 2452.380 0.900 2522.980 2.500 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2140.065 3399.745 2140.235 3401.955 ;
        RECT 2173.645 3399.065 2173.815 3399.915 ;
        RECT 2221.485 3399.065 2221.655 3400.595 ;
        RECT 2428.485 3399.575 2428.655 3400.595 ;
        RECT 2428.025 3399.405 2428.655 3399.575 ;
        RECT 2532.445 3399.405 2532.615 3400.595 ;
        RECT 2646.065 3399.405 2646.235 3400.595 ;
        RECT 2788.665 3400.425 2788.835 3402.295 ;
        RECT 7.045 52.445 7.215 61.795 ;
        RECT 8.885 61.625 9.055 99.875 ;
        RECT 25.905 6.885 26.075 7.735 ;
      LAYER mcon ;
        RECT 2788.665 3402.125 2788.835 3402.295 ;
        RECT 2140.065 3401.785 2140.235 3401.955 ;
        RECT 2221.485 3400.425 2221.655 3400.595 ;
        RECT 2173.645 3399.745 2173.815 3399.915 ;
        RECT 2428.485 3400.425 2428.655 3400.595 ;
        RECT 2532.445 3400.425 2532.615 3400.595 ;
        RECT 2646.065 3400.425 2646.235 3400.595 ;
        RECT 8.885 99.705 9.055 99.875 ;
        RECT 7.045 61.625 7.215 61.795 ;
        RECT 25.905 7.565 26.075 7.735 ;
      LAYER met1 ;
        RECT 2788.605 3402.280 2788.895 3402.325 ;
        RECT 2796.870 3402.280 2797.190 3402.340 ;
        RECT 2788.605 3402.140 2797.190 3402.280 ;
        RECT 2788.605 3402.095 2788.895 3402.140 ;
        RECT 2796.870 3402.080 2797.190 3402.140 ;
        RECT 2117.910 3401.940 2118.230 3402.000 ;
        RECT 2140.005 3401.940 2140.295 3401.985 ;
        RECT 2117.910 3401.800 2140.295 3401.940 ;
        RECT 2117.910 3401.740 2118.230 3401.800 ;
        RECT 2140.005 3401.755 2140.295 3401.800 ;
        RECT 2221.425 3400.580 2221.715 3400.625 ;
        RECT 2428.425 3400.580 2428.715 3400.625 ;
        RECT 2532.385 3400.580 2532.675 3400.625 ;
        RECT 2221.425 3400.440 2347.680 3400.580 ;
        RECT 2221.425 3400.395 2221.715 3400.440 ;
        RECT 2140.005 3399.900 2140.295 3399.945 ;
        RECT 2173.585 3399.900 2173.875 3399.945 ;
        RECT 2140.005 3399.760 2173.875 3399.900 ;
        RECT 2140.005 3399.715 2140.295 3399.760 ;
        RECT 2173.585 3399.715 2173.875 3399.760 ;
        RECT 2347.540 3399.560 2347.680 3400.440 ;
        RECT 2428.425 3400.440 2532.675 3400.580 ;
        RECT 2428.425 3400.395 2428.715 3400.440 ;
        RECT 2532.385 3400.395 2532.675 3400.440 ;
        RECT 2646.005 3400.580 2646.295 3400.625 ;
        RECT 2788.605 3400.580 2788.895 3400.625 ;
        RECT 2646.005 3400.440 2788.895 3400.580 ;
        RECT 2646.005 3400.395 2646.295 3400.440 ;
        RECT 2788.605 3400.395 2788.895 3400.440 ;
        RECT 2427.965 3399.560 2428.255 3399.605 ;
        RECT 2347.540 3399.420 2428.255 3399.560 ;
        RECT 2427.965 3399.375 2428.255 3399.420 ;
        RECT 2532.385 3399.560 2532.675 3399.605 ;
        RECT 2646.005 3399.560 2646.295 3399.605 ;
        RECT 2532.385 3399.420 2646.295 3399.560 ;
        RECT 2532.385 3399.375 2532.675 3399.420 ;
        RECT 2646.005 3399.375 2646.295 3399.420 ;
        RECT 2173.585 3399.220 2173.875 3399.265 ;
        RECT 2221.425 3399.220 2221.715 3399.265 ;
        RECT 2173.585 3399.080 2221.715 3399.220 ;
        RECT 2173.585 3399.035 2173.875 3399.080 ;
        RECT 2221.425 3399.035 2221.715 3399.080 ;
        RECT 6.970 99.860 7.290 99.920 ;
        RECT 8.825 99.860 9.115 99.905 ;
        RECT 6.970 99.720 9.115 99.860 ;
        RECT 6.970 99.660 7.290 99.720 ;
        RECT 8.825 99.675 9.115 99.720 ;
        RECT 6.985 61.780 7.275 61.825 ;
        RECT 8.825 61.780 9.115 61.825 ;
        RECT 6.985 61.640 9.115 61.780 ;
        RECT 6.985 61.595 7.275 61.640 ;
        RECT 8.825 61.595 9.115 61.640 ;
        RECT 4.210 52.600 4.530 52.660 ;
        RECT 6.985 52.600 7.275 52.645 ;
        RECT 4.210 52.460 7.275 52.600 ;
        RECT 4.210 52.400 4.530 52.460 ;
        RECT 6.985 52.415 7.275 52.460 ;
        RECT 91.610 8.400 91.930 8.460 ;
        RECT 51.680 8.260 91.930 8.400 ;
        RECT 25.845 7.720 26.135 7.765 ;
        RECT 51.680 7.720 51.820 8.260 ;
        RECT 91.610 8.200 91.930 8.260 ;
        RECT 25.845 7.580 51.820 7.720 ;
        RECT 25.845 7.535 26.135 7.580 ;
        RECT 4.670 7.040 4.990 7.100 ;
        RECT 25.845 7.040 26.135 7.085 ;
        RECT 4.670 6.900 26.135 7.040 ;
        RECT 4.670 6.840 4.990 6.900 ;
        RECT 25.845 6.855 26.135 6.900 ;
      LAYER via ;
        RECT 2796.900 3402.080 2797.160 3402.340 ;
        RECT 2117.940 3401.740 2118.200 3402.000 ;
        RECT 7.000 99.660 7.260 99.920 ;
        RECT 4.240 52.400 4.500 52.660 ;
        RECT 91.640 8.200 91.900 8.460 ;
        RECT 4.700 6.840 4.960 7.100 ;
      LAYER met2 ;
        RECT 2117.410 3401.770 2117.690 3405.000 ;
        RECT 2796.890 3402.875 2797.170 3403.245 ;
        RECT 2796.960 3402.370 2797.100 3402.875 ;
        RECT 2796.900 3402.050 2797.160 3402.370 ;
        RECT 2117.940 3401.770 2118.200 3402.030 ;
        RECT 2117.410 3401.710 2118.200 3401.770 ;
        RECT 2117.410 3401.630 2118.140 3401.710 ;
        RECT 2117.410 3401.000 2117.690 3401.630 ;
        RECT 6.990 100.115 7.270 100.485 ;
        RECT 7.060 99.950 7.200 100.115 ;
        RECT 7.000 99.630 7.260 99.950 ;
        RECT 4.240 52.370 4.500 52.690 ;
        RECT 4.300 50.730 4.440 52.370 ;
        RECT 4.300 50.590 4.900 50.730 ;
        RECT 4.760 7.130 4.900 50.590 ;
        RECT 91.640 8.170 91.900 8.490 ;
        RECT 4.700 6.810 4.960 7.130 ;
        RECT 91.700 2.400 91.840 8.170 ;
        RECT 91.490 -4.800 92.050 2.400 ;
      LAYER via2 ;
        RECT 2796.890 3402.920 2797.170 3403.200 ;
        RECT 6.990 100.160 7.270 100.440 ;
      LAYER met3 ;
        RECT 2796.865 3403.210 2797.195 3403.225 ;
        RECT 2809.950 3403.210 2810.330 3403.220 ;
        RECT 2796.865 3402.910 2810.330 3403.210 ;
        RECT 2796.865 3402.895 2797.195 3402.910 ;
        RECT 2809.950 3402.900 2810.330 3402.910 ;
        RECT 6.965 100.450 7.295 100.465 ;
        RECT 7.630 100.450 8.010 100.460 ;
        RECT 6.965 100.150 8.010 100.450 ;
        RECT 6.965 100.135 7.295 100.150 ;
        RECT 7.630 100.140 8.010 100.150 ;
      LAYER via3 ;
        RECT 2809.980 3402.900 2810.300 3403.220 ;
        RECT 7.660 100.140 7.980 100.460 ;
      LAYER met4 ;
        RECT 2809.975 3402.895 2810.305 3403.225 ;
        RECT 2809.990 175.690 2810.290 3402.895 ;
        RECT 2798.510 174.510 2799.690 175.690 ;
        RECT 2809.550 174.510 2810.730 175.690 ;
        RECT 2798.950 124.690 2799.250 174.510 ;
        RECT 7.230 123.510 8.410 124.690 ;
        RECT 2798.510 123.510 2799.690 124.690 ;
        RECT 7.670 100.465 7.970 123.510 ;
        RECT 7.655 100.135 7.985 100.465 ;
      LAYER met5 ;
        RECT 2798.300 174.300 2810.940 175.900 ;
        RECT 7.020 123.300 2799.900 124.900 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 5.665 1210.145 5.835 1307.555 ;
        RECT 7.505 1107.465 7.675 1190.935 ;
        RECT 3.365 110.245 3.535 167.875 ;
        RECT 3.825 60.265 3.995 92.395 ;
      LAYER mcon ;
        RECT 5.665 1307.385 5.835 1307.555 ;
        RECT 7.505 1190.765 7.675 1190.935 ;
        RECT 3.365 167.705 3.535 167.875 ;
        RECT 3.825 92.225 3.995 92.395 ;
      LAYER met1 ;
        RECT 5.590 1307.540 5.910 1307.600 ;
        RECT 5.395 1307.400 5.910 1307.540 ;
        RECT 5.590 1307.340 5.910 1307.400 ;
        RECT 5.605 1210.300 5.895 1210.345 ;
        RECT 8.810 1210.300 9.130 1210.360 ;
        RECT 5.605 1210.160 9.130 1210.300 ;
        RECT 5.605 1210.115 5.895 1210.160 ;
        RECT 8.810 1210.100 9.130 1210.160 ;
        RECT 7.445 1190.920 7.735 1190.965 ;
        RECT 8.810 1190.920 9.130 1190.980 ;
        RECT 7.445 1190.780 9.130 1190.920 ;
        RECT 7.445 1190.735 7.735 1190.780 ;
        RECT 8.810 1190.720 9.130 1190.780 ;
        RECT 6.970 1107.620 7.290 1107.680 ;
        RECT 7.445 1107.620 7.735 1107.665 ;
        RECT 6.970 1107.480 7.735 1107.620 ;
        RECT 6.970 1107.420 7.290 1107.480 ;
        RECT 7.445 1107.435 7.735 1107.480 ;
        RECT 6.510 977.740 6.830 977.800 ;
        RECT 7.430 977.740 7.750 977.800 ;
        RECT 6.510 977.600 7.750 977.740 ;
        RECT 6.510 977.540 6.830 977.600 ;
        RECT 7.430 977.540 7.750 977.600 ;
        RECT 0.990 872.340 1.310 872.400 ;
        RECT 7.430 872.340 7.750 872.400 ;
        RECT 0.990 872.200 7.750 872.340 ;
        RECT 0.990 872.140 1.310 872.200 ;
        RECT 7.430 872.140 7.750 872.200 ;
        RECT 0.990 692.820 1.310 692.880 ;
        RECT 3.290 692.820 3.610 692.880 ;
        RECT 0.990 692.680 3.610 692.820 ;
        RECT 0.990 692.620 1.310 692.680 ;
        RECT 3.290 692.620 3.610 692.680 ;
        RECT 3.290 167.860 3.610 167.920 ;
        RECT 3.095 167.720 3.610 167.860 ;
        RECT 3.290 167.660 3.610 167.720 ;
        RECT 3.305 110.400 3.595 110.445 ;
        RECT 9.730 110.400 10.050 110.460 ;
        RECT 3.305 110.260 10.050 110.400 ;
        RECT 3.305 110.215 3.595 110.260 ;
        RECT 9.730 110.200 10.050 110.260 ;
        RECT 3.765 92.380 4.055 92.425 ;
        RECT 9.730 92.380 10.050 92.440 ;
        RECT 3.765 92.240 10.050 92.380 ;
        RECT 3.765 92.195 4.055 92.240 ;
        RECT 9.730 92.180 10.050 92.240 ;
        RECT 3.765 60.420 4.055 60.465 ;
        RECT 6.510 60.420 6.830 60.480 ;
        RECT 3.765 60.280 6.830 60.420 ;
        RECT 3.765 60.235 4.055 60.280 ;
        RECT 6.510 60.220 6.830 60.280 ;
        RECT 568.630 3.980 568.950 4.040 ;
        RECT 602.670 3.980 602.990 4.040 ;
        RECT 568.630 3.840 602.990 3.980 ;
        RECT 568.630 3.780 568.950 3.840 ;
        RECT 602.670 3.780 602.990 3.840 ;
        RECT 513.430 3.640 513.750 3.700 ;
        RECT 539.190 3.640 539.510 3.700 ;
        RECT 513.430 3.500 539.510 3.640 ;
        RECT 513.430 3.440 513.750 3.500 ;
        RECT 539.190 3.440 539.510 3.500 ;
      LAYER via ;
        RECT 5.620 1307.340 5.880 1307.600 ;
        RECT 8.840 1210.100 9.100 1210.360 ;
        RECT 8.840 1190.720 9.100 1190.980 ;
        RECT 7.000 1107.420 7.260 1107.680 ;
        RECT 6.540 977.540 6.800 977.800 ;
        RECT 7.460 977.540 7.720 977.800 ;
        RECT 1.020 872.140 1.280 872.400 ;
        RECT 7.460 872.140 7.720 872.400 ;
        RECT 1.020 692.620 1.280 692.880 ;
        RECT 3.320 692.620 3.580 692.880 ;
        RECT 3.320 167.660 3.580 167.920 ;
        RECT 9.760 110.200 10.020 110.460 ;
        RECT 9.760 92.180 10.020 92.440 ;
        RECT 6.540 60.220 6.800 60.480 ;
        RECT 568.660 3.780 568.920 4.040 ;
        RECT 602.700 3.780 602.960 4.040 ;
        RECT 513.460 3.440 513.720 3.700 ;
        RECT 539.220 3.440 539.480 3.700 ;
      LAYER met2 ;
        RECT 5.610 3347.115 5.890 3347.485 ;
        RECT 5.680 1307.630 5.820 3347.115 ;
        RECT 5.620 1307.310 5.880 1307.630 ;
        RECT 8.840 1210.070 9.100 1210.390 ;
        RECT 8.900 1191.010 9.040 1210.070 ;
        RECT 8.840 1190.690 9.100 1191.010 ;
        RECT 7.000 1107.565 7.260 1107.710 ;
        RECT 6.990 1107.195 7.270 1107.565 ;
        RECT 6.530 1072.515 6.810 1072.885 ;
        RECT 6.600 977.830 6.740 1072.515 ;
        RECT 6.540 977.510 6.800 977.830 ;
        RECT 7.460 977.510 7.720 977.830 ;
        RECT 7.520 872.430 7.660 977.510 ;
        RECT 1.020 872.110 1.280 872.430 ;
        RECT 7.460 872.110 7.720 872.430 ;
        RECT 1.080 692.910 1.220 872.110 ;
        RECT 1.020 692.590 1.280 692.910 ;
        RECT 3.320 692.590 3.580 692.910 ;
        RECT 3.380 167.950 3.520 692.590 ;
        RECT 3.320 167.630 3.580 167.950 ;
        RECT 9.760 110.170 10.020 110.490 ;
        RECT 9.820 98.330 9.960 110.170 ;
        RECT 9.820 98.190 10.420 98.330 ;
        RECT 10.280 92.890 10.420 98.190 ;
        RECT 9.820 92.750 10.420 92.890 ;
        RECT 9.820 92.470 9.960 92.750 ;
        RECT 9.760 92.150 10.020 92.470 ;
        RECT 6.540 60.190 6.800 60.510 ;
        RECT 6.600 51.410 6.740 60.190 ;
        RECT 6.140 51.270 6.740 51.410 ;
        RECT 6.140 22.285 6.280 51.270 ;
        RECT 6.070 21.915 6.350 22.285 ;
        RECT 568.660 3.925 568.920 4.070 ;
        RECT 602.700 3.980 602.960 4.070 ;
        RECT 513.450 3.555 513.730 3.925 ;
        RECT 539.210 3.555 539.490 3.925 ;
        RECT 568.650 3.555 568.930 3.925 ;
        RECT 602.700 3.840 603.360 3.980 ;
        RECT 602.700 3.750 602.960 3.840 ;
        RECT 513.460 3.410 513.720 3.555 ;
        RECT 539.220 3.410 539.480 3.555 ;
        RECT 603.220 2.400 603.360 3.840 ;
        RECT 603.010 -4.800 603.570 2.400 ;
      LAYER via2 ;
        RECT 5.610 3347.160 5.890 3347.440 ;
        RECT 6.990 1107.240 7.270 1107.520 ;
        RECT 6.530 1072.560 6.810 1072.840 ;
        RECT 6.070 21.960 6.350 22.240 ;
        RECT 513.450 3.600 513.730 3.880 ;
        RECT 539.210 3.600 539.490 3.880 ;
        RECT 568.650 3.600 568.930 3.880 ;
      LAYER met3 ;
        RECT 5.000 3347.920 9.000 3348.520 ;
        RECT 5.830 3347.465 6.130 3347.920 ;
        RECT 5.585 3347.150 6.130 3347.465 ;
        RECT 5.585 3347.135 5.915 3347.150 ;
        RECT 6.965 1107.540 7.295 1107.545 ;
        RECT 6.710 1107.530 7.295 1107.540 ;
        RECT 6.510 1107.230 7.295 1107.530 ;
        RECT 6.710 1107.220 7.295 1107.230 ;
        RECT 6.965 1107.215 7.295 1107.220 ;
        RECT 6.505 1072.860 6.835 1072.865 ;
        RECT 6.505 1072.850 7.090 1072.860 ;
        RECT 6.280 1072.550 7.090 1072.850 ;
        RECT 6.505 1072.540 7.090 1072.550 ;
        RECT 6.505 1072.535 6.835 1072.540 ;
        RECT 6.045 22.250 6.375 22.265 ;
        RECT 6.710 22.250 7.090 22.260 ;
        RECT 6.045 21.950 7.090 22.250 ;
        RECT 6.045 21.935 6.375 21.950 ;
        RECT 6.710 21.940 7.090 21.950 ;
        RECT 458.660 9.030 459.920 9.255 ;
        RECT 458.660 9.020 459.040 9.030 ;
        RECT 459.620 8.650 459.920 9.030 ;
        RECT 463.950 8.650 464.330 8.660 ;
        RECT 459.620 8.350 464.330 8.650 ;
        RECT 463.950 8.340 464.330 8.350 ;
        RECT 511.790 3.890 512.170 3.900 ;
        RECT 513.425 3.890 513.755 3.905 ;
        RECT 511.790 3.590 513.755 3.890 ;
        RECT 511.790 3.580 512.170 3.590 ;
        RECT 513.425 3.575 513.755 3.590 ;
        RECT 539.185 3.890 539.515 3.905 ;
        RECT 557.790 3.890 558.170 3.900 ;
        RECT 539.185 3.590 558.170 3.890 ;
        RECT 539.185 3.575 539.515 3.590 ;
        RECT 557.790 3.580 558.170 3.590 ;
        RECT 558.710 3.890 559.090 3.900 ;
        RECT 568.625 3.890 568.955 3.905 ;
        RECT 558.710 3.590 568.955 3.890 ;
        RECT 558.710 3.580 559.090 3.590 ;
        RECT 568.625 3.575 568.955 3.590 ;
      LAYER via3 ;
        RECT 6.740 1107.220 7.060 1107.540 ;
        RECT 6.740 1072.540 7.060 1072.860 ;
        RECT 6.740 21.940 7.060 22.260 ;
        RECT 458.690 9.020 459.010 9.255 ;
        RECT 463.980 8.340 464.300 8.660 ;
        RECT 511.820 3.580 512.140 3.900 ;
        RECT 557.820 3.580 558.140 3.900 ;
        RECT 558.740 3.580 559.060 3.900 ;
      LAYER met4 ;
        RECT 6.735 1107.215 7.065 1107.545 ;
        RECT 6.750 1072.865 7.050 1107.215 ;
        RECT 6.735 1072.535 7.065 1072.865 ;
        RECT 6.310 21.510 7.490 22.690 ;
        RECT 381.670 14.710 382.850 15.890 ;
        RECT 411.110 14.710 412.290 15.890 ;
        RECT 457.110 14.710 458.290 15.890 ;
        RECT 382.110 12.050 382.410 14.710 ;
        RECT 382.110 11.750 383.330 12.050 ;
        RECT 383.030 7.970 383.330 11.750 ;
        RECT 411.550 9.330 411.850 14.710 ;
        RECT 408.790 9.030 411.850 9.330 ;
        RECT 457.550 9.330 457.850 14.710 ;
        RECT 458.685 9.330 459.015 9.345 ;
        RECT 457.550 9.030 459.015 9.330 ;
        RECT 408.790 8.650 409.090 9.030 ;
        RECT 458.685 9.015 459.015 9.030 ;
        RECT 384.870 8.350 409.090 8.650 ;
        RECT 384.870 7.970 385.170 8.350 ;
        RECT 463.975 8.335 464.305 8.665 ;
        RECT 383.030 7.670 385.170 7.970 ;
        RECT 463.990 7.970 464.290 8.335 ;
        RECT 463.990 7.670 472.570 7.970 ;
        RECT 472.270 3.890 472.570 7.670 ;
        RECT 511.815 3.890 512.145 3.905 ;
        RECT 472.270 3.590 512.145 3.890 ;
        RECT 511.815 3.575 512.145 3.590 ;
        RECT 557.815 3.890 558.145 3.905 ;
        RECT 558.735 3.890 559.065 3.905 ;
        RECT 557.815 3.590 559.065 3.890 ;
        RECT 557.815 3.575 558.145 3.590 ;
        RECT 558.735 3.575 559.065 3.590 ;
      LAYER met5 ;
        RECT 6.100 21.300 169.390 22.900 ;
        RECT 167.790 19.500 169.390 21.300 ;
        RECT 177.220 21.300 383.060 22.900 ;
        RECT 177.220 19.500 178.820 21.300 ;
        RECT 167.790 17.900 178.820 19.500 ;
        RECT 381.460 14.500 383.060 21.300 ;
        RECT 410.900 14.500 458.500 16.100 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 917.845 9.265 950.215 9.435 ;
        RECT 850.225 8.415 850.395 9.095 ;
        RECT 917.845 8.925 918.015 9.265 ;
        RECT 871.385 8.585 877.075 8.755 ;
        RECT 871.385 8.415 871.555 8.585 ;
        RECT 704.405 8.245 705.495 8.415 ;
        RECT 850.225 8.245 871.555 8.415 ;
        RECT 705.325 7.905 705.495 8.245 ;
        RECT 950.045 6.885 950.215 9.265 ;
        RECT 952.345 7.565 953.895 7.735 ;
        RECT 952.345 6.885 952.515 7.565 ;
        RECT 953.725 7.395 953.895 7.565 ;
        RECT 958.325 7.565 983.795 7.735 ;
        RECT 953.725 7.225 955.735 7.395 ;
        RECT 958.325 7.225 958.495 7.565 ;
        RECT 983.625 6.375 983.795 7.565 ;
        RECT 995.125 6.885 996.215 7.055 ;
        RECT 983.625 6.205 984.715 6.375 ;
        RECT 984.545 2.975 984.715 6.205 ;
        RECT 985.465 2.975 985.635 3.315 ;
        RECT 995.125 3.145 995.295 6.885 ;
        RECT 996.045 6.545 996.215 6.885 ;
        RECT 1192.925 6.545 1195.855 6.715 ;
        RECT 1122.085 3.485 1123.175 3.655 ;
        RECT 1122.085 3.145 1122.255 3.485 ;
        RECT 1123.005 3.315 1123.175 3.485 ;
        RECT 1125.765 3.315 1125.935 3.655 ;
        RECT 1123.005 3.145 1125.935 3.315 ;
        RECT 984.545 2.805 985.635 2.975 ;
        RECT 1157.965 2.975 1158.135 3.315 ;
        RECT 1160.265 2.975 1160.435 3.995 ;
        RECT 1164.405 3.825 1167.335 3.995 ;
        RECT 1192.005 3.655 1192.175 3.995 ;
        RECT 1192.925 3.655 1193.095 6.545 ;
        RECT 1195.685 6.205 1195.855 6.545 ;
        RECT 1192.005 3.485 1193.095 3.655 ;
        RECT 1157.965 2.805 1160.435 2.975 ;
      LAYER mcon ;
        RECT 850.225 8.925 850.395 9.095 ;
        RECT 876.905 8.585 877.075 8.755 ;
        RECT 955.565 7.225 955.735 7.395 ;
        RECT 1160.265 3.825 1160.435 3.995 ;
        RECT 1167.165 3.825 1167.335 3.995 ;
        RECT 1192.005 3.825 1192.175 3.995 ;
        RECT 985.465 3.145 985.635 3.315 ;
        RECT 1125.765 3.485 1125.935 3.655 ;
        RECT 1157.965 3.145 1158.135 3.315 ;
      LAYER met1 ;
        RECT 850.165 9.080 850.455 9.125 ;
        RECT 917.785 9.080 918.075 9.125 ;
        RECT 786.760 8.940 850.455 9.080 ;
        RECT 694.670 8.740 694.990 8.800 ;
        RECT 783.910 8.740 784.230 8.800 ;
        RECT 786.760 8.740 786.900 8.940 ;
        RECT 850.165 8.895 850.455 8.940 ;
        RECT 878.300 8.940 918.075 9.080 ;
        RECT 694.670 8.600 702.260 8.740 ;
        RECT 694.670 8.540 694.990 8.600 ;
        RECT 702.120 8.400 702.260 8.600 ;
        RECT 783.910 8.600 786.900 8.740 ;
        RECT 876.845 8.740 877.135 8.785 ;
        RECT 878.300 8.740 878.440 8.940 ;
        RECT 917.785 8.895 918.075 8.940 ;
        RECT 876.845 8.600 878.440 8.740 ;
        RECT 783.910 8.540 784.230 8.600 ;
        RECT 876.845 8.555 877.135 8.600 ;
        RECT 704.345 8.400 704.635 8.445 ;
        RECT 702.120 8.260 704.635 8.400 ;
        RECT 704.345 8.215 704.635 8.260 ;
        RECT 705.265 8.060 705.555 8.105 ;
        RECT 723.650 8.060 723.970 8.120 ;
        RECT 705.265 7.920 723.970 8.060 ;
        RECT 705.265 7.875 705.555 7.920 ;
        RECT 723.650 7.860 723.970 7.920 ;
        RECT 955.505 7.380 955.795 7.425 ;
        RECT 956.410 7.380 956.730 7.440 ;
        RECT 955.505 7.240 956.730 7.380 ;
        RECT 955.505 7.195 955.795 7.240 ;
        RECT 956.410 7.180 956.730 7.240 ;
        RECT 958.250 7.380 958.570 7.440 ;
        RECT 1401.230 7.380 1401.550 7.440 ;
        RECT 1408.590 7.380 1408.910 7.440 ;
        RECT 958.250 7.240 958.765 7.380 ;
        RECT 1401.230 7.240 1408.910 7.380 ;
        RECT 958.250 7.180 958.570 7.240 ;
        RECT 1401.230 7.180 1401.550 7.240 ;
        RECT 1408.590 7.180 1408.910 7.240 ;
        RECT 949.985 7.040 950.275 7.085 ;
        RECT 952.285 7.040 952.575 7.085 ;
        RECT 949.985 6.900 952.575 7.040 ;
        RECT 949.985 6.855 950.275 6.900 ;
        RECT 952.285 6.855 952.575 6.900 ;
        RECT 995.970 6.700 996.290 6.760 ;
        RECT 1014.830 6.700 1015.150 6.760 ;
        RECT 1055.770 6.700 1056.090 6.760 ;
        RECT 995.970 6.560 996.485 6.700 ;
        RECT 1014.830 6.560 1056.090 6.700 ;
        RECT 995.970 6.500 996.290 6.560 ;
        RECT 1014.830 6.500 1015.150 6.560 ;
        RECT 1055.770 6.500 1056.090 6.560 ;
        RECT 1195.610 6.360 1195.930 6.420 ;
        RECT 1195.610 6.220 1196.125 6.360 ;
        RECT 1195.610 6.160 1195.930 6.220 ;
        RECT 1069.110 3.980 1069.430 4.040 ;
        RECT 1096.710 3.980 1097.030 4.040 ;
        RECT 1069.110 3.840 1097.030 3.980 ;
        RECT 1069.110 3.780 1069.430 3.840 ;
        RECT 1096.710 3.780 1097.030 3.840 ;
        RECT 1160.205 3.980 1160.495 4.025 ;
        RECT 1164.345 3.980 1164.635 4.025 ;
        RECT 1160.205 3.840 1164.635 3.980 ;
        RECT 1160.205 3.795 1160.495 3.840 ;
        RECT 1164.345 3.795 1164.635 3.840 ;
        RECT 1167.105 3.980 1167.395 4.025 ;
        RECT 1191.945 3.980 1192.235 4.025 ;
        RECT 1167.105 3.840 1192.235 3.980 ;
        RECT 1167.105 3.795 1167.395 3.840 ;
        RECT 1191.945 3.795 1192.235 3.840 ;
        RECT 1125.705 3.640 1125.995 3.685 ;
        RECT 1125.705 3.500 1158.120 3.640 ;
        RECT 1125.705 3.455 1125.995 3.500 ;
        RECT 985.405 3.300 985.695 3.345 ;
        RECT 995.065 3.300 995.355 3.345 ;
        RECT 985.405 3.160 995.355 3.300 ;
        RECT 985.405 3.115 985.695 3.160 ;
        RECT 995.065 3.115 995.355 3.160 ;
        RECT 1122.010 3.300 1122.330 3.360 ;
        RECT 1157.980 3.345 1158.120 3.500 ;
        RECT 1122.010 3.160 1122.525 3.300 ;
        RECT 1122.010 3.100 1122.330 3.160 ;
        RECT 1157.905 3.115 1158.195 3.345 ;
        RECT 1208.490 2.280 1208.810 2.340 ;
        RECT 1236.090 2.280 1236.410 2.340 ;
        RECT 1208.490 2.140 1236.410 2.280 ;
        RECT 1208.490 2.080 1208.810 2.140 ;
        RECT 1236.090 2.080 1236.410 2.140 ;
      LAYER via ;
        RECT 694.700 8.540 694.960 8.800 ;
        RECT 783.940 8.540 784.200 8.800 ;
        RECT 723.680 7.860 723.940 8.120 ;
        RECT 956.440 7.180 956.700 7.440 ;
        RECT 958.280 7.180 958.540 7.440 ;
        RECT 1401.260 7.180 1401.520 7.440 ;
        RECT 1408.620 7.180 1408.880 7.440 ;
        RECT 996.000 6.500 996.260 6.760 ;
        RECT 1014.860 6.500 1015.120 6.760 ;
        RECT 1055.800 6.500 1056.060 6.760 ;
        RECT 1195.640 6.160 1195.900 6.420 ;
        RECT 1069.140 3.780 1069.400 4.040 ;
        RECT 1096.740 3.780 1097.000 4.040 ;
        RECT 1122.040 3.100 1122.300 3.360 ;
        RECT 1208.520 2.080 1208.780 2.340 ;
        RECT 1236.120 2.080 1236.380 2.340 ;
      LAYER met2 ;
        RECT 694.700 8.510 694.960 8.830 ;
        RECT 783.940 8.740 784.200 8.830 ;
        RECT 771.580 8.685 784.200 8.740 ;
        RECT 771.510 8.600 784.200 8.685 ;
        RECT 676.820 4.180 681.100 4.320 ;
        RECT 676.820 3.245 676.960 4.180 ;
        RECT 680.960 3.810 681.100 4.180 ;
        RECT 694.760 3.810 694.900 8.510 ;
        RECT 771.510 8.315 771.790 8.600 ;
        RECT 783.940 8.510 784.200 8.600 ;
        RECT 723.680 8.060 723.940 8.150 ;
        RECT 723.680 7.920 724.340 8.060 ;
        RECT 723.680 7.830 723.940 7.920 ;
        RECT 724.200 7.890 724.340 7.920 ;
        RECT 725.050 7.890 725.330 8.005 ;
        RECT 724.200 7.750 725.330 7.890 ;
        RECT 725.050 7.635 725.330 7.750 ;
        RECT 729.190 7.890 729.470 8.005 ;
        RECT 737.010 7.890 737.290 8.005 ;
        RECT 729.190 7.750 737.290 7.890 ;
        RECT 729.190 7.635 729.470 7.750 ;
        RECT 737.010 7.635 737.290 7.750 ;
        RECT 743.450 7.635 743.730 8.005 ;
        RECT 1251.360 7.750 1254.260 7.890 ;
        RECT 743.520 6.645 743.660 7.635 ;
        RECT 956.440 7.380 956.700 7.470 ;
        RECT 958.280 7.380 958.540 7.470 ;
        RECT 956.440 7.240 958.540 7.380 ;
        RECT 956.440 7.150 956.700 7.240 ;
        RECT 958.280 7.150 958.540 7.240 ;
        RECT 1244.850 7.210 1245.130 7.325 ;
        RECT 1195.700 7.070 1197.220 7.210 ;
        RECT 996.000 6.700 996.260 6.790 ;
        RECT 1014.860 6.700 1015.120 6.790 ;
        RECT 743.450 6.275 743.730 6.645 ;
        RECT 996.000 6.560 1015.120 6.700 ;
        RECT 996.000 6.470 996.260 6.560 ;
        RECT 1014.860 6.470 1015.120 6.560 ;
        RECT 1055.800 6.470 1056.060 6.790 ;
        RECT 1055.860 5.170 1056.000 6.470 ;
        RECT 1195.700 6.450 1195.840 7.070 ;
        RECT 1195.640 6.130 1195.900 6.450 ;
        RECT 1055.860 5.030 1069.340 5.170 ;
        RECT 1069.200 4.070 1069.340 5.030 ;
        RECT 680.960 3.670 694.900 3.810 ;
        RECT 1069.140 3.750 1069.400 4.070 ;
        RECT 1096.740 3.750 1097.000 4.070 ;
        RECT 1096.800 3.245 1096.940 3.750 ;
        RECT 1122.030 3.555 1122.310 3.925 ;
        RECT 1197.080 3.810 1197.220 7.070 ;
        RECT 1236.180 7.070 1245.130 7.210 ;
        RECT 1197.080 3.670 1207.800 3.810 ;
        RECT 1207.660 3.640 1207.800 3.670 ;
        RECT 1122.100 3.390 1122.240 3.555 ;
        RECT 1207.660 3.500 1208.720 3.640 ;
        RECT 621.090 2.875 621.370 3.245 ;
        RECT 676.750 2.875 677.030 3.245 ;
        RECT 1096.730 2.875 1097.010 3.245 ;
        RECT 1122.040 3.070 1122.300 3.390 ;
        RECT 621.160 2.400 621.300 2.875 ;
        RECT 620.950 -4.800 621.510 2.400 ;
        RECT 1208.580 2.370 1208.720 3.500 ;
        RECT 1236.180 2.370 1236.320 7.070 ;
        RECT 1244.850 6.955 1245.130 7.070 ;
        RECT 1249.910 7.210 1250.190 7.325 ;
        RECT 1251.360 7.210 1251.500 7.750 ;
        RECT 1249.910 7.070 1251.500 7.210 ;
        RECT 1254.120 7.210 1254.260 7.750 ;
        RECT 1257.730 7.210 1258.010 7.325 ;
        RECT 1254.120 7.070 1258.010 7.210 ;
        RECT 1401.260 7.150 1401.520 7.470 ;
        RECT 1408.620 7.325 1408.880 7.470 ;
        RECT 1249.910 6.955 1250.190 7.070 ;
        RECT 1257.730 6.955 1258.010 7.070 ;
        RECT 1401.320 6.020 1401.460 7.150 ;
        RECT 1408.610 6.955 1408.890 7.325 ;
        RECT 1426.550 7.210 1426.830 7.325 ;
        RECT 1429.770 7.210 1430.050 7.325 ;
        RECT 1426.550 7.070 1430.050 7.210 ;
        RECT 1426.550 6.955 1426.830 7.070 ;
        RECT 1429.770 6.955 1430.050 7.070 ;
        RECT 2782.170 7.210 2782.450 7.325 ;
        RECT 2783.490 7.210 2783.770 9.000 ;
        RECT 2782.170 7.070 2783.770 7.210 ;
        RECT 2782.170 6.955 2782.450 7.070 ;
        RECT 1401.320 5.880 1401.920 6.020 ;
        RECT 1266.470 4.915 1266.750 5.285 ;
        RECT 1266.540 3.300 1266.680 4.915 ;
        RECT 1291.770 3.810 1292.050 3.925 ;
        RECT 1280.340 3.670 1292.050 3.810 ;
        RECT 1280.340 3.300 1280.480 3.670 ;
        RECT 1291.770 3.555 1292.050 3.670 ;
        RECT 1401.250 3.810 1401.530 3.925 ;
        RECT 1401.780 3.810 1401.920 5.880 ;
        RECT 2783.490 5.000 2783.770 7.070 ;
        RECT 1401.250 3.670 1401.920 3.810 ;
        RECT 1401.250 3.555 1401.530 3.670 ;
        RECT 1266.540 3.160 1280.480 3.300 ;
        RECT 1208.520 2.050 1208.780 2.370 ;
        RECT 1236.120 2.050 1236.380 2.370 ;
      LAYER via2 ;
        RECT 771.510 8.360 771.790 8.640 ;
        RECT 725.050 7.680 725.330 7.960 ;
        RECT 729.190 7.680 729.470 7.960 ;
        RECT 737.010 7.680 737.290 7.960 ;
        RECT 743.450 7.680 743.730 7.960 ;
        RECT 743.450 6.320 743.730 6.600 ;
        RECT 1122.030 3.600 1122.310 3.880 ;
        RECT 621.090 2.920 621.370 3.200 ;
        RECT 676.750 2.920 677.030 3.200 ;
        RECT 1096.730 2.920 1097.010 3.200 ;
        RECT 1244.850 7.000 1245.130 7.280 ;
        RECT 1249.910 7.000 1250.190 7.280 ;
        RECT 1257.730 7.000 1258.010 7.280 ;
        RECT 1408.610 7.000 1408.890 7.280 ;
        RECT 1426.550 7.000 1426.830 7.280 ;
        RECT 1429.770 7.000 1430.050 7.280 ;
        RECT 2782.170 7.000 2782.450 7.280 ;
        RECT 1266.470 4.960 1266.750 5.240 ;
        RECT 1291.770 3.600 1292.050 3.880 ;
        RECT 1401.250 3.600 1401.530 3.880 ;
      LAYER met3 ;
        RECT 771.485 8.650 771.815 8.665 ;
        RECT 763.910 8.350 771.815 8.650 ;
        RECT 725.025 7.970 725.355 7.985 ;
        RECT 729.165 7.970 729.495 7.985 ;
        RECT 725.025 7.670 729.495 7.970 ;
        RECT 725.025 7.655 725.355 7.670 ;
        RECT 729.165 7.655 729.495 7.670 ;
        RECT 736.985 7.970 737.315 7.985 ;
        RECT 739.030 7.970 739.410 7.980 ;
        RECT 736.985 7.670 739.410 7.970 ;
        RECT 736.985 7.655 737.315 7.670 ;
        RECT 739.030 7.660 739.410 7.670 ;
        RECT 743.425 7.970 743.755 7.985 ;
        RECT 763.910 7.970 764.210 8.350 ;
        RECT 771.485 8.335 771.815 8.350 ;
        RECT 743.425 7.670 764.210 7.970 ;
        RECT 743.425 7.655 743.755 7.670 ;
        RECT 1244.825 7.290 1245.155 7.305 ;
        RECT 1249.885 7.290 1250.215 7.305 ;
        RECT 1244.825 6.990 1250.215 7.290 ;
        RECT 1244.825 6.975 1245.155 6.990 ;
        RECT 1249.885 6.975 1250.215 6.990 ;
        RECT 1257.705 7.290 1258.035 7.305 ;
        RECT 1408.585 7.290 1408.915 7.305 ;
        RECT 1426.525 7.290 1426.855 7.305 ;
        RECT 1257.705 6.990 1264.690 7.290 ;
        RECT 1257.705 6.975 1258.035 6.990 ;
        RECT 740.870 6.610 741.250 6.620 ;
        RECT 743.425 6.610 743.755 6.625 ;
        RECT 740.870 6.310 743.755 6.610 ;
        RECT 740.870 6.300 741.250 6.310 ;
        RECT 743.425 6.295 743.755 6.310 ;
        RECT 1264.390 5.250 1264.690 6.990 ;
        RECT 1408.585 6.990 1426.855 7.290 ;
        RECT 1408.585 6.975 1408.915 6.990 ;
        RECT 1426.525 6.975 1426.855 6.990 ;
        RECT 1429.745 7.290 1430.075 7.305 ;
        RECT 2782.145 7.290 2782.475 7.305 ;
        RECT 1429.745 6.990 2782.475 7.290 ;
        RECT 1429.745 6.975 1430.075 6.990 ;
        RECT 2782.145 6.975 2782.475 6.990 ;
        RECT 1266.445 5.250 1266.775 5.265 ;
        RECT 1264.390 4.950 1266.775 5.250 ;
        RECT 1266.445 4.935 1266.775 4.950 ;
        RECT 1122.005 3.890 1122.335 3.905 ;
        RECT 1106.150 3.590 1122.335 3.890 ;
        RECT 621.065 3.210 621.395 3.225 ;
        RECT 676.725 3.210 677.055 3.225 ;
        RECT 621.065 3.040 647.600 3.210 ;
        RECT 648.910 3.040 677.055 3.210 ;
        RECT 621.065 2.910 677.055 3.040 ;
        RECT 621.065 2.895 621.395 2.910 ;
        RECT 647.300 2.740 649.210 2.910 ;
        RECT 676.725 2.895 677.055 2.910 ;
        RECT 1096.705 3.210 1097.035 3.225 ;
        RECT 1106.150 3.210 1106.450 3.590 ;
        RECT 1122.005 3.575 1122.335 3.590 ;
        RECT 1291.745 3.890 1292.075 3.905 ;
        RECT 1301.150 3.890 1301.530 3.900 ;
        RECT 1291.745 3.590 1301.530 3.890 ;
        RECT 1291.745 3.575 1292.075 3.590 ;
        RECT 1301.150 3.580 1301.530 3.590 ;
        RECT 1400.510 3.890 1400.890 3.900 ;
        RECT 1401.225 3.890 1401.555 3.905 ;
        RECT 1400.510 3.590 1401.555 3.890 ;
        RECT 1400.510 3.580 1400.890 3.590 ;
        RECT 1401.225 3.575 1401.555 3.590 ;
        RECT 1096.705 2.910 1106.450 3.210 ;
        RECT 1096.705 2.895 1097.035 2.910 ;
      LAYER via3 ;
        RECT 739.060 7.660 739.380 7.980 ;
        RECT 740.900 6.300 741.220 6.620 ;
        RECT 1301.180 3.580 1301.500 3.900 ;
        RECT 1400.540 3.580 1400.860 3.900 ;
      LAYER met4 ;
        RECT 739.055 7.970 739.385 7.985 ;
        RECT 739.055 7.670 741.210 7.970 ;
        RECT 739.055 7.655 739.385 7.670 ;
        RECT 740.910 6.625 741.210 7.670 ;
        RECT 1315.910 6.990 1337.370 7.290 ;
        RECT 740.895 6.295 741.225 6.625 ;
        RECT 1301.190 4.950 1305.170 5.250 ;
        RECT 1301.190 3.905 1301.490 4.950 ;
        RECT 1301.175 3.575 1301.505 3.905 ;
        RECT 1304.870 1.850 1305.170 4.950 ;
        RECT 1315.910 1.850 1316.210 6.990 ;
        RECT 1331.110 3.210 1332.290 3.650 ;
        RECT 1337.070 3.210 1337.370 6.990 ;
        RECT 1400.535 3.575 1400.865 3.905 ;
        RECT 1331.110 2.910 1337.370 3.210 ;
        RECT 1331.110 2.470 1332.290 2.910 ;
        RECT 1400.550 2.290 1400.850 3.575 ;
        RECT 1304.870 1.550 1316.210 1.850 ;
        RECT 1400.110 1.110 1401.290 2.290 ;
      LAYER met5 ;
        RECT 1330.900 2.500 1332.500 3.860 ;
        RECT 1330.900 0.900 1401.500 2.500 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 9.345 2204.645 9.515 2245.955 ;
        RECT 9.345 1969.705 9.515 2028.015 ;
        RECT 8.885 1728.305 9.055 1791.375 ;
        RECT 8.885 1259.105 9.055 1307.555 ;
        RECT 8.425 1189.745 8.595 1211.335 ;
        RECT 9.345 880.855 9.515 898.195 ;
        RECT 8.885 880.685 9.515 880.855 ;
        RECT 8.885 797.725 9.055 880.685 ;
        RECT 2.905 707.965 3.075 714.935 ;
        RECT 9.345 362.185 9.515 465.715 ;
        RECT 7.505 80.325 7.675 108.035 ;
      LAYER mcon ;
        RECT 9.345 2245.785 9.515 2245.955 ;
        RECT 9.345 2027.845 9.515 2028.015 ;
        RECT 8.885 1791.205 9.055 1791.375 ;
        RECT 8.885 1307.385 9.055 1307.555 ;
        RECT 8.425 1211.165 8.595 1211.335 ;
        RECT 9.345 898.025 9.515 898.195 ;
        RECT 2.905 714.765 3.075 714.935 ;
        RECT 9.345 465.545 9.515 465.715 ;
        RECT 7.505 107.865 7.675 108.035 ;
      LAYER met1 ;
        RECT 6.970 2299.320 7.290 2299.380 ;
        RECT 9.270 2299.320 9.590 2299.380 ;
        RECT 6.970 2299.180 9.590 2299.320 ;
        RECT 6.970 2299.120 7.290 2299.180 ;
        RECT 9.270 2299.120 9.590 2299.180 ;
        RECT 9.270 2245.940 9.590 2246.000 ;
        RECT 9.075 2245.800 9.590 2245.940 ;
        RECT 9.270 2245.740 9.590 2245.800 ;
        RECT 9.270 2204.800 9.590 2204.860 ;
        RECT 9.075 2204.660 9.590 2204.800 ;
        RECT 9.270 2204.600 9.590 2204.660 ;
        RECT 9.270 2074.720 9.590 2074.980 ;
        RECT 9.360 2073.960 9.500 2074.720 ;
        RECT 9.270 2073.700 9.590 2073.960 ;
        RECT 9.270 2028.000 9.590 2028.060 ;
        RECT 9.075 2027.860 9.590 2028.000 ;
        RECT 9.270 2027.800 9.590 2027.860 ;
        RECT 9.270 1969.860 9.590 1969.920 ;
        RECT 9.075 1969.720 9.590 1969.860 ;
        RECT 9.270 1969.660 9.590 1969.720 ;
        RECT 8.825 1791.360 9.115 1791.405 ;
        RECT 9.270 1791.360 9.590 1791.420 ;
        RECT 8.825 1791.220 9.590 1791.360 ;
        RECT 8.825 1791.175 9.115 1791.220 ;
        RECT 9.270 1791.160 9.590 1791.220 ;
        RECT 8.825 1728.460 9.115 1728.505 ;
        RECT 9.270 1728.460 9.590 1728.520 ;
        RECT 8.825 1728.320 9.590 1728.460 ;
        RECT 8.825 1728.275 9.115 1728.320 ;
        RECT 9.270 1728.260 9.590 1728.320 ;
        RECT 8.825 1307.540 9.115 1307.585 ;
        RECT 9.270 1307.540 9.590 1307.600 ;
        RECT 8.825 1307.400 9.590 1307.540 ;
        RECT 8.825 1307.355 9.115 1307.400 ;
        RECT 9.270 1307.340 9.590 1307.400 ;
        RECT 8.825 1259.260 9.115 1259.305 ;
        RECT 9.270 1259.260 9.590 1259.320 ;
        RECT 8.825 1259.120 9.590 1259.260 ;
        RECT 8.825 1259.075 9.115 1259.120 ;
        RECT 9.270 1259.060 9.590 1259.120 ;
        RECT 8.365 1211.320 8.655 1211.365 ;
        RECT 9.270 1211.320 9.590 1211.380 ;
        RECT 8.365 1211.180 9.590 1211.320 ;
        RECT 8.365 1211.135 8.655 1211.180 ;
        RECT 9.270 1211.120 9.590 1211.180 ;
        RECT 8.365 1189.900 8.655 1189.945 ;
        RECT 9.270 1189.900 9.590 1189.960 ;
        RECT 8.365 1189.760 9.590 1189.900 ;
        RECT 8.365 1189.715 8.655 1189.760 ;
        RECT 9.270 1189.700 9.590 1189.760 ;
        RECT 9.270 898.180 9.590 898.240 ;
        RECT 9.075 898.040 9.590 898.180 ;
        RECT 9.270 897.980 9.590 898.040 ;
        RECT 5.130 797.880 5.450 797.940 ;
        RECT 8.825 797.880 9.115 797.925 ;
        RECT 5.130 797.740 9.115 797.880 ;
        RECT 5.130 797.680 5.450 797.740 ;
        RECT 8.825 797.695 9.115 797.740 ;
        RECT 2.845 714.920 3.135 714.965 ;
        RECT 5.130 714.920 5.450 714.980 ;
        RECT 2.845 714.780 5.450 714.920 ;
        RECT 2.845 714.735 3.135 714.780 ;
        RECT 5.130 714.720 5.450 714.780 ;
        RECT 2.830 708.120 3.150 708.180 ;
        RECT 2.635 707.980 3.150 708.120 ;
        RECT 2.830 707.920 3.150 707.980 ;
        RECT 2.830 465.700 3.150 465.760 ;
        RECT 9.285 465.700 9.575 465.745 ;
        RECT 2.830 465.560 9.575 465.700 ;
        RECT 2.830 465.500 3.150 465.560 ;
        RECT 9.285 465.515 9.575 465.560 ;
        RECT 9.270 362.340 9.590 362.400 ;
        RECT 9.075 362.200 9.590 362.340 ;
        RECT 9.270 362.140 9.590 362.200 ;
        RECT 6.510 192.680 6.830 192.740 ;
        RECT 9.270 192.680 9.590 192.740 ;
        RECT 6.510 192.540 9.590 192.680 ;
        RECT 6.510 192.480 6.830 192.540 ;
        RECT 9.270 192.480 9.590 192.540 ;
        RECT 6.510 108.020 6.830 108.080 ;
        RECT 7.445 108.020 7.735 108.065 ;
        RECT 6.510 107.880 7.735 108.020 ;
        RECT 6.510 107.820 6.830 107.880 ;
        RECT 7.445 107.835 7.735 107.880 ;
        RECT 7.445 80.480 7.735 80.525 ;
        RECT 9.270 80.480 9.590 80.540 ;
        RECT 7.445 80.340 9.590 80.480 ;
        RECT 7.445 80.295 7.735 80.340 ;
        RECT 9.270 80.280 9.590 80.340 ;
      LAYER via ;
        RECT 7.000 2299.120 7.260 2299.380 ;
        RECT 9.300 2299.120 9.560 2299.380 ;
        RECT 9.300 2245.740 9.560 2246.000 ;
        RECT 9.300 2204.600 9.560 2204.860 ;
        RECT 9.300 2074.720 9.560 2074.980 ;
        RECT 9.300 2073.700 9.560 2073.960 ;
        RECT 9.300 2027.800 9.560 2028.060 ;
        RECT 9.300 1969.660 9.560 1969.920 ;
        RECT 9.300 1791.160 9.560 1791.420 ;
        RECT 9.300 1728.260 9.560 1728.520 ;
        RECT 9.300 1307.340 9.560 1307.600 ;
        RECT 9.300 1259.060 9.560 1259.320 ;
        RECT 9.300 1211.120 9.560 1211.380 ;
        RECT 9.300 1189.700 9.560 1189.960 ;
        RECT 9.300 897.980 9.560 898.240 ;
        RECT 5.160 797.680 5.420 797.940 ;
        RECT 5.160 714.720 5.420 714.980 ;
        RECT 2.860 707.920 3.120 708.180 ;
        RECT 2.860 465.500 3.120 465.760 ;
        RECT 9.300 362.140 9.560 362.400 ;
        RECT 6.540 192.480 6.800 192.740 ;
        RECT 9.300 192.480 9.560 192.740 ;
        RECT 6.540 107.820 6.800 108.080 ;
        RECT 9.300 80.280 9.560 80.540 ;
      LAYER met2 ;
        RECT 6.990 2325.075 7.270 2325.445 ;
        RECT 7.060 2299.410 7.200 2325.075 ;
        RECT 7.000 2299.090 7.260 2299.410 ;
        RECT 9.300 2299.090 9.560 2299.410 ;
        RECT 9.360 2246.030 9.500 2299.090 ;
        RECT 9.300 2245.710 9.560 2246.030 ;
        RECT 9.300 2204.570 9.560 2204.890 ;
        RECT 9.360 2075.010 9.500 2204.570 ;
        RECT 9.300 2074.690 9.560 2075.010 ;
        RECT 9.300 2073.670 9.560 2073.990 ;
        RECT 9.360 2028.090 9.500 2073.670 ;
        RECT 9.300 2027.770 9.560 2028.090 ;
        RECT 9.300 1969.630 9.560 1969.950 ;
        RECT 9.360 1791.450 9.500 1969.630 ;
        RECT 9.300 1791.130 9.560 1791.450 ;
        RECT 9.300 1728.230 9.560 1728.550 ;
        RECT 9.360 1682.050 9.500 1728.230 ;
        RECT 8.900 1681.910 9.500 1682.050 ;
        RECT 8.900 1667.090 9.040 1681.910 ;
        RECT 8.900 1666.950 9.500 1667.090 ;
        RECT 9.360 1307.630 9.500 1666.950 ;
        RECT 9.300 1307.310 9.560 1307.630 ;
        RECT 9.300 1259.030 9.560 1259.350 ;
        RECT 9.360 1211.410 9.500 1259.030 ;
        RECT 9.300 1211.090 9.560 1211.410 ;
        RECT 9.300 1189.670 9.560 1189.990 ;
        RECT 9.360 898.270 9.500 1189.670 ;
        RECT 9.300 897.950 9.560 898.270 ;
        RECT 5.160 797.650 5.420 797.970 ;
        RECT 5.220 715.010 5.360 797.650 ;
        RECT 5.160 714.690 5.420 715.010 ;
        RECT 2.860 707.890 3.120 708.210 ;
        RECT 2.920 465.790 3.060 707.890 ;
        RECT 2.860 465.470 3.120 465.790 ;
        RECT 9.300 362.110 9.560 362.430 ;
        RECT 9.360 192.770 9.500 362.110 ;
        RECT 6.540 192.450 6.800 192.770 ;
        RECT 9.300 192.450 9.560 192.770 ;
        RECT 6.600 108.110 6.740 192.450 ;
        RECT 6.540 107.790 6.800 108.110 ;
        RECT 9.300 80.250 9.560 80.570 ;
        RECT 9.360 74.530 9.500 80.250 ;
        RECT 8.900 74.390 9.500 74.530 ;
        RECT 8.900 4.605 9.040 74.390 ;
        RECT 8.830 4.235 9.110 4.605 ;
        RECT 115.550 3.555 115.830 3.925 ;
        RECT 115.620 2.400 115.760 3.555 ;
        RECT 115.410 -4.800 115.970 2.400 ;
      LAYER via2 ;
        RECT 6.990 2325.120 7.270 2325.400 ;
        RECT 8.830 4.280 9.110 4.560 ;
        RECT 115.550 3.600 115.830 3.880 ;
      LAYER met3 ;
        RECT 5.000 2327.920 9.000 2328.520 ;
        RECT 6.750 2325.425 7.050 2327.920 ;
        RECT 6.750 2325.110 7.295 2325.425 ;
        RECT 6.965 2325.095 7.295 2325.110 ;
        RECT 8.805 4.570 9.135 4.585 ;
        RECT 8.805 4.270 52.130 4.570 ;
        RECT 8.805 4.255 9.135 4.270 ;
        RECT 51.830 3.890 52.130 4.270 ;
        RECT 115.525 3.890 115.855 3.905 ;
        RECT 51.830 3.590 115.855 3.890 ;
        RECT 115.525 3.575 115.855 3.590 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1314.825 15.385 1342.135 15.555 ;
        RECT 745.345 7.395 745.515 8.075 ;
        RECT 761.905 7.735 762.075 9.095 ;
        RECT 760.525 7.565 762.075 7.735 ;
        RECT 766.505 7.565 766.675 9.095 ;
        RECT 784.905 8.585 787.375 8.755 ;
        RECT 784.905 7.905 785.075 8.585 ;
        RECT 1312.065 7.735 1312.235 8.075 ;
        RECT 1314.825 7.735 1314.995 15.385 ;
        RECT 1312.065 7.565 1314.995 7.735 ;
        RECT 745.345 7.225 746.895 7.395 ;
        RECT 459.225 6.035 459.395 6.375 ;
        RECT 487.285 6.205 502.175 6.375 ;
        RECT 503.385 6.205 504.015 6.375 ;
        RECT 459.225 5.865 459.855 6.035 ;
        RECT 459.685 5.185 459.855 5.865 ;
        RECT 487.285 4.335 487.455 6.205 ;
        RECT 469.805 3.995 469.975 4.335 ;
        RECT 482.225 3.995 482.395 4.335 ;
        RECT 484.985 4.165 487.455 4.335 ;
        RECT 469.805 3.825 482.395 3.995 ;
        RECT 830.445 3.145 830.615 3.995 ;
      LAYER mcon ;
        RECT 1341.965 15.385 1342.135 15.555 ;
        RECT 761.905 8.925 762.075 9.095 ;
        RECT 745.345 7.905 745.515 8.075 ;
        RECT 766.505 8.925 766.675 9.095 ;
        RECT 787.205 8.585 787.375 8.755 ;
        RECT 1312.065 7.905 1312.235 8.075 ;
        RECT 746.725 7.225 746.895 7.395 ;
        RECT 459.225 6.205 459.395 6.375 ;
        RECT 502.005 6.205 502.175 6.375 ;
        RECT 503.845 6.205 504.015 6.375 ;
        RECT 469.805 4.165 469.975 4.335 ;
        RECT 482.225 4.165 482.395 4.335 ;
        RECT 830.445 3.825 830.615 3.995 ;
      LAYER met1 ;
        RECT 761.845 9.080 762.135 9.125 ;
        RECT 766.445 9.080 766.735 9.125 ;
        RECT 761.845 8.940 766.735 9.080 ;
        RECT 761.845 8.895 762.135 8.940 ;
        RECT 766.445 8.895 766.735 8.940 ;
        RECT 787.145 8.740 787.435 8.785 ;
        RECT 787.145 8.600 788.740 8.740 ;
        RECT 787.145 8.555 787.435 8.600 ;
        RECT 788.600 8.400 788.740 8.600 ;
        RECT 794.490 8.400 794.810 8.460 ;
        RECT 788.600 8.260 794.810 8.400 ;
        RECT 794.490 8.200 794.810 8.260 ;
        RECT 744.810 8.060 745.130 8.120 ;
        RECT 745.285 8.060 745.575 8.105 ;
        RECT 784.845 8.060 785.135 8.105 ;
        RECT 744.810 7.920 745.575 8.060 ;
        RECT 744.810 7.860 745.130 7.920 ;
        RECT 745.285 7.875 745.575 7.920 ;
        RECT 768.360 7.920 785.135 8.060 ;
        RECT 759.990 7.720 760.310 7.780 ;
        RECT 760.465 7.720 760.755 7.765 ;
        RECT 759.990 7.580 760.755 7.720 ;
        RECT 759.990 7.520 760.310 7.580 ;
        RECT 760.465 7.535 760.755 7.580 ;
        RECT 766.445 7.720 766.735 7.765 ;
        RECT 768.360 7.720 768.500 7.920 ;
        RECT 784.845 7.875 785.135 7.920 ;
        RECT 1311.530 8.060 1311.850 8.120 ;
        RECT 1312.005 8.060 1312.295 8.105 ;
        RECT 1311.530 7.920 1312.295 8.060 ;
        RECT 1311.530 7.860 1311.850 7.920 ;
        RECT 1312.005 7.875 1312.295 7.920 ;
        RECT 766.445 7.580 768.500 7.720 ;
        RECT 766.445 7.535 766.735 7.580 ;
        RECT 746.665 7.380 746.955 7.425 ;
        RECT 747.110 7.380 747.430 7.440 ;
        RECT 746.665 7.240 747.430 7.380 ;
        RECT 746.665 7.195 746.955 7.240 ;
        RECT 747.110 7.180 747.430 7.240 ;
        RECT 1024.030 7.380 1024.350 7.440 ;
        RECT 1056.690 7.380 1057.010 7.440 ;
        RECT 1024.030 7.240 1057.010 7.380 ;
        RECT 1024.030 7.180 1024.350 7.240 ;
        RECT 1056.690 7.180 1057.010 7.240 ;
        RECT 409.010 7.040 409.330 7.100 ;
        RECT 409.010 6.900 416.600 7.040 ;
        RECT 409.010 6.840 409.330 6.900 ;
        RECT 416.460 6.360 416.600 6.900 ;
        RECT 957.330 6.700 957.650 6.760 ;
        RECT 976.190 6.700 976.510 6.760 ;
        RECT 957.330 6.560 976.510 6.700 ;
        RECT 957.330 6.500 957.650 6.560 ;
        RECT 976.190 6.500 976.510 6.560 ;
        RECT 459.165 6.360 459.455 6.405 ;
        RECT 416.460 6.220 430.860 6.360 ;
        RECT 430.720 6.020 430.860 6.220 ;
        RECT 439.000 6.220 459.455 6.360 ;
        RECT 439.000 6.020 439.140 6.220 ;
        RECT 459.165 6.175 459.455 6.220 ;
        RECT 501.945 6.360 502.235 6.405 ;
        RECT 503.325 6.360 503.615 6.405 ;
        RECT 501.945 6.220 503.615 6.360 ;
        RECT 501.945 6.175 502.235 6.220 ;
        RECT 503.325 6.175 503.615 6.220 ;
        RECT 503.785 6.360 504.075 6.405 ;
        RECT 509.750 6.360 510.070 6.420 ;
        RECT 503.785 6.220 510.070 6.360 ;
        RECT 503.785 6.175 504.075 6.220 ;
        RECT 509.750 6.160 510.070 6.220 ;
        RECT 534.130 6.360 534.450 6.420 ;
        RECT 552.070 6.360 552.390 6.420 ;
        RECT 534.130 6.220 552.390 6.360 ;
        RECT 534.130 6.160 534.450 6.220 ;
        RECT 552.070 6.160 552.390 6.220 ;
        RECT 430.720 5.880 439.140 6.020 ;
        RECT 1190.090 6.020 1190.410 6.080 ;
        RECT 1191.930 6.020 1192.250 6.080 ;
        RECT 1190.090 5.880 1192.250 6.020 ;
        RECT 1190.090 5.820 1190.410 5.880 ;
        RECT 1191.930 5.820 1192.250 5.880 ;
        RECT 459.625 5.340 459.915 5.385 ;
        RECT 460.070 5.340 460.390 5.400 ;
        RECT 459.625 5.200 460.390 5.340 ;
        RECT 459.625 5.155 459.915 5.200 ;
        RECT 460.070 5.140 460.390 5.200 ;
        RECT 467.430 4.320 467.750 4.380 ;
        RECT 469.745 4.320 470.035 4.365 ;
        RECT 467.430 4.180 470.035 4.320 ;
        RECT 467.430 4.120 467.750 4.180 ;
        RECT 469.745 4.135 470.035 4.180 ;
        RECT 482.165 4.320 482.455 4.365 ;
        RECT 484.925 4.320 485.215 4.365 ;
        RECT 482.165 4.180 485.215 4.320 ;
        RECT 482.165 4.135 482.455 4.180 ;
        RECT 484.925 4.135 485.215 4.180 ;
        RECT 830.385 3.980 830.675 4.025 ;
        RECT 847.390 3.980 847.710 4.040 ;
        RECT 830.385 3.840 847.710 3.980 ;
        RECT 830.385 3.795 830.675 3.840 ;
        RECT 847.390 3.780 847.710 3.840 ;
        RECT 815.650 3.300 815.970 3.360 ;
        RECT 830.385 3.300 830.675 3.345 ;
        RECT 815.650 3.160 830.675 3.300 ;
        RECT 815.650 3.100 815.970 3.160 ;
        RECT 830.385 3.115 830.675 3.160 ;
        RECT 1208.950 2.620 1209.270 2.680 ;
        RECT 1232.870 2.620 1233.190 2.680 ;
        RECT 1208.950 2.480 1233.190 2.620 ;
        RECT 1208.950 2.420 1209.270 2.480 ;
        RECT 1232.870 2.420 1233.190 2.480 ;
      LAYER via ;
        RECT 794.520 8.200 794.780 8.460 ;
        RECT 744.840 7.860 745.100 8.120 ;
        RECT 760.020 7.520 760.280 7.780 ;
        RECT 1311.560 7.860 1311.820 8.120 ;
        RECT 747.140 7.180 747.400 7.440 ;
        RECT 1024.060 7.180 1024.320 7.440 ;
        RECT 1056.720 7.180 1056.980 7.440 ;
        RECT 409.040 6.840 409.300 7.100 ;
        RECT 957.360 6.500 957.620 6.760 ;
        RECT 976.220 6.500 976.480 6.760 ;
        RECT 509.780 6.160 510.040 6.420 ;
        RECT 534.160 6.160 534.420 6.420 ;
        RECT 552.100 6.160 552.360 6.420 ;
        RECT 1190.120 5.820 1190.380 6.080 ;
        RECT 1191.960 5.820 1192.220 6.080 ;
        RECT 460.100 5.140 460.360 5.400 ;
        RECT 467.460 4.120 467.720 4.380 ;
        RECT 847.420 3.780 847.680 4.040 ;
        RECT 815.680 3.100 815.940 3.360 ;
        RECT 1208.980 2.420 1209.240 2.680 ;
        RECT 1232.900 2.420 1233.160 2.680 ;
      LAYER met2 ;
        RECT 1341.920 15.340 1342.180 15.600 ;
        RECT 509.840 8.260 518.260 8.400 ;
        RECT 157.410 6.955 157.690 7.325 ;
        RECT 157.480 2.400 157.620 6.955 ;
        RECT 409.040 6.810 409.300 7.130 ;
        RECT 409.100 3.810 409.240 6.810 ;
        RECT 509.840 6.450 509.980 8.260 ;
        RECT 518.120 7.040 518.260 8.260 ;
        RECT 794.520 8.170 794.780 8.490 ;
        RECT 698.900 7.920 702.720 8.060 ;
        RECT 558.600 7.580 560.580 7.720 ;
        RECT 518.120 6.900 534.360 7.040 ;
        RECT 534.220 6.450 534.360 6.900 ;
        RECT 558.600 6.530 558.740 7.580 ;
        RECT 509.780 6.130 510.040 6.450 ;
        RECT 534.160 6.130 534.420 6.450 ;
        RECT 552.100 6.130 552.360 6.450 ;
        RECT 556.300 6.390 558.740 6.530 ;
        RECT 461.540 5.710 464.900 5.850 ;
        RECT 460.100 5.170 460.360 5.430 ;
        RECT 461.540 5.170 461.680 5.710 ;
        RECT 460.100 5.110 461.680 5.170 ;
        RECT 460.160 5.030 461.680 5.110 ;
        RECT 396.220 3.670 409.240 3.810 ;
        RECT 396.220 2.565 396.360 3.670 ;
        RECT 464.760 3.300 464.900 5.710 ;
        RECT 552.160 5.340 552.300 6.130 ;
        RECT 556.300 5.340 556.440 6.390 ;
        RECT 560.440 5.850 560.580 7.580 ;
        RECT 698.900 5.965 699.040 7.920 ;
        RECT 563.130 5.850 563.410 5.965 ;
        RECT 560.440 5.710 563.410 5.850 ;
        RECT 563.130 5.595 563.410 5.710 ;
        RECT 698.830 5.595 699.110 5.965 ;
        RECT 702.580 5.850 702.720 7.920 ;
        RECT 744.840 7.830 745.100 8.150 ;
        RECT 726.500 6.560 738.600 6.700 ;
        RECT 726.500 5.965 726.640 6.560 ;
        RECT 706.650 5.850 706.930 5.965 ;
        RECT 702.580 5.710 706.930 5.850 ;
        RECT 706.650 5.595 706.930 5.710 ;
        RECT 726.430 5.595 726.710 5.965 ;
        RECT 552.160 5.200 556.440 5.340 ;
        RECT 618.790 5.170 619.070 5.285 ;
        RECT 618.400 5.030 619.070 5.170 ;
        RECT 467.460 4.320 467.720 4.410 ;
        RECT 465.680 4.180 467.720 4.320 ;
        RECT 465.680 3.300 465.820 4.180 ;
        RECT 467.460 4.090 467.720 4.180 ;
        RECT 618.400 3.980 618.540 5.030 ;
        RECT 618.790 4.915 619.070 5.030 ;
        RECT 738.460 4.320 738.600 6.560 ;
        RECT 744.900 5.850 745.040 7.830 ;
        RECT 760.020 7.720 760.280 7.810 ;
        RECT 754.100 7.580 760.280 7.720 ;
        RECT 747.140 7.210 747.400 7.470 ;
        RECT 754.100 7.210 754.240 7.580 ;
        RECT 760.020 7.490 760.280 7.580 ;
        RECT 747.140 7.150 754.240 7.210 ;
        RECT 747.200 7.070 754.240 7.150 ;
        RECT 743.980 5.710 745.040 5.850 ;
        RECT 743.980 4.320 744.120 5.710 ;
        RECT 738.460 4.180 744.120 4.320 ;
        RECT 464.760 3.160 465.820 3.300 ;
        RECT 617.940 3.840 618.540 3.980 ;
        RECT 794.580 3.980 794.720 8.170 ;
        RECT 979.890 7.890 980.170 8.005 ;
        RECT 979.040 7.750 980.170 7.890 ;
        RECT 957.360 6.700 957.620 6.790 ;
        RECT 955.580 6.645 957.620 6.700 ;
        RECT 955.510 6.560 957.620 6.645 ;
        RECT 955.510 6.275 955.790 6.560 ;
        RECT 957.360 6.470 957.620 6.560 ;
        RECT 976.220 6.470 976.480 6.790 ;
        RECT 796.420 4.860 807.140 5.000 ;
        RECT 796.420 3.980 796.560 4.860 ;
        RECT 794.580 3.840 796.560 3.980 ;
        RECT 157.270 -4.800 157.830 2.400 ;
        RECT 396.150 2.195 396.430 2.565 ;
        RECT 617.940 1.770 618.080 3.840 ;
        RECT 619.710 3.130 619.990 3.245 ;
        RECT 619.320 2.990 619.990 3.130 ;
        RECT 619.320 1.770 619.460 2.990 ;
        RECT 619.710 2.875 619.990 2.990 ;
        RECT 807.000 1.885 807.140 4.860 ;
        RECT 976.280 4.490 976.420 6.470 ;
        RECT 979.040 4.490 979.180 7.750 ;
        RECT 979.890 7.635 980.170 7.750 ;
        RECT 1024.050 7.635 1024.330 8.005 ;
        RECT 1056.710 7.635 1056.990 8.005 ;
        RECT 1311.560 7.830 1311.820 8.150 ;
        RECT 1024.120 7.470 1024.260 7.635 ;
        RECT 1056.780 7.470 1056.920 7.635 ;
        RECT 1024.060 7.150 1024.320 7.470 ;
        RECT 1056.720 7.150 1056.980 7.470 ;
        RECT 1127.090 6.955 1127.370 7.325 ;
        RECT 1271.070 6.955 1271.350 7.325 ;
        RECT 1127.160 5.170 1127.300 6.955 ;
        RECT 1162.510 6.275 1162.790 6.645 ;
        RECT 1190.110 6.275 1190.390 6.645 ;
        RECT 1253.130 6.530 1253.410 6.645 ;
        RECT 1250.900 6.390 1253.410 6.530 ;
        RECT 1127.160 5.030 1158.120 5.170 ;
        RECT 847.480 4.350 849.920 4.490 ;
        RECT 976.280 4.350 979.180 4.490 ;
        RECT 1157.980 4.490 1158.120 5.030 ;
        RECT 1157.980 4.350 1159.040 4.490 ;
        RECT 847.480 4.070 847.620 4.350 ;
        RECT 847.420 3.750 847.680 4.070 ;
        RECT 815.680 3.070 815.940 3.390 ;
        RECT 849.780 3.130 849.920 4.350 ;
        RECT 1158.900 3.980 1159.040 4.350 ;
        RECT 1162.580 3.980 1162.720 6.275 ;
        RECT 1190.180 6.110 1190.320 6.275 ;
        RECT 1190.120 5.790 1190.380 6.110 ;
        RECT 1191.960 5.790 1192.220 6.110 ;
        RECT 1158.900 3.840 1162.720 3.980 ;
        RECT 1192.020 3.925 1192.160 5.790 ;
        RECT 1232.960 5.030 1234.480 5.170 ;
        RECT 1191.950 3.555 1192.230 3.925 ;
        RECT 1195.630 3.555 1195.910 3.925 ;
        RECT 850.170 3.130 850.450 3.245 ;
        RECT 815.740 1.885 815.880 3.070 ;
        RECT 849.780 2.990 850.450 3.130 ;
        RECT 1195.700 3.130 1195.840 3.555 ;
        RECT 1195.700 2.990 1207.800 3.130 ;
        RECT 850.170 2.875 850.450 2.990 ;
        RECT 617.940 1.630 619.460 1.770 ;
        RECT 806.930 1.515 807.210 1.885 ;
        RECT 815.670 1.515 815.950 1.885 ;
        RECT 1207.660 1.770 1207.800 2.990 ;
        RECT 1232.960 2.710 1233.100 5.030 ;
        RECT 1234.340 4.490 1234.480 5.030 ;
        RECT 1250.900 4.605 1251.040 6.390 ;
        RECT 1253.130 6.275 1253.410 6.390 ;
        RECT 1269.230 6.275 1269.510 6.645 ;
        RECT 1269.300 5.850 1269.440 6.275 ;
        RECT 1271.140 5.850 1271.280 6.955 ;
        RECT 1269.300 5.710 1271.280 5.850 ;
        RECT 1311.620 5.285 1311.760 7.830 ;
        RECT 1311.550 4.915 1311.830 5.285 ;
        RECT 1234.730 4.490 1235.010 4.605 ;
        RECT 1234.340 4.350 1235.010 4.490 ;
        RECT 1234.730 4.235 1235.010 4.350 ;
        RECT 1250.830 4.235 1251.110 4.605 ;
        RECT 1208.980 2.390 1209.240 2.710 ;
        RECT 1232.900 2.390 1233.160 2.710 ;
        RECT 1209.040 1.770 1209.180 2.390 ;
        RECT 1207.660 1.630 1209.180 1.770 ;
      LAYER via2 ;
        RECT 157.410 7.000 157.690 7.280 ;
        RECT 563.130 5.640 563.410 5.920 ;
        RECT 698.830 5.640 699.110 5.920 ;
        RECT 706.650 5.640 706.930 5.920 ;
        RECT 726.430 5.640 726.710 5.920 ;
        RECT 618.790 4.960 619.070 5.240 ;
        RECT 955.510 6.320 955.790 6.600 ;
        RECT 396.150 2.240 396.430 2.520 ;
        RECT 619.710 2.920 619.990 3.200 ;
        RECT 979.890 7.680 980.170 7.960 ;
        RECT 1024.050 7.680 1024.330 7.960 ;
        RECT 1056.710 7.680 1056.990 7.960 ;
        RECT 1127.090 7.000 1127.370 7.280 ;
        RECT 1271.070 7.000 1271.350 7.280 ;
        RECT 1162.510 6.320 1162.790 6.600 ;
        RECT 1190.110 6.320 1190.390 6.600 ;
        RECT 1191.950 3.600 1192.230 3.880 ;
        RECT 1195.630 3.600 1195.910 3.880 ;
        RECT 850.170 2.920 850.450 3.200 ;
        RECT 806.930 1.560 807.210 1.840 ;
        RECT 815.670 1.560 815.950 1.840 ;
        RECT 1253.130 6.320 1253.410 6.600 ;
        RECT 1269.230 6.320 1269.510 6.600 ;
        RECT 1311.550 4.960 1311.830 5.240 ;
        RECT 1234.730 4.280 1235.010 4.560 ;
        RECT 1250.830 4.280 1251.110 4.560 ;
      LAYER met3 ;
        RECT 1308.510 8.650 1308.890 8.660 ;
        RECT 1291.070 8.350 1308.890 8.650 ;
        RECT 979.865 7.970 980.195 7.985 ;
        RECT 1024.025 7.980 1024.355 7.985 ;
        RECT 985.590 7.970 985.970 7.980 ;
        RECT 979.865 7.670 985.970 7.970 ;
        RECT 979.865 7.655 980.195 7.670 ;
        RECT 985.590 7.660 985.970 7.670 ;
        RECT 1015.950 7.970 1016.330 7.980 ;
        RECT 1021.470 7.970 1021.850 7.980 ;
        RECT 1015.950 7.670 1021.850 7.970 ;
        RECT 1015.950 7.660 1016.330 7.670 ;
        RECT 1021.470 7.660 1021.850 7.670 ;
        RECT 1024.025 7.970 1024.610 7.980 ;
        RECT 1056.685 7.970 1057.015 7.985 ;
        RECT 1291.070 7.970 1291.370 8.350 ;
        RECT 1308.510 8.340 1308.890 8.350 ;
        RECT 1024.025 7.670 1024.810 7.970 ;
        RECT 1056.685 7.670 1123.700 7.970 ;
        RECT 1024.025 7.660 1024.610 7.670 ;
        RECT 1024.025 7.655 1024.355 7.660 ;
        RECT 1056.685 7.655 1057.015 7.670 ;
        RECT 157.385 7.290 157.715 7.305 ;
        RECT 195.310 7.290 195.690 7.300 ;
        RECT 157.385 6.990 195.690 7.290 ;
        RECT 1123.400 7.290 1123.700 7.670 ;
        RECT 1284.630 7.670 1291.370 7.970 ;
        RECT 1127.065 7.290 1127.395 7.305 ;
        RECT 1123.400 6.990 1127.395 7.290 ;
        RECT 157.385 6.975 157.715 6.990 ;
        RECT 195.310 6.980 195.690 6.990 ;
        RECT 1127.065 6.975 1127.395 6.990 ;
        RECT 1271.045 7.290 1271.375 7.305 ;
        RECT 1284.630 7.290 1284.930 7.670 ;
        RECT 1271.045 6.990 1284.930 7.290 ;
        RECT 1271.045 6.975 1271.375 6.990 ;
        RECT 948.790 6.610 949.170 6.620 ;
        RECT 955.485 6.610 955.815 6.625 ;
        RECT 948.790 6.310 955.815 6.610 ;
        RECT 948.790 6.300 949.170 6.310 ;
        RECT 955.485 6.295 955.815 6.310 ;
        RECT 1162.485 6.610 1162.815 6.625 ;
        RECT 1190.085 6.610 1190.415 6.625 ;
        RECT 1162.485 6.310 1190.415 6.610 ;
        RECT 1162.485 6.295 1162.815 6.310 ;
        RECT 1190.085 6.295 1190.415 6.310 ;
        RECT 1253.105 6.610 1253.435 6.625 ;
        RECT 1256.070 6.610 1256.450 6.620 ;
        RECT 1253.105 6.310 1256.450 6.610 ;
        RECT 1253.105 6.295 1253.435 6.310 ;
        RECT 1256.070 6.300 1256.450 6.310 ;
        RECT 1265.270 6.610 1265.650 6.620 ;
        RECT 1269.205 6.610 1269.535 6.625 ;
        RECT 1265.270 6.310 1269.535 6.610 ;
        RECT 1265.270 6.300 1265.650 6.310 ;
        RECT 1269.205 6.295 1269.535 6.310 ;
        RECT 563.105 5.930 563.435 5.945 ;
        RECT 601.030 5.930 601.410 5.940 ;
        RECT 563.105 5.630 601.410 5.930 ;
        RECT 563.105 5.615 563.435 5.630 ;
        RECT 601.030 5.620 601.410 5.630 ;
        RECT 697.860 5.930 698.240 5.940 ;
        RECT 698.805 5.930 699.135 5.945 ;
        RECT 697.860 5.630 699.135 5.930 ;
        RECT 697.860 5.620 698.240 5.630 ;
        RECT 698.805 5.615 699.135 5.630 ;
        RECT 706.625 5.930 706.955 5.945 ;
        RECT 726.405 5.930 726.735 5.945 ;
        RECT 706.625 5.630 726.735 5.930 ;
        RECT 706.625 5.615 706.955 5.630 ;
        RECT 726.405 5.615 726.735 5.630 ;
        RECT 618.765 5.260 619.095 5.265 ;
        RECT 1311.525 5.260 1311.855 5.265 ;
        RECT 618.510 5.250 619.095 5.260 ;
        RECT 1311.270 5.250 1311.855 5.260 ;
        RECT 618.510 4.950 619.320 5.250 ;
        RECT 1311.070 4.950 1311.855 5.250 ;
        RECT 618.510 4.940 619.095 4.950 ;
        RECT 1311.270 4.940 1311.855 4.950 ;
        RECT 618.765 4.935 619.095 4.940 ;
        RECT 1311.525 4.935 1311.855 4.940 ;
        RECT 1234.705 4.570 1235.035 4.585 ;
        RECT 1250.805 4.570 1251.135 4.585 ;
        RECT 1234.705 4.270 1251.135 4.570 ;
        RECT 1234.705 4.255 1235.035 4.270 ;
        RECT 1250.805 4.255 1251.135 4.270 ;
        RECT 652.550 3.890 652.930 3.900 ;
        RECT 674.630 3.890 675.010 3.900 ;
        RECT 652.550 3.590 675.010 3.890 ;
        RECT 652.550 3.580 652.930 3.590 ;
        RECT 674.630 3.580 675.010 3.590 ;
        RECT 681.070 3.890 681.450 3.900 ;
        RECT 688.430 3.890 688.810 3.900 ;
        RECT 681.070 3.590 688.810 3.890 ;
        RECT 681.070 3.580 681.450 3.590 ;
        RECT 688.430 3.580 688.810 3.590 ;
        RECT 1191.925 3.890 1192.255 3.905 ;
        RECT 1195.605 3.890 1195.935 3.905 ;
        RECT 1191.925 3.590 1195.935 3.890 ;
        RECT 1191.925 3.575 1192.255 3.590 ;
        RECT 1195.605 3.575 1195.935 3.590 ;
        RECT 619.685 3.210 620.015 3.225 ;
        RECT 620.350 3.210 620.730 3.220 ;
        RECT 619.685 2.910 620.730 3.210 ;
        RECT 619.685 2.895 620.015 2.910 ;
        RECT 620.350 2.900 620.730 2.910 ;
        RECT 850.145 3.210 850.475 3.225 ;
        RECT 875.190 3.210 875.570 3.220 ;
        RECT 850.145 2.910 875.570 3.210 ;
        RECT 850.145 2.895 850.475 2.910 ;
        RECT 875.190 2.900 875.570 2.910 ;
        RECT 393.110 2.530 393.490 2.540 ;
        RECT 396.125 2.530 396.455 2.545 ;
        RECT 393.110 2.230 396.455 2.530 ;
        RECT 393.110 2.220 393.490 2.230 ;
        RECT 396.125 2.215 396.455 2.230 ;
        RECT 806.905 1.850 807.235 1.865 ;
        RECT 815.645 1.850 815.975 1.865 ;
        RECT 806.905 1.550 815.975 1.850 ;
        RECT 806.905 1.535 807.235 1.550 ;
        RECT 815.645 1.535 815.975 1.550 ;
      LAYER via3 ;
        RECT 985.620 7.660 985.940 7.980 ;
        RECT 1015.980 7.660 1016.300 7.980 ;
        RECT 1021.500 7.660 1021.820 7.980 ;
        RECT 1024.260 7.660 1024.580 7.980 ;
        RECT 1308.540 8.340 1308.860 8.660 ;
        RECT 195.340 6.980 195.660 7.300 ;
        RECT 948.820 6.300 949.140 6.620 ;
        RECT 1256.100 6.300 1256.420 6.620 ;
        RECT 1265.300 6.300 1265.620 6.620 ;
        RECT 601.060 5.620 601.380 5.940 ;
        RECT 697.890 5.620 698.210 5.940 ;
        RECT 618.540 4.940 618.860 5.260 ;
        RECT 1311.300 4.940 1311.620 5.260 ;
        RECT 652.580 3.580 652.900 3.900 ;
        RECT 674.660 3.580 674.980 3.900 ;
        RECT 681.100 3.580 681.420 3.900 ;
        RECT 688.460 3.580 688.780 3.900 ;
        RECT 620.380 2.900 620.700 3.220 ;
        RECT 875.220 2.900 875.540 3.220 ;
        RECT 393.140 2.220 393.460 2.540 ;
      LAYER met4 ;
        RECT 985.630 8.350 1003.410 8.650 ;
        RECT 985.630 7.985 985.930 8.350 ;
        RECT 985.615 7.655 985.945 7.985 ;
        RECT 195.335 6.975 195.665 7.305 ;
        RECT 1003.110 7.290 1003.410 8.350 ;
        RECT 1308.535 8.335 1308.865 8.665 ;
        RECT 1015.975 7.655 1016.305 7.985 ;
        RECT 1021.495 7.655 1021.825 7.985 ;
        RECT 1024.255 7.655 1024.585 7.985 ;
        RECT 1015.990 7.290 1016.290 7.655 ;
        RECT 1003.110 6.990 1016.290 7.290 ;
        RECT 1021.510 7.290 1021.810 7.655 ;
        RECT 1024.270 7.290 1024.570 7.655 ;
        RECT 1021.510 6.990 1024.570 7.290 ;
        RECT 1308.550 7.290 1308.850 8.335 ;
        RECT 1308.550 6.990 1315.290 7.290 ;
        RECT 195.350 5.690 195.650 6.975 ;
        RECT 948.815 6.610 949.145 6.625 ;
        RECT 919.390 6.310 949.145 6.610 ;
        RECT 601.055 5.930 601.385 5.945 ;
        RECT 697.885 5.930 698.215 5.945 ;
        RECT 919.390 5.930 919.690 6.310 ;
        RECT 948.815 6.295 949.145 6.310 ;
        RECT 1256.095 6.610 1256.425 6.625 ;
        RECT 1265.295 6.610 1265.625 6.625 ;
        RECT 1256.095 6.310 1265.625 6.610 ;
        RECT 1256.095 6.295 1256.425 6.310 ;
        RECT 1265.295 6.295 1265.625 6.310 ;
        RECT 194.910 4.510 196.090 5.690 ;
        RECT 601.055 5.630 618.850 5.930 ;
        RECT 601.055 5.615 601.385 5.630 ;
        RECT 618.550 5.265 618.850 5.630 ;
        RECT 697.670 5.615 698.215 5.930 ;
        RECT 905.590 5.630 919.690 5.930 ;
        RECT 618.535 4.935 618.865 5.265 ;
        RECT 697.670 5.250 697.970 5.615 ;
        RECT 905.590 5.250 905.890 5.630 ;
        RECT 689.390 4.950 697.970 5.250 ;
        RECT 875.230 4.950 877.370 5.250 ;
        RECT 621.540 3.590 622.530 3.890 ;
        RECT 620.375 3.210 620.705 3.225 ;
        RECT 621.540 3.210 621.840 3.590 ;
        RECT 367.390 2.910 381.490 3.210 ;
        RECT 367.390 2.290 367.690 2.910 ;
        RECT 381.190 2.530 381.490 2.910 ;
        RECT 620.375 2.910 621.840 3.210 ;
        RECT 622.230 3.210 622.530 3.590 ;
        RECT 652.575 3.575 652.905 3.905 ;
        RECT 674.655 3.575 674.985 3.905 ;
        RECT 681.095 3.890 681.425 3.905 ;
        RECT 678.350 3.590 681.425 3.890 ;
        RECT 652.590 3.210 652.890 3.575 ;
        RECT 622.230 2.910 652.890 3.210 ;
        RECT 674.670 3.210 674.970 3.575 ;
        RECT 674.670 2.910 675.200 3.210 ;
        RECT 620.375 2.895 620.705 2.910 ;
        RECT 393.135 2.530 393.465 2.545 ;
        RECT 366.950 1.110 368.130 2.290 ;
        RECT 381.190 2.230 393.465 2.530 ;
        RECT 674.900 2.530 675.200 2.910 ;
        RECT 678.350 2.530 678.650 3.590 ;
        RECT 681.095 3.575 681.425 3.590 ;
        RECT 688.455 3.890 688.785 3.905 ;
        RECT 689.390 3.890 689.690 4.950 ;
        RECT 688.455 3.590 689.690 3.890 ;
        RECT 688.455 3.575 688.785 3.590 ;
        RECT 875.230 3.225 875.530 4.950 ;
        RECT 877.070 4.570 877.370 4.950 ;
        RECT 882.590 4.950 905.890 5.250 ;
        RECT 1311.295 5.250 1311.625 5.265 ;
        RECT 1314.990 5.250 1315.290 6.990 ;
        RECT 1311.295 4.950 1315.290 5.250 ;
        RECT 882.590 4.570 882.890 4.950 ;
        RECT 1311.295 4.935 1311.625 4.950 ;
        RECT 877.070 4.270 882.890 4.570 ;
        RECT 875.215 2.895 875.545 3.225 ;
        RECT 674.900 2.230 678.650 2.530 ;
        RECT 393.135 2.215 393.465 2.230 ;
      LAYER met5 ;
        RECT 194.700 4.300 231.260 5.900 ;
        RECT 229.660 2.500 231.260 4.300 ;
        RECT 229.660 0.900 368.340 2.500 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 5.205 705.585 5.375 751.315 ;
        RECT 7.505 751.145 7.675 781.915 ;
        RECT 7.505 631.125 7.675 673.115 ;
        RECT 27.745 8.245 27.915 9.095 ;
        RECT 50.745 7.395 50.915 8.415 ;
        RECT 50.745 7.225 53.215 7.395 ;
        RECT 64.545 6.715 64.715 7.395 ;
        RECT 64.545 6.545 66.095 6.715 ;
      LAYER mcon ;
        RECT 7.505 781.745 7.675 781.915 ;
        RECT 5.205 751.145 5.375 751.315 ;
        RECT 7.505 672.945 7.675 673.115 ;
        RECT 27.745 8.925 27.915 9.095 ;
        RECT 50.745 8.245 50.915 8.415 ;
        RECT 53.045 7.225 53.215 7.395 ;
        RECT 64.545 7.225 64.715 7.395 ;
        RECT 65.925 6.545 66.095 6.715 ;
      LAYER met1 ;
        RECT 7.445 781.900 7.735 781.945 ;
        RECT 7.890 781.900 8.210 781.960 ;
        RECT 7.445 781.760 8.210 781.900 ;
        RECT 7.445 781.715 7.735 781.760 ;
        RECT 7.890 781.700 8.210 781.760 ;
        RECT 5.145 751.300 5.435 751.345 ;
        RECT 7.445 751.300 7.735 751.345 ;
        RECT 5.145 751.160 7.735 751.300 ;
        RECT 5.145 751.115 5.435 751.160 ;
        RECT 7.445 751.115 7.735 751.160 ;
        RECT 5.145 705.740 5.435 705.785 ;
        RECT 9.270 705.740 9.590 705.800 ;
        RECT 5.145 705.600 9.590 705.740 ;
        RECT 5.145 705.555 5.435 705.600 ;
        RECT 9.270 705.540 9.590 705.600 ;
        RECT 7.445 673.100 7.735 673.145 ;
        RECT 9.270 673.100 9.590 673.160 ;
        RECT 7.445 672.960 9.590 673.100 ;
        RECT 7.445 672.915 7.735 672.960 ;
        RECT 9.270 672.900 9.590 672.960 ;
        RECT 7.445 631.280 7.735 631.325 ;
        RECT 7.890 631.280 8.210 631.340 ;
        RECT 7.445 631.140 8.210 631.280 ;
        RECT 7.445 631.095 7.735 631.140 ;
        RECT 7.890 631.080 8.210 631.140 ;
        RECT 7.430 9.080 7.750 9.140 ;
        RECT 27.685 9.080 27.975 9.125 ;
        RECT 7.430 8.940 27.975 9.080 ;
        RECT 7.430 8.880 7.750 8.940 ;
        RECT 27.685 8.895 27.975 8.940 ;
        RECT 27.685 8.400 27.975 8.445 ;
        RECT 50.685 8.400 50.975 8.445 ;
        RECT 27.685 8.260 50.975 8.400 ;
        RECT 27.685 8.215 27.975 8.260 ;
        RECT 50.685 8.215 50.975 8.260 ;
        RECT 52.985 7.380 53.275 7.425 ;
        RECT 64.485 7.380 64.775 7.425 ;
        RECT 52.985 7.240 64.775 7.380 ;
        RECT 52.985 7.195 53.275 7.240 ;
        RECT 64.485 7.195 64.775 7.240 ;
        RECT 65.865 6.700 66.155 6.745 ;
        RECT 72.290 6.700 72.610 6.760 ;
        RECT 65.865 6.560 72.610 6.700 ;
        RECT 65.865 6.515 66.155 6.560 ;
        RECT 72.290 6.500 72.610 6.560 ;
      LAYER via ;
        RECT 7.920 781.700 8.180 781.960 ;
        RECT 9.300 705.540 9.560 705.800 ;
        RECT 9.300 672.900 9.560 673.160 ;
        RECT 7.920 631.080 8.180 631.340 ;
        RECT 7.460 8.880 7.720 9.140 ;
        RECT 72.320 6.500 72.580 6.760 ;
      LAYER met2 ;
        RECT 7.910 2438.635 8.190 2439.005 ;
        RECT 7.980 781.990 8.120 2438.635 ;
        RECT 7.920 781.670 8.180 781.990 ;
        RECT 9.300 705.510 9.560 705.830 ;
        RECT 9.360 673.190 9.500 705.510 ;
        RECT 9.300 672.870 9.560 673.190 ;
        RECT 7.920 631.050 8.180 631.370 ;
        RECT 7.980 52.090 8.120 631.050 ;
        RECT 7.520 51.950 8.120 52.090 ;
        RECT 7.520 9.170 7.660 51.950 ;
        RECT 7.460 8.850 7.720 9.170 ;
        RECT 72.320 6.470 72.580 6.790 ;
        RECT 72.380 4.605 72.520 6.470 ;
        RECT 72.310 4.235 72.590 4.605 ;
        RECT 174.890 4.235 175.170 4.605 ;
        RECT 174.960 2.400 175.100 4.235 ;
        RECT 174.750 -4.800 175.310 2.400 ;
      LAYER via2 ;
        RECT 7.910 2438.680 8.190 2438.960 ;
        RECT 72.310 4.280 72.590 4.560 ;
        RECT 174.890 4.280 175.170 4.560 ;
      LAYER met3 ;
        RECT 5.000 2441.480 9.000 2442.080 ;
        RECT 7.670 2438.985 7.970 2441.480 ;
        RECT 7.670 2438.670 8.215 2438.985 ;
        RECT 7.885 2438.655 8.215 2438.670 ;
        RECT 72.285 4.570 72.615 4.585 ;
        RECT 95.950 4.570 96.330 4.580 ;
        RECT 72.285 4.270 96.330 4.570 ;
        RECT 72.285 4.255 72.615 4.270 ;
        RECT 95.950 4.260 96.330 4.270 ;
        RECT 141.030 4.570 141.410 4.580 ;
        RECT 174.865 4.570 175.195 4.585 ;
        RECT 141.030 4.270 175.195 4.570 ;
        RECT 141.030 4.260 141.410 4.270 ;
        RECT 174.865 4.255 175.195 4.270 ;
      LAYER via3 ;
        RECT 95.980 4.260 96.300 4.580 ;
        RECT 141.060 4.260 141.380 4.580 ;
      LAYER met4 ;
        RECT 95.550 4.510 96.730 5.690 ;
        RECT 140.630 4.510 141.810 5.690 ;
        RECT 95.975 4.255 96.305 4.510 ;
        RECT 141.055 4.255 141.385 4.510 ;
      LAYER via4 ;
        RECT 95.550 4.510 96.730 5.690 ;
        RECT 140.630 4.510 141.810 5.690 ;
      LAYER met5 ;
        RECT 95.340 4.300 142.020 5.900 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 317.545 0.935 317.715 1.275 ;
        RECT 318.465 0.935 318.635 4.335 ;
        RECT 488.665 3.485 492.515 3.655 ;
        RECT 478.545 1.615 478.715 2.295 ;
        RECT 488.665 1.615 488.835 3.485 ;
        RECT 478.545 1.445 488.835 1.615 ;
        RECT 492.345 1.615 492.515 3.485 ;
        RECT 513.045 2.805 515.975 2.975 ;
        RECT 554.445 2.805 554.615 4.335 ;
        RECT 559.045 4.165 559.675 4.335 ;
        RECT 559.505 3.995 559.675 4.165 ;
        RECT 559.505 3.825 560.135 3.995 ;
        RECT 513.045 1.955 513.215 2.805 ;
        RECT 505.225 1.785 513.215 1.955 ;
        RECT 505.225 1.615 505.395 1.785 ;
        RECT 492.345 1.445 505.395 1.615 ;
        RECT 317.545 0.765 318.635 0.935 ;
      LAYER mcon ;
        RECT 318.465 4.165 318.635 4.335 ;
        RECT 317.545 1.105 317.715 1.275 ;
        RECT 554.445 4.165 554.615 4.335 ;
        RECT 478.545 2.125 478.715 2.295 ;
        RECT 559.965 3.825 560.135 3.995 ;
        RECT 515.805 2.805 515.975 2.975 ;
      LAYER met1 ;
        RECT 239.730 6.360 240.050 6.420 ;
        RECT 243.410 6.360 243.730 6.420 ;
        RECT 239.730 6.220 243.730 6.360 ;
        RECT 239.730 6.160 240.050 6.220 ;
        RECT 243.410 6.160 243.730 6.220 ;
        RECT 417.750 5.680 418.070 5.740 ;
        RECT 417.750 5.540 460.760 5.680 ;
        RECT 417.750 5.480 418.070 5.540 ;
        RECT 460.620 5.340 460.760 5.540 ;
        RECT 463.750 5.340 464.070 5.400 ;
        RECT 460.620 5.200 464.070 5.340 ;
        RECT 463.750 5.140 464.070 5.200 ;
        RECT 318.405 4.320 318.695 4.365 ;
        RECT 318.850 4.320 319.170 4.380 ;
        RECT 318.405 4.180 319.170 4.320 ;
        RECT 318.405 4.135 318.695 4.180 ;
        RECT 318.850 4.120 319.170 4.180 ;
        RECT 384.170 4.320 384.490 4.380 ;
        RECT 412.690 4.320 413.010 4.380 ;
        RECT 384.170 4.180 413.010 4.320 ;
        RECT 384.170 4.120 384.490 4.180 ;
        RECT 412.690 4.120 413.010 4.180 ;
        RECT 554.385 4.320 554.675 4.365 ;
        RECT 558.985 4.320 559.275 4.365 ;
        RECT 554.385 4.180 559.275 4.320 ;
        RECT 554.385 4.135 554.675 4.180 ;
        RECT 558.985 4.135 559.275 4.180 ;
        RECT 559.905 3.980 560.195 4.025 ;
        RECT 561.730 3.980 562.050 4.040 ;
        RECT 559.905 3.840 562.050 3.980 ;
        RECT 559.905 3.795 560.195 3.840 ;
        RECT 561.730 3.780 562.050 3.840 ;
        RECT 515.745 2.960 516.035 3.005 ;
        RECT 554.385 2.960 554.675 3.005 ;
        RECT 515.745 2.820 554.675 2.960 ;
        RECT 515.745 2.775 516.035 2.820 ;
        RECT 554.385 2.775 554.675 2.820 ;
        RECT 463.750 2.280 464.070 2.340 ;
        RECT 478.485 2.280 478.775 2.325 ;
        RECT 463.750 2.140 478.775 2.280 ;
        RECT 463.750 2.080 464.070 2.140 ;
        RECT 478.485 2.095 478.775 2.140 ;
        RECT 305.050 1.260 305.370 1.320 ;
        RECT 317.485 1.260 317.775 1.305 ;
        RECT 305.050 1.120 317.775 1.260 ;
        RECT 305.050 1.060 305.370 1.120 ;
        RECT 317.485 1.075 317.775 1.120 ;
      LAYER via ;
        RECT 239.760 6.160 240.020 6.420 ;
        RECT 243.440 6.160 243.700 6.420 ;
        RECT 417.780 5.480 418.040 5.740 ;
        RECT 463.780 5.140 464.040 5.400 ;
        RECT 318.880 4.120 319.140 4.380 ;
        RECT 384.200 4.120 384.460 4.380 ;
        RECT 412.720 4.120 412.980 4.380 ;
        RECT 561.760 3.780 562.020 4.040 ;
        RECT 463.780 2.080 464.040 2.340 ;
        RECT 305.080 1.060 305.340 1.320 ;
      LAYER met2 ;
        RECT 275.170 8.315 275.450 8.685 ;
        RECT 368.550 8.400 368.830 8.685 ;
        RECT 378.280 8.430 382.100 8.570 ;
        RECT 368.550 8.315 377.500 8.400 ;
        RECT 243.430 7.635 243.710 8.005 ;
        RECT 243.500 6.450 243.640 7.635 ;
        RECT 275.240 7.325 275.380 8.315 ;
        RECT 368.620 8.260 377.500 8.315 ;
        RECT 305.070 7.635 305.350 8.005 ;
        RECT 377.360 7.890 377.500 8.260 ;
        RECT 378.280 7.890 378.420 8.430 ;
        RECT 381.960 8.400 382.100 8.430 ;
        RECT 381.960 8.260 386.240 8.400 ;
        RECT 377.360 7.750 378.420 7.890 ;
        RECT 275.170 6.955 275.450 7.325 ;
        RECT 239.760 6.130 240.020 6.450 ;
        RECT 243.440 6.130 243.700 6.450 ;
        RECT 239.820 4.605 239.960 6.130 ;
        RECT 192.830 4.235 193.110 4.605 ;
        RECT 239.750 4.235 240.030 4.605 ;
        RECT 192.900 2.400 193.040 4.235 ;
        RECT 192.690 -4.800 193.250 2.400 ;
        RECT 305.140 1.350 305.280 7.635 ;
        RECT 386.100 7.210 386.240 8.260 ;
        RECT 382.880 7.070 386.240 7.210 ;
        RECT 319.330 5.850 319.610 5.965 ;
        RECT 318.940 5.710 319.610 5.850 ;
        RECT 318.940 4.410 319.080 5.710 ;
        RECT 319.330 5.595 319.610 5.710 ;
        RECT 318.880 4.090 319.140 4.410 ;
        RECT 382.880 4.320 383.020 7.070 ;
        RECT 417.780 5.680 418.040 5.770 ;
        RECT 417.380 5.540 418.040 5.680 ;
        RECT 413.240 5.030 414.300 5.170 ;
        RECT 413.240 4.490 413.380 5.030 ;
        RECT 414.160 4.660 414.300 5.030 ;
        RECT 417.380 4.660 417.520 5.540 ;
        RECT 417.780 5.450 418.040 5.540 ;
        RECT 463.780 5.110 464.040 5.430 ;
        RECT 414.160 4.520 417.520 4.660 ;
        RECT 412.780 4.410 413.380 4.490 ;
        RECT 384.200 4.320 384.460 4.410 ;
        RECT 382.880 4.180 384.460 4.320 ;
        RECT 384.200 4.090 384.460 4.180 ;
        RECT 412.720 4.350 413.380 4.410 ;
        RECT 412.720 4.090 412.980 4.350 ;
        RECT 463.840 2.370 463.980 5.110 ;
        RECT 561.760 3.980 562.020 4.070 ;
        RECT 561.760 3.840 563.340 3.980 ;
        RECT 561.760 3.750 562.020 3.840 ;
        RECT 463.780 2.050 464.040 2.370 ;
        RECT 305.080 1.030 305.340 1.350 ;
        RECT 563.200 0.525 563.340 3.840 ;
        RECT 563.130 0.155 563.410 0.525 ;
      LAYER via2 ;
        RECT 275.170 8.360 275.450 8.640 ;
        RECT 368.550 8.360 368.830 8.640 ;
        RECT 243.430 7.680 243.710 7.960 ;
        RECT 305.070 7.680 305.350 7.960 ;
        RECT 275.170 7.000 275.450 7.280 ;
        RECT 192.830 4.280 193.110 4.560 ;
        RECT 239.750 4.280 240.030 4.560 ;
        RECT 319.330 5.640 319.610 5.920 ;
        RECT 563.130 0.200 563.410 0.480 ;
      LAYER met3 ;
        RECT 275.145 8.650 275.475 8.665 ;
        RECT 245.950 8.350 275.475 8.650 ;
        RECT 243.405 7.970 243.735 7.985 ;
        RECT 245.950 7.970 246.250 8.350 ;
        RECT 275.145 8.335 275.475 8.350 ;
        RECT 325.030 8.650 325.410 8.660 ;
        RECT 343.430 8.650 343.810 8.660 ;
        RECT 325.030 8.350 343.810 8.650 ;
        RECT 325.030 8.340 325.410 8.350 ;
        RECT 343.430 8.340 343.810 8.350 ;
        RECT 362.750 8.650 363.130 8.660 ;
        RECT 368.525 8.650 368.855 8.665 ;
        RECT 362.750 8.350 368.855 8.650 ;
        RECT 362.750 8.340 363.130 8.350 ;
        RECT 368.525 8.335 368.855 8.350 ;
        RECT 772.150 8.650 772.530 8.660 ;
        RECT 780.430 8.650 780.810 8.660 ;
        RECT 772.150 8.350 780.810 8.650 ;
        RECT 772.150 8.340 772.530 8.350 ;
        RECT 780.430 8.340 780.810 8.350 ;
        RECT 243.405 7.670 246.250 7.970 ;
        RECT 292.830 7.970 293.210 7.980 ;
        RECT 305.045 7.970 305.375 7.985 ;
        RECT 292.830 7.670 305.375 7.970 ;
        RECT 243.405 7.655 243.735 7.670 ;
        RECT 292.830 7.660 293.210 7.670 ;
        RECT 305.045 7.655 305.375 7.670 ;
        RECT 275.145 7.290 275.475 7.305 ;
        RECT 281.790 7.290 282.170 7.300 ;
        RECT 275.145 6.990 282.170 7.290 ;
        RECT 275.145 6.975 275.475 6.990 ;
        RECT 281.790 6.980 282.170 6.990 ;
        RECT 319.305 5.930 319.635 5.945 ;
        RECT 323.190 5.930 323.570 5.940 ;
        RECT 319.305 5.630 323.570 5.930 ;
        RECT 319.305 5.615 319.635 5.630 ;
        RECT 323.190 5.620 323.570 5.630 ;
        RECT 192.805 4.570 193.135 4.585 ;
        RECT 239.725 4.570 240.055 4.585 ;
        RECT 192.805 4.270 240.055 4.570 ;
        RECT 192.805 4.255 193.135 4.270 ;
        RECT 239.725 4.255 240.055 4.270 ;
        RECT 583.550 0.860 583.930 1.180 ;
        RECT 563.105 0.490 563.435 0.505 ;
        RECT 583.590 0.490 583.890 0.860 ;
        RECT 563.105 0.190 583.890 0.490 ;
        RECT 563.105 0.175 563.435 0.190 ;
      LAYER via3 ;
        RECT 325.060 8.340 325.380 8.660 ;
        RECT 343.460 8.340 343.780 8.660 ;
        RECT 362.780 8.340 363.100 8.660 ;
        RECT 772.180 8.340 772.500 8.660 ;
        RECT 780.460 8.340 780.780 8.660 ;
        RECT 292.860 7.660 293.180 7.980 ;
        RECT 281.820 6.980 282.140 7.300 ;
        RECT 323.220 5.620 323.540 5.940 ;
        RECT 583.580 0.860 583.900 1.180 ;
      LAYER met4 ;
        RECT 889.280 18.110 890.460 19.290 ;
        RECT 635.590 14.710 636.770 15.890 ;
        RECT 771.750 14.710 772.930 15.890 ;
        RECT 780.030 14.710 781.210 15.890 ;
        RECT 636.030 12.050 636.330 14.710 ;
        RECT 633.500 11.750 636.330 12.050 ;
        RECT 325.055 8.650 325.385 8.665 ;
        RECT 323.230 8.350 325.385 8.650 ;
        RECT 292.855 7.970 293.185 7.985 ;
        RECT 281.830 7.670 293.185 7.970 ;
        RECT 281.830 7.305 282.130 7.670 ;
        RECT 292.855 7.655 293.185 7.670 ;
        RECT 281.815 6.975 282.145 7.305 ;
        RECT 323.230 5.945 323.530 8.350 ;
        RECT 325.055 8.335 325.385 8.350 ;
        RECT 343.455 8.650 343.785 8.665 ;
        RECT 362.775 8.650 363.105 8.665 ;
        RECT 343.455 8.350 363.105 8.650 ;
        RECT 343.455 8.335 343.785 8.350 ;
        RECT 362.775 8.335 363.105 8.350 ;
        RECT 633.500 7.290 633.800 11.750 ;
        RECT 772.190 8.665 772.490 14.710 ;
        RECT 780.470 8.665 780.770 14.710 ;
        RECT 772.175 8.335 772.505 8.665 ;
        RECT 780.455 8.335 780.785 8.665 ;
        RECT 633.500 6.990 635.410 7.290 ;
        RECT 621.310 6.310 628.050 6.610 ;
        RECT 323.215 5.615 323.545 5.945 ;
        RECT 621.310 4.570 621.610 6.310 ;
        RECT 627.750 5.250 628.050 6.310 ;
        RECT 635.110 5.250 635.410 6.990 ;
        RECT 627.750 4.950 635.410 5.250 ;
        RECT 620.390 4.270 621.610 4.570 ;
        RECT 620.390 3.890 620.690 4.270 ;
        RECT 615.790 3.590 620.690 3.890 ;
        RECT 583.575 1.170 583.905 1.185 ;
        RECT 615.790 1.170 616.090 3.590 ;
        RECT 583.575 0.870 616.090 1.170 ;
        RECT 583.575 0.855 583.905 0.870 ;
      LAYER met5 ;
        RECT 674.940 21.300 763.710 22.900 ;
        RECT 674.940 16.100 676.540 21.300 ;
        RECT 762.110 19.500 763.710 21.300 ;
        RECT 762.110 17.900 773.140 19.500 ;
        RECT 635.380 14.500 676.540 16.100 ;
        RECT 771.540 14.500 773.140 17.900 ;
        RECT 779.820 17.900 890.670 19.500 ;
        RECT 779.820 14.500 781.420 17.900 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 8.425 914.345 8.595 978.435 ;
        RECT 7.505 818.295 7.675 878.135 ;
        RECT 7.045 818.125 7.675 818.295 ;
        RECT 7.045 796.705 7.215 818.125 ;
        RECT 7.045 144.925 7.215 196.775 ;
        RECT 4.745 118.745 4.915 144.415 ;
        RECT 131.245 6.545 131.415 8.755 ;
        RECT 171.725 5.525 171.895 6.715 ;
        RECT 191.965 4.165 192.135 5.695 ;
        RECT 28.665 1.275 28.835 1.955 ;
        RECT 48.445 1.445 48.615 2.975 ;
        RECT 52.125 1.785 52.295 2.975 ;
        RECT 71.445 1.785 71.615 2.975 ;
        RECT 28.205 1.105 28.835 1.275 ;
      LAYER mcon ;
        RECT 8.425 978.265 8.595 978.435 ;
        RECT 7.505 877.965 7.675 878.135 ;
        RECT 7.045 196.605 7.215 196.775 ;
        RECT 4.745 144.245 4.915 144.415 ;
        RECT 131.245 8.585 131.415 8.755 ;
        RECT 171.725 6.545 171.895 6.715 ;
        RECT 191.965 5.525 192.135 5.695 ;
        RECT 48.445 2.805 48.615 2.975 ;
        RECT 28.665 1.785 28.835 1.955 ;
        RECT 52.125 2.805 52.295 2.975 ;
        RECT 71.445 2.805 71.615 2.975 ;
      LAYER met1 ;
        RECT 7.430 978.420 7.750 978.480 ;
        RECT 8.365 978.420 8.655 978.465 ;
        RECT 7.430 978.280 8.655 978.420 ;
        RECT 7.430 978.220 7.750 978.280 ;
        RECT 8.365 978.235 8.655 978.280 ;
        RECT 6.050 914.500 6.370 914.560 ;
        RECT 8.365 914.500 8.655 914.545 ;
        RECT 6.050 914.360 8.655 914.500 ;
        RECT 6.050 914.300 6.370 914.360 ;
        RECT 8.365 914.315 8.655 914.360 ;
        RECT 6.050 878.120 6.370 878.180 ;
        RECT 7.445 878.120 7.735 878.165 ;
        RECT 6.050 877.980 7.735 878.120 ;
        RECT 6.050 877.920 6.370 877.980 ;
        RECT 7.445 877.935 7.735 877.980 ;
        RECT 6.985 796.860 7.275 796.905 ;
        RECT 7.430 796.860 7.750 796.920 ;
        RECT 6.985 796.720 7.750 796.860 ;
        RECT 6.985 796.675 7.275 796.720 ;
        RECT 7.430 796.660 7.750 796.720 ;
        RECT 6.985 196.760 7.275 196.805 ;
        RECT 7.430 196.760 7.750 196.820 ;
        RECT 6.985 196.620 7.750 196.760 ;
        RECT 6.985 196.575 7.275 196.620 ;
        RECT 7.430 196.560 7.750 196.620 ;
        RECT 6.985 145.080 7.275 145.125 ;
        RECT 6.985 144.940 7.660 145.080 ;
        RECT 6.985 144.895 7.275 144.940 ;
        RECT 4.685 144.400 4.975 144.445 ;
        RECT 7.520 144.400 7.660 144.940 ;
        RECT 4.685 144.260 7.660 144.400 ;
        RECT 4.685 144.215 4.975 144.260 ;
        RECT 4.685 118.900 4.975 118.945 ;
        RECT 7.430 118.900 7.750 118.960 ;
        RECT 4.685 118.760 7.750 118.900 ;
        RECT 4.685 118.715 4.975 118.760 ;
        RECT 7.430 118.700 7.750 118.760 ;
        RECT 110.930 8.740 111.250 8.800 ;
        RECT 131.185 8.740 131.475 8.785 ;
        RECT 110.930 8.600 131.475 8.740 ;
        RECT 110.930 8.540 111.250 8.600 ;
        RECT 131.185 8.555 131.475 8.600 ;
        RECT 131.185 6.700 131.475 6.745 ;
        RECT 171.665 6.700 171.955 6.745 ;
        RECT 131.185 6.560 171.955 6.700 ;
        RECT 131.185 6.515 131.475 6.560 ;
        RECT 171.665 6.515 171.955 6.560 ;
        RECT 171.665 5.680 171.955 5.725 ;
        RECT 191.905 5.680 192.195 5.725 ;
        RECT 171.665 5.540 192.195 5.680 ;
        RECT 171.665 5.495 171.955 5.540 ;
        RECT 191.905 5.495 192.195 5.540 ;
        RECT 191.905 4.320 192.195 4.365 ;
        RECT 210.750 4.320 211.070 4.380 ;
        RECT 191.905 4.180 211.070 4.320 ;
        RECT 191.905 4.135 192.195 4.180 ;
        RECT 210.750 4.120 211.070 4.180 ;
        RECT 48.385 2.960 48.675 3.005 ;
        RECT 52.065 2.960 52.355 3.005 ;
        RECT 48.385 2.820 52.355 2.960 ;
        RECT 48.385 2.775 48.675 2.820 ;
        RECT 52.065 2.775 52.355 2.820 ;
        RECT 71.385 2.960 71.675 3.005 ;
        RECT 110.930 2.960 111.250 3.020 ;
        RECT 71.385 2.820 111.250 2.960 ;
        RECT 71.385 2.775 71.675 2.820 ;
        RECT 110.930 2.760 111.250 2.820 ;
        RECT 28.605 1.755 28.895 1.985 ;
        RECT 52.065 1.940 52.355 1.985 ;
        RECT 71.385 1.940 71.675 1.985 ;
        RECT 52.065 1.800 71.675 1.940 ;
        RECT 52.065 1.755 52.355 1.800 ;
        RECT 71.385 1.755 71.675 1.800 ;
        RECT 28.680 1.600 28.820 1.755 ;
        RECT 48.385 1.600 48.675 1.645 ;
        RECT 28.680 1.460 48.675 1.600 ;
        RECT 48.385 1.415 48.675 1.460 ;
        RECT 6.970 1.260 7.290 1.320 ;
        RECT 28.145 1.260 28.435 1.305 ;
        RECT 6.970 1.120 28.435 1.260 ;
        RECT 6.970 1.060 7.290 1.120 ;
        RECT 28.145 1.075 28.435 1.120 ;
      LAYER via ;
        RECT 7.460 978.220 7.720 978.480 ;
        RECT 6.080 914.300 6.340 914.560 ;
        RECT 6.080 877.920 6.340 878.180 ;
        RECT 7.460 796.660 7.720 796.920 ;
        RECT 7.460 196.560 7.720 196.820 ;
        RECT 7.460 118.700 7.720 118.960 ;
        RECT 110.960 8.540 111.220 8.800 ;
        RECT 210.780 4.120 211.040 4.380 ;
        RECT 110.960 2.760 111.220 3.020 ;
        RECT 7.000 1.060 7.260 1.320 ;
      LAYER met2 ;
        RECT 7.450 2552.875 7.730 2553.245 ;
        RECT 7.520 978.510 7.660 2552.875 ;
        RECT 7.460 978.190 7.720 978.510 ;
        RECT 6.080 914.270 6.340 914.590 ;
        RECT 6.140 878.210 6.280 914.270 ;
        RECT 6.080 877.890 6.340 878.210 ;
        RECT 7.460 796.630 7.720 796.950 ;
        RECT 7.520 714.410 7.660 796.630 ;
        RECT 7.520 714.270 8.120 714.410 ;
        RECT 7.980 672.250 8.120 714.270 ;
        RECT 7.980 672.110 8.580 672.250 ;
        RECT 8.440 662.050 8.580 672.110 ;
        RECT 7.520 661.910 8.580 662.050 ;
        RECT 7.520 196.850 7.660 661.910 ;
        RECT 7.460 196.530 7.720 196.850 ;
        RECT 7.460 118.670 7.720 118.990 ;
        RECT 7.520 79.290 7.660 118.670 ;
        RECT 7.060 79.150 7.660 79.290 ;
        RECT 7.060 1.350 7.200 79.150 ;
        RECT 110.960 8.510 111.220 8.830 ;
        RECT 111.020 3.050 111.160 8.510 ;
        RECT 210.780 4.090 211.040 4.410 ;
        RECT 110.960 2.730 111.220 3.050 ;
        RECT 210.840 2.400 210.980 4.090 ;
        RECT 7.000 1.030 7.260 1.350 ;
        RECT 210.630 -4.800 211.190 2.400 ;
      LAYER via2 ;
        RECT 7.450 2552.920 7.730 2553.200 ;
      LAYER met3 ;
        RECT 5.000 2554.360 9.000 2554.960 ;
        RECT 7.670 2553.225 7.970 2554.360 ;
        RECT 7.425 2552.910 7.970 2553.225 ;
        RECT 7.425 2552.895 7.755 2552.910 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 394.290 7.040 394.610 7.100 ;
        RECT 406.710 7.040 407.030 7.100 ;
        RECT 394.290 6.900 407.030 7.040 ;
        RECT 394.290 6.840 394.610 6.900 ;
        RECT 406.710 6.840 407.030 6.900 ;
      LAYER via ;
        RECT 394.320 6.840 394.580 7.100 ;
        RECT 406.740 6.840 407.000 7.100 ;
      LAYER met2 ;
        RECT 392.080 8.260 393.600 8.400 ;
        RECT 392.080 8.005 392.220 8.260 ;
        RECT 385.570 7.890 385.850 8.005 ;
        RECT 381.960 7.750 385.850 7.890 ;
        RECT 50.300 2.990 51.360 3.130 ;
        RECT 50.300 2.400 50.440 2.990 ;
        RECT 50.090 -4.800 50.650 2.400 ;
        RECT 51.220 0.525 51.360 2.990 ;
        RECT 378.670 2.195 378.950 2.565 ;
        RECT 378.740 1.770 378.880 2.195 ;
        RECT 381.960 1.770 382.100 7.750 ;
        RECT 385.570 7.635 385.850 7.750 ;
        RECT 392.010 7.635 392.290 8.005 ;
        RECT 393.460 7.040 393.600 8.260 ;
        RECT 408.510 7.210 408.790 9.000 ;
        RECT 406.800 7.130 408.790 7.210 ;
        RECT 394.320 7.040 394.580 7.130 ;
        RECT 393.460 6.900 394.580 7.040 ;
        RECT 394.320 6.810 394.580 6.900 ;
        RECT 406.740 7.070 408.790 7.130 ;
        RECT 406.740 6.810 407.000 7.070 ;
        RECT 408.510 5.000 408.790 7.070 ;
        RECT 378.740 1.630 382.100 1.770 ;
        RECT 51.150 0.155 51.430 0.525 ;
      LAYER via2 ;
        RECT 378.670 2.240 378.950 2.520 ;
        RECT 385.570 7.680 385.850 7.960 ;
        RECT 392.010 7.680 392.290 7.960 ;
        RECT 51.150 0.200 51.430 0.480 ;
      LAYER met3 ;
        RECT 385.545 7.970 385.875 7.985 ;
        RECT 391.985 7.970 392.315 7.985 ;
        RECT 385.545 7.670 392.315 7.970 ;
        RECT 385.545 7.655 385.875 7.670 ;
        RECT 391.985 7.655 392.315 7.670 ;
        RECT 371.030 2.530 371.410 2.540 ;
        RECT 378.645 2.530 378.975 2.545 ;
        RECT 371.030 2.230 378.975 2.530 ;
        RECT 371.030 2.220 371.410 2.230 ;
        RECT 378.645 2.215 378.975 2.230 ;
        RECT 369.190 1.170 369.570 1.180 ;
        RECT 368.310 0.870 369.570 1.170 ;
        RECT 51.125 0.490 51.455 0.505 ;
        RECT 368.310 0.490 368.610 0.870 ;
        RECT 369.190 0.860 369.570 0.870 ;
        RECT 51.125 0.190 368.610 0.490 ;
        RECT 51.125 0.175 51.455 0.190 ;
      LAYER via3 ;
        RECT 371.060 2.220 371.380 2.540 ;
        RECT 369.220 0.860 369.540 1.180 ;
      LAYER met4 ;
        RECT 371.055 2.530 371.385 2.545 ;
        RECT 369.230 2.230 371.385 2.530 ;
        RECT 369.230 1.185 369.530 2.230 ;
        RECT 371.055 2.215 371.385 2.230 ;
        RECT 369.215 0.855 369.545 1.185 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 621.605 15.215 621.775 15.555 ;
        RECT 628.045 15.385 634.195 15.555 ;
        RECT 628.045 15.215 628.215 15.385 ;
        RECT 621.605 15.045 629.135 15.215 ;
        RECT 628.045 13.855 628.215 15.045 ;
        RECT 613.325 13.685 628.215 13.855 ;
        RECT 579.285 9.605 581.755 9.775 ;
        RECT 508.905 6.885 510.455 7.055 ;
        RECT 508.905 6.715 509.075 6.885 ;
        RECT 336.865 5.185 344.855 5.355 ;
        RECT 336.865 1.275 337.035 5.185 ;
        RECT 364.925 4.505 365.095 5.355 ;
        RECT 377.345 4.845 380.275 5.015 ;
        RECT 377.345 4.505 377.515 4.845 ;
        RECT 380.105 4.165 380.275 4.845 ;
        RECT 383.785 4.165 383.955 6.715 ;
        RECT 415.525 6.375 415.695 6.715 ;
        RECT 483.145 6.545 509.075 6.715 ;
        RECT 415.525 6.205 417.075 6.375 ;
        RECT 416.905 4.165 417.075 6.205 ;
        RECT 483.145 5.355 483.315 6.545 ;
        RECT 529.605 5.525 529.775 7.055 ;
        RECT 579.285 5.525 579.455 9.605 ;
        RECT 581.585 9.435 581.755 9.605 ;
        RECT 581.585 9.265 612.115 9.435 ;
        RECT 611.945 6.035 612.115 9.265 ;
        RECT 613.325 7.225 613.495 13.685 ;
        RECT 628.965 12.835 629.135 15.045 ;
        RECT 624.365 12.665 629.595 12.835 ;
        RECT 622.065 8.245 623.615 8.415 ;
        RECT 610.105 5.865 612.115 6.035 ;
        RECT 467.045 5.185 483.315 5.355 ;
        RECT 467.045 4.165 467.215 5.185 ;
        RECT 610.105 2.975 610.275 5.865 ;
        RECT 622.065 2.975 622.235 8.245 ;
        RECT 624.365 3.995 624.535 12.665 ;
        RECT 628.965 11.135 629.135 12.665 ;
        RECT 626.205 10.965 629.135 11.135 ;
        RECT 626.205 6.035 626.375 10.965 ;
        RECT 629.425 10.795 629.595 12.665 ;
        RECT 634.025 11.815 634.195 15.385 ;
        RECT 710.845 12.325 737.235 12.495 ;
        RECT 710.845 12.155 711.015 12.325 ;
        RECT 662.545 11.985 711.015 12.155 ;
        RECT 737.065 12.155 737.235 12.325 ;
        RECT 737.065 11.985 780.935 12.155 ;
        RECT 662.545 11.815 662.715 11.985 ;
        RECT 634.025 11.645 662.715 11.815 ;
        RECT 780.765 11.815 780.935 11.985 ;
        RECT 780.765 11.645 801.175 11.815 ;
        RECT 801.005 11.475 801.175 11.645 ;
        RECT 780.765 11.305 787.375 11.475 ;
        RECT 648.745 10.965 649.835 11.135 ;
        RECT 648.745 10.795 648.915 10.965 ;
        RECT 629.425 10.625 648.915 10.795 ;
        RECT 649.665 10.795 649.835 10.965 ;
        RECT 649.665 10.625 695.835 10.795 ;
        RECT 695.665 10.115 695.835 10.625 ;
        RECT 739.365 10.625 772.655 10.795 ;
        RECT 695.665 9.945 718.835 10.115 ;
        RECT 642.305 9.265 671.915 9.435 ;
        RECT 628.505 7.905 628.675 9.095 ;
        RECT 642.305 8.925 642.475 9.265 ;
        RECT 671.745 8.925 671.915 9.265 ;
        RECT 718.665 9.095 718.835 9.945 ;
        RECT 724.185 9.605 734.475 9.775 ;
        RECT 703.025 8.925 708.715 9.095 ;
        RECT 718.665 8.925 723.435 9.095 ;
        RECT 629.425 8.245 630.975 8.415 ;
        RECT 628.045 6.035 628.215 7.395 ;
        RECT 629.425 7.225 629.595 8.245 ;
        RECT 630.805 7.055 630.975 8.245 ;
        RECT 641.385 7.055 641.555 8.755 ;
        RECT 703.025 8.415 703.195 8.925 ;
        RECT 708.545 8.585 708.715 8.925 ;
        RECT 692.445 7.735 692.615 8.415 ;
        RECT 701.645 8.245 703.195 8.415 ;
        RECT 723.265 8.075 723.435 8.925 ;
        RECT 724.185 8.585 724.355 9.605 ;
        RECT 734.305 9.435 734.475 9.605 ;
        RECT 734.305 9.265 736.315 9.435 ;
        RECT 736.145 8.925 736.315 9.265 ;
        RECT 739.365 8.925 739.535 10.625 ;
        RECT 745.805 9.265 751.955 9.435 ;
        RECT 745.805 8.925 745.975 9.265 ;
        RECT 751.785 8.925 751.955 9.265 ;
        RECT 744.425 8.585 745.055 8.755 ;
        RECT 723.265 7.905 724.355 8.075 ;
        RECT 744.425 7.905 744.595 8.585 ;
        RECT 692.445 7.565 705.955 7.735 ;
        RECT 757.305 7.565 757.475 9.095 ;
        RECT 772.485 8.925 772.655 10.625 ;
        RECT 780.765 8.925 780.935 11.305 ;
        RECT 787.205 10.795 787.375 11.305 ;
        RECT 789.045 11.305 797.955 11.475 ;
        RECT 801.005 11.305 808.995 11.475 ;
        RECT 789.045 10.795 789.215 11.305 ;
        RECT 797.785 11.135 797.955 11.305 ;
        RECT 797.785 10.965 806.235 11.135 ;
        RECT 787.205 10.625 789.215 10.795 ;
        RECT 806.065 10.115 806.235 10.965 ;
        RECT 806.065 9.945 808.535 10.115 ;
        RECT 808.365 8.585 808.535 9.945 ;
        RECT 630.805 6.885 641.555 7.055 ;
        RECT 626.205 5.865 628.215 6.035 ;
        RECT 705.785 4.505 705.955 7.565 ;
        RECT 759.605 7.055 759.775 7.735 ;
        RECT 759.605 6.885 763.455 7.055 ;
        RECT 763.285 6.035 763.455 6.885 ;
        RECT 762.365 5.865 763.455 6.035 ;
        RECT 739.825 5.355 739.995 5.695 ;
        RECT 739.825 5.185 740.915 5.355 ;
        RECT 711.765 4.335 711.935 4.675 ;
        RECT 716.365 4.335 716.535 4.675 ;
        RECT 762.365 4.505 762.535 5.865 ;
        RECT 711.765 4.165 716.535 4.335 ;
        RECT 622.525 3.825 624.535 3.995 ;
        RECT 622.525 3.145 622.695 3.825 ;
        RECT 610.105 2.805 622.235 2.975 ;
        RECT 791.345 2.975 791.515 5.695 ;
        RECT 795.945 2.975 796.115 7.735 ;
        RECT 808.825 6.205 808.995 11.305 ;
        RECT 884.725 6.885 888.115 7.055 ;
        RECT 889.785 6.885 889.955 8.075 ;
        RECT 1454.205 7.905 1455.295 8.075 ;
        RECT 884.725 6.205 884.895 6.885 ;
        RECT 973.045 6.545 976.895 6.715 ;
        RECT 899.905 4.165 900.535 4.335 ;
        RECT 791.345 2.805 796.115 2.975 ;
        RECT 887.025 2.295 887.195 3.315 ;
        RECT 899.905 2.295 900.075 4.165 ;
        RECT 919.685 3.485 920.315 3.655 ;
        RECT 920.145 2.635 920.315 3.485 ;
        RECT 973.045 3.315 973.215 6.545 ;
        RECT 983.165 6.035 983.335 6.715 ;
        RECT 983.165 5.865 984.255 6.035 ;
        RECT 956.485 3.145 973.215 3.315 ;
        RECT 956.485 2.975 956.655 3.145 ;
        RECT 952.805 2.805 956.655 2.975 ;
        RECT 952.805 2.635 952.975 2.805 ;
        RECT 920.145 2.465 952.975 2.635 ;
        RECT 984.085 2.635 984.255 5.865 ;
        RECT 1437.185 3.655 1437.355 4.335 ;
        RECT 1453.285 3.655 1453.455 6.035 ;
        RECT 1454.205 5.865 1454.375 7.905 ;
        RECT 1090.805 3.485 1098.795 3.655 ;
        RECT 996.505 3.145 1022.435 3.315 ;
        RECT 984.085 2.465 992.995 2.635 ;
        RECT 887.025 2.125 900.075 2.295 ;
        RECT 992.825 1.955 992.995 2.465 ;
        RECT 992.825 1.785 993.455 1.955 ;
        RECT 996.505 1.785 996.675 3.145 ;
        RECT 1090.805 2.635 1090.975 3.485 ;
        RECT 1098.625 2.975 1098.795 3.485 ;
        RECT 1127.605 3.485 1159.055 3.655 ;
        RECT 1437.185 3.485 1453.455 3.655 ;
        RECT 1098.625 2.805 1111.215 2.975 ;
        RECT 1089.425 2.465 1090.975 2.635 ;
        RECT 1111.045 2.635 1111.215 2.805 ;
        RECT 1127.605 2.635 1127.775 3.485 ;
        RECT 1111.045 2.465 1127.775 2.635 ;
        RECT 336.405 1.105 337.035 1.275 ;
      LAYER mcon ;
        RECT 621.605 15.385 621.775 15.555 ;
        RECT 510.285 6.885 510.455 7.055 ;
        RECT 529.605 6.885 529.775 7.055 ;
        RECT 383.785 6.545 383.955 6.715 ;
        RECT 344.685 5.185 344.855 5.355 ;
        RECT 364.925 5.185 365.095 5.355 ;
        RECT 415.525 6.545 415.695 6.715 ;
        RECT 623.445 8.245 623.615 8.415 ;
        RECT 628.505 8.925 628.675 9.095 ;
        RECT 641.385 8.585 641.555 8.755 ;
        RECT 628.045 7.225 628.215 7.395 ;
        RECT 692.445 8.245 692.615 8.415 ;
        RECT 757.305 8.925 757.475 9.095 ;
        RECT 744.885 8.585 745.055 8.755 ;
        RECT 724.185 7.905 724.355 8.075 ;
        RECT 759.605 7.565 759.775 7.735 ;
        RECT 795.945 7.565 796.115 7.735 ;
        RECT 739.825 5.525 739.995 5.695 ;
        RECT 740.745 5.185 740.915 5.355 ;
        RECT 711.765 4.505 711.935 4.675 ;
        RECT 716.365 4.505 716.535 4.675 ;
        RECT 791.345 5.525 791.515 5.695 ;
        RECT 889.785 7.905 889.955 8.075 ;
        RECT 887.945 6.885 888.115 7.055 ;
        RECT 1455.125 7.905 1455.295 8.075 ;
        RECT 976.725 6.545 976.895 6.715 ;
        RECT 983.165 6.545 983.335 6.715 ;
        RECT 900.365 4.165 900.535 4.335 ;
        RECT 887.025 3.145 887.195 3.315 ;
        RECT 1453.285 5.865 1453.455 6.035 ;
        RECT 1437.185 4.165 1437.355 4.335 ;
        RECT 1022.265 3.145 1022.435 3.315 ;
        RECT 1158.885 3.485 1159.055 3.655 ;
        RECT 993.285 1.785 993.455 1.955 ;
      LAYER met1 ;
        RECT 628.445 9.080 628.735 9.125 ;
        RECT 642.245 9.080 642.535 9.125 ;
        RECT 628.445 8.940 642.535 9.080 ;
        RECT 628.445 8.895 628.735 8.940 ;
        RECT 642.245 8.895 642.535 8.940 ;
        RECT 671.685 9.080 671.975 9.125 ;
        RECT 736.085 9.080 736.375 9.125 ;
        RECT 739.305 9.080 739.595 9.125 ;
        RECT 671.685 8.940 672.820 9.080 ;
        RECT 671.685 8.895 671.975 8.940 ;
        RECT 641.310 8.740 641.630 8.800 ;
        RECT 641.115 8.600 641.630 8.740 ;
        RECT 672.680 8.740 672.820 8.940 ;
        RECT 736.085 8.940 739.595 9.080 ;
        RECT 736.085 8.895 736.375 8.940 ;
        RECT 739.305 8.895 739.595 8.940 ;
        RECT 745.745 8.895 746.035 9.125 ;
        RECT 751.725 9.080 752.015 9.125 ;
        RECT 757.245 9.080 757.535 9.125 ;
        RECT 751.725 8.940 757.535 9.080 ;
        RECT 751.725 8.895 752.015 8.940 ;
        RECT 757.245 8.895 757.535 8.940 ;
        RECT 772.425 9.080 772.715 9.125 ;
        RECT 780.705 9.080 780.995 9.125 ;
        RECT 772.425 8.940 780.995 9.080 ;
        RECT 772.425 8.895 772.715 8.940 ;
        RECT 780.705 8.895 780.995 8.940 ;
        RECT 708.485 8.740 708.775 8.785 ;
        RECT 724.125 8.740 724.415 8.785 ;
        RECT 672.680 8.600 694.440 8.740 ;
        RECT 641.310 8.540 641.630 8.600 ;
        RECT 623.385 8.400 623.675 8.445 ;
        RECT 691.910 8.400 692.230 8.460 ;
        RECT 692.385 8.400 692.675 8.445 ;
        RECT 623.385 8.260 627.280 8.400 ;
        RECT 623.385 8.215 623.675 8.260 ;
        RECT 627.140 8.060 627.280 8.260 ;
        RECT 691.910 8.260 692.675 8.400 ;
        RECT 694.300 8.400 694.440 8.600 ;
        RECT 708.485 8.600 724.415 8.740 ;
        RECT 708.485 8.555 708.775 8.600 ;
        RECT 724.125 8.555 724.415 8.600 ;
        RECT 744.825 8.740 745.115 8.785 ;
        RECT 745.820 8.740 745.960 8.895 ;
        RECT 744.825 8.600 745.960 8.740 ;
        RECT 808.305 8.740 808.595 8.785 ;
        RECT 847.390 8.740 847.710 8.800 ;
        RECT 808.305 8.600 847.710 8.740 ;
        RECT 744.825 8.555 745.115 8.600 ;
        RECT 808.305 8.555 808.595 8.600 ;
        RECT 847.390 8.540 847.710 8.600 ;
        RECT 871.310 8.740 871.630 8.800 ;
        RECT 876.370 8.740 876.690 8.800 ;
        RECT 871.310 8.600 876.690 8.740 ;
        RECT 871.310 8.540 871.630 8.600 ;
        RECT 876.370 8.540 876.690 8.600 ;
        RECT 1764.630 8.740 1764.950 8.800 ;
        RECT 1831.790 8.740 1832.110 8.800 ;
        RECT 1764.630 8.600 1832.110 8.740 ;
        RECT 1764.630 8.540 1764.950 8.600 ;
        RECT 1831.790 8.540 1832.110 8.600 ;
        RECT 701.585 8.400 701.875 8.445 ;
        RECT 694.300 8.260 701.875 8.400 ;
        RECT 691.910 8.200 692.230 8.260 ;
        RECT 692.385 8.215 692.675 8.260 ;
        RECT 701.585 8.215 701.875 8.260 ;
        RECT 1573.730 8.400 1574.050 8.460 ;
        RECT 1598.570 8.400 1598.890 8.460 ;
        RECT 1573.730 8.260 1598.890 8.400 ;
        RECT 1573.730 8.200 1574.050 8.260 ;
        RECT 1598.570 8.200 1598.890 8.260 ;
        RECT 628.445 8.060 628.735 8.105 ;
        RECT 627.140 7.920 628.735 8.060 ;
        RECT 628.445 7.875 628.735 7.920 ;
        RECT 724.125 8.060 724.415 8.105 ;
        RECT 744.365 8.060 744.655 8.105 ;
        RECT 724.125 7.920 744.655 8.060 ;
        RECT 724.125 7.875 724.415 7.920 ;
        RECT 744.365 7.875 744.655 7.920 ;
        RECT 889.725 8.060 890.015 8.105 ;
        RECT 893.390 8.060 893.710 8.120 ;
        RECT 889.725 7.920 893.710 8.060 ;
        RECT 889.725 7.875 890.015 7.920 ;
        RECT 893.390 7.860 893.710 7.920 ;
        RECT 1455.065 8.060 1455.355 8.105 ;
        RECT 1468.390 8.060 1468.710 8.120 ;
        RECT 1455.065 7.920 1468.710 8.060 ;
        RECT 1455.065 7.875 1455.355 7.920 ;
        RECT 1468.390 7.860 1468.710 7.920 ;
        RECT 757.245 7.720 757.535 7.765 ;
        RECT 759.545 7.720 759.835 7.765 ;
        RECT 757.245 7.580 759.835 7.720 ;
        RECT 757.245 7.535 757.535 7.580 ;
        RECT 759.545 7.535 759.835 7.580 ;
        RECT 795.885 7.720 796.175 7.765 ;
        RECT 801.390 7.720 801.710 7.780 ;
        RECT 795.885 7.580 801.710 7.720 ;
        RECT 795.885 7.535 796.175 7.580 ;
        RECT 801.390 7.520 801.710 7.580 ;
        RECT 613.265 7.380 613.555 7.425 ;
        RECT 611.040 7.240 613.555 7.380 ;
        RECT 510.225 7.040 510.515 7.085 ;
        RECT 529.545 7.040 529.835 7.085 ;
        RECT 510.225 6.900 529.835 7.040 ;
        RECT 510.225 6.855 510.515 6.900 ;
        RECT 529.545 6.855 529.835 6.900 ;
        RECT 610.030 7.040 610.350 7.100 ;
        RECT 611.040 7.040 611.180 7.240 ;
        RECT 613.265 7.195 613.555 7.240 ;
        RECT 627.985 7.380 628.275 7.425 ;
        RECT 629.365 7.380 629.655 7.425 ;
        RECT 627.985 7.240 629.655 7.380 ;
        RECT 627.985 7.195 628.275 7.240 ;
        RECT 629.365 7.195 629.655 7.240 ;
        RECT 846.930 7.380 847.250 7.440 ;
        RECT 857.510 7.380 857.830 7.440 ;
        RECT 846.930 7.240 857.830 7.380 ;
        RECT 846.930 7.180 847.250 7.240 ;
        RECT 857.510 7.180 857.830 7.240 ;
        RECT 1328.090 7.380 1328.410 7.440 ;
        RECT 1343.270 7.380 1343.590 7.440 ;
        RECT 1328.090 7.240 1343.590 7.380 ;
        RECT 1328.090 7.180 1328.410 7.240 ;
        RECT 1343.270 7.180 1343.590 7.240 ;
        RECT 1469.770 7.380 1470.090 7.440 ;
        RECT 1473.910 7.380 1474.230 7.440 ;
        RECT 1469.770 7.240 1474.230 7.380 ;
        RECT 1469.770 7.180 1470.090 7.240 ;
        RECT 1473.910 7.180 1474.230 7.240 ;
        RECT 610.030 6.900 611.180 7.040 ;
        RECT 887.885 7.040 888.175 7.085 ;
        RECT 889.725 7.040 890.015 7.085 ;
        RECT 887.885 6.900 890.015 7.040 ;
        RECT 610.030 6.840 610.350 6.900 ;
        RECT 887.885 6.855 888.175 6.900 ;
        RECT 889.725 6.855 890.015 6.900 ;
        RECT 383.725 6.700 384.015 6.745 ;
        RECT 415.465 6.700 415.755 6.745 ;
        RECT 383.725 6.560 415.755 6.700 ;
        RECT 383.725 6.515 384.015 6.560 ;
        RECT 415.465 6.515 415.755 6.560 ;
        RECT 976.665 6.700 976.955 6.745 ;
        RECT 983.105 6.700 983.395 6.745 ;
        RECT 976.665 6.560 983.395 6.700 ;
        RECT 976.665 6.515 976.955 6.560 ;
        RECT 983.105 6.515 983.395 6.560 ;
        RECT 808.765 6.360 809.055 6.405 ;
        RECT 811.510 6.360 811.830 6.420 ;
        RECT 808.765 6.220 811.830 6.360 ;
        RECT 808.765 6.175 809.055 6.220 ;
        RECT 811.510 6.160 811.830 6.220 ;
        RECT 880.050 6.360 880.370 6.420 ;
        RECT 884.665 6.360 884.955 6.405 ;
        RECT 880.050 6.220 884.955 6.360 ;
        RECT 880.050 6.160 880.370 6.220 ;
        RECT 884.665 6.175 884.955 6.220 ;
        RECT 1270.590 6.360 1270.910 6.420 ;
        RECT 1282.550 6.360 1282.870 6.420 ;
        RECT 1270.590 6.220 1282.870 6.360 ;
        RECT 1270.590 6.160 1270.910 6.220 ;
        RECT 1282.550 6.160 1282.870 6.220 ;
        RECT 1353.850 6.020 1354.170 6.080 ;
        RECT 1399.390 6.020 1399.710 6.080 ;
        RECT 1353.850 5.880 1399.710 6.020 ;
        RECT 1353.850 5.820 1354.170 5.880 ;
        RECT 1399.390 5.820 1399.710 5.880 ;
        RECT 1453.225 6.020 1453.515 6.065 ;
        RECT 1454.145 6.020 1454.435 6.065 ;
        RECT 1453.225 5.880 1454.435 6.020 ;
        RECT 1453.225 5.835 1453.515 5.880 ;
        RECT 1454.145 5.835 1454.435 5.880 ;
        RECT 529.545 5.680 529.835 5.725 ;
        RECT 579.225 5.680 579.515 5.725 ;
        RECT 739.765 5.680 740.055 5.725 ;
        RECT 529.545 5.540 579.515 5.680 ;
        RECT 529.545 5.495 529.835 5.540 ;
        RECT 579.225 5.495 579.515 5.540 ;
        RECT 738.460 5.540 740.055 5.680 ;
        RECT 344.625 5.340 344.915 5.385 ;
        RECT 364.865 5.340 365.155 5.385 ;
        RECT 344.625 5.200 365.155 5.340 ;
        RECT 344.625 5.155 344.915 5.200 ;
        RECT 364.865 5.155 365.155 5.200 ;
        RECT 737.450 5.340 737.770 5.400 ;
        RECT 738.460 5.340 738.600 5.540 ;
        RECT 739.765 5.495 740.055 5.540 ;
        RECT 787.590 5.680 787.910 5.740 ;
        RECT 791.285 5.680 791.575 5.725 ;
        RECT 787.590 5.540 791.575 5.680 ;
        RECT 787.590 5.480 787.910 5.540 ;
        RECT 791.285 5.495 791.575 5.540 ;
        RECT 737.450 5.200 738.600 5.340 ;
        RECT 740.685 5.340 740.975 5.385 ;
        RECT 744.350 5.340 744.670 5.400 ;
        RECT 740.685 5.200 744.670 5.340 ;
        RECT 737.450 5.140 737.770 5.200 ;
        RECT 740.685 5.155 740.975 5.200 ;
        RECT 744.350 5.140 744.670 5.200 ;
        RECT 730.550 5.000 730.870 5.060 ;
        RECT 728.340 4.860 730.870 5.000 ;
        RECT 364.865 4.660 365.155 4.705 ;
        RECT 377.285 4.660 377.575 4.705 ;
        RECT 364.865 4.520 377.575 4.660 ;
        RECT 364.865 4.475 365.155 4.520 ;
        RECT 377.285 4.475 377.575 4.520 ;
        RECT 705.725 4.660 706.015 4.705 ;
        RECT 711.705 4.660 711.995 4.705 ;
        RECT 705.725 4.520 711.995 4.660 ;
        RECT 705.725 4.475 706.015 4.520 ;
        RECT 711.705 4.475 711.995 4.520 ;
        RECT 716.305 4.660 716.595 4.705 ;
        RECT 728.340 4.660 728.480 4.860 ;
        RECT 730.550 4.800 730.870 4.860 ;
        RECT 716.305 4.520 728.480 4.660 ;
        RECT 762.305 4.660 762.595 4.705 ;
        RECT 770.570 4.660 770.890 4.720 ;
        RECT 762.305 4.520 770.890 4.660 ;
        RECT 716.305 4.475 716.595 4.520 ;
        RECT 762.305 4.475 762.595 4.520 ;
        RECT 770.570 4.460 770.890 4.520 ;
        RECT 380.045 4.320 380.335 4.365 ;
        RECT 383.725 4.320 384.015 4.365 ;
        RECT 380.045 4.180 384.015 4.320 ;
        RECT 380.045 4.135 380.335 4.180 ;
        RECT 383.725 4.135 384.015 4.180 ;
        RECT 416.845 4.320 417.135 4.365 ;
        RECT 419.130 4.320 419.450 4.380 ;
        RECT 416.845 4.180 419.450 4.320 ;
        RECT 416.845 4.135 417.135 4.180 ;
        RECT 419.130 4.120 419.450 4.180 ;
        RECT 439.370 4.320 439.690 4.380 ;
        RECT 466.985 4.320 467.275 4.365 ;
        RECT 439.370 4.180 467.275 4.320 ;
        RECT 439.370 4.120 439.690 4.180 ;
        RECT 466.985 4.135 467.275 4.180 ;
        RECT 898.450 4.320 898.770 4.380 ;
        RECT 900.305 4.320 900.595 4.365 ;
        RECT 898.450 4.180 900.595 4.320 ;
        RECT 898.450 4.120 898.770 4.180 ;
        RECT 900.305 4.135 900.595 4.180 ;
        RECT 1431.130 4.320 1431.450 4.380 ;
        RECT 1437.125 4.320 1437.415 4.365 ;
        RECT 1431.130 4.180 1437.415 4.320 ;
        RECT 1431.130 4.120 1431.450 4.180 ;
        RECT 1437.125 4.135 1437.415 4.180 ;
        RECT 901.210 3.640 901.530 3.700 ;
        RECT 919.625 3.640 919.915 3.685 ;
        RECT 901.210 3.500 919.915 3.640 ;
        RECT 901.210 3.440 901.530 3.500 ;
        RECT 919.625 3.455 919.915 3.500 ;
        RECT 1158.825 3.640 1159.115 3.685 ;
        RECT 1158.825 3.500 1166.400 3.640 ;
        RECT 1158.825 3.455 1159.115 3.500 ;
        RECT 610.950 3.300 611.270 3.360 ;
        RECT 622.465 3.300 622.755 3.345 ;
        RECT 610.950 3.160 622.755 3.300 ;
        RECT 610.950 3.100 611.270 3.160 ;
        RECT 622.465 3.115 622.755 3.160 ;
        RECT 885.570 3.300 885.890 3.360 ;
        RECT 886.965 3.300 887.255 3.345 ;
        RECT 885.570 3.160 887.255 3.300 ;
        RECT 885.570 3.100 885.890 3.160 ;
        RECT 886.965 3.115 887.255 3.160 ;
        RECT 1022.205 3.300 1022.495 3.345 ;
        RECT 1038.750 3.300 1039.070 3.360 ;
        RECT 1022.205 3.160 1039.070 3.300 ;
        RECT 1166.260 3.300 1166.400 3.500 ;
        RECT 1259.550 3.300 1259.870 3.360 ;
        RECT 1166.260 3.160 1259.870 3.300 ;
        RECT 1022.205 3.115 1022.495 3.160 ;
        RECT 1038.750 3.100 1039.070 3.160 ;
        RECT 1259.550 3.100 1259.870 3.160 ;
        RECT 1088.890 2.620 1089.210 2.680 ;
        RECT 1089.365 2.620 1089.655 2.665 ;
        RECT 1088.890 2.480 1089.655 2.620 ;
        RECT 1088.890 2.420 1089.210 2.480 ;
        RECT 1089.365 2.435 1089.655 2.480 ;
        RECT 1314.750 2.280 1315.070 2.340 ;
        RECT 1324.410 2.280 1324.730 2.340 ;
        RECT 1314.750 2.140 1324.730 2.280 ;
        RECT 1314.750 2.080 1315.070 2.140 ;
        RECT 1324.410 2.080 1324.730 2.140 ;
        RECT 1401.690 2.280 1402.010 2.340 ;
        RECT 1407.670 2.280 1407.990 2.340 ;
        RECT 1401.690 2.140 1407.990 2.280 ;
        RECT 1401.690 2.080 1402.010 2.140 ;
        RECT 1407.670 2.080 1407.990 2.140 ;
        RECT 1427.910 2.280 1428.230 2.340 ;
        RECT 1428.370 2.280 1428.690 2.340 ;
        RECT 1427.910 2.140 1428.690 2.280 ;
        RECT 1427.910 2.080 1428.230 2.140 ;
        RECT 1428.370 2.080 1428.690 2.140 ;
        RECT 993.225 1.940 993.515 1.985 ;
        RECT 996.445 1.940 996.735 1.985 ;
        RECT 993.225 1.800 996.735 1.940 ;
        RECT 993.225 1.755 993.515 1.800 ;
        RECT 996.445 1.755 996.735 1.800 ;
        RECT 334.950 1.260 335.270 1.320 ;
        RECT 336.345 1.260 336.635 1.305 ;
        RECT 334.950 1.120 336.635 1.260 ;
        RECT 334.950 1.060 335.270 1.120 ;
        RECT 336.345 1.075 336.635 1.120 ;
        RECT 423.270 0.920 423.590 0.980 ;
        RECT 438.450 0.920 438.770 0.980 ;
        RECT 423.270 0.780 438.770 0.920 ;
        RECT 423.270 0.720 423.590 0.780 ;
        RECT 438.450 0.720 438.770 0.780 ;
      LAYER via ;
        RECT 641.340 8.540 641.600 8.800 ;
        RECT 691.940 8.200 692.200 8.460 ;
        RECT 847.420 8.540 847.680 8.800 ;
        RECT 871.340 8.540 871.600 8.800 ;
        RECT 876.400 8.540 876.660 8.800 ;
        RECT 1764.660 8.540 1764.920 8.800 ;
        RECT 1831.820 8.540 1832.080 8.800 ;
        RECT 1573.760 8.200 1574.020 8.460 ;
        RECT 1598.600 8.200 1598.860 8.460 ;
        RECT 893.420 7.860 893.680 8.120 ;
        RECT 1468.420 7.860 1468.680 8.120 ;
        RECT 801.420 7.520 801.680 7.780 ;
        RECT 610.060 6.840 610.320 7.100 ;
        RECT 846.960 7.180 847.220 7.440 ;
        RECT 857.540 7.180 857.800 7.440 ;
        RECT 1328.120 7.180 1328.380 7.440 ;
        RECT 1343.300 7.180 1343.560 7.440 ;
        RECT 1469.800 7.180 1470.060 7.440 ;
        RECT 1473.940 7.180 1474.200 7.440 ;
        RECT 811.540 6.160 811.800 6.420 ;
        RECT 880.080 6.160 880.340 6.420 ;
        RECT 1270.620 6.160 1270.880 6.420 ;
        RECT 1282.580 6.160 1282.840 6.420 ;
        RECT 1353.880 5.820 1354.140 6.080 ;
        RECT 1399.420 5.820 1399.680 6.080 ;
        RECT 737.480 5.140 737.740 5.400 ;
        RECT 787.620 5.480 787.880 5.740 ;
        RECT 744.380 5.140 744.640 5.400 ;
        RECT 730.580 4.800 730.840 5.060 ;
        RECT 770.600 4.460 770.860 4.720 ;
        RECT 419.160 4.120 419.420 4.380 ;
        RECT 439.400 4.120 439.660 4.380 ;
        RECT 898.480 4.120 898.740 4.380 ;
        RECT 1431.160 4.120 1431.420 4.380 ;
        RECT 901.240 3.440 901.500 3.700 ;
        RECT 610.980 3.100 611.240 3.360 ;
        RECT 885.600 3.100 885.860 3.360 ;
        RECT 1038.780 3.100 1039.040 3.360 ;
        RECT 1259.580 3.100 1259.840 3.360 ;
        RECT 1088.920 2.420 1089.180 2.680 ;
        RECT 1314.780 2.080 1315.040 2.340 ;
        RECT 1324.440 2.080 1324.700 2.340 ;
        RECT 1401.720 2.080 1401.980 2.340 ;
        RECT 1407.700 2.080 1407.960 2.340 ;
        RECT 1427.940 2.080 1428.200 2.340 ;
        RECT 1428.400 2.080 1428.660 2.340 ;
        RECT 334.980 1.060 335.240 1.320 ;
        RECT 423.300 0.720 423.560 0.980 ;
        RECT 438.480 0.720 438.740 0.980 ;
      LAYER met2 ;
        RECT 621.560 15.340 621.820 15.600 ;
        RECT 641.340 8.685 641.600 8.830 ;
        RECT 641.330 8.315 641.610 8.685 ;
        RECT 691.930 8.315 692.210 8.685 ;
        RECT 745.750 8.315 746.030 8.685 ;
        RECT 847.420 8.510 847.680 8.830 ;
        RECT 871.340 8.740 871.600 8.830 ;
        RECT 857.600 8.600 871.600 8.740 ;
        RECT 691.940 8.170 692.200 8.315 ;
        RECT 609.590 7.635 609.870 8.005 ;
        RECT 609.660 7.040 609.800 7.635 ;
        RECT 610.060 7.040 610.320 7.130 ;
        RECT 609.660 6.900 610.320 7.040 ;
        RECT 610.060 6.810 610.320 6.900 ;
        RECT 730.640 5.710 733.540 5.850 ;
        RECT 730.640 5.090 730.780 5.710 ;
        RECT 733.400 5.340 733.540 5.710 ;
        RECT 737.480 5.340 737.740 5.430 ;
        RECT 733.400 5.200 737.740 5.340 ;
        RECT 737.480 5.110 737.740 5.200 ;
        RECT 744.380 5.340 744.640 5.430 ;
        RECT 745.820 5.340 745.960 8.315 ;
        RECT 801.410 7.635 801.690 8.005 ;
        RECT 801.420 7.490 801.680 7.635 ;
        RECT 811.600 7.580 819.100 7.720 ;
        RECT 770.590 6.275 770.870 6.645 ;
        RECT 787.610 6.275 787.890 6.645 ;
        RECT 811.600 6.450 811.740 7.580 ;
        RECT 818.960 6.645 819.100 7.580 ;
        RECT 844.720 7.580 846.700 7.720 ;
        RECT 844.720 6.645 844.860 7.580 ;
        RECT 744.380 5.200 745.960 5.340 ;
        RECT 744.380 5.110 744.640 5.200 ;
        RECT 730.580 4.770 730.840 5.090 ;
        RECT 770.660 4.750 770.800 6.275 ;
        RECT 787.680 5.770 787.820 6.275 ;
        RECT 811.540 6.130 811.800 6.450 ;
        RECT 818.890 6.275 819.170 6.645 ;
        RECT 844.650 6.275 844.930 6.645 ;
        RECT 787.620 5.450 787.880 5.770 ;
        RECT 846.560 5.340 846.700 7.580 ;
        RECT 846.960 7.150 847.220 7.470 ;
        RECT 847.480 7.210 847.620 8.510 ;
        RECT 857.600 7.470 857.740 8.600 ;
        RECT 871.340 8.510 871.600 8.600 ;
        RECT 876.400 8.740 876.660 8.830 ;
        RECT 876.400 8.600 877.060 8.740 ;
        RECT 876.400 8.510 876.660 8.600 ;
        RECT 876.920 7.720 877.060 8.600 ;
        RECT 883.230 7.720 883.510 9.000 ;
        RECT 954.590 8.315 954.870 8.685 ;
        RECT 961.030 8.570 961.310 8.685 ;
        RECT 961.030 8.430 961.700 8.570 ;
        RECT 961.030 8.315 961.310 8.430 ;
        RECT 893.420 7.830 893.680 8.150 ;
        RECT 876.920 7.580 886.260 7.720 ;
        RECT 847.020 5.965 847.160 7.150 ;
        RECT 847.480 7.070 854.520 7.210 ;
        RECT 857.540 7.150 857.800 7.470 ;
        RECT 853.850 6.530 854.130 6.645 ;
        RECT 852.540 6.390 854.130 6.530 ;
        RECT 852.540 5.965 852.680 6.390 ;
        RECT 853.850 6.275 854.130 6.390 ;
        RECT 846.950 5.595 847.230 5.965 ;
        RECT 847.870 5.850 848.150 5.965 ;
        RECT 847.480 5.710 848.150 5.850 ;
        RECT 847.480 5.340 847.620 5.710 ;
        RECT 847.870 5.595 848.150 5.710 ;
        RECT 852.470 5.595 852.750 5.965 ;
        RECT 846.560 5.200 847.620 5.340 ;
        RECT 854.380 5.170 854.520 7.070 ;
        RECT 869.030 6.360 869.310 6.645 ;
        RECT 880.080 6.360 880.340 6.450 ;
        RECT 869.030 6.275 880.340 6.360 ;
        RECT 869.100 6.220 880.340 6.275 ;
        RECT 880.080 6.130 880.340 6.220 ;
        RECT 866.270 5.850 866.550 5.965 ;
        RECT 881.450 5.850 881.730 5.965 ;
        RECT 866.270 5.710 881.730 5.850 ;
        RECT 866.270 5.595 866.550 5.710 ;
        RECT 881.450 5.595 881.730 5.710 ;
        RECT 883.230 5.170 883.510 7.580 ;
        RECT 885.590 5.595 885.870 5.965 ;
        RECT 854.380 5.030 883.510 5.170 ;
        RECT 883.230 5.000 883.510 5.030 ;
        RECT 419.220 4.410 421.200 4.490 ;
        RECT 770.600 4.430 770.860 4.750 ;
        RECT 419.160 4.350 421.200 4.410 ;
        RECT 419.160 4.090 419.420 4.350 ;
        RECT 421.060 3.130 421.200 4.350 ;
        RECT 439.400 4.090 439.660 4.410 ;
        RECT 252.700 2.990 253.760 3.130 ;
        RECT 252.700 2.400 252.840 2.990 ;
        RECT 253.620 2.565 253.760 2.990 ;
        RECT 288.120 2.990 289.180 3.130 ;
        RECT 421.060 2.990 423.500 3.130 ;
        RECT 252.490 -4.800 253.050 2.400 ;
        RECT 253.550 2.195 253.830 2.565 ;
        RECT 288.120 2.400 288.260 2.990 ;
        RECT 287.910 -4.800 288.470 2.400 ;
        RECT 289.040 1.205 289.180 2.990 ;
        RECT 333.660 1.630 335.180 1.770 ;
        RECT 333.660 1.205 333.800 1.630 ;
        RECT 335.040 1.350 335.180 1.630 ;
        RECT 288.970 0.835 289.250 1.205 ;
        RECT 333.590 0.835 333.870 1.205 ;
        RECT 334.980 1.030 335.240 1.350 ;
        RECT 423.360 1.010 423.500 2.990 ;
        RECT 439.460 1.090 439.600 4.090 ;
        RECT 885.660 3.390 885.800 5.595 ;
        RECT 610.980 3.300 611.240 3.390 ;
        RECT 609.200 3.160 611.240 3.300 ;
        RECT 609.200 2.400 609.340 3.160 ;
        RECT 610.980 3.070 611.240 3.160 ;
        RECT 885.600 3.070 885.860 3.390 ;
        RECT 886.120 3.130 886.260 7.580 ;
        RECT 893.480 7.325 893.620 7.830 ;
        RECT 954.660 7.325 954.800 8.315 ;
        RECT 961.560 7.890 961.700 8.430 ;
        RECT 978.450 7.890 978.730 9.000 ;
        RECT 961.560 7.750 978.730 7.890 ;
        RECT 893.410 6.955 893.690 7.325 ;
        RECT 918.710 7.040 918.990 7.325 ;
        RECT 921.930 7.040 922.210 7.325 ;
        RECT 918.710 6.955 922.210 7.040 ;
        RECT 954.590 6.955 954.870 7.325 ;
        RECT 918.780 6.900 922.140 6.955 ;
        RECT 898.470 6.275 898.750 6.645 ;
        RECT 901.230 6.275 901.510 6.645 ;
        RECT 898.540 4.410 898.680 6.275 ;
        RECT 898.480 4.090 898.740 4.410 ;
        RECT 901.300 3.730 901.440 6.275 ;
        RECT 978.450 5.000 978.730 7.750 ;
        RECT 1128.470 7.635 1128.750 8.005 ;
        RECT 1128.540 6.530 1128.680 7.635 ;
        RECT 1128.930 6.530 1129.210 6.645 ;
        RECT 1128.540 6.390 1129.210 6.530 ;
        RECT 1128.930 6.275 1129.210 6.390 ;
        RECT 1263.190 5.170 1263.470 9.000 ;
        RECT 1764.660 8.510 1764.920 8.830 ;
        RECT 1831.820 8.570 1832.080 8.830 ;
        RECT 1833.590 8.570 1833.870 9.000 ;
        RECT 1831.820 8.510 1833.870 8.570 ;
        RECT 1475.380 8.260 1478.740 8.400 ;
        RECT 1468.420 8.060 1468.680 8.150 ;
        RECT 1468.420 7.920 1470.000 8.060 ;
        RECT 1343.820 7.750 1353.620 7.890 ;
        RECT 1468.420 7.830 1468.680 7.920 ;
        RECT 1270.150 7.210 1270.430 7.325 ;
        RECT 1270.150 7.070 1270.820 7.210 ;
        RECT 1328.120 7.150 1328.380 7.470 ;
        RECT 1343.300 7.380 1343.560 7.470 ;
        RECT 1343.820 7.380 1343.960 7.750 ;
        RECT 1343.300 7.240 1343.960 7.380 ;
        RECT 1353.480 7.380 1353.620 7.750 ;
        RECT 1469.860 7.470 1470.000 7.920 ;
        RECT 1475.380 7.890 1475.520 8.260 ;
        RECT 1474.000 7.750 1475.520 7.890 ;
        RECT 1478.600 7.890 1478.740 8.260 ;
        RECT 1573.760 8.170 1574.020 8.490 ;
        RECT 1598.600 8.170 1598.860 8.490 ;
        RECT 1478.990 7.890 1479.270 8.005 ;
        RECT 1478.600 7.750 1479.270 7.890 ;
        RECT 1474.000 7.470 1474.140 7.750 ;
        RECT 1478.990 7.635 1479.270 7.750 ;
        RECT 1353.480 7.240 1354.080 7.380 ;
        RECT 1343.300 7.150 1343.560 7.240 ;
        RECT 1270.150 6.955 1270.430 7.070 ;
        RECT 1270.680 6.450 1270.820 7.070 ;
        RECT 1270.620 6.130 1270.880 6.450 ;
        RECT 1282.570 6.275 1282.850 6.645 ;
        RECT 1306.030 6.275 1306.310 6.645 ;
        RECT 1282.580 6.130 1282.840 6.275 ;
        RECT 1306.100 6.020 1306.240 6.275 ;
        RECT 1306.100 5.880 1309.460 6.020 ;
        RECT 1260.560 5.030 1263.470 5.170 ;
        RECT 1041.600 4.350 1047.260 4.490 ;
        RECT 901.240 3.410 901.500 3.730 ;
        RECT 886.970 3.130 887.250 3.245 ;
        RECT 886.120 2.990 887.250 3.130 ;
        RECT 1038.780 3.070 1039.040 3.390 ;
        RECT 886.970 2.875 887.250 2.990 ;
        RECT 1038.840 2.450 1038.980 3.070 ;
        RECT 1041.600 2.450 1041.740 4.350 ;
        RECT 1047.120 3.980 1047.260 4.350 ;
        RECT 1047.120 3.840 1057.840 3.980 ;
        RECT 438.540 1.010 439.600 1.090 ;
        RECT 423.300 0.690 423.560 1.010 ;
        RECT 438.480 0.950 439.600 1.010 ;
        RECT 438.480 0.690 438.740 0.950 ;
        RECT 608.990 -4.800 609.550 2.400 ;
        RECT 1038.840 2.310 1041.740 2.450 ;
        RECT 1057.700 1.770 1057.840 3.840 ;
        RECT 1076.030 3.130 1076.310 3.245 ;
        RECT 1060.460 2.990 1068.420 3.130 ;
        RECT 1060.460 1.770 1060.600 2.990 ;
        RECT 1068.280 2.620 1068.420 2.990 ;
        RECT 1071.040 2.990 1074.400 3.130 ;
        RECT 1071.040 2.620 1071.180 2.990 ;
        RECT 1068.280 2.480 1071.180 2.620 ;
        RECT 1074.260 2.620 1074.400 2.990 ;
        RECT 1075.640 2.990 1076.310 3.130 ;
        RECT 1075.640 2.620 1075.780 2.990 ;
        RECT 1076.030 2.875 1076.310 2.990 ;
        RECT 1088.910 2.875 1089.190 3.245 ;
        RECT 1259.580 3.070 1259.840 3.390 ;
        RECT 1088.980 2.710 1089.120 2.875 ;
        RECT 1074.260 2.480 1075.780 2.620 ;
        RECT 1088.920 2.390 1089.180 2.710 ;
        RECT 1259.640 2.620 1259.780 3.070 ;
        RECT 1260.560 2.620 1260.700 5.030 ;
        RECT 1263.190 5.000 1263.470 5.030 ;
        RECT 1309.320 3.925 1309.460 5.880 ;
        RECT 1309.250 3.555 1309.530 3.925 ;
        RECT 1313.390 3.555 1313.670 3.925 ;
        RECT 1259.640 2.480 1260.700 2.620 ;
        RECT 1057.700 1.630 1060.600 1.770 ;
        RECT 1313.460 1.770 1313.600 3.555 ;
        RECT 1314.780 2.050 1315.040 2.370 ;
        RECT 1324.440 2.050 1324.700 2.370 ;
        RECT 1314.840 1.770 1314.980 2.050 ;
        RECT 1313.460 1.630 1314.980 1.770 ;
        RECT 1324.500 1.770 1324.640 2.050 ;
        RECT 1328.180 1.940 1328.320 7.150 ;
        RECT 1353.940 6.110 1354.080 7.240 ;
        RECT 1469.800 7.150 1470.060 7.470 ;
        RECT 1473.940 7.150 1474.200 7.470 ;
        RECT 1353.880 5.790 1354.140 6.110 ;
        RECT 1399.420 5.850 1399.680 6.110 ;
        RECT 1399.420 5.790 1400.080 5.850 ;
        RECT 1399.480 5.710 1400.080 5.790 ;
        RECT 1399.940 3.810 1400.080 5.710 ;
        RECT 1573.820 4.605 1573.960 8.170 ;
        RECT 1598.660 8.005 1598.800 8.170 ;
        RECT 1764.720 8.005 1764.860 8.510 ;
        RECT 1831.880 8.430 1833.870 8.510 ;
        RECT 1598.590 7.635 1598.870 8.005 ;
        RECT 1764.650 7.635 1764.930 8.005 ;
        RECT 1833.590 5.000 1833.870 8.430 ;
        RECT 1431.160 4.320 1431.420 4.410 ;
        RECT 1429.380 4.180 1431.420 4.320 ;
        RECT 1573.750 4.235 1574.030 4.605 ;
        RECT 1399.940 3.670 1401.000 3.810 ;
        RECT 1400.860 3.300 1401.000 3.670 ;
        RECT 1410.450 3.555 1410.730 3.925 ;
        RECT 1426.550 3.555 1426.830 3.925 ;
        RECT 1400.860 3.160 1401.920 3.300 ;
        RECT 1401.780 2.370 1401.920 3.160 ;
        RECT 1410.520 2.450 1410.660 3.555 ;
        RECT 1426.620 3.130 1426.760 3.555 ;
        RECT 1429.380 3.130 1429.520 4.180 ;
        RECT 1431.160 4.090 1431.420 4.180 ;
        RECT 1426.620 2.990 1428.140 3.130 ;
        RECT 1407.760 2.370 1410.660 2.450 ;
        RECT 1428.000 2.370 1428.140 2.990 ;
        RECT 1428.460 2.990 1429.520 3.130 ;
        RECT 1428.460 2.370 1428.600 2.990 ;
        RECT 1401.720 2.050 1401.980 2.370 ;
        RECT 1407.700 2.310 1410.660 2.370 ;
        RECT 1407.700 2.050 1407.960 2.310 ;
        RECT 1427.940 2.050 1428.200 2.370 ;
        RECT 1428.400 2.050 1428.660 2.370 ;
        RECT 1325.420 1.800 1328.320 1.940 ;
        RECT 1325.420 1.770 1325.560 1.800 ;
        RECT 1324.500 1.630 1325.560 1.770 ;
      LAYER via2 ;
        RECT 641.330 8.360 641.610 8.640 ;
        RECT 691.930 8.360 692.210 8.640 ;
        RECT 745.750 8.360 746.030 8.640 ;
        RECT 609.590 7.680 609.870 7.960 ;
        RECT 801.410 7.680 801.690 7.960 ;
        RECT 770.590 6.320 770.870 6.600 ;
        RECT 787.610 6.320 787.890 6.600 ;
        RECT 818.890 6.320 819.170 6.600 ;
        RECT 844.650 6.320 844.930 6.600 ;
        RECT 954.590 8.360 954.870 8.640 ;
        RECT 961.030 8.360 961.310 8.640 ;
        RECT 853.850 6.320 854.130 6.600 ;
        RECT 846.950 5.640 847.230 5.920 ;
        RECT 847.870 5.640 848.150 5.920 ;
        RECT 852.470 5.640 852.750 5.920 ;
        RECT 869.030 6.320 869.310 6.600 ;
        RECT 866.270 5.640 866.550 5.920 ;
        RECT 881.450 5.640 881.730 5.920 ;
        RECT 885.590 5.640 885.870 5.920 ;
        RECT 253.550 2.240 253.830 2.520 ;
        RECT 288.970 0.880 289.250 1.160 ;
        RECT 333.590 0.880 333.870 1.160 ;
        RECT 893.410 7.000 893.690 7.280 ;
        RECT 918.710 7.000 918.990 7.280 ;
        RECT 921.930 7.000 922.210 7.280 ;
        RECT 954.590 7.000 954.870 7.280 ;
        RECT 898.470 6.320 898.750 6.600 ;
        RECT 901.230 6.320 901.510 6.600 ;
        RECT 1128.470 7.680 1128.750 7.960 ;
        RECT 1128.930 6.320 1129.210 6.600 ;
        RECT 1270.150 7.000 1270.430 7.280 ;
        RECT 1478.990 7.680 1479.270 7.960 ;
        RECT 1282.570 6.320 1282.850 6.600 ;
        RECT 1306.030 6.320 1306.310 6.600 ;
        RECT 886.970 2.920 887.250 3.200 ;
        RECT 1076.030 2.920 1076.310 3.200 ;
        RECT 1088.910 2.920 1089.190 3.200 ;
        RECT 1309.250 3.600 1309.530 3.880 ;
        RECT 1313.390 3.600 1313.670 3.880 ;
        RECT 1598.590 7.680 1598.870 7.960 ;
        RECT 1764.650 7.680 1764.930 7.960 ;
        RECT 1573.750 4.280 1574.030 4.560 ;
        RECT 1410.450 3.600 1410.730 3.880 ;
        RECT 1426.550 3.600 1426.830 3.880 ;
      LAYER met3 ;
        RECT 376.550 8.650 376.930 8.660 ;
        RECT 369.230 8.350 376.930 8.650 ;
        RECT 366.430 7.970 366.810 7.980 ;
        RECT 369.230 7.970 369.530 8.350 ;
        RECT 376.550 8.340 376.930 8.350 ;
        RECT 380.230 8.650 380.610 8.660 ;
        RECT 383.910 8.650 384.290 8.660 ;
        RECT 380.230 8.350 384.290 8.650 ;
        RECT 380.230 8.340 380.610 8.350 ;
        RECT 383.910 8.340 384.290 8.350 ;
        RECT 477.750 8.650 478.130 8.660 ;
        RECT 501.670 8.650 502.050 8.660 ;
        RECT 477.750 8.350 502.050 8.650 ;
        RECT 477.750 8.340 478.130 8.350 ;
        RECT 501.670 8.340 502.050 8.350 ;
        RECT 641.305 8.650 641.635 8.665 ;
        RECT 644.270 8.650 644.650 8.660 ;
        RECT 641.305 8.350 644.650 8.650 ;
        RECT 641.305 8.335 641.635 8.350 ;
        RECT 644.270 8.340 644.650 8.350 ;
        RECT 681.990 8.650 682.370 8.660 ;
        RECT 691.905 8.650 692.235 8.665 ;
        RECT 681.990 8.350 692.235 8.650 ;
        RECT 681.990 8.340 682.370 8.350 ;
        RECT 691.905 8.335 692.235 8.350 ;
        RECT 745.725 8.650 746.055 8.665 ;
        RECT 761.110 8.650 761.490 8.660 ;
        RECT 745.725 8.350 761.490 8.650 ;
        RECT 745.725 8.335 746.055 8.350 ;
        RECT 761.110 8.340 761.490 8.350 ;
        RECT 834.710 8.650 835.090 8.660 ;
        RECT 844.830 8.650 845.210 8.660 ;
        RECT 834.710 8.350 845.210 8.650 ;
        RECT 834.710 8.340 835.090 8.350 ;
        RECT 844.830 8.340 845.210 8.350 ;
        RECT 954.565 8.650 954.895 8.665 ;
        RECT 961.005 8.650 961.335 8.665 ;
        RECT 954.565 8.350 961.335 8.650 ;
        RECT 954.565 8.335 954.895 8.350 ;
        RECT 961.005 8.335 961.335 8.350 ;
        RECT 609.565 7.970 609.895 7.985 ;
        RECT 366.430 7.670 369.530 7.970 ;
        RECT 603.830 7.670 609.895 7.970 ;
        RECT 366.430 7.660 366.810 7.670 ;
        RECT 603.830 7.300 604.130 7.670 ;
        RECT 609.565 7.655 609.895 7.670 ;
        RECT 789.630 7.970 790.010 7.980 ;
        RECT 800.670 7.970 801.050 7.980 ;
        RECT 789.630 7.670 801.050 7.970 ;
        RECT 789.630 7.660 790.010 7.670 ;
        RECT 800.670 7.660 801.050 7.670 ;
        RECT 801.385 7.970 801.715 7.985 ;
        RECT 805.270 7.970 805.650 7.980 ;
        RECT 801.385 7.670 805.650 7.970 ;
        RECT 801.385 7.655 801.715 7.670 ;
        RECT 805.270 7.660 805.650 7.670 ;
        RECT 1124.510 7.970 1124.890 7.980 ;
        RECT 1128.445 7.970 1128.775 7.985 ;
        RECT 1124.510 7.670 1128.775 7.970 ;
        RECT 1124.510 7.660 1124.890 7.670 ;
        RECT 1128.445 7.655 1128.775 7.670 ;
        RECT 1266.190 7.970 1266.570 7.980 ;
        RECT 1478.965 7.970 1479.295 7.985 ;
        RECT 1480.550 7.970 1480.930 7.980 ;
        RECT 1266.190 7.670 1268.370 7.970 ;
        RECT 1266.190 7.660 1266.570 7.670 ;
        RECT 603.790 6.980 604.170 7.300 ;
        RECT 893.385 7.290 893.715 7.305 ;
        RECT 918.685 7.290 919.015 7.305 ;
        RECT 893.385 6.990 919.015 7.290 ;
        RECT 893.385 6.975 893.715 6.990 ;
        RECT 918.685 6.975 919.015 6.990 ;
        RECT 921.905 7.290 922.235 7.305 ;
        RECT 954.565 7.290 954.895 7.305 ;
        RECT 921.905 6.990 954.895 7.290 ;
        RECT 1268.070 7.290 1268.370 7.670 ;
        RECT 1478.965 7.670 1480.930 7.970 ;
        RECT 1478.965 7.655 1479.295 7.670 ;
        RECT 1480.550 7.660 1480.930 7.670 ;
        RECT 1598.565 7.970 1598.895 7.985 ;
        RECT 1764.625 7.970 1764.955 7.985 ;
        RECT 1598.565 7.670 1764.955 7.970 ;
        RECT 1598.565 7.655 1598.895 7.670 ;
        RECT 1764.625 7.655 1764.955 7.670 ;
        RECT 1270.125 7.290 1270.455 7.305 ;
        RECT 1268.070 6.990 1270.455 7.290 ;
        RECT 921.905 6.975 922.235 6.990 ;
        RECT 954.565 6.975 954.895 6.990 ;
        RECT 1270.125 6.975 1270.455 6.990 ;
        RECT 770.565 6.610 770.895 6.625 ;
        RECT 787.585 6.610 787.915 6.625 ;
        RECT 770.565 6.310 787.915 6.610 ;
        RECT 770.565 6.295 770.895 6.310 ;
        RECT 787.585 6.295 787.915 6.310 ;
        RECT 818.865 6.610 819.195 6.625 ;
        RECT 844.625 6.610 844.955 6.625 ;
        RECT 818.865 6.310 844.955 6.610 ;
        RECT 818.865 6.295 819.195 6.310 ;
        RECT 844.625 6.295 844.955 6.310 ;
        RECT 850.350 6.610 850.730 6.620 ;
        RECT 853.825 6.610 854.155 6.625 ;
        RECT 869.005 6.610 869.335 6.625 ;
        RECT 850.350 6.310 853.450 6.610 ;
        RECT 850.350 6.300 850.730 6.310 ;
        RECT 558.940 5.930 559.320 5.940 ;
        RECT 562.390 5.930 562.770 5.940 ;
        RECT 558.940 5.630 562.770 5.930 ;
        RECT 558.940 5.620 559.320 5.630 ;
        RECT 562.390 5.620 562.770 5.630 ;
        RECT 843.910 5.930 844.290 5.940 ;
        RECT 846.925 5.930 847.255 5.945 ;
        RECT 843.910 5.630 847.255 5.930 ;
        RECT 843.910 5.620 844.290 5.630 ;
        RECT 846.925 5.615 847.255 5.630 ;
        RECT 847.845 5.930 848.175 5.945 ;
        RECT 852.445 5.930 852.775 5.945 ;
        RECT 847.845 5.630 852.775 5.930 ;
        RECT 853.150 5.930 853.450 6.310 ;
        RECT 853.825 6.310 869.335 6.610 ;
        RECT 853.825 6.295 854.155 6.310 ;
        RECT 869.005 6.295 869.335 6.310 ;
        RECT 898.445 6.610 898.775 6.625 ;
        RECT 901.205 6.610 901.535 6.625 ;
        RECT 898.445 6.310 901.535 6.610 ;
        RECT 898.445 6.295 898.775 6.310 ;
        RECT 901.205 6.295 901.535 6.310 ;
        RECT 1128.905 6.610 1129.235 6.625 ;
        RECT 1135.550 6.610 1135.930 6.620 ;
        RECT 1128.905 6.310 1135.930 6.610 ;
        RECT 1128.905 6.295 1129.235 6.310 ;
        RECT 1135.550 6.300 1135.930 6.310 ;
        RECT 1282.545 6.610 1282.875 6.625 ;
        RECT 1306.005 6.610 1306.335 6.625 ;
        RECT 1282.545 6.310 1306.335 6.610 ;
        RECT 1282.545 6.295 1282.875 6.310 ;
        RECT 1306.005 6.295 1306.335 6.310 ;
        RECT 866.245 5.930 866.575 5.945 ;
        RECT 853.150 5.630 866.575 5.930 ;
        RECT 847.845 5.615 848.175 5.630 ;
        RECT 852.445 5.615 852.775 5.630 ;
        RECT 866.245 5.615 866.575 5.630 ;
        RECT 881.425 5.930 881.755 5.945 ;
        RECT 885.565 5.930 885.895 5.945 ;
        RECT 881.425 5.630 885.895 5.930 ;
        RECT 881.425 5.615 881.755 5.630 ;
        RECT 885.565 5.615 885.895 5.630 ;
        RECT 922.110 5.250 922.490 5.260 ;
        RECT 948.790 5.250 949.170 5.260 ;
        RECT 922.110 4.950 949.170 5.250 ;
        RECT 922.110 4.940 922.490 4.950 ;
        RECT 948.790 4.940 949.170 4.950 ;
        RECT 1549.550 4.570 1549.930 4.580 ;
        RECT 1573.725 4.570 1574.055 4.585 ;
        RECT 1549.550 4.270 1574.055 4.570 ;
        RECT 1549.550 4.260 1549.930 4.270 ;
        RECT 1573.725 4.255 1574.055 4.270 ;
        RECT 1309.225 3.890 1309.555 3.905 ;
        RECT 1313.365 3.890 1313.695 3.905 ;
        RECT 1309.225 3.590 1313.695 3.890 ;
        RECT 1309.225 3.575 1309.555 3.590 ;
        RECT 1313.365 3.575 1313.695 3.590 ;
        RECT 1410.425 3.890 1410.755 3.905 ;
        RECT 1426.525 3.890 1426.855 3.905 ;
        RECT 1410.425 3.590 1426.855 3.890 ;
        RECT 1410.425 3.575 1410.755 3.590 ;
        RECT 1426.525 3.575 1426.855 3.590 ;
        RECT 886.945 3.210 887.275 3.225 ;
        RECT 888.990 3.210 889.370 3.220 ;
        RECT 886.945 2.910 889.370 3.210 ;
        RECT 886.945 2.895 887.275 2.910 ;
        RECT 888.990 2.900 889.370 2.910 ;
        RECT 1039.870 3.210 1040.250 3.220 ;
        RECT 1051.830 3.210 1052.210 3.220 ;
        RECT 1039.870 2.910 1052.210 3.210 ;
        RECT 1039.870 2.900 1040.250 2.910 ;
        RECT 1051.830 2.900 1052.210 2.910 ;
        RECT 1076.005 3.210 1076.335 3.225 ;
        RECT 1088.885 3.210 1089.215 3.225 ;
        RECT 1076.005 2.910 1089.215 3.210 ;
        RECT 1076.005 2.895 1076.335 2.910 ;
        RECT 1088.885 2.895 1089.215 2.910 ;
        RECT 253.525 2.530 253.855 2.545 ;
        RECT 957.070 2.530 957.450 2.540 ;
        RECT 985.590 2.530 985.970 2.540 ;
        RECT 253.525 2.230 326.290 2.530 ;
        RECT 253.525 2.215 253.855 2.230 ;
        RECT 288.945 1.170 289.275 1.185 ;
        RECT 305.710 1.170 306.090 1.180 ;
        RECT 288.945 0.870 306.090 1.170 ;
        RECT 325.990 1.170 326.290 2.230 ;
        RECT 957.070 2.230 985.970 2.530 ;
        RECT 957.070 2.220 957.450 2.230 ;
        RECT 985.590 2.220 985.970 2.230 ;
        RECT 333.565 1.170 333.895 1.185 ;
        RECT 325.990 0.870 333.895 1.170 ;
        RECT 288.945 0.855 289.275 0.870 ;
        RECT 305.710 0.860 306.090 0.870 ;
        RECT 333.565 0.855 333.895 0.870 ;
      LAYER via3 ;
        RECT 366.460 7.660 366.780 7.980 ;
        RECT 376.580 8.340 376.900 8.660 ;
        RECT 380.260 8.340 380.580 8.660 ;
        RECT 383.940 8.340 384.260 8.660 ;
        RECT 477.780 8.340 478.100 8.660 ;
        RECT 501.700 8.340 502.020 8.660 ;
        RECT 644.300 8.340 644.620 8.660 ;
        RECT 682.020 8.340 682.340 8.660 ;
        RECT 761.140 8.340 761.460 8.660 ;
        RECT 834.740 8.340 835.060 8.660 ;
        RECT 844.860 8.340 845.180 8.660 ;
        RECT 789.660 7.660 789.980 7.980 ;
        RECT 800.700 7.660 801.020 7.980 ;
        RECT 805.300 7.660 805.620 7.980 ;
        RECT 1124.540 7.660 1124.860 7.980 ;
        RECT 1266.220 7.660 1266.540 7.980 ;
        RECT 603.820 6.980 604.140 7.300 ;
        RECT 1480.580 7.660 1480.900 7.980 ;
        RECT 850.380 6.300 850.700 6.620 ;
        RECT 558.970 5.620 559.290 5.940 ;
        RECT 562.420 5.620 562.740 5.940 ;
        RECT 843.940 5.620 844.260 5.940 ;
        RECT 1135.580 6.300 1135.900 6.620 ;
        RECT 922.140 4.940 922.460 5.260 ;
        RECT 948.820 4.940 949.140 5.260 ;
        RECT 1549.580 4.260 1549.900 4.580 ;
        RECT 889.020 2.900 889.340 3.220 ;
        RECT 1039.900 2.900 1040.220 3.220 ;
        RECT 1051.860 2.900 1052.180 3.220 ;
        RECT 305.740 0.860 306.060 1.180 ;
        RECT 957.100 2.220 957.420 2.540 ;
        RECT 985.620 2.220 985.940 2.540 ;
      LAYER met4 ;
        RECT 392.710 14.710 393.890 15.890 ;
        RECT 473.670 14.710 474.850 15.890 ;
        RECT 1143.430 14.710 1144.610 15.890 ;
        RECT 1266.710 14.710 1267.890 15.890 ;
        RECT 325.990 11.750 339.170 12.050 ;
        RECT 325.990 5.930 326.290 11.750 ;
        RECT 338.870 9.330 339.170 11.750 ;
        RECT 383.950 11.750 387.930 12.050 ;
        RECT 338.870 9.030 366.770 9.330 ;
        RECT 366.470 7.985 366.770 9.030 ;
        RECT 383.950 8.665 384.250 11.750 ;
        RECT 387.630 9.330 387.930 11.750 ;
        RECT 393.150 9.330 393.450 14.710 ;
        RECT 474.110 12.050 474.410 14.710 ;
        RECT 474.110 11.750 476.250 12.050 ;
        RECT 387.630 9.030 393.450 9.330 ;
        RECT 376.575 8.650 376.905 8.665 ;
        RECT 380.255 8.650 380.585 8.665 ;
        RECT 376.575 8.350 380.585 8.650 ;
        RECT 376.575 8.335 376.905 8.350 ;
        RECT 380.255 8.335 380.585 8.350 ;
        RECT 383.935 8.335 384.265 8.665 ;
        RECT 366.455 7.655 366.785 7.985 ;
        RECT 475.950 7.970 476.250 11.750 ;
        RECT 477.775 8.335 478.105 8.665 ;
        RECT 501.695 8.650 502.025 8.665 ;
        RECT 644.295 8.650 644.625 8.665 ;
        RECT 501.695 8.350 513.050 8.650 ;
        RECT 501.695 8.335 502.025 8.350 ;
        RECT 477.790 7.970 478.090 8.335 ;
        RECT 475.950 7.670 478.090 7.970 ;
        RECT 512.750 6.610 513.050 8.350 ;
        RECT 644.295 8.350 669.450 8.650 ;
        RECT 644.295 8.335 644.625 8.350 ;
        RECT 603.815 7.290 604.145 7.305 ;
        RECT 515.510 6.990 546.170 7.290 ;
        RECT 515.510 6.610 515.810 6.990 ;
        RECT 512.750 6.310 515.810 6.610 ;
        RECT 325.070 5.630 326.290 5.930 ;
        RECT 325.070 1.850 325.370 5.630 ;
        RECT 545.870 5.250 546.170 6.990 ;
        RECT 562.430 6.990 604.145 7.290 ;
        RECT 562.430 5.945 562.730 6.990 ;
        RECT 603.815 6.975 604.145 6.990 ;
        RECT 558.965 5.930 559.295 5.945 ;
        RECT 558.750 5.615 559.295 5.930 ;
        RECT 562.415 5.615 562.745 5.945 ;
        RECT 669.150 5.930 669.450 8.350 ;
        RECT 682.015 8.335 682.345 8.665 ;
        RECT 761.135 8.650 761.465 8.665 ;
        RECT 834.735 8.650 835.065 8.665 ;
        RECT 761.135 8.350 762.370 8.650 ;
        RECT 761.135 8.335 761.465 8.350 ;
        RECT 682.030 5.930 682.330 8.335 ;
        RECT 762.070 7.290 762.370 8.350 ;
        RECT 800.710 8.350 835.065 8.650 ;
        RECT 800.710 7.985 801.010 8.350 ;
        RECT 834.735 8.335 835.065 8.350 ;
        RECT 844.855 8.335 845.185 8.665 ;
        RECT 1143.870 8.650 1144.170 14.710 ;
        RECT 1267.150 12.050 1267.450 14.710 ;
        RECT 1057.390 8.350 1079.770 8.650 ;
        RECT 789.655 7.970 789.985 7.985 ;
        RECT 775.870 7.670 789.985 7.970 ;
        RECT 775.870 7.290 776.170 7.670 ;
        RECT 789.655 7.655 789.985 7.670 ;
        RECT 800.695 7.655 801.025 7.985 ;
        RECT 805.295 7.970 805.625 7.985 ;
        RECT 805.295 7.670 833.210 7.970 ;
        RECT 805.295 7.655 805.625 7.670 ;
        RECT 762.070 6.990 776.170 7.290 ;
        RECT 669.150 5.630 682.330 5.930 ;
        RECT 832.910 5.930 833.210 7.670 ;
        RECT 843.935 5.930 844.265 5.945 ;
        RECT 832.910 5.630 844.265 5.930 ;
        RECT 844.870 5.930 845.170 8.335 ;
        RECT 850.375 6.295 850.705 6.625 ;
        RECT 1057.390 6.610 1057.690 8.350 ;
        RECT 1079.470 7.970 1079.770 8.350 ;
        RECT 1084.990 8.350 1093.570 8.650 ;
        RECT 1084.990 7.970 1085.290 8.350 ;
        RECT 1079.470 7.670 1085.290 7.970 ;
        RECT 1051.870 6.310 1057.690 6.610 ;
        RECT 850.390 5.930 850.690 6.295 ;
        RECT 844.870 5.630 850.690 5.930 ;
        RECT 843.935 5.615 844.265 5.630 ;
        RECT 558.750 5.250 559.050 5.615 ;
        RECT 545.870 4.950 559.050 5.250 ;
        RECT 922.135 4.935 922.465 5.265 ;
        RECT 948.815 5.250 949.145 5.265 ;
        RECT 948.815 4.950 952.810 5.250 ;
        RECT 948.815 4.935 949.145 4.950 ;
        RECT 922.150 4.570 922.450 4.935 ;
        RECT 889.030 4.270 922.450 4.570 ;
        RECT 889.030 3.225 889.330 4.270 ;
        RECT 889.015 2.895 889.345 3.225 ;
        RECT 952.510 3.210 952.810 4.950 ;
        RECT 1051.870 3.225 1052.170 6.310 ;
        RECT 1093.270 5.250 1093.570 8.350 ;
        RECT 1135.590 8.350 1144.170 8.650 ;
        RECT 1266.230 11.750 1267.450 12.050 ;
        RECT 1480.590 11.750 1486.410 12.050 ;
        RECT 1124.535 7.970 1124.865 7.985 ;
        RECT 1104.310 7.670 1124.865 7.970 ;
        RECT 1104.310 5.250 1104.610 7.670 ;
        RECT 1124.535 7.655 1124.865 7.670 ;
        RECT 1135.590 6.625 1135.890 8.350 ;
        RECT 1266.230 7.985 1266.530 11.750 ;
        RECT 1480.590 7.985 1480.890 11.750 ;
        RECT 1266.215 7.655 1266.545 7.985 ;
        RECT 1480.575 7.655 1480.905 7.985 ;
        RECT 1135.575 6.295 1135.905 6.625 ;
        RECT 1093.270 4.950 1104.610 5.250 ;
        RECT 952.510 2.910 957.410 3.210 ;
        RECT 957.110 2.545 957.410 2.910 ;
        RECT 985.630 2.910 992.140 3.210 ;
        RECT 985.630 2.545 985.930 2.910 ;
        RECT 957.095 2.215 957.425 2.545 ;
        RECT 985.615 2.215 985.945 2.545 ;
        RECT 991.840 2.530 992.140 2.910 ;
        RECT 1039.895 2.895 1040.225 3.225 ;
        RECT 1051.855 2.895 1052.185 3.225 ;
        RECT 1039.910 2.530 1040.210 2.895 ;
        RECT 991.840 2.230 1040.210 2.530 ;
        RECT 317.710 1.550 325.370 1.850 ;
        RECT 1486.110 1.850 1486.410 11.750 ;
        RECT 1499.910 6.310 1519.530 6.610 ;
        RECT 1499.910 1.850 1500.210 6.310 ;
        RECT 1519.230 5.250 1519.530 6.310 ;
        RECT 1519.230 4.950 1549.890 5.250 ;
        RECT 1549.590 4.585 1549.890 4.950 ;
        RECT 1549.575 4.255 1549.905 4.585 ;
        RECT 1486.110 1.550 1500.210 1.850 ;
        RECT 305.735 1.170 306.065 1.185 ;
        RECT 317.710 1.170 318.010 1.550 ;
        RECT 305.735 0.870 318.010 1.170 ;
        RECT 305.735 0.855 306.065 0.870 ;
      LAYER met5 ;
        RECT 392.500 21.300 400.540 22.900 ;
        RECT 392.500 14.500 394.100 21.300 ;
        RECT 398.940 19.500 400.540 21.300 ;
        RECT 398.940 17.900 475.060 19.500 ;
        RECT 473.460 14.500 475.060 17.900 ;
        RECT 1143.220 14.500 1268.100 16.100 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 727.865 7.565 728.955 7.735 ;
        RECT 727.865 7.225 728.035 7.565 ;
        RECT 415.985 6.545 417.075 6.715 ;
        RECT 420.585 4.165 420.755 7.055 ;
        RECT 439.445 6.545 460.315 6.715 ;
        RECT 439.445 5.865 439.615 6.545 ;
        RECT 460.145 5.695 460.315 6.545 ;
        RECT 728.785 6.035 728.955 7.565 ;
        RECT 728.785 5.865 741.375 6.035 ;
        RECT 460.145 5.525 461.695 5.695 ;
        RECT 463.365 5.015 463.535 5.695 ;
        RECT 741.205 5.355 741.375 5.865 ;
        RECT 746.725 5.525 748.735 5.695 ;
        RECT 741.205 5.185 745.055 5.355 ;
        RECT 746.725 5.185 746.895 5.525 ;
        RECT 463.365 4.845 465.375 5.015 ;
        RECT 465.205 1.955 465.375 4.845 ;
        RECT 956.025 3.995 956.195 8.755 ;
        RECT 984.085 6.545 984.255 8.415 ;
        RECT 985.925 6.545 992.995 6.715 ;
        RECT 950.965 3.655 951.135 3.995 ;
        RECT 952.345 3.825 956.195 3.995 ;
        RECT 952.345 3.655 952.515 3.825 ;
        RECT 487.285 2.295 487.455 3.655 ;
        RECT 479.005 2.125 483.775 2.295 ;
        RECT 485.905 2.125 487.455 2.295 ;
        RECT 465.205 1.785 471.815 1.955 ;
        RECT 479.005 1.785 479.175 2.125 ;
        RECT 500.625 1.955 500.795 3.655 ;
        RECT 950.965 3.485 952.515 3.655 ;
        RECT 511.205 3.145 512.295 3.315 ;
        RECT 995.585 3.145 995.755 6.715 ;
        RECT 511.205 2.295 511.375 3.145 ;
        RECT 512.125 2.805 512.295 3.145 ;
        RECT 504.765 2.125 511.375 2.295 ;
        RECT 504.765 1.955 504.935 2.125 ;
        RECT 500.625 1.785 504.935 1.955 ;
      LAYER mcon ;
        RECT 956.025 8.585 956.195 8.755 ;
        RECT 420.585 6.885 420.755 7.055 ;
        RECT 416.905 6.545 417.075 6.715 ;
        RECT 461.525 5.525 461.695 5.695 ;
        RECT 463.365 5.525 463.535 5.695 ;
        RECT 748.565 5.525 748.735 5.695 ;
        RECT 744.885 5.185 745.055 5.355 ;
        RECT 984.085 8.245 984.255 8.415 ;
        RECT 992.825 6.545 992.995 6.715 ;
        RECT 995.585 6.545 995.755 6.715 ;
        RECT 950.965 3.825 951.135 3.995 ;
        RECT 487.285 3.485 487.455 3.655 ;
        RECT 483.605 2.125 483.775 2.295 ;
        RECT 500.625 3.485 500.795 3.655 ;
        RECT 471.645 1.785 471.815 1.955 ;
      LAYER met1 ;
        RECT 727.790 8.740 728.110 8.800 ;
        RECT 729.170 8.740 729.490 8.800 ;
        RECT 955.950 8.740 956.270 8.800 ;
        RECT 727.790 8.600 729.490 8.740 ;
        RECT 955.755 8.600 956.270 8.740 ;
        RECT 727.790 8.540 728.110 8.600 ;
        RECT 729.170 8.540 729.490 8.600 ;
        RECT 955.950 8.540 956.270 8.600 ;
        RECT 958.710 8.740 959.030 8.800 ;
        RECT 958.710 8.600 984.240 8.740 ;
        RECT 958.710 8.540 959.030 8.600 ;
        RECT 984.100 8.445 984.240 8.600 ;
        RECT 984.025 8.215 984.315 8.445 ;
        RECT 727.790 7.380 728.110 7.440 ;
        RECT 727.595 7.240 728.110 7.380 ;
        RECT 727.790 7.180 728.110 7.240 ;
        RECT 420.525 7.040 420.815 7.085 ;
        RECT 416.920 6.900 420.815 7.040 ;
        RECT 416.920 6.745 417.060 6.900 ;
        RECT 420.525 6.855 420.815 6.900 ;
        RECT 836.810 7.040 837.130 7.100 ;
        RECT 846.010 7.040 846.330 7.100 ;
        RECT 836.810 6.900 846.330 7.040 ;
        RECT 836.810 6.840 837.130 6.900 ;
        RECT 846.010 6.840 846.330 6.900 ;
        RECT 415.925 6.515 416.215 6.745 ;
        RECT 416.845 6.515 417.135 6.745 ;
        RECT 984.025 6.700 984.315 6.745 ;
        RECT 985.865 6.700 986.155 6.745 ;
        RECT 984.025 6.560 986.155 6.700 ;
        RECT 984.025 6.515 984.315 6.560 ;
        RECT 985.865 6.515 986.155 6.560 ;
        RECT 992.765 6.700 993.055 6.745 ;
        RECT 995.525 6.700 995.815 6.745 ;
        RECT 992.765 6.560 995.815 6.700 ;
        RECT 992.765 6.515 993.055 6.560 ;
        RECT 995.525 6.515 995.815 6.560 ;
        RECT 416.000 6.360 416.140 6.515 ;
        RECT 414.620 6.220 416.140 6.360 ;
        RECT 414.620 5.680 414.760 6.220 ;
        RECT 439.370 6.020 439.690 6.080 ;
        RECT 439.370 5.880 439.885 6.020 ;
        RECT 439.370 5.820 439.690 5.880 ;
        RECT 415.910 5.680 416.230 5.740 ;
        RECT 414.620 5.540 416.230 5.680 ;
        RECT 415.910 5.480 416.230 5.540 ;
        RECT 461.465 5.680 461.755 5.725 ;
        RECT 463.305 5.680 463.595 5.725 ;
        RECT 461.465 5.540 463.595 5.680 ;
        RECT 461.465 5.495 461.755 5.540 ;
        RECT 463.305 5.495 463.595 5.540 ;
        RECT 748.505 5.680 748.795 5.725 ;
        RECT 749.870 5.680 750.190 5.740 ;
        RECT 748.505 5.540 750.190 5.680 ;
        RECT 748.505 5.495 748.795 5.540 ;
        RECT 749.870 5.480 750.190 5.540 ;
        RECT 744.825 5.340 745.115 5.385 ;
        RECT 746.665 5.340 746.955 5.385 ;
        RECT 744.825 5.200 746.955 5.340 ;
        RECT 744.825 5.155 745.115 5.200 ;
        RECT 746.665 5.155 746.955 5.200 ;
        RECT 420.525 4.320 420.815 4.365 ;
        RECT 423.730 4.320 424.050 4.380 ;
        RECT 420.525 4.180 424.050 4.320 ;
        RECT 420.525 4.135 420.815 4.180 ;
        RECT 423.730 4.120 424.050 4.180 ;
        RECT 918.690 3.980 919.010 4.040 ;
        RECT 950.905 3.980 951.195 4.025 ;
        RECT 918.690 3.840 951.195 3.980 ;
        RECT 918.690 3.780 919.010 3.840 ;
        RECT 950.905 3.795 951.195 3.840 ;
        RECT 487.225 3.640 487.515 3.685 ;
        RECT 500.565 3.640 500.855 3.685 ;
        RECT 487.225 3.500 500.855 3.640 ;
        RECT 487.225 3.455 487.515 3.500 ;
        RECT 500.565 3.455 500.855 3.500 ;
        RECT 995.525 3.300 995.815 3.345 ;
        RECT 1021.730 3.300 1022.050 3.360 ;
        RECT 995.525 3.160 1022.050 3.300 ;
        RECT 995.525 3.115 995.815 3.160 ;
        RECT 1021.730 3.100 1022.050 3.160 ;
        RECT 512.065 2.960 512.355 3.005 ;
        RECT 515.270 2.960 515.590 3.020 ;
        RECT 512.065 2.820 515.590 2.960 ;
        RECT 512.065 2.775 512.355 2.820 ;
        RECT 515.270 2.760 515.590 2.820 ;
        RECT 483.545 2.280 483.835 2.325 ;
        RECT 485.845 2.280 486.135 2.325 ;
        RECT 483.545 2.140 486.135 2.280 ;
        RECT 483.545 2.095 483.835 2.140 ;
        RECT 485.845 2.095 486.135 2.140 ;
        RECT 471.585 1.940 471.875 1.985 ;
        RECT 478.945 1.940 479.235 1.985 ;
        RECT 471.585 1.800 479.235 1.940 ;
        RECT 471.585 1.755 471.875 1.800 ;
        RECT 478.945 1.755 479.235 1.800 ;
      LAYER via ;
        RECT 727.820 8.540 728.080 8.800 ;
        RECT 729.200 8.540 729.460 8.800 ;
        RECT 955.980 8.540 956.240 8.800 ;
        RECT 958.740 8.540 959.000 8.800 ;
        RECT 727.820 7.180 728.080 7.440 ;
        RECT 836.840 6.840 837.100 7.100 ;
        RECT 846.040 6.840 846.300 7.100 ;
        RECT 439.400 5.820 439.660 6.080 ;
        RECT 415.940 5.480 416.200 5.740 ;
        RECT 749.900 5.480 750.160 5.740 ;
        RECT 423.760 4.120 424.020 4.380 ;
        RECT 918.720 3.780 918.980 4.040 ;
        RECT 1021.760 3.100 1022.020 3.360 ;
        RECT 515.300 2.760 515.560 3.020 ;
      LAYER met2 ;
        RECT 344.170 8.570 344.450 8.685 ;
        RECT 327.680 8.430 344.450 8.570 ;
        RECT 322.160 8.260 323.220 8.400 ;
        RECT 306.060 2.990 307.120 3.130 ;
        RECT 306.060 2.400 306.200 2.990 ;
        RECT 305.850 -4.800 306.410 2.400 ;
        RECT 306.980 1.205 307.120 2.990 ;
        RECT 322.160 1.205 322.300 8.260 ;
        RECT 323.080 7.210 323.220 8.260 ;
        RECT 327.680 7.210 327.820 8.430 ;
        RECT 344.170 8.315 344.450 8.430 ;
        RECT 362.110 8.400 362.390 8.685 ;
        RECT 727.820 8.510 728.080 8.830 ;
        RECT 729.200 8.685 729.460 8.830 ;
        RECT 955.980 8.740 956.240 8.830 ;
        RECT 958.740 8.740 959.000 8.830 ;
        RECT 362.110 8.315 366.000 8.400 ;
        RECT 362.180 8.260 366.000 8.315 ;
        RECT 365.860 7.890 366.000 8.260 ;
        RECT 365.860 7.750 368.760 7.890 ;
        RECT 323.080 7.070 327.820 7.210 ;
        RECT 368.620 7.210 368.760 7.750 ;
        RECT 727.880 7.470 728.020 8.510 ;
        RECT 729.190 8.315 729.470 8.685 ;
        RECT 955.980 8.600 959.000 8.740 ;
        RECT 798.260 8.430 807.140 8.570 ;
        RECT 955.980 8.510 956.240 8.600 ;
        RECT 958.740 8.510 959.000 8.600 ;
        RECT 369.930 7.210 370.210 7.325 ;
        RECT 368.620 7.070 370.210 7.210 ;
        RECT 369.930 6.955 370.210 7.070 ;
        RECT 415.930 7.210 416.210 7.325 ;
        RECT 415.930 7.070 416.600 7.210 ;
        RECT 727.820 7.150 728.080 7.470 ;
        RECT 798.260 7.325 798.400 8.430 ;
        RECT 415.930 6.955 416.210 7.070 ;
        RECT 415.940 5.680 416.200 5.770 ;
        RECT 416.460 5.680 416.600 7.070 ;
        RECT 798.190 6.955 798.470 7.325 ;
        RECT 415.940 5.540 416.600 5.680 ;
        RECT 423.820 6.390 425.340 6.530 ;
        RECT 415.940 5.450 416.200 5.540 ;
        RECT 423.820 4.410 423.960 6.390 ;
        RECT 425.200 5.170 425.340 6.390 ;
        RECT 515.290 6.275 515.570 6.645 ;
        RECT 439.400 6.020 439.660 6.110 ;
        RECT 432.100 5.880 439.660 6.020 ;
        RECT 432.100 5.170 432.240 5.880 ;
        RECT 439.400 5.790 439.660 5.880 ;
        RECT 425.200 5.030 432.240 5.170 ;
        RECT 423.760 4.090 424.020 4.410 ;
        RECT 515.360 3.050 515.500 6.275 ;
        RECT 754.490 5.850 754.770 5.965 ;
        RECT 749.960 5.770 754.770 5.850 ;
        RECT 749.900 5.710 754.770 5.770 ;
        RECT 807.000 5.850 807.140 8.430 ;
        RECT 888.350 7.890 888.630 8.005 ;
        RECT 888.350 7.750 892.240 7.890 ;
        RECT 888.350 7.635 888.630 7.750 ;
        RECT 836.840 6.810 837.100 7.130 ;
        RECT 846.030 6.955 846.310 7.325 ;
        RECT 846.040 6.810 846.300 6.955 ;
        RECT 807.000 5.710 817.260 5.850 ;
        RECT 749.900 5.450 750.160 5.710 ;
        RECT 754.490 5.595 754.770 5.710 ;
        RECT 817.120 4.660 817.260 5.710 ;
        RECT 817.120 4.520 831.520 4.660 ;
        RECT 515.300 2.730 515.560 3.050 ;
        RECT 831.380 2.620 831.520 4.520 ;
        RECT 836.900 3.300 837.040 6.810 ;
        RECT 892.100 5.170 892.240 7.750 ;
        RECT 896.630 5.595 896.910 5.965 ;
        RECT 903.990 5.595 904.270 5.965 ;
        RECT 896.700 5.170 896.840 5.595 ;
        RECT 892.100 5.030 896.840 5.170 ;
        RECT 904.060 3.980 904.200 5.595 ;
        RECT 1025.830 5.170 1026.110 9.000 ;
        RECT 1021.820 5.030 1026.110 5.170 ;
        RECT 918.720 3.980 918.980 4.070 ;
        RECT 904.060 3.840 918.980 3.980 ;
        RECT 918.720 3.750 918.980 3.840 ;
        RECT 1021.820 3.390 1021.960 5.030 ;
        RECT 1025.830 5.000 1026.110 5.030 ;
        RECT 833.680 3.160 837.040 3.300 ;
        RECT 833.680 2.620 833.820 3.160 ;
        RECT 1021.760 3.070 1022.020 3.390 ;
        RECT 831.380 2.480 833.820 2.620 ;
        RECT 306.910 0.835 307.190 1.205 ;
        RECT 322.090 0.835 322.370 1.205 ;
      LAYER via2 ;
        RECT 344.170 8.360 344.450 8.640 ;
        RECT 362.110 8.360 362.390 8.640 ;
        RECT 729.190 8.360 729.470 8.640 ;
        RECT 369.930 7.000 370.210 7.280 ;
        RECT 415.930 7.000 416.210 7.280 ;
        RECT 798.190 7.000 798.470 7.280 ;
        RECT 515.290 6.320 515.570 6.600 ;
        RECT 754.490 5.640 754.770 5.920 ;
        RECT 888.350 7.680 888.630 7.960 ;
        RECT 846.030 7.000 846.310 7.280 ;
        RECT 896.630 5.640 896.910 5.920 ;
        RECT 903.990 5.640 904.270 5.920 ;
        RECT 306.910 0.880 307.190 1.160 ;
        RECT 322.090 0.880 322.370 1.160 ;
      LAYER met3 ;
        RECT 344.145 8.650 344.475 8.665 ;
        RECT 362.085 8.650 362.415 8.665 ;
        RECT 729.165 8.660 729.495 8.665 ;
        RECT 344.145 8.350 362.415 8.650 ;
        RECT 344.145 8.335 344.475 8.350 ;
        RECT 362.085 8.335 362.415 8.350 ;
        RECT 728.910 8.650 729.495 8.660 ;
        RECT 728.910 8.350 729.720 8.650 ;
        RECT 728.910 8.340 729.495 8.350 ;
        RECT 729.165 8.335 729.495 8.340 ;
        RECT 888.325 7.970 888.655 7.985 ;
        RECT 866.030 7.670 888.655 7.970 ;
        RECT 369.905 7.290 370.235 7.305 ;
        RECT 415.905 7.290 416.235 7.305 ;
        RECT 369.905 6.990 416.235 7.290 ;
        RECT 369.905 6.975 370.235 6.990 ;
        RECT 415.905 6.975 416.235 6.990 ;
        RECT 796.990 7.290 797.370 7.300 ;
        RECT 798.165 7.290 798.495 7.305 ;
        RECT 796.990 6.990 798.495 7.290 ;
        RECT 796.990 6.980 797.370 6.990 ;
        RECT 798.165 6.975 798.495 6.990 ;
        RECT 846.005 7.290 846.335 7.305 ;
        RECT 866.030 7.290 866.330 7.670 ;
        RECT 888.325 7.655 888.655 7.670 ;
        RECT 846.005 6.990 866.330 7.290 ;
        RECT 846.005 6.975 846.335 6.990 ;
        RECT 515.265 6.610 515.595 6.625 ;
        RECT 516.390 6.610 516.770 6.620 ;
        RECT 515.265 6.310 516.770 6.610 ;
        RECT 515.265 6.295 515.595 6.310 ;
        RECT 516.390 6.300 516.770 6.310 ;
        RECT 754.465 5.930 754.795 5.945 ;
        RECT 756.510 5.930 756.890 5.940 ;
        RECT 754.465 5.630 756.890 5.930 ;
        RECT 754.465 5.615 754.795 5.630 ;
        RECT 756.510 5.620 756.890 5.630 ;
        RECT 896.605 5.930 896.935 5.945 ;
        RECT 903.965 5.930 904.295 5.945 ;
        RECT 896.605 5.630 904.295 5.930 ;
        RECT 896.605 5.615 896.935 5.630 ;
        RECT 903.965 5.615 904.295 5.630 ;
        RECT 306.885 1.170 307.215 1.185 ;
        RECT 322.065 1.170 322.395 1.185 ;
        RECT 306.885 0.870 322.395 1.170 ;
        RECT 306.885 0.855 307.215 0.870 ;
        RECT 322.065 0.855 322.395 0.870 ;
        RECT 584.470 0.490 584.850 0.500 ;
        RECT 597.350 0.490 597.730 0.500 ;
        RECT 584.470 0.190 597.730 0.490 ;
        RECT 584.470 0.180 584.850 0.190 ;
        RECT 597.350 0.180 597.730 0.190 ;
      LAYER via3 ;
        RECT 728.940 8.340 729.260 8.660 ;
        RECT 797.020 6.980 797.340 7.300 ;
        RECT 516.420 6.300 516.740 6.620 ;
        RECT 756.540 5.620 756.860 5.940 ;
        RECT 584.500 0.180 584.820 0.500 ;
        RECT 597.380 0.180 597.700 0.500 ;
      LAYER met4 ;
        RECT 709.630 9.030 726.490 9.330 ;
        RECT 709.630 7.970 709.930 9.030 ;
        RECT 726.190 8.650 726.490 9.030 ;
        RECT 728.935 8.650 729.265 8.665 ;
        RECT 726.190 8.350 729.265 8.650 ;
        RECT 728.935 8.335 729.265 8.350 ;
        RECT 705.030 7.670 709.930 7.970 ;
        RECT 516.415 6.610 516.745 6.625 ;
        RECT 516.415 6.310 538.810 6.610 ;
        RECT 516.415 6.295 516.745 6.310 ;
        RECT 538.510 5.250 538.810 6.310 ;
        RECT 537.590 4.950 538.810 5.250 ;
        RECT 537.590 3.210 537.890 4.950 ;
        RECT 705.030 3.890 705.330 7.670 ;
        RECT 797.015 6.975 797.345 7.305 ;
        RECT 756.535 5.615 756.865 5.945 ;
        RECT 797.030 5.690 797.330 6.975 ;
        RECT 756.550 5.250 756.850 5.615 ;
        RECT 757.260 5.250 758.440 5.690 ;
        RECT 756.550 4.950 758.440 5.250 ;
        RECT 757.260 4.510 758.440 4.950 ;
        RECT 796.590 4.510 797.770 5.690 ;
        RECT 696.750 3.590 705.330 3.890 ;
        RECT 537.590 2.910 539.730 3.210 ;
        RECT 539.430 1.170 539.730 2.910 ;
        RECT 696.750 1.850 697.050 3.590 ;
        RECT 675.590 1.550 697.050 1.850 ;
        RECT 539.430 0.870 566.410 1.170 ;
        RECT 566.110 0.490 566.410 0.870 ;
        RECT 584.495 0.490 584.825 0.505 ;
        RECT 566.110 0.190 584.825 0.490 ;
        RECT 584.495 0.175 584.825 0.190 ;
        RECT 597.375 0.490 597.705 0.505 ;
        RECT 675.590 0.490 675.890 1.550 ;
        RECT 597.375 0.190 675.890 0.490 ;
        RECT 597.375 0.175 597.705 0.190 ;
      LAYER met5 ;
        RECT 757.050 4.300 797.980 5.900 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 555.365 8.245 557.835 8.415 ;
        RECT 362.625 6.885 364.635 7.055 ;
        RECT 393.905 6.885 407.415 7.055 ;
        RECT 346.985 0.765 347.155 4.675 ;
        RECT 362.625 0.765 362.795 6.885 ;
        RECT 364.465 6.545 364.635 6.885 ;
        RECT 408.625 0.255 408.795 7.055 ;
        RECT 421.045 0.255 421.215 7.055 ;
        RECT 553.985 4.165 554.155 7.395 ;
        RECT 555.365 7.225 555.535 8.245 ;
        RECT 557.665 6.885 557.835 8.245 ;
        RECT 582.505 5.185 582.675 8.075 ;
        RECT 756.845 5.355 757.015 7.055 ;
        RECT 758.225 5.355 758.395 8.075 ;
        RECT 766.045 7.395 766.215 7.735 ;
        RECT 766.045 7.225 769.435 7.395 ;
        RECT 769.265 7.055 769.435 7.225 ;
        RECT 769.265 6.885 775.415 7.055 ;
        RECT 775.245 6.205 775.415 6.885 ;
        RECT 756.845 5.185 758.395 5.355 ;
        RECT 1071.485 4.675 1071.655 6.715 ;
        RECT 1068.725 4.505 1071.655 4.675 ;
        RECT 1068.725 3.825 1068.895 4.505 ;
        RECT 408.625 0.085 421.215 0.255 ;
      LAYER mcon ;
        RECT 553.985 7.225 554.155 7.395 ;
        RECT 407.245 6.885 407.415 7.055 ;
        RECT 408.625 6.885 408.795 7.055 ;
        RECT 346.985 4.505 347.155 4.675 ;
        RECT 421.045 6.885 421.215 7.055 ;
        RECT 582.505 7.905 582.675 8.075 ;
        RECT 758.225 7.905 758.395 8.075 ;
        RECT 756.845 6.885 757.015 7.055 ;
        RECT 766.045 7.565 766.215 7.735 ;
        RECT 1071.485 6.545 1071.655 6.715 ;
      LAYER met1 ;
        RECT 575.990 8.060 576.310 8.120 ;
        RECT 582.445 8.060 582.735 8.105 ;
        RECT 575.990 7.920 582.735 8.060 ;
        RECT 575.990 7.860 576.310 7.920 ;
        RECT 582.445 7.875 582.735 7.920 ;
        RECT 758.165 8.060 758.455 8.105 ;
        RECT 758.165 7.920 761.140 8.060 ;
        RECT 758.165 7.875 758.455 7.920 ;
        RECT 761.000 7.720 761.140 7.920 ;
        RECT 765.985 7.720 766.275 7.765 ;
        RECT 761.000 7.580 766.275 7.720 ;
        RECT 765.985 7.535 766.275 7.580 ;
        RECT 553.925 7.380 554.215 7.425 ;
        RECT 555.305 7.380 555.595 7.425 ;
        RECT 553.925 7.240 555.595 7.380 ;
        RECT 553.925 7.195 554.215 7.240 ;
        RECT 555.305 7.195 555.595 7.240 ;
        RECT 393.845 7.040 394.135 7.085 ;
        RECT 374.600 6.900 394.135 7.040 ;
        RECT 364.405 6.700 364.695 6.745 ;
        RECT 374.600 6.700 374.740 6.900 ;
        RECT 393.845 6.855 394.135 6.900 ;
        RECT 407.185 7.040 407.475 7.085 ;
        RECT 408.565 7.040 408.855 7.085 ;
        RECT 407.185 6.900 408.855 7.040 ;
        RECT 407.185 6.855 407.475 6.900 ;
        RECT 408.565 6.855 408.855 6.900 ;
        RECT 420.985 7.040 421.275 7.085 ;
        RECT 428.330 7.040 428.650 7.100 ;
        RECT 420.985 6.900 428.650 7.040 ;
        RECT 420.985 6.855 421.275 6.900 ;
        RECT 428.330 6.840 428.650 6.900 ;
        RECT 557.605 7.040 557.895 7.085 ;
        RECT 575.990 7.040 576.310 7.100 ;
        RECT 557.605 6.900 576.310 7.040 ;
        RECT 557.605 6.855 557.895 6.900 ;
        RECT 575.990 6.840 576.310 6.900 ;
        RECT 744.350 7.040 744.670 7.100 ;
        RECT 756.785 7.040 757.075 7.085 ;
        RECT 744.350 6.900 757.075 7.040 ;
        RECT 744.350 6.840 744.670 6.900 ;
        RECT 756.785 6.855 757.075 6.900 ;
        RECT 834.050 7.040 834.370 7.100 ;
        RECT 836.350 7.040 836.670 7.100 ;
        RECT 834.050 6.900 836.670 7.040 ;
        RECT 834.050 6.840 834.370 6.900 ;
        RECT 836.350 6.840 836.670 6.900 ;
        RECT 364.405 6.560 374.740 6.700 ;
        RECT 1071.425 6.700 1071.715 6.745 ;
        RECT 1071.870 6.700 1072.190 6.760 ;
        RECT 1071.425 6.560 1072.190 6.700 ;
        RECT 364.405 6.515 364.695 6.560 ;
        RECT 1071.425 6.515 1071.715 6.560 ;
        RECT 1071.870 6.500 1072.190 6.560 ;
        RECT 775.185 6.360 775.475 6.405 ;
        RECT 782.070 6.360 782.390 6.420 ;
        RECT 775.185 6.220 782.390 6.360 ;
        RECT 775.185 6.175 775.475 6.220 ;
        RECT 782.070 6.160 782.390 6.220 ;
        RECT 787.130 6.360 787.450 6.420 ;
        RECT 790.810 6.360 791.130 6.420 ;
        RECT 787.130 6.220 791.130 6.360 ;
        RECT 787.130 6.160 787.450 6.220 ;
        RECT 790.810 6.160 791.130 6.220 ;
        RECT 333.570 5.340 333.890 5.400 ;
        RECT 344.150 5.340 344.470 5.400 ;
        RECT 333.570 5.200 344.470 5.340 ;
        RECT 333.570 5.140 333.890 5.200 ;
        RECT 344.150 5.140 344.470 5.200 ;
        RECT 582.445 5.340 582.735 5.385 ;
        RECT 605.890 5.340 606.210 5.400 ;
        RECT 582.445 5.200 606.210 5.340 ;
        RECT 582.445 5.155 582.735 5.200 ;
        RECT 605.890 5.140 606.210 5.200 ;
        RECT 344.610 4.660 344.930 4.720 ;
        RECT 346.925 4.660 347.215 4.705 ;
        RECT 344.610 4.520 347.215 4.660 ;
        RECT 344.610 4.460 344.930 4.520 ;
        RECT 346.925 4.475 347.215 4.520 ;
        RECT 550.230 4.320 550.550 4.380 ;
        RECT 553.925 4.320 554.215 4.365 ;
        RECT 550.230 4.180 554.215 4.320 ;
        RECT 550.230 4.120 550.550 4.180 ;
        RECT 553.925 4.135 554.215 4.180 ;
        RECT 1041.050 3.980 1041.370 4.040 ;
        RECT 1068.665 3.980 1068.955 4.025 ;
        RECT 1041.050 3.840 1068.955 3.980 ;
        RECT 1041.050 3.780 1041.370 3.840 ;
        RECT 1068.665 3.795 1068.955 3.840 ;
        RECT 346.925 0.920 347.215 0.965 ;
        RECT 362.565 0.920 362.855 0.965 ;
        RECT 346.925 0.780 362.855 0.920 ;
        RECT 346.925 0.735 347.215 0.780 ;
        RECT 362.565 0.735 362.855 0.780 ;
      LAYER via ;
        RECT 576.020 7.860 576.280 8.120 ;
        RECT 428.360 6.840 428.620 7.100 ;
        RECT 576.020 6.840 576.280 7.100 ;
        RECT 744.380 6.840 744.640 7.100 ;
        RECT 834.080 6.840 834.340 7.100 ;
        RECT 836.380 6.840 836.640 7.100 ;
        RECT 1071.900 6.500 1072.160 6.760 ;
        RECT 782.100 6.160 782.360 6.420 ;
        RECT 787.160 6.160 787.420 6.420 ;
        RECT 790.840 6.160 791.100 6.420 ;
        RECT 333.600 5.140 333.860 5.400 ;
        RECT 344.180 5.140 344.440 5.400 ;
        RECT 605.920 5.140 606.180 5.400 ;
        RECT 344.640 4.460 344.900 4.720 ;
        RECT 550.260 4.120 550.520 4.380 ;
        RECT 1041.080 3.780 1041.340 4.040 ;
      LAYER met2 ;
        RECT 794.970 8.315 795.250 8.685 ;
        RECT 834.070 8.315 834.350 8.685 ;
        RECT 576.020 7.830 576.280 8.150 ;
        RECT 576.080 7.130 576.220 7.830 ;
        RECT 795.040 7.325 795.180 8.315 ;
        RECT 428.360 6.810 428.620 7.130 ;
        RECT 576.020 6.810 576.280 7.130 ;
        RECT 744.380 6.810 744.640 7.130 ;
        RECT 790.830 6.955 791.110 7.325 ;
        RECT 794.970 6.955 795.250 7.325 ;
        RECT 834.140 7.130 834.280 8.315 ;
        RECT 836.440 7.580 837.500 7.720 ;
        RECT 836.440 7.130 836.580 7.580 ;
        RECT 428.420 6.020 428.560 6.810 ;
        RECT 744.440 6.645 744.580 6.810 ;
        RECT 430.190 6.530 430.470 6.645 ;
        RECT 429.800 6.390 430.470 6.530 ;
        RECT 429.800 6.020 429.940 6.390 ;
        RECT 430.190 6.275 430.470 6.390 ;
        RECT 744.370 6.275 744.650 6.645 ;
        RECT 790.900 6.450 791.040 6.955 ;
        RECT 834.080 6.810 834.340 7.130 ;
        RECT 836.380 6.810 836.640 7.130 ;
        RECT 782.100 6.360 782.360 6.450 ;
        RECT 787.160 6.360 787.420 6.450 ;
        RECT 782.100 6.220 787.420 6.360 ;
        RECT 782.100 6.130 782.360 6.220 ;
        RECT 787.160 6.130 787.420 6.220 ;
        RECT 790.840 6.130 791.100 6.450 ;
        RECT 323.930 5.595 324.210 5.965 ;
        RECT 333.590 5.595 333.870 5.965 ;
        RECT 428.420 5.880 429.940 6.020 ;
        RECT 536.910 5.680 537.190 5.965 ;
        RECT 536.910 5.595 545.860 5.680 ;
        RECT 324.000 2.400 324.140 5.595 ;
        RECT 333.660 5.430 333.800 5.595 ;
        RECT 536.980 5.540 545.860 5.595 ;
        RECT 333.600 5.110 333.860 5.430 ;
        RECT 344.180 5.170 344.440 5.430 ;
        RECT 344.180 5.110 344.840 5.170 ;
        RECT 344.240 5.030 344.840 5.110 ;
        RECT 344.700 4.750 344.840 5.030 ;
        RECT 344.640 4.430 344.900 4.750 ;
        RECT 545.720 4.660 545.860 5.540 ;
        RECT 605.920 5.110 606.180 5.430 ;
        RECT 546.640 4.860 550.460 5.000 ;
        RECT 546.640 4.660 546.780 4.860 ;
        RECT 460.550 4.490 460.830 4.605 ;
        RECT 545.720 4.520 546.780 4.660 ;
        RECT 460.550 4.350 461.680 4.490 ;
        RECT 550.320 4.410 550.460 4.860 ;
        RECT 460.550 4.235 460.830 4.350 ;
        RECT 323.790 -4.800 324.350 2.400 ;
        RECT 461.540 1.090 461.680 4.350 ;
        RECT 550.260 4.090 550.520 4.410 ;
        RECT 466.140 3.500 467.660 3.640 ;
        RECT 466.140 2.960 466.280 3.500 ;
        RECT 464.300 2.820 466.280 2.960 ;
        RECT 464.300 1.090 464.440 2.820 ;
        RECT 461.540 0.950 464.440 1.090 ;
        RECT 467.520 0.410 467.660 3.500 ;
        RECT 605.980 3.245 606.120 5.110 ;
        RECT 644.090 4.915 644.370 5.285 ;
        RECT 644.160 4.490 644.300 4.915 ;
        RECT 622.080 4.350 644.300 4.490 ;
        RECT 622.080 4.320 622.220 4.350 ;
        RECT 618.860 4.180 622.220 4.320 ;
        RECT 618.860 3.245 619.000 4.180 ;
        RECT 837.360 3.300 837.500 7.580 ;
        RECT 1040.150 6.275 1040.430 6.645 ;
        RECT 1071.900 6.530 1072.160 6.790 ;
        RECT 1073.210 6.530 1073.490 9.000 ;
        RECT 1071.900 6.470 1073.490 6.530 ;
        RECT 1071.960 6.390 1073.490 6.470 ;
        RECT 1040.220 3.980 1040.360 6.275 ;
        RECT 1073.210 5.000 1073.490 6.390 ;
        RECT 1041.080 3.980 1041.340 4.070 ;
        RECT 1040.220 3.840 1041.340 3.980 ;
        RECT 1041.080 3.750 1041.340 3.840 ;
        RECT 605.910 2.875 606.190 3.245 ;
        RECT 618.790 2.875 619.070 3.245 ;
        RECT 837.360 3.160 848.080 3.300 ;
        RECT 847.940 2.620 848.080 3.160 ;
        RECT 849.250 3.130 849.530 3.245 ;
        RECT 848.860 2.990 849.530 3.130 ;
        RECT 848.860 2.620 849.000 2.990 ;
        RECT 849.250 2.875 849.530 2.990 ;
        RECT 847.940 2.480 849.000 2.620 ;
        RECT 468.830 1.090 469.110 1.205 ;
        RECT 468.440 0.950 469.110 1.090 ;
        RECT 468.440 0.410 468.580 0.950 ;
        RECT 468.830 0.835 469.110 0.950 ;
        RECT 467.520 0.270 468.580 0.410 ;
      LAYER via2 ;
        RECT 794.970 8.360 795.250 8.640 ;
        RECT 834.070 8.360 834.350 8.640 ;
        RECT 790.830 7.000 791.110 7.280 ;
        RECT 794.970 7.000 795.250 7.280 ;
        RECT 430.190 6.320 430.470 6.600 ;
        RECT 744.370 6.320 744.650 6.600 ;
        RECT 323.930 5.640 324.210 5.920 ;
        RECT 333.590 5.640 333.870 5.920 ;
        RECT 536.910 5.640 537.190 5.920 ;
        RECT 460.550 4.280 460.830 4.560 ;
        RECT 644.090 4.960 644.370 5.240 ;
        RECT 1040.150 6.320 1040.430 6.600 ;
        RECT 605.910 2.920 606.190 3.200 ;
        RECT 618.790 2.920 619.070 3.200 ;
        RECT 849.250 2.920 849.530 3.200 ;
        RECT 468.830 0.880 469.110 1.160 ;
      LAYER met3 ;
        RECT 794.945 8.650 795.275 8.665 ;
        RECT 834.045 8.650 834.375 8.665 ;
        RECT 794.945 8.350 834.375 8.650 ;
        RECT 794.945 8.335 795.275 8.350 ;
        RECT 834.045 8.335 834.375 8.350 ;
        RECT 790.805 7.290 791.135 7.305 ;
        RECT 794.945 7.290 795.275 7.305 ;
        RECT 790.805 6.990 795.275 7.290 ;
        RECT 790.805 6.975 791.135 6.990 ;
        RECT 794.945 6.975 795.275 6.990 ;
        RECT 430.165 6.610 430.495 6.625 ;
        RECT 454.750 6.610 455.130 6.620 ;
        RECT 430.165 6.310 455.130 6.610 ;
        RECT 430.165 6.295 430.495 6.310 ;
        RECT 454.750 6.300 455.130 6.310 ;
        RECT 744.345 6.295 744.675 6.625 ;
        RECT 956.150 6.610 956.530 6.620 ;
        RECT 1040.125 6.610 1040.455 6.625 ;
        RECT 956.150 6.310 1040.455 6.610 ;
        RECT 956.150 6.300 956.530 6.310 ;
        RECT 1040.125 6.295 1040.455 6.310 ;
        RECT 323.905 5.930 324.235 5.945 ;
        RECT 333.565 5.930 333.895 5.945 ;
        RECT 323.905 5.630 333.895 5.930 ;
        RECT 323.905 5.615 324.235 5.630 ;
        RECT 333.565 5.615 333.895 5.630 ;
        RECT 535.710 5.930 536.090 5.940 ;
        RECT 536.885 5.930 537.215 5.945 ;
        RECT 535.710 5.630 537.215 5.930 ;
        RECT 535.710 5.620 536.090 5.630 ;
        RECT 536.885 5.615 537.215 5.630 ;
        RECT 743.630 5.930 744.010 5.940 ;
        RECT 744.360 5.930 744.660 6.295 ;
        RECT 743.630 5.630 744.660 5.930 ;
        RECT 743.630 5.620 744.010 5.630 ;
        RECT 644.065 5.250 644.395 5.265 ;
        RECT 644.065 4.950 649.210 5.250 ;
        RECT 644.065 4.935 644.395 4.950 ;
        RECT 460.525 4.570 460.855 4.585 ;
        RECT 459.390 4.270 460.855 4.570 ;
        RECT 459.390 3.900 459.690 4.270 ;
        RECT 460.525 4.255 460.855 4.270 ;
        RECT 459.350 3.580 459.730 3.900 ;
        RECT 648.910 3.890 649.210 4.950 ;
        RECT 651.630 3.890 652.010 3.900 ;
        RECT 648.910 3.590 652.010 3.890 ;
        RECT 651.630 3.580 652.010 3.590 ;
        RECT 605.885 3.210 606.215 3.225 ;
        RECT 618.765 3.210 619.095 3.225 ;
        RECT 849.225 3.220 849.555 3.225 ;
        RECT 605.885 2.910 619.095 3.210 ;
        RECT 605.885 2.895 606.215 2.910 ;
        RECT 618.765 2.895 619.095 2.910 ;
        RECT 677.390 3.210 677.770 3.220 ;
        RECT 699.470 3.210 699.850 3.220 ;
        RECT 849.225 3.210 849.810 3.220 ;
        RECT 677.390 2.910 699.850 3.210 ;
        RECT 849.000 2.910 849.810 3.210 ;
        RECT 677.390 2.900 677.770 2.910 ;
        RECT 699.470 2.900 699.850 2.910 ;
        RECT 849.225 2.900 849.810 2.910 ;
        RECT 877.030 3.210 877.410 3.220 ;
        RECT 886.230 3.210 886.610 3.220 ;
        RECT 877.030 2.910 886.610 3.210 ;
        RECT 877.030 2.900 877.410 2.910 ;
        RECT 886.230 2.900 886.610 2.910 ;
        RECT 849.225 2.895 849.555 2.900 ;
        RECT 468.805 1.170 469.135 1.185 ;
        RECT 469.470 1.170 469.850 1.180 ;
        RECT 468.805 0.870 469.850 1.170 ;
        RECT 468.805 0.855 469.135 0.870 ;
        RECT 469.470 0.860 469.850 0.870 ;
      LAYER via3 ;
        RECT 454.780 6.300 455.100 6.620 ;
        RECT 956.180 6.300 956.500 6.620 ;
        RECT 535.740 5.620 536.060 5.940 ;
        RECT 743.660 5.620 743.980 5.940 ;
        RECT 459.380 3.580 459.700 3.900 ;
        RECT 651.660 3.580 651.980 3.900 ;
        RECT 677.420 2.900 677.740 3.220 ;
        RECT 699.500 2.900 699.820 3.220 ;
        RECT 849.460 2.900 849.780 3.220 ;
        RECT 877.060 2.900 877.380 3.220 ;
        RECT 886.260 2.900 886.580 3.220 ;
        RECT 469.500 0.860 469.820 1.180 ;
      LAYER met4 ;
        RECT 454.775 6.295 455.105 6.625 ;
        RECT 956.175 6.610 956.505 6.625 ;
        RECT 949.750 6.310 956.505 6.610 ;
        RECT 454.790 3.890 455.090 6.295 ;
        RECT 535.735 5.930 536.065 5.945 ;
        RECT 524.710 5.630 536.065 5.930 ;
        RECT 524.710 5.250 525.010 5.630 ;
        RECT 535.735 5.615 536.065 5.630 ;
        RECT 743.655 5.615 743.985 5.945 ;
        RECT 949.750 5.930 950.050 6.310 ;
        RECT 956.175 6.295 956.505 6.310 ;
        RECT 923.070 5.630 950.050 5.930 ;
        RECT 523.790 4.950 525.010 5.250 ;
        RECT 459.375 3.890 459.705 3.905 ;
        RECT 454.790 3.590 459.705 3.890 ;
        RECT 459.375 3.575 459.705 3.590 ;
        RECT 523.790 3.210 524.090 4.950 ;
        RECT 651.670 4.270 675.890 4.570 ;
        RECT 651.670 3.905 651.970 4.270 ;
        RECT 651.655 3.575 651.985 3.905 ;
        RECT 675.590 3.210 675.890 4.270 ;
        RECT 677.415 3.210 677.745 3.225 ;
        RECT 523.790 2.910 524.320 3.210 ;
        RECT 675.590 2.910 677.745 3.210 ;
        RECT 469.070 1.110 470.250 2.290 ;
        RECT 518.750 1.110 519.930 2.290 ;
        RECT 469.495 0.855 469.825 1.110 ;
        RECT 519.190 0.490 519.490 1.110 ;
        RECT 524.020 0.490 524.320 2.910 ;
        RECT 677.415 2.895 677.745 2.910 ;
        RECT 699.495 2.895 699.825 3.225 ;
        RECT 699.510 2.530 699.810 2.895 ;
        RECT 743.670 2.530 743.970 5.615 ;
        RECT 923.070 3.890 923.370 5.630 ;
        RECT 849.455 2.895 849.785 3.225 ;
        RECT 699.510 2.230 743.970 2.530 ;
        RECT 849.470 2.290 849.770 2.895 ;
        RECT 876.630 2.470 877.810 3.650 ;
        RECT 889.950 3.590 923.370 3.890 ;
        RECT 886.255 2.895 886.585 3.225 ;
        RECT 849.030 1.110 850.210 2.290 ;
        RECT 886.270 1.850 886.570 2.895 ;
        RECT 889.950 1.850 890.250 3.590 ;
        RECT 886.270 1.550 890.250 1.850 ;
        RECT 519.190 0.190 524.320 0.490 ;
      LAYER via4 ;
        RECT 469.070 1.110 470.250 2.290 ;
      LAYER met5 ;
        RECT 874.580 2.500 878.020 3.860 ;
        RECT 468.860 0.900 520.140 2.500 ;
        RECT 848.820 2.260 878.020 2.500 ;
        RECT 848.820 0.900 876.180 2.260 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 507.525 8.585 512.295 8.755 ;
        RECT 429.785 7.565 432.255 7.735 ;
        RECT 429.785 6.885 429.955 7.565 ;
        RECT 432.085 4.165 432.255 7.565 ;
        RECT 438.985 7.225 463.995 7.395 ;
        RECT 507.525 7.225 507.695 8.585 ;
        RECT 512.125 8.415 512.295 8.585 ;
        RECT 512.125 8.245 519.195 8.415 ;
        RECT 519.025 7.565 519.195 8.245 ;
        RECT 438.985 4.165 439.155 7.225 ;
        RECT 521.785 5.695 521.955 7.735 ;
        RECT 953.265 6.545 953.435 7.395 ;
        RECT 521.785 5.525 524.715 5.695 ;
        RECT 532.825 4.165 536.675 4.335 ;
        RECT 1074.705 3.825 1076.715 3.995 ;
        RECT 1119.325 3.825 1119.495 5.695 ;
        RECT 1074.705 3.145 1074.875 3.825 ;
        RECT 1076.545 3.315 1076.715 3.825 ;
        RECT 1076.545 3.145 1088.675 3.315 ;
      LAYER mcon ;
        RECT 521.785 7.565 521.955 7.735 ;
        RECT 463.825 7.225 463.995 7.395 ;
        RECT 953.265 7.225 953.435 7.395 ;
        RECT 524.545 5.525 524.715 5.695 ;
        RECT 1119.325 5.525 1119.495 5.695 ;
        RECT 536.505 4.165 536.675 4.335 ;
        RECT 1088.505 3.145 1088.675 3.315 ;
      LAYER met1 ;
        RECT 518.965 7.720 519.255 7.765 ;
        RECT 521.725 7.720 522.015 7.765 ;
        RECT 518.965 7.580 522.015 7.720 ;
        RECT 518.965 7.535 519.255 7.580 ;
        RECT 521.725 7.535 522.015 7.580 ;
        RECT 463.765 7.380 464.055 7.425 ;
        RECT 507.465 7.380 507.755 7.425 ;
        RECT 463.765 7.240 507.755 7.380 ;
        RECT 463.765 7.195 464.055 7.240 ;
        RECT 507.465 7.195 507.755 7.240 ;
        RECT 629.810 7.380 630.130 7.440 ;
        RECT 639.930 7.380 640.250 7.440 ;
        RECT 629.810 7.240 640.250 7.380 ;
        RECT 629.810 7.180 630.130 7.240 ;
        RECT 639.930 7.180 640.250 7.240 ;
        RECT 953.205 7.380 953.495 7.425 ;
        RECT 955.030 7.380 955.350 7.440 ;
        RECT 953.205 7.240 955.350 7.380 ;
        RECT 953.205 7.195 953.495 7.240 ;
        RECT 955.030 7.180 955.350 7.240 ;
        RECT 429.250 7.040 429.570 7.100 ;
        RECT 429.725 7.040 430.015 7.085 ;
        RECT 429.250 6.900 430.015 7.040 ;
        RECT 429.250 6.840 429.570 6.900 ;
        RECT 429.725 6.855 430.015 6.900 ;
        RECT 950.890 6.700 951.210 6.760 ;
        RECT 953.205 6.700 953.495 6.745 ;
        RECT 950.890 6.560 953.495 6.700 ;
        RECT 950.890 6.500 951.210 6.560 ;
        RECT 953.205 6.515 953.495 6.560 ;
        RECT 524.485 5.680 524.775 5.725 ;
        RECT 529.070 5.680 529.390 5.740 ;
        RECT 524.485 5.540 529.390 5.680 ;
        RECT 524.485 5.495 524.775 5.540 ;
        RECT 529.070 5.480 529.390 5.540 ;
        RECT 1119.250 5.680 1119.570 5.740 ;
        RECT 1119.250 5.540 1119.765 5.680 ;
        RECT 1119.250 5.480 1119.570 5.540 ;
        RECT 432.025 4.320 432.315 4.365 ;
        RECT 438.925 4.320 439.215 4.365 ;
        RECT 432.025 4.180 439.215 4.320 ;
        RECT 432.025 4.135 432.315 4.180 ;
        RECT 438.925 4.135 439.215 4.180 ;
        RECT 532.290 4.320 532.610 4.380 ;
        RECT 532.765 4.320 533.055 4.365 ;
        RECT 532.290 4.180 533.055 4.320 ;
        RECT 532.290 4.120 532.610 4.180 ;
        RECT 532.765 4.135 533.055 4.180 ;
        RECT 536.445 4.320 536.735 4.365 ;
        RECT 544.250 4.320 544.570 4.380 ;
        RECT 536.445 4.180 544.570 4.320 ;
        RECT 536.445 4.135 536.735 4.180 ;
        RECT 544.250 4.120 544.570 4.180 ;
        RECT 1097.170 3.980 1097.490 4.040 ;
        RECT 1119.265 3.980 1119.555 4.025 ;
        RECT 1097.170 3.840 1119.555 3.980 ;
        RECT 1097.170 3.780 1097.490 3.840 ;
        RECT 1119.265 3.795 1119.555 3.840 ;
        RECT 1070.490 3.300 1070.810 3.360 ;
        RECT 1074.645 3.300 1074.935 3.345 ;
        RECT 1070.490 3.160 1074.935 3.300 ;
        RECT 1070.490 3.100 1070.810 3.160 ;
        RECT 1074.645 3.115 1074.935 3.160 ;
        RECT 1088.445 3.300 1088.735 3.345 ;
        RECT 1097.170 3.300 1097.490 3.360 ;
        RECT 1088.445 3.160 1097.490 3.300 ;
        RECT 1088.445 3.115 1088.735 3.160 ;
        RECT 1097.170 3.100 1097.490 3.160 ;
        RECT 1015.750 2.280 1016.070 2.340 ;
        RECT 1059.910 2.280 1060.230 2.340 ;
        RECT 1015.750 2.140 1060.230 2.280 ;
        RECT 1015.750 2.080 1016.070 2.140 ;
        RECT 1059.910 2.080 1060.230 2.140 ;
      LAYER via ;
        RECT 629.840 7.180 630.100 7.440 ;
        RECT 639.960 7.180 640.220 7.440 ;
        RECT 955.060 7.180 955.320 7.440 ;
        RECT 429.280 6.840 429.540 7.100 ;
        RECT 950.920 6.500 951.180 6.760 ;
        RECT 529.100 5.480 529.360 5.740 ;
        RECT 1119.280 5.480 1119.540 5.740 ;
        RECT 532.320 4.120 532.580 4.380 ;
        RECT 544.280 4.120 544.540 4.380 ;
        RECT 1097.200 3.780 1097.460 4.040 ;
        RECT 1070.520 3.100 1070.780 3.360 ;
        RECT 1097.200 3.100 1097.460 3.360 ;
        RECT 1015.780 2.080 1016.040 2.340 ;
        RECT 1059.940 2.080 1060.200 2.340 ;
      LAYER met2 ;
        RECT 563.660 8.600 585.420 8.740 ;
        RECT 370.390 7.635 370.670 8.005 ;
        RECT 376.830 7.635 377.110 8.005 ;
        RECT 370.460 6.530 370.600 7.635 ;
        RECT 365.860 6.390 370.600 6.530 ;
        RECT 365.860 3.810 366.000 6.390 ;
        RECT 376.900 4.660 377.040 7.635 ;
        RECT 429.280 6.810 429.540 7.130 ;
        RECT 429.340 6.645 429.480 6.810 ;
        RECT 429.270 6.275 429.550 6.645 ;
        RECT 529.100 5.680 529.360 5.770 ;
        RECT 529.100 5.540 532.520 5.680 ;
        RECT 529.100 5.450 529.360 5.540 ;
        RECT 376.900 4.520 379.800 4.660 ;
        RECT 363.100 3.670 366.000 3.810 ;
        RECT 341.480 2.990 342.540 3.130 ;
        RECT 341.480 2.400 341.620 2.990 ;
        RECT 342.400 2.565 342.540 2.990 ;
        RECT 363.100 2.565 363.240 3.670 ;
        RECT 379.660 2.565 379.800 4.520 ;
        RECT 532.380 4.410 532.520 5.540 ;
        RECT 563.660 5.340 563.800 8.600 ;
        RECT 585.280 6.645 585.420 8.600 ;
        RECT 611.430 8.570 611.710 8.685 ;
        RECT 609.200 8.430 611.710 8.570 ;
        RECT 609.200 6.645 609.340 8.430 ;
        RECT 611.430 8.315 611.710 8.430 ;
        RECT 621.550 8.570 621.830 8.685 ;
        RECT 621.550 8.430 622.220 8.570 ;
        RECT 621.550 8.315 621.830 8.430 ;
        RECT 622.080 6.700 622.220 8.430 ;
        RECT 676.750 8.315 677.030 8.685 ;
        RECT 983.570 8.315 983.850 8.685 ;
        RECT 676.820 8.060 676.960 8.315 ;
        RECT 639.950 7.635 640.230 8.005 ;
        RECT 676.820 7.920 677.880 8.060 ;
        RECT 640.020 7.470 640.160 7.635 ;
        RECT 629.840 7.150 630.100 7.470 ;
        RECT 639.960 7.150 640.220 7.470 ;
        RECT 677.740 7.325 677.880 7.920 ;
        RECT 629.900 6.700 630.040 7.150 ;
        RECT 677.670 6.955 677.950 7.325 ;
        RECT 955.060 7.150 955.320 7.470 ;
        RECT 950.920 6.700 951.180 6.790 ;
        RECT 585.210 6.275 585.490 6.645 ;
        RECT 609.130 6.275 609.410 6.645 ;
        RECT 622.080 6.560 630.040 6.700 ;
        RECT 948.150 6.530 948.430 6.645 ;
        RECT 950.060 6.560 951.180 6.700 ;
        RECT 950.060 6.530 950.200 6.560 ;
        RECT 948.150 6.390 950.200 6.530 ;
        RECT 950.920 6.470 951.180 6.560 ;
        RECT 948.150 6.275 948.430 6.390 ;
        RECT 955.120 5.850 955.260 7.150 ;
        RECT 983.640 5.965 983.780 8.315 ;
        RECT 1001.510 7.210 1001.790 7.325 ;
        RECT 1001.510 7.070 1015.980 7.210 ;
        RECT 1001.510 6.955 1001.790 7.070 ;
        RECT 957.810 5.850 958.090 5.965 ;
        RECT 955.120 5.710 958.090 5.850 ;
        RECT 957.810 5.595 958.090 5.710 ;
        RECT 983.570 5.595 983.850 5.965 ;
        RECT 559.980 5.200 563.800 5.340 ;
        RECT 532.320 4.090 532.580 4.410 ;
        RECT 544.280 4.320 544.540 4.410 ;
        RECT 544.280 4.180 544.940 4.320 ;
        RECT 544.280 4.090 544.540 4.180 ;
        RECT 341.270 -4.800 341.830 2.400 ;
        RECT 342.330 2.195 342.610 2.565 ;
        RECT 363.030 2.195 363.310 2.565 ;
        RECT 379.590 2.195 379.870 2.565 ;
        RECT 544.800 1.205 544.940 4.180 ;
        RECT 544.730 0.835 545.010 1.205 ;
        RECT 558.530 1.090 558.810 1.205 ;
        RECT 559.980 1.090 560.120 5.200 ;
        RECT 1015.840 2.370 1015.980 7.070 ;
        RECT 1119.280 5.450 1119.540 5.770 ;
        RECT 1119.340 5.170 1119.480 5.450 ;
        RECT 1121.050 5.170 1121.330 9.000 ;
        RECT 1119.340 5.030 1121.330 5.170 ;
        RECT 1121.050 5.000 1121.330 5.030 ;
        RECT 1060.460 4.350 1068.880 4.490 ;
        RECT 1060.460 3.640 1060.600 4.350 ;
        RECT 1060.000 3.500 1060.600 3.640 ;
        RECT 1060.000 2.370 1060.140 3.500 ;
        RECT 1068.740 3.300 1068.880 4.350 ;
        RECT 1097.200 3.750 1097.460 4.070 ;
        RECT 1097.260 3.390 1097.400 3.750 ;
        RECT 1070.520 3.300 1070.780 3.390 ;
        RECT 1068.740 3.160 1070.780 3.300 ;
        RECT 1070.520 3.070 1070.780 3.160 ;
        RECT 1097.200 3.070 1097.460 3.390 ;
        RECT 1015.780 2.050 1016.040 2.370 ;
        RECT 1059.940 2.050 1060.200 2.370 ;
        RECT 558.530 0.950 560.120 1.090 ;
        RECT 558.530 0.835 558.810 0.950 ;
      LAYER via2 ;
        RECT 370.390 7.680 370.670 7.960 ;
        RECT 376.830 7.680 377.110 7.960 ;
        RECT 429.270 6.320 429.550 6.600 ;
        RECT 611.430 8.360 611.710 8.640 ;
        RECT 621.550 8.360 621.830 8.640 ;
        RECT 676.750 8.360 677.030 8.640 ;
        RECT 983.570 8.360 983.850 8.640 ;
        RECT 639.950 7.680 640.230 7.960 ;
        RECT 677.670 7.000 677.950 7.280 ;
        RECT 585.210 6.320 585.490 6.600 ;
        RECT 609.130 6.320 609.410 6.600 ;
        RECT 948.150 6.320 948.430 6.600 ;
        RECT 1001.510 7.000 1001.790 7.280 ;
        RECT 957.810 5.640 958.090 5.920 ;
        RECT 983.570 5.640 983.850 5.920 ;
        RECT 342.330 2.240 342.610 2.520 ;
        RECT 363.030 2.240 363.310 2.520 ;
        RECT 379.590 2.240 379.870 2.520 ;
        RECT 544.730 0.880 545.010 1.160 ;
        RECT 558.530 0.880 558.810 1.160 ;
      LAYER met3 ;
        RECT 611.405 8.650 611.735 8.665 ;
        RECT 621.525 8.650 621.855 8.665 ;
        RECT 676.725 8.660 677.055 8.665 ;
        RECT 611.405 8.350 621.855 8.650 ;
        RECT 611.405 8.335 611.735 8.350 ;
        RECT 621.525 8.335 621.855 8.350 ;
        RECT 676.470 8.650 677.055 8.660 ;
        RECT 879.790 8.650 880.170 8.660 ;
        RECT 890.830 8.650 891.210 8.660 ;
        RECT 676.470 8.350 677.280 8.650 ;
        RECT 879.790 8.350 891.210 8.650 ;
        RECT 676.470 8.340 677.055 8.350 ;
        RECT 879.790 8.340 880.170 8.350 ;
        RECT 890.830 8.340 891.210 8.350 ;
        RECT 983.545 8.650 983.875 8.665 ;
        RECT 983.545 8.350 993.060 8.650 ;
        RECT 676.725 8.335 677.055 8.340 ;
        RECT 983.545 8.335 983.875 8.350 ;
        RECT 370.365 7.970 370.695 7.985 ;
        RECT 376.805 7.970 377.135 7.985 ;
        RECT 370.365 7.670 377.135 7.970 ;
        RECT 370.365 7.655 370.695 7.670 ;
        RECT 376.805 7.655 377.135 7.670 ;
        RECT 639.925 7.970 640.255 7.985 ;
        RECT 642.430 7.970 642.810 7.980 ;
        RECT 639.925 7.670 642.810 7.970 ;
        RECT 639.925 7.655 640.255 7.670 ;
        RECT 642.430 7.660 642.810 7.670 ;
        RECT 858.630 7.970 859.010 7.980 ;
        RECT 865.070 7.970 865.450 7.980 ;
        RECT 858.630 7.670 865.450 7.970 ;
        RECT 858.630 7.660 859.010 7.670 ;
        RECT 865.070 7.660 865.450 7.670 ;
        RECT 891.750 7.970 892.130 7.980 ;
        RECT 898.190 7.970 898.570 7.980 ;
        RECT 891.750 7.670 898.570 7.970 ;
        RECT 891.750 7.660 892.130 7.670 ;
        RECT 898.190 7.660 898.570 7.670 ;
        RECT 909.230 7.970 909.610 7.980 ;
        RECT 992.760 7.970 993.060 8.350 ;
        RECT 909.230 7.670 919.920 7.970 ;
        RECT 992.760 7.670 995.130 7.970 ;
        RECT 909.230 7.660 909.610 7.670 ;
        RECT 677.645 7.290 677.975 7.305 ;
        RECT 682.910 7.290 683.290 7.300 ;
        RECT 677.645 6.990 683.290 7.290 ;
        RECT 677.645 6.975 677.975 6.990 ;
        RECT 682.910 6.980 683.290 6.990 ;
        RECT 416.110 6.610 416.490 6.620 ;
        RECT 429.245 6.610 429.575 6.625 ;
        RECT 416.110 6.310 429.575 6.610 ;
        RECT 416.110 6.300 416.490 6.310 ;
        RECT 429.245 6.295 429.575 6.310 ;
        RECT 585.185 6.610 585.515 6.625 ;
        RECT 609.105 6.610 609.435 6.625 ;
        RECT 585.185 6.310 609.435 6.610 ;
        RECT 585.185 6.295 585.515 6.310 ;
        RECT 609.105 6.295 609.435 6.310 ;
        RECT 869.670 6.610 870.050 6.620 ;
        RECT 879.790 6.610 880.170 6.620 ;
        RECT 869.670 6.310 880.170 6.610 ;
        RECT 919.620 6.610 919.920 7.670 ;
        RECT 994.830 7.290 995.130 7.670 ;
        RECT 1001.485 7.290 1001.815 7.305 ;
        RECT 994.830 6.990 1001.815 7.290 ;
        RECT 1001.485 6.975 1001.815 6.990 ;
        RECT 948.125 6.610 948.455 6.625 ;
        RECT 919.620 6.310 948.455 6.610 ;
        RECT 869.670 6.300 870.050 6.310 ;
        RECT 879.790 6.300 880.170 6.310 ;
        RECT 948.125 6.295 948.455 6.310 ;
        RECT 699.470 5.930 699.850 5.940 ;
        RECT 705.910 5.930 706.290 5.940 ;
        RECT 699.470 5.630 706.290 5.930 ;
        RECT 699.470 5.620 699.850 5.630 ;
        RECT 705.910 5.620 706.290 5.630 ;
        RECT 957.785 5.930 958.115 5.945 ;
        RECT 983.545 5.930 983.875 5.945 ;
        RECT 957.785 5.630 983.875 5.930 ;
        RECT 957.785 5.615 958.115 5.630 ;
        RECT 983.545 5.615 983.875 5.630 ;
        RECT 721.550 3.890 721.930 3.900 ;
        RECT 727.990 3.890 728.370 3.900 ;
        RECT 721.550 3.590 728.370 3.890 ;
        RECT 721.550 3.580 721.930 3.590 ;
        RECT 727.990 3.580 728.370 3.590 ;
        RECT 342.305 2.530 342.635 2.545 ;
        RECT 363.005 2.530 363.335 2.545 ;
        RECT 342.305 2.230 363.335 2.530 ;
        RECT 342.305 2.215 342.635 2.230 ;
        RECT 363.005 2.215 363.335 2.230 ;
        RECT 379.565 2.530 379.895 2.545 ;
        RECT 380.230 2.530 380.610 2.540 ;
        RECT 379.565 2.230 380.610 2.530 ;
        RECT 379.565 2.215 379.895 2.230 ;
        RECT 380.230 2.220 380.610 2.230 ;
        RECT 544.705 1.170 545.035 1.185 ;
        RECT 558.505 1.170 558.835 1.185 ;
        RECT 544.705 0.870 558.835 1.170 ;
        RECT 544.705 0.855 545.035 0.870 ;
        RECT 558.505 0.855 558.835 0.870 ;
      LAYER via3 ;
        RECT 676.500 8.340 676.820 8.660 ;
        RECT 879.820 8.340 880.140 8.660 ;
        RECT 890.860 8.340 891.180 8.660 ;
        RECT 642.460 7.660 642.780 7.980 ;
        RECT 858.660 7.660 858.980 7.980 ;
        RECT 865.100 7.660 865.420 7.980 ;
        RECT 891.780 7.660 892.100 7.980 ;
        RECT 898.220 7.660 898.540 7.980 ;
        RECT 909.260 7.660 909.580 7.980 ;
        RECT 682.940 6.980 683.260 7.300 ;
        RECT 416.140 6.300 416.460 6.620 ;
        RECT 869.700 6.300 870.020 6.620 ;
        RECT 879.820 6.300 880.140 6.620 ;
        RECT 699.500 5.620 699.820 5.940 ;
        RECT 705.940 5.620 706.260 5.940 ;
        RECT 721.580 3.580 721.900 3.900 ;
        RECT 728.020 3.580 728.340 3.900 ;
        RECT 380.260 2.220 380.580 2.540 ;
      LAYER met4 ;
        RECT 793.350 11.750 851.610 12.050 ;
        RECT 642.470 9.030 670.370 9.330 ;
        RECT 642.470 7.985 642.770 9.030 ;
        RECT 670.070 8.650 670.370 9.030 ;
        RECT 676.495 8.650 676.825 8.665 ;
        RECT 670.070 8.350 676.825 8.650 ;
        RECT 676.495 8.335 676.825 8.350 ;
        RECT 642.455 7.655 642.785 7.985 ;
        RECT 394.070 6.990 416.450 7.290 ;
        RECT 380.255 2.215 380.585 2.545 ;
        RECT 380.270 1.850 380.570 2.215 ;
        RECT 394.070 1.850 394.370 6.990 ;
        RECT 416.150 6.625 416.450 6.990 ;
        RECT 682.935 6.975 683.265 7.305 ;
        RECT 745.510 6.990 760.530 7.290 ;
        RECT 416.135 6.295 416.465 6.625 ;
        RECT 682.950 3.210 683.250 6.975 ;
        RECT 742.750 6.310 744.890 6.610 ;
        RECT 699.495 5.930 699.825 5.945 ;
        RECT 698.590 5.630 699.825 5.930 ;
        RECT 698.590 4.570 698.890 5.630 ;
        RECT 699.495 5.615 699.825 5.630 ;
        RECT 705.935 5.615 706.265 5.945 ;
        RECT 690.310 4.270 698.890 4.570 ;
        RECT 690.310 3.210 690.610 4.270 ;
        RECT 705.950 3.890 706.250 5.615 ;
        RECT 721.575 3.890 721.905 3.905 ;
        RECT 705.950 3.590 721.905 3.890 ;
        RECT 721.575 3.575 721.905 3.590 ;
        RECT 728.015 3.575 728.345 3.905 ;
        RECT 682.950 2.910 690.610 3.210 ;
        RECT 728.030 3.210 728.330 3.575 ;
        RECT 742.750 3.210 743.050 6.310 ;
        RECT 728.030 2.910 743.050 3.210 ;
        RECT 744.590 3.210 744.890 6.310 ;
        RECT 745.510 3.210 745.810 6.990 ;
        RECT 760.230 4.570 760.530 6.990 ;
        RECT 793.350 5.250 793.650 11.750 ;
        RECT 851.310 9.330 851.610 11.750 ;
        RECT 851.310 9.030 857.130 9.330 ;
        RECT 856.830 7.970 857.130 9.030 ;
        RECT 879.815 8.335 880.145 8.665 ;
        RECT 890.855 8.650 891.185 8.665 ;
        RECT 890.855 8.350 892.090 8.650 ;
        RECT 890.855 8.335 891.185 8.350 ;
        RECT 858.655 7.970 858.985 7.985 ;
        RECT 856.830 7.670 858.985 7.970 ;
        RECT 858.655 7.655 858.985 7.670 ;
        RECT 865.095 7.655 865.425 7.985 ;
        RECT 865.110 6.610 865.410 7.655 ;
        RECT 879.830 6.625 880.130 8.335 ;
        RECT 891.790 7.985 892.090 8.350 ;
        RECT 891.775 7.655 892.105 7.985 ;
        RECT 898.215 7.970 898.545 7.985 ;
        RECT 909.255 7.970 909.585 7.985 ;
        RECT 898.215 7.670 909.585 7.970 ;
        RECT 898.215 7.655 898.545 7.670 ;
        RECT 909.255 7.655 909.585 7.670 ;
        RECT 869.695 6.610 870.025 6.625 ;
        RECT 865.110 6.310 870.025 6.610 ;
        RECT 869.695 6.295 870.025 6.310 ;
        RECT 879.815 6.295 880.145 6.625 ;
        RECT 762.990 4.950 793.650 5.250 ;
        RECT 762.990 4.570 763.290 4.950 ;
        RECT 760.230 4.270 763.290 4.570 ;
        RECT 744.590 2.910 745.810 3.210 ;
        RECT 380.270 1.550 394.370 1.850 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 197.485 3.825 197.655 6.375 ;
        RECT 290.865 1.105 291.035 7.395 ;
        RECT 327.665 7.225 327.835 9.095 ;
        RECT 334.105 5.865 334.275 7.395 ;
        RECT 381.485 5.865 381.655 7.395 ;
        RECT 438.525 6.375 438.695 7.395 ;
        RECT 530.065 6.885 530.235 9.095 ;
        RECT 643.225 7.225 643.395 8.415 ;
        RECT 751.325 7.735 751.495 9.095 ;
        RECT 1103.225 8.245 1104.775 8.415 ;
        RECT 1089.885 7.905 1102.015 8.075 ;
        RECT 1103.225 7.905 1103.395 8.245 ;
        RECT 1104.605 7.905 1104.775 8.245 ;
        RECT 1158.425 8.075 1158.595 9.095 ;
        RECT 1160.725 8.245 1160.895 9.095 ;
        RECT 751.325 7.565 752.875 7.735 ;
        RECT 752.705 7.225 752.875 7.565 ;
        RECT 437.145 6.205 438.695 6.375 ;
        RECT 414.145 5.865 415.235 6.035 ;
        RECT 424.265 4.165 424.435 6.035 ;
        RECT 429.325 3.995 429.495 4.335 ;
        RECT 437.145 3.995 437.315 6.205 ;
        RECT 1089.885 6.035 1090.055 7.905 ;
        RECT 1110.125 7.395 1110.295 8.075 ;
        RECT 1126.225 7.905 1158.595 8.075 ;
        RECT 1126.225 7.395 1126.395 7.905 ;
        RECT 1110.125 7.225 1126.395 7.395 ;
        RECT 429.325 3.825 437.315 3.995 ;
        RECT 1088.965 5.865 1090.055 6.035 ;
        RECT 1062.745 2.295 1062.915 3.315 ;
        RECT 1088.965 2.295 1089.135 5.865 ;
        RECT 1062.745 2.125 1089.135 2.295 ;
      LAYER mcon ;
        RECT 327.665 8.925 327.835 9.095 ;
        RECT 530.065 8.925 530.235 9.095 ;
        RECT 290.865 7.225 291.035 7.395 ;
        RECT 334.105 7.225 334.275 7.395 ;
        RECT 197.485 6.205 197.655 6.375 ;
        RECT 381.485 7.225 381.655 7.395 ;
        RECT 438.525 7.225 438.695 7.395 ;
        RECT 751.325 8.925 751.495 9.095 ;
        RECT 643.225 8.245 643.395 8.415 ;
        RECT 1158.425 8.925 1158.595 9.095 ;
        RECT 1101.845 7.905 1102.015 8.075 ;
        RECT 1160.725 8.925 1160.895 9.095 ;
        RECT 1110.125 7.905 1110.295 8.075 ;
        RECT 415.065 5.865 415.235 6.035 ;
        RECT 424.265 5.865 424.435 6.035 ;
        RECT 429.325 4.165 429.495 4.335 ;
        RECT 1062.745 3.145 1062.915 3.315 ;
      LAYER met1 ;
        RECT 327.605 9.080 327.895 9.125 ;
        RECT 530.005 9.080 530.295 9.125 ;
        RECT 751.265 9.080 751.555 9.125 ;
        RECT 327.605 8.940 530.295 9.080 ;
        RECT 327.605 8.895 327.895 8.940 ;
        RECT 530.005 8.895 530.295 8.940 ;
        RECT 746.280 8.940 751.555 9.080 ;
        RECT 746.280 8.800 746.420 8.940 ;
        RECT 751.265 8.895 751.555 8.940 ;
        RECT 1158.365 9.080 1158.655 9.125 ;
        RECT 1160.665 9.080 1160.955 9.125 ;
        RECT 1158.365 8.940 1160.955 9.080 ;
        RECT 1158.365 8.895 1158.655 8.940 ;
        RECT 1160.665 8.895 1160.955 8.940 ;
        RECT 643.240 8.600 647.520 8.740 ;
        RECT 643.240 8.445 643.380 8.600 ;
        RECT 643.165 8.215 643.455 8.445 ;
        RECT 647.380 8.400 647.520 8.600 ;
        RECT 746.190 8.540 746.510 8.800 ;
        RECT 1167.550 8.740 1167.870 8.800 ;
        RECT 1163.960 8.600 1167.870 8.740 ;
        RECT 672.590 8.400 672.910 8.460 ;
        RECT 647.380 8.260 672.910 8.400 ;
        RECT 672.590 8.200 672.910 8.260 ;
        RECT 1160.665 8.400 1160.955 8.445 ;
        RECT 1163.960 8.400 1164.100 8.600 ;
        RECT 1167.550 8.540 1167.870 8.600 ;
        RECT 1160.665 8.260 1164.100 8.400 ;
        RECT 1160.665 8.215 1160.955 8.260 ;
        RECT 1101.785 8.060 1102.075 8.105 ;
        RECT 1103.165 8.060 1103.455 8.105 ;
        RECT 1101.785 7.920 1103.455 8.060 ;
        RECT 1101.785 7.875 1102.075 7.920 ;
        RECT 1103.165 7.875 1103.455 7.920 ;
        RECT 1104.545 8.060 1104.835 8.105 ;
        RECT 1110.065 8.060 1110.355 8.105 ;
        RECT 1104.545 7.920 1110.355 8.060 ;
        RECT 1104.545 7.875 1104.835 7.920 ;
        RECT 1110.065 7.875 1110.355 7.920 ;
        RECT 290.805 7.380 291.095 7.425 ;
        RECT 303.670 7.380 303.990 7.440 ;
        RECT 327.605 7.380 327.895 7.425 ;
        RECT 290.805 7.240 303.990 7.380 ;
        RECT 290.805 7.195 291.095 7.240 ;
        RECT 303.670 7.180 303.990 7.240 ;
        RECT 311.120 7.240 327.895 7.380 ;
        RECT 311.120 7.040 311.260 7.240 ;
        RECT 327.605 7.195 327.895 7.240 ;
        RECT 334.045 7.380 334.335 7.425 ;
        RECT 381.425 7.380 381.715 7.425 ;
        RECT 334.045 7.240 381.715 7.380 ;
        RECT 334.045 7.195 334.335 7.240 ;
        RECT 381.425 7.195 381.715 7.240 ;
        RECT 438.465 7.380 438.755 7.425 ;
        RECT 642.230 7.380 642.550 7.440 ;
        RECT 643.165 7.380 643.455 7.425 ;
        RECT 746.190 7.380 746.510 7.440 ;
        RECT 438.465 7.240 463.520 7.380 ;
        RECT 438.465 7.195 438.755 7.240 ;
        RECT 274.780 6.900 311.260 7.040 ;
        RECT 359.330 7.040 359.650 7.100 ;
        RECT 372.210 7.040 372.530 7.100 ;
        RECT 359.330 6.900 372.530 7.040 ;
        RECT 463.380 7.040 463.520 7.240 ;
        RECT 642.230 7.240 643.455 7.380 ;
        RECT 642.230 7.180 642.550 7.240 ;
        RECT 643.165 7.195 643.455 7.240 ;
        RECT 737.540 7.240 746.510 7.380 ;
        RECT 530.005 7.040 530.295 7.085 ;
        RECT 549.310 7.040 549.630 7.100 ;
        RECT 463.380 6.900 463.980 7.040 ;
        RECT 274.780 6.700 274.920 6.900 ;
        RECT 359.330 6.840 359.650 6.900 ;
        RECT 372.210 6.840 372.530 6.900 ;
        RECT 235.680 6.560 274.920 6.700 ;
        RECT 197.425 6.360 197.715 6.405 ;
        RECT 235.680 6.360 235.820 6.560 ;
        RECT 197.425 6.220 235.820 6.360 ;
        RECT 463.840 6.360 463.980 6.900 ;
        RECT 530.005 6.900 549.630 7.040 ;
        RECT 530.005 6.855 530.295 6.900 ;
        RECT 549.310 6.840 549.630 6.900 ;
        RECT 725.950 7.040 726.270 7.100 ;
        RECT 737.540 7.040 737.680 7.240 ;
        RECT 746.190 7.180 746.510 7.240 ;
        RECT 752.645 7.380 752.935 7.425 ;
        RECT 762.750 7.380 763.070 7.440 ;
        RECT 752.645 7.240 763.070 7.380 ;
        RECT 752.645 7.195 752.935 7.240 ;
        RECT 762.750 7.180 763.070 7.240 ;
        RECT 725.950 6.900 737.680 7.040 ;
        RECT 725.950 6.840 726.270 6.900 ;
        RECT 501.470 6.360 501.790 6.420 ;
        RECT 463.840 6.220 501.790 6.360 ;
        RECT 197.425 6.175 197.715 6.220 ;
        RECT 501.470 6.160 501.790 6.220 ;
        RECT 552.990 6.360 553.310 6.420 ;
        RECT 555.750 6.360 556.070 6.420 ;
        RECT 552.990 6.220 556.070 6.360 ;
        RECT 552.990 6.160 553.310 6.220 ;
        RECT 555.750 6.160 556.070 6.220 ;
        RECT 317.930 6.020 318.250 6.080 ;
        RECT 334.045 6.020 334.335 6.065 ;
        RECT 317.930 5.880 334.335 6.020 ;
        RECT 317.930 5.820 318.250 5.880 ;
        RECT 334.045 5.835 334.335 5.880 ;
        RECT 381.425 6.020 381.715 6.065 ;
        RECT 414.085 6.020 414.375 6.065 ;
        RECT 381.425 5.880 414.375 6.020 ;
        RECT 381.425 5.835 381.715 5.880 ;
        RECT 414.085 5.835 414.375 5.880 ;
        RECT 415.005 6.020 415.295 6.065 ;
        RECT 424.205 6.020 424.495 6.065 ;
        RECT 415.005 5.880 424.495 6.020 ;
        RECT 415.005 5.835 415.295 5.880 ;
        RECT 424.205 5.835 424.495 5.880 ;
        RECT 424.205 4.320 424.495 4.365 ;
        RECT 429.265 4.320 429.555 4.365 ;
        RECT 424.205 4.180 429.555 4.320 ;
        RECT 424.205 4.135 424.495 4.180 ;
        RECT 429.265 4.135 429.555 4.180 ;
        RECT 190.970 3.980 191.290 4.040 ;
        RECT 197.425 3.980 197.715 4.025 ;
        RECT 190.970 3.840 197.715 3.980 ;
        RECT 190.970 3.780 191.290 3.840 ;
        RECT 197.425 3.795 197.715 3.840 ;
        RECT 1039.210 3.300 1039.530 3.360 ;
        RECT 1062.685 3.300 1062.975 3.345 ;
        RECT 1039.210 3.160 1062.975 3.300 ;
        RECT 1039.210 3.100 1039.530 3.160 ;
        RECT 1062.685 3.115 1062.975 3.160 ;
        RECT 278.370 1.260 278.690 1.320 ;
        RECT 290.805 1.260 291.095 1.305 ;
        RECT 278.370 1.120 291.095 1.260 ;
        RECT 278.370 1.060 278.690 1.120 ;
        RECT 290.805 1.075 291.095 1.120 ;
      LAYER via ;
        RECT 746.220 8.540 746.480 8.800 ;
        RECT 672.620 8.200 672.880 8.460 ;
        RECT 1167.580 8.540 1167.840 8.800 ;
        RECT 303.700 7.180 303.960 7.440 ;
        RECT 359.360 6.840 359.620 7.100 ;
        RECT 372.240 6.840 372.500 7.100 ;
        RECT 642.260 7.180 642.520 7.440 ;
        RECT 549.340 6.840 549.600 7.100 ;
        RECT 725.980 6.840 726.240 7.100 ;
        RECT 746.220 7.180 746.480 7.440 ;
        RECT 762.780 7.180 763.040 7.440 ;
        RECT 501.500 6.160 501.760 6.420 ;
        RECT 553.020 6.160 553.280 6.420 ;
        RECT 555.780 6.160 556.040 6.420 ;
        RECT 317.960 5.820 318.220 6.080 ;
        RECT 191.000 3.780 191.260 4.040 ;
        RECT 1039.240 3.100 1039.500 3.360 ;
        RECT 278.400 1.060 278.660 1.320 ;
      LAYER met2 ;
        RECT 503.270 7.720 503.550 9.000 ;
        RECT 504.780 8.600 538.040 8.740 ;
        RECT 504.780 8.570 504.920 8.600 ;
        RECT 504.320 8.430 504.920 8.570 ;
        RECT 504.320 7.720 504.460 8.430 ;
        RECT 537.900 7.890 538.040 8.600 ;
        RECT 537.900 7.750 545.400 7.890 ;
        RECT 501.100 7.580 504.460 7.720 ;
        RECT 545.260 7.720 545.400 7.750 ;
        RECT 545.260 7.580 546.780 7.720 ;
        RECT 303.700 7.150 303.960 7.470 ;
        RECT 303.760 5.965 303.900 7.150 ;
        RECT 359.360 6.810 359.620 7.130 ;
        RECT 372.240 6.810 372.500 7.130 ;
        RECT 303.690 5.595 303.970 5.965 ;
        RECT 316.570 5.595 316.850 5.965 ;
        RECT 317.960 5.790 318.220 6.110 ;
        RECT 316.640 4.660 316.780 5.595 ;
        RECT 318.020 4.660 318.160 5.790 ;
        RECT 316.640 4.520 318.160 4.660 ;
        RECT 191.000 3.925 191.260 4.070 ;
        RECT 121.530 3.555 121.810 3.925 ;
        RECT 190.990 3.555 191.270 3.925 ;
        RECT 247.570 3.555 247.850 3.925 ;
        RECT 278.390 3.555 278.670 3.925 ;
        RECT 97.680 2.820 98.740 2.960 ;
        RECT 97.680 2.400 97.820 2.820 ;
        RECT 97.470 -4.800 98.030 2.400 ;
        RECT 98.600 1.205 98.740 2.820 ;
        RECT 121.600 2.400 121.740 3.555 ;
        RECT 98.530 0.835 98.810 1.205 ;
        RECT 121.390 -4.800 121.950 2.400 ;
        RECT 247.640 1.205 247.780 3.555 ;
        RECT 278.460 1.350 278.600 3.555 ;
        RECT 359.420 2.400 359.560 6.810 ;
        RECT 372.300 5.285 372.440 6.810 ;
        RECT 501.100 6.645 501.240 7.580 ;
        RECT 489.530 6.530 489.810 6.645 ;
        RECT 489.140 6.390 489.810 6.530 ;
        RECT 372.230 4.915 372.510 5.285 ;
        RECT 247.570 0.835 247.850 1.205 ;
        RECT 278.400 1.030 278.660 1.350 ;
        RECT 359.210 -4.800 359.770 2.400 ;
        RECT 489.140 1.205 489.280 6.390 ;
        RECT 489.530 6.275 489.810 6.390 ;
        RECT 501.030 6.275 501.310 6.645 ;
        RECT 503.270 6.530 503.550 7.580 ;
        RECT 501.560 6.450 503.550 6.530 ;
        RECT 501.500 6.390 503.550 6.450 ;
        RECT 501.500 6.130 501.760 6.390 ;
        RECT 503.270 5.000 503.550 6.390 ;
        RECT 546.640 5.850 546.780 7.580 ;
        RECT 550.650 7.210 550.930 9.000 ;
        RECT 672.620 8.400 672.880 8.490 ;
        RECT 672.620 8.260 675.120 8.400 ;
        RECT 721.830 8.315 722.110 8.685 ;
        RECT 746.220 8.510 746.480 8.830 ;
        RECT 1167.580 8.570 1167.840 8.830 ;
        RECT 1168.430 8.570 1168.710 9.000 ;
        RECT 1167.580 8.510 1168.710 8.570 ;
        RECT 672.620 8.170 672.880 8.260 ;
        RECT 556.230 7.890 556.510 8.005 ;
        RECT 549.400 7.130 550.930 7.210 ;
        RECT 549.340 7.070 550.930 7.130 ;
        RECT 549.340 6.810 549.600 7.070 ;
        RECT 550.650 5.850 550.930 7.070 ;
        RECT 555.840 7.750 556.510 7.890 ;
        RECT 551.240 6.900 553.220 7.040 ;
        RECT 551.240 5.850 551.380 6.900 ;
        RECT 553.080 6.450 553.220 6.900 ;
        RECT 555.840 6.450 555.980 7.750 ;
        RECT 556.230 7.635 556.510 7.750 ;
        RECT 639.030 7.635 639.310 8.005 ;
        RECT 674.980 7.890 675.120 8.260 ;
        RECT 675.370 7.890 675.650 8.005 ;
        RECT 674.980 7.750 675.650 7.890 ;
        RECT 675.370 7.635 675.650 7.750 ;
        RECT 682.730 7.635 683.010 8.005 ;
        RECT 721.900 7.720 722.040 8.315 ;
        RECT 639.100 6.700 639.240 7.635 ;
        RECT 642.260 7.150 642.520 7.470 ;
        RECT 682.800 7.210 682.940 7.635 ;
        RECT 721.900 7.580 722.500 7.720 ;
        RECT 722.360 7.380 722.500 7.580 ;
        RECT 746.280 7.470 746.420 8.510 ;
        RECT 1167.640 8.430 1168.710 8.510 ;
        RECT 684.570 7.210 684.850 7.325 ;
        RECT 722.360 7.240 725.260 7.380 ;
        RECT 642.320 6.700 642.460 7.150 ;
        RECT 682.800 7.070 684.850 7.210 ;
        RECT 684.570 6.955 684.850 7.070 ;
        RECT 639.100 6.560 642.460 6.700 ;
        RECT 725.120 6.530 725.260 7.240 ;
        RECT 746.220 7.150 746.480 7.470 ;
        RECT 762.780 7.150 763.040 7.470 ;
        RECT 725.980 6.810 726.240 7.130 ;
        RECT 726.040 6.530 726.180 6.810 ;
        RECT 762.840 6.645 762.980 7.150 ;
        RECT 553.020 6.130 553.280 6.450 ;
        RECT 555.780 6.130 556.040 6.450 ;
        RECT 725.120 6.390 726.180 6.530 ;
        RECT 762.770 6.275 763.050 6.645 ;
        RECT 546.640 5.710 551.380 5.850 ;
        RECT 550.650 5.000 550.930 5.710 ;
        RECT 1168.430 5.000 1168.710 8.430 ;
        RECT 1039.240 3.245 1039.500 3.390 ;
        RECT 1039.230 2.875 1039.510 3.245 ;
        RECT 489.070 0.835 489.350 1.205 ;
      LAYER via2 ;
        RECT 303.690 5.640 303.970 5.920 ;
        RECT 316.570 5.640 316.850 5.920 ;
        RECT 121.530 3.600 121.810 3.880 ;
        RECT 190.990 3.600 191.270 3.880 ;
        RECT 247.570 3.600 247.850 3.880 ;
        RECT 278.390 3.600 278.670 3.880 ;
        RECT 98.530 0.880 98.810 1.160 ;
        RECT 372.230 4.960 372.510 5.240 ;
        RECT 247.570 0.880 247.850 1.160 ;
        RECT 489.530 6.320 489.810 6.600 ;
        RECT 501.030 6.320 501.310 6.600 ;
        RECT 721.830 8.360 722.110 8.640 ;
        RECT 556.230 7.680 556.510 7.960 ;
        RECT 639.030 7.680 639.310 7.960 ;
        RECT 675.370 7.680 675.650 7.960 ;
        RECT 682.730 7.680 683.010 7.960 ;
        RECT 684.570 7.000 684.850 7.280 ;
        RECT 762.770 6.320 763.050 6.600 ;
        RECT 1039.230 2.920 1039.510 3.200 ;
        RECT 489.070 0.880 489.350 1.160 ;
      LAYER met3 ;
        RECT 603.790 8.650 604.170 8.660 ;
        RECT 696.710 8.650 697.090 8.660 ;
        RECT 704.990 8.650 705.370 8.660 ;
        RECT 603.790 8.350 610.800 8.650 ;
        RECT 603.790 8.340 604.170 8.350 ;
        RECT 556.205 7.980 556.535 7.985 ;
        RECT 555.950 7.970 556.535 7.980 ;
        RECT 610.500 7.970 610.800 8.350 ;
        RECT 696.710 8.350 705.370 8.650 ;
        RECT 696.710 8.340 697.090 8.350 ;
        RECT 704.990 8.340 705.370 8.350 ;
        RECT 708.670 8.650 709.050 8.660 ;
        RECT 721.805 8.650 722.135 8.665 ;
        RECT 708.670 8.350 722.135 8.650 ;
        RECT 708.670 8.340 709.050 8.350 ;
        RECT 721.805 8.335 722.135 8.350 ;
        RECT 639.005 7.970 639.335 7.985 ;
        RECT 555.950 7.670 556.760 7.970 ;
        RECT 610.500 7.670 639.335 7.970 ;
        RECT 555.950 7.660 556.535 7.670 ;
        RECT 556.205 7.655 556.535 7.660 ;
        RECT 639.005 7.655 639.335 7.670 ;
        RECT 675.345 7.970 675.675 7.985 ;
        RECT 682.705 7.970 683.035 7.985 ;
        RECT 675.345 7.670 683.035 7.970 ;
        RECT 675.345 7.655 675.675 7.670 ;
        RECT 682.705 7.655 683.035 7.670 ;
        RECT 684.545 7.290 684.875 7.305 ;
        RECT 693.030 7.290 693.410 7.300 ;
        RECT 684.545 6.990 693.410 7.290 ;
        RECT 684.545 6.975 684.875 6.990 ;
        RECT 693.030 6.980 693.410 6.990 ;
        RECT 489.505 6.610 489.835 6.625 ;
        RECT 501.005 6.610 501.335 6.625 ;
        RECT 489.505 6.310 501.335 6.610 ;
        RECT 489.505 6.295 489.835 6.310 ;
        RECT 501.005 6.295 501.335 6.310 ;
        RECT 762.745 6.610 763.075 6.625 ;
        RECT 769.390 6.610 769.770 6.620 ;
        RECT 762.745 6.310 769.770 6.610 ;
        RECT 762.745 6.295 763.075 6.310 ;
        RECT 769.390 6.300 769.770 6.310 ;
        RECT 303.665 5.930 303.995 5.945 ;
        RECT 316.545 5.930 316.875 5.945 ;
        RECT 303.665 5.630 316.875 5.930 ;
        RECT 303.665 5.615 303.995 5.630 ;
        RECT 316.545 5.615 316.875 5.630 ;
        RECT 411.510 5.620 411.890 5.940 ;
        RECT 413.350 5.930 413.730 5.940 ;
        RECT 452.910 5.930 453.290 5.940 ;
        RECT 413.350 5.630 453.290 5.930 ;
        RECT 413.350 5.620 413.730 5.630 ;
        RECT 452.910 5.620 453.290 5.630 ;
        RECT 372.205 5.250 372.535 5.265 ;
        RECT 411.550 5.250 411.850 5.620 ;
        RECT 372.205 4.950 411.850 5.250 ;
        RECT 372.205 4.935 372.535 4.950 ;
        RECT 989.270 4.260 989.650 4.580 ;
        RECT 121.505 3.890 121.835 3.905 ;
        RECT 190.965 3.890 191.295 3.905 ;
        RECT 121.505 3.590 191.295 3.890 ;
        RECT 121.505 3.575 121.835 3.590 ;
        RECT 190.965 3.575 191.295 3.590 ;
        RECT 247.545 3.890 247.875 3.905 ;
        RECT 278.365 3.890 278.695 3.905 ;
        RECT 247.545 3.590 278.695 3.890 ;
        RECT 989.310 3.890 989.610 4.260 ;
        RECT 992.030 3.890 992.410 3.900 ;
        RECT 989.310 3.590 992.410 3.890 ;
        RECT 247.545 3.575 247.875 3.590 ;
        RECT 278.365 3.575 278.695 3.590 ;
        RECT 992.030 3.580 992.410 3.590 ;
        RECT 1026.070 3.210 1026.450 3.220 ;
        RECT 1039.205 3.210 1039.535 3.225 ;
        RECT 1026.070 2.910 1039.535 3.210 ;
        RECT 1026.070 2.900 1026.450 2.910 ;
        RECT 1039.205 2.895 1039.535 2.910 ;
        RECT 98.505 1.170 98.835 1.185 ;
        RECT 247.545 1.170 247.875 1.185 ;
        RECT 98.505 0.870 247.875 1.170 ;
        RECT 98.505 0.855 98.835 0.870 ;
        RECT 247.545 0.855 247.875 0.870 ;
        RECT 471.310 1.170 471.690 1.180 ;
        RECT 489.045 1.170 489.375 1.185 ;
        RECT 471.310 0.870 489.375 1.170 ;
        RECT 471.310 0.860 471.690 0.870 ;
        RECT 489.045 0.855 489.375 0.870 ;
      LAYER via3 ;
        RECT 603.820 8.340 604.140 8.660 ;
        RECT 555.980 7.660 556.300 7.980 ;
        RECT 696.740 8.340 697.060 8.660 ;
        RECT 705.020 8.340 705.340 8.660 ;
        RECT 708.700 8.340 709.020 8.660 ;
        RECT 693.060 6.980 693.380 7.300 ;
        RECT 769.420 6.300 769.740 6.620 ;
        RECT 411.540 5.620 411.860 5.940 ;
        RECT 413.380 5.620 413.700 5.940 ;
        RECT 452.940 5.620 453.260 5.940 ;
        RECT 989.300 4.260 989.620 4.580 ;
        RECT 992.060 3.580 992.380 3.900 ;
        RECT 1026.100 2.900 1026.420 3.220 ;
        RECT 471.340 0.860 471.660 1.180 ;
      LAYER met4 ;
        RECT 790.150 14.710 791.330 15.890 ;
        RECT 970.470 14.710 971.650 15.890 ;
        RECT 555.990 9.030 559.050 9.330 ;
        RECT 555.990 7.985 556.290 9.030 ;
        RECT 558.750 8.650 559.050 9.030 ;
        RECT 603.815 8.650 604.145 8.665 ;
        RECT 696.735 8.650 697.065 8.665 ;
        RECT 558.750 8.350 604.145 8.650 ;
        RECT 603.815 8.335 604.145 8.350 ;
        RECT 693.070 8.350 697.065 8.650 ;
        RECT 555.975 7.655 556.305 7.985 ;
        RECT 693.070 7.305 693.370 8.350 ;
        RECT 696.735 8.335 697.065 8.350 ;
        RECT 705.015 8.650 705.345 8.665 ;
        RECT 708.695 8.650 709.025 8.665 ;
        RECT 705.015 8.350 709.025 8.650 ;
        RECT 705.015 8.335 705.345 8.350 ;
        RECT 708.695 8.335 709.025 8.350 ;
        RECT 452.950 6.990 471.650 7.290 ;
        RECT 452.950 5.945 453.250 6.990 ;
        RECT 411.535 5.930 411.865 5.945 ;
        RECT 413.375 5.930 413.705 5.945 ;
        RECT 411.535 5.630 413.705 5.930 ;
        RECT 411.535 5.615 411.865 5.630 ;
        RECT 413.375 5.615 413.705 5.630 ;
        RECT 452.935 5.615 453.265 5.945 ;
        RECT 471.350 1.185 471.650 6.990 ;
        RECT 693.055 6.975 693.385 7.305 ;
        RECT 769.415 6.610 769.745 6.625 ;
        RECT 790.590 6.610 790.890 14.710 ;
        RECT 769.415 6.310 790.890 6.610 ;
        RECT 970.910 6.610 971.210 14.710 ;
        RECT 970.910 6.310 988.690 6.610 ;
        RECT 769.415 6.295 769.745 6.310 ;
        RECT 988.390 4.570 988.690 6.310 ;
        RECT 989.295 4.570 989.625 4.585 ;
        RECT 988.390 4.270 989.625 4.570 ;
        RECT 989.295 4.255 989.625 4.270 ;
        RECT 992.070 4.270 1024.340 4.570 ;
        RECT 992.070 3.905 992.370 4.270 ;
        RECT 992.055 3.575 992.385 3.905 ;
        RECT 1024.040 3.210 1024.340 4.270 ;
        RECT 1026.095 3.210 1026.425 3.225 ;
        RECT 1024.040 2.910 1026.425 3.210 ;
        RECT 1026.095 2.895 1026.425 2.910 ;
        RECT 471.335 0.855 471.665 1.185 ;
      LAYER met5 ;
        RECT 892.750 17.900 971.860 19.500 ;
        RECT 892.750 16.100 894.350 17.900 ;
        RECT 789.940 14.500 894.350 16.100 ;
        RECT 970.260 14.500 971.860 17.900 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 415.065 5.525 416.615 5.695 ;
        RECT 415.065 3.825 415.235 5.525 ;
      LAYER mcon ;
        RECT 416.445 5.525 416.615 5.695 ;
      LAYER met1 ;
        RECT 416.385 5.680 416.675 5.725 ;
        RECT 416.830 5.680 417.150 5.740 ;
        RECT 416.385 5.540 417.150 5.680 ;
        RECT 416.385 5.495 416.675 5.540 ;
        RECT 416.830 5.480 417.150 5.540 ;
        RECT 395.210 3.980 395.530 4.040 ;
        RECT 415.005 3.980 415.295 4.025 ;
        RECT 395.210 3.840 415.295 3.980 ;
        RECT 395.210 3.780 395.530 3.840 ;
        RECT 415.005 3.795 415.295 3.840 ;
      LAYER via ;
        RECT 416.860 5.480 417.120 5.740 ;
        RECT 395.240 3.780 395.500 4.040 ;
      LAYER met2 ;
        RECT 416.850 6.955 417.130 7.325 ;
        RECT 416.920 5.770 417.060 6.955 ;
        RECT 416.860 5.450 417.120 5.770 ;
        RECT 395.240 3.750 395.500 4.070 ;
        RECT 395.300 2.400 395.440 3.750 ;
        RECT 395.090 -4.800 395.650 2.400 ;
      LAYER via2 ;
        RECT 416.850 7.000 417.130 7.280 ;
      LAYER met3 ;
        RECT 464.870 8.650 465.250 8.660 ;
        RECT 472.230 8.650 472.610 8.660 ;
        RECT 464.870 8.350 472.610 8.650 ;
        RECT 464.870 8.340 465.250 8.350 ;
        RECT 472.230 8.340 472.610 8.350 ;
        RECT 474.070 7.970 474.450 7.980 ;
        RECT 478.670 7.970 479.050 7.980 ;
        RECT 474.070 7.670 479.050 7.970 ;
        RECT 474.070 7.660 474.450 7.670 ;
        RECT 478.670 7.660 479.050 7.670 ;
        RECT 416.825 7.300 417.155 7.305 ;
        RECT 416.825 7.290 417.410 7.300 ;
        RECT 416.600 6.990 417.410 7.290 ;
        RECT 416.825 6.980 417.410 6.990 ;
        RECT 416.825 6.975 417.155 6.980 ;
        RECT 428.070 1.170 428.450 1.180 ;
        RECT 436.350 1.170 436.730 1.180 ;
        RECT 428.070 0.870 436.730 1.170 ;
        RECT 428.070 0.860 428.450 0.870 ;
        RECT 436.350 0.860 436.730 0.870 ;
      LAYER via3 ;
        RECT 464.900 8.340 465.220 8.660 ;
        RECT 472.260 8.340 472.580 8.660 ;
        RECT 474.100 7.660 474.420 7.980 ;
        RECT 478.700 7.660 479.020 7.980 ;
        RECT 417.060 6.980 417.380 7.300 ;
        RECT 428.100 0.860 428.420 1.180 ;
        RECT 436.380 0.860 436.700 1.180 ;
      LAYER met4 ;
        RECT 621.100 18.110 622.280 19.290 ;
        RECT 483.790 14.710 484.970 15.890 ;
        RECT 484.230 9.330 484.530 14.710 ;
        RECT 463.070 9.030 465.210 9.330 ;
        RECT 463.070 7.970 463.370 9.030 ;
        RECT 464.910 8.665 465.210 9.030 ;
        RECT 478.710 9.030 484.530 9.330 ;
        RECT 464.895 8.335 465.225 8.665 ;
        RECT 472.255 8.650 472.585 8.665 ;
        RECT 472.255 8.350 474.410 8.650 ;
        RECT 472.255 8.335 472.585 8.350 ;
        RECT 474.110 7.985 474.410 8.350 ;
        RECT 478.710 7.985 479.010 9.030 ;
        RECT 417.070 7.670 428.410 7.970 ;
        RECT 417.070 7.305 417.370 7.670 ;
        RECT 417.055 6.975 417.385 7.305 ;
        RECT 428.110 1.185 428.410 7.670 ;
        RECT 443.750 7.670 463.370 7.970 ;
        RECT 443.750 3.890 444.050 7.670 ;
        RECT 474.095 7.655 474.425 7.985 ;
        RECT 478.695 7.655 479.025 7.985 ;
        RECT 436.390 3.590 444.050 3.890 ;
        RECT 436.390 1.185 436.690 3.590 ;
        RECT 428.095 0.855 428.425 1.185 ;
        RECT 436.375 0.855 436.705 1.185 ;
      LAYER met5 ;
        RECT 483.580 17.900 622.490 19.500 ;
        RECT 483.580 14.500 485.180 17.900 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 125.725 5.865 125.895 8.415 ;
        RECT 196.105 6.885 197.195 7.055 ;
        RECT 196.105 5.865 196.275 6.885 ;
        RECT 244.405 6.205 244.575 7.055 ;
        RECT 317.545 5.695 317.715 6.035 ;
        RECT 317.545 5.525 319.095 5.695 ;
        RECT 318.925 4.335 319.095 5.525 ;
        RECT 344.225 4.845 347.615 5.015 ;
        RECT 324.905 4.335 325.075 4.675 ;
        RECT 344.225 4.505 344.395 4.845 ;
        RECT 347.445 4.505 347.615 4.845 ;
        RECT 318.925 4.165 325.075 4.335 ;
        RECT 352.965 0.595 353.135 4.675 ;
        RECT 702.565 3.315 702.735 4.675 ;
        RECT 725.105 3.485 749.655 3.655 ;
        RECT 725.105 3.315 725.275 3.485 ;
        RECT 702.565 3.145 725.275 3.315 ;
        RECT 749.485 2.805 749.655 3.485 ;
        RECT 766.965 3.145 767.135 3.995 ;
        RECT 363.085 0.595 363.255 0.935 ;
        RECT 352.965 0.425 363.255 0.595 ;
        RECT 382.405 0.595 382.575 0.935 ;
        RECT 383.325 0.595 383.495 1.955 ;
        RECT 382.405 0.425 383.495 0.595 ;
      LAYER mcon ;
        RECT 125.725 8.245 125.895 8.415 ;
        RECT 197.025 6.885 197.195 7.055 ;
        RECT 244.405 6.885 244.575 7.055 ;
        RECT 317.545 5.865 317.715 6.035 ;
        RECT 324.905 4.505 325.075 4.675 ;
        RECT 352.965 4.505 353.135 4.675 ;
        RECT 702.565 4.505 702.735 4.675 ;
        RECT 766.965 3.825 767.135 3.995 ;
        RECT 383.325 1.785 383.495 1.955 ;
        RECT 363.085 0.765 363.255 0.935 ;
        RECT 382.405 0.765 382.575 0.935 ;
      LAYER met1 ;
        RECT 96.670 8.400 96.990 8.460 ;
        RECT 125.665 8.400 125.955 8.445 ;
        RECT 96.670 8.260 125.955 8.400 ;
        RECT 96.670 8.200 96.990 8.260 ;
        RECT 125.665 8.215 125.955 8.260 ;
        RECT 196.965 7.040 197.255 7.085 ;
        RECT 244.345 7.040 244.635 7.085 ;
        RECT 196.965 6.900 244.635 7.040 ;
        RECT 196.965 6.855 197.255 6.900 ;
        RECT 244.345 6.855 244.635 6.900 ;
        RECT 431.550 6.700 431.870 6.760 ;
        RECT 434.310 6.700 434.630 6.760 ;
        RECT 431.550 6.560 434.630 6.700 ;
        RECT 431.550 6.500 431.870 6.560 ;
        RECT 434.310 6.500 434.630 6.560 ;
        RECT 244.345 6.360 244.635 6.405 ;
        RECT 459.610 6.360 459.930 6.420 ;
        RECT 462.830 6.360 463.150 6.420 ;
        RECT 244.345 6.220 317.240 6.360 ;
        RECT 244.345 6.175 244.635 6.220 ;
        RECT 125.665 6.020 125.955 6.065 ;
        RECT 196.045 6.020 196.335 6.065 ;
        RECT 125.665 5.880 196.335 6.020 ;
        RECT 317.100 6.020 317.240 6.220 ;
        RECT 459.610 6.220 463.150 6.360 ;
        RECT 459.610 6.160 459.930 6.220 ;
        RECT 462.830 6.160 463.150 6.220 ;
        RECT 317.485 6.020 317.775 6.065 ;
        RECT 317.100 5.880 317.775 6.020 ;
        RECT 125.665 5.835 125.955 5.880 ;
        RECT 196.045 5.835 196.335 5.880 ;
        RECT 317.485 5.835 317.775 5.880 ;
        RECT 324.845 4.660 325.135 4.705 ;
        RECT 344.165 4.660 344.455 4.705 ;
        RECT 324.845 4.520 344.455 4.660 ;
        RECT 324.845 4.475 325.135 4.520 ;
        RECT 344.165 4.475 344.455 4.520 ;
        RECT 347.385 4.660 347.675 4.705 ;
        RECT 352.905 4.660 353.195 4.705 ;
        RECT 347.385 4.520 353.195 4.660 ;
        RECT 347.385 4.475 347.675 4.520 ;
        RECT 352.905 4.475 353.195 4.520 ;
        RECT 702.490 4.660 702.810 4.720 ;
        RECT 702.490 4.520 703.005 4.660 ;
        RECT 702.490 4.460 702.810 4.520 ;
        RECT 413.610 4.320 413.930 4.380 ;
        RECT 413.610 4.180 415.680 4.320 ;
        RECT 413.610 4.120 413.930 4.180 ;
        RECT 415.540 3.980 415.680 4.180 ;
        RECT 766.980 4.180 785.060 4.320 ;
        RECT 418.210 3.980 418.530 4.040 ;
        RECT 766.980 4.025 767.120 4.180 ;
        RECT 415.540 3.840 418.530 3.980 ;
        RECT 418.210 3.780 418.530 3.840 ;
        RECT 766.905 3.795 767.195 4.025 ;
        RECT 784.920 3.640 785.060 4.180 ;
        RECT 784.920 3.500 785.520 3.640 ;
        RECT 766.905 3.300 767.195 3.345 ;
        RECT 751.800 3.160 767.195 3.300 ;
        RECT 785.380 3.300 785.520 3.500 ;
        RECT 786.670 3.300 786.990 3.360 ;
        RECT 785.380 3.160 786.990 3.300 ;
        RECT 749.425 2.960 749.715 3.005 ;
        RECT 751.800 2.960 751.940 3.160 ;
        RECT 766.905 3.115 767.195 3.160 ;
        RECT 786.670 3.100 786.990 3.160 ;
        RECT 749.425 2.820 751.940 2.960 ;
        RECT 749.425 2.775 749.715 2.820 ;
        RECT 383.265 1.940 383.555 1.985 ;
        RECT 447.650 1.940 447.970 2.000 ;
        RECT 383.265 1.800 447.970 1.940 ;
        RECT 383.265 1.755 383.555 1.800 ;
        RECT 447.650 1.740 447.970 1.800 ;
        RECT 363.025 0.920 363.315 0.965 ;
        RECT 382.345 0.920 382.635 0.965 ;
        RECT 363.025 0.780 382.635 0.920 ;
        RECT 363.025 0.735 363.315 0.780 ;
        RECT 382.345 0.735 382.635 0.780 ;
      LAYER via ;
        RECT 96.700 8.200 96.960 8.460 ;
        RECT 431.580 6.500 431.840 6.760 ;
        RECT 434.340 6.500 434.600 6.760 ;
        RECT 459.640 6.160 459.900 6.420 ;
        RECT 462.860 6.160 463.120 6.420 ;
        RECT 702.520 4.460 702.780 4.720 ;
        RECT 413.640 4.120 413.900 4.380 ;
        RECT 418.240 3.780 418.500 4.040 ;
        RECT 786.700 3.100 786.960 3.360 ;
        RECT 447.680 1.740 447.940 2.000 ;
      LAYER met2 ;
        RECT 96.700 8.170 96.960 8.490 ;
        RECT 418.690 8.315 418.970 8.685 ;
        RECT 428.350 8.570 428.630 8.685 ;
        RECT 428.350 8.430 430.860 8.570 ;
        RECT 428.350 8.315 428.630 8.430 ;
        RECT 74.220 2.990 75.280 3.130 ;
        RECT 74.220 2.400 74.360 2.990 ;
        RECT 74.010 -4.800 74.570 2.400 ;
        RECT 75.140 1.205 75.280 2.990 ;
        RECT 96.760 1.205 96.900 8.170 ;
        RECT 413.640 4.090 413.900 4.410 ;
        RECT 413.700 3.640 413.840 4.090 ;
        RECT 418.240 3.980 418.500 4.070 ;
        RECT 418.760 3.980 418.900 8.315 ;
        RECT 430.720 6.700 430.860 8.430 ;
        RECT 434.400 7.070 435.920 7.210 ;
        RECT 434.400 6.790 434.540 7.070 ;
        RECT 435.780 7.040 435.920 7.070 ;
        RECT 455.890 7.040 456.170 9.000 ;
        RECT 463.770 7.635 464.050 8.005 ;
        RECT 463.840 7.040 463.980 7.635 ;
        RECT 435.780 6.900 456.620 7.040 ;
        RECT 431.580 6.700 431.840 6.790 ;
        RECT 430.720 6.560 431.840 6.700 ;
        RECT 431.580 6.470 431.840 6.560 ;
        RECT 434.340 6.470 434.600 6.790 ;
        RECT 455.890 5.170 456.170 6.900 ;
        RECT 456.480 6.360 456.620 6.900 ;
        RECT 462.920 6.900 463.980 7.040 ;
        RECT 462.920 6.450 463.060 6.900 ;
        RECT 459.640 6.360 459.900 6.450 ;
        RECT 456.480 6.220 459.900 6.360 ;
        RECT 459.640 6.130 459.900 6.220 ;
        RECT 462.860 6.130 463.120 6.450 ;
        RECT 418.240 3.840 418.900 3.980 ;
        RECT 447.740 5.030 456.170 5.170 ;
        RECT 418.240 3.750 418.500 3.840 ;
        RECT 413.240 3.500 413.840 3.640 ;
        RECT 413.240 2.400 413.380 3.500 ;
        RECT 75.070 0.835 75.350 1.205 ;
        RECT 96.690 0.835 96.970 1.205 ;
        RECT 413.030 -4.800 413.590 2.400 ;
        RECT 447.740 2.030 447.880 5.030 ;
        RECT 455.890 5.000 456.170 5.030 ;
        RECT 1309.710 5.170 1309.990 5.285 ;
        RECT 1311.030 5.170 1311.310 9.000 ;
        RECT 1309.710 5.030 1311.310 5.170 ;
        RECT 1309.710 4.915 1309.990 5.030 ;
        RECT 1311.030 5.000 1311.310 5.030 ;
        RECT 702.520 4.660 702.780 4.750 ;
        RECT 700.740 4.520 702.780 4.660 ;
        RECT 680.430 3.555 680.710 3.925 ;
        RECT 680.500 3.300 680.640 3.555 ;
        RECT 680.500 3.160 699.960 3.300 ;
        RECT 699.820 2.450 699.960 3.160 ;
        RECT 700.740 2.450 700.880 4.520 ;
        RECT 702.520 4.430 702.780 4.520 ;
        RECT 786.700 3.070 786.960 3.390 ;
        RECT 790.370 3.130 790.650 3.245 ;
        RECT 699.820 2.310 700.880 2.450 ;
        RECT 447.680 1.710 447.940 2.030 ;
        RECT 786.760 1.885 786.900 3.070 ;
        RECT 789.980 2.990 790.650 3.130 ;
        RECT 789.980 1.940 790.120 2.990 ;
        RECT 790.370 2.875 790.650 2.990 ;
        RECT 789.060 1.885 790.120 1.940 ;
        RECT 786.690 1.515 786.970 1.885 ;
        RECT 788.990 1.800 790.120 1.885 ;
        RECT 788.990 1.515 789.270 1.800 ;
      LAYER via2 ;
        RECT 418.690 8.360 418.970 8.640 ;
        RECT 428.350 8.360 428.630 8.640 ;
        RECT 463.770 7.680 464.050 7.960 ;
        RECT 75.070 0.880 75.350 1.160 ;
        RECT 96.690 0.880 96.970 1.160 ;
        RECT 1309.710 4.960 1309.990 5.240 ;
        RECT 680.430 3.600 680.710 3.880 ;
        RECT 790.370 2.920 790.650 3.200 ;
        RECT 786.690 1.560 786.970 1.840 ;
        RECT 788.990 1.560 789.270 1.840 ;
      LAYER met3 ;
        RECT 418.665 8.650 418.995 8.665 ;
        RECT 428.325 8.650 428.655 8.665 ;
        RECT 476.830 8.650 477.210 8.660 ;
        RECT 418.665 8.350 428.655 8.650 ;
        RECT 418.665 8.335 418.995 8.350 ;
        RECT 428.325 8.335 428.655 8.350 ;
        RECT 473.190 8.350 477.210 8.650 ;
        RECT 463.745 7.970 464.075 7.985 ;
        RECT 473.190 7.970 473.490 8.350 ;
        RECT 476.830 8.340 477.210 8.350 ;
        RECT 463.745 7.670 473.490 7.970 ;
        RECT 463.745 7.655 464.075 7.670 ;
        RECT 1279.990 5.250 1280.370 5.260 ;
        RECT 1309.685 5.250 1310.015 5.265 ;
        RECT 1279.990 4.950 1310.015 5.250 ;
        RECT 1279.990 4.940 1280.370 4.950 ;
        RECT 1309.685 4.935 1310.015 4.950 ;
        RECT 676.470 3.890 676.850 3.900 ;
        RECT 680.405 3.890 680.735 3.905 ;
        RECT 676.470 3.590 680.735 3.890 ;
        RECT 676.470 3.580 676.850 3.590 ;
        RECT 680.405 3.575 680.735 3.590 ;
        RECT 808.030 3.580 808.410 3.900 ;
        RECT 790.345 3.210 790.675 3.225 ;
        RECT 808.070 3.210 808.370 3.580 ;
        RECT 790.345 2.910 808.370 3.210 ;
        RECT 790.345 2.895 790.675 2.910 ;
        RECT 786.665 1.850 786.995 1.865 ;
        RECT 788.965 1.850 789.295 1.865 ;
        RECT 786.665 1.550 789.295 1.850 ;
        RECT 786.665 1.535 786.995 1.550 ;
        RECT 788.965 1.535 789.295 1.550 ;
        RECT 75.045 1.170 75.375 1.185 ;
        RECT 96.665 1.170 96.995 1.185 ;
        RECT 75.045 0.870 96.995 1.170 ;
        RECT 75.045 0.855 75.375 0.870 ;
        RECT 96.665 0.855 96.995 0.870 ;
      LAYER via3 ;
        RECT 476.860 8.340 477.180 8.660 ;
        RECT 1280.020 4.940 1280.340 5.260 ;
        RECT 676.500 3.580 676.820 3.900 ;
        RECT 808.060 3.580 808.380 3.900 ;
      LAYER met4 ;
        RECT 478.270 14.710 479.450 15.890 ;
        RECT 630.070 14.710 631.250 15.890 ;
        RECT 478.710 12.050 479.010 14.710 ;
        RECT 476.870 11.750 479.010 12.050 ;
        RECT 630.510 12.050 630.810 14.710 ;
        RECT 630.510 11.750 632.650 12.050 ;
        RECT 476.870 8.665 477.170 11.750 ;
        RECT 632.350 9.090 632.650 11.750 ;
        RECT 476.855 8.335 477.185 8.665 ;
        RECT 631.910 7.910 633.090 9.090 ;
        RECT 635.590 7.910 636.770 9.090 ;
        RECT 636.030 7.290 636.330 7.910 ;
        RECT 636.030 6.990 658.410 7.290 ;
        RECT 658.110 5.250 658.410 6.990 ;
        RECT 658.110 4.950 676.810 5.250 ;
        RECT 676.510 3.905 676.810 4.950 ;
        RECT 811.310 4.570 812.490 5.690 ;
        RECT 808.070 4.510 812.490 4.570 ;
        RECT 1205.070 5.250 1206.250 5.690 ;
        RECT 1210.590 5.250 1211.770 5.690 ;
        RECT 1205.070 4.950 1211.770 5.250 ;
        RECT 1205.070 4.510 1206.250 4.950 ;
        RECT 1210.590 4.510 1211.770 4.950 ;
        RECT 1274.070 5.250 1275.250 5.690 ;
        RECT 1280.015 5.250 1280.345 5.265 ;
        RECT 1274.070 4.950 1280.345 5.250 ;
        RECT 1274.070 4.510 1275.250 4.950 ;
        RECT 1280.015 4.935 1280.345 4.950 ;
        RECT 808.070 4.270 812.050 4.510 ;
        RECT 808.070 3.905 808.370 4.270 ;
        RECT 676.495 3.575 676.825 3.905 ;
        RECT 808.055 3.575 808.385 3.905 ;
      LAYER via4 ;
        RECT 811.310 4.510 812.490 5.690 ;
      LAYER met5 ;
        RECT 479.900 21.300 631.460 22.900 ;
        RECT 479.900 19.500 481.500 21.300 ;
        RECT 478.980 17.900 481.500 19.500 ;
        RECT 478.980 16.100 480.580 17.900 ;
        RECT 478.060 14.500 480.580 16.100 ;
        RECT 629.860 14.500 631.460 21.300 ;
        RECT 631.700 7.700 636.980 9.300 ;
        RECT 870.900 5.900 881.470 7.260 ;
        RECT 1005.220 5.900 1015.100 6.580 ;
        RECT 811.100 5.660 1206.460 5.900 ;
        RECT 811.100 4.300 872.500 5.660 ;
        RECT 879.870 4.980 1206.460 5.660 ;
        RECT 879.870 4.300 1006.820 4.980 ;
        RECT 1013.500 4.300 1206.460 4.980 ;
        RECT 1210.380 4.980 1275.460 6.580 ;
        RECT 1210.380 4.300 1211.980 4.980 ;
        RECT 1273.860 4.300 1275.460 4.980 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2850.765 1945.225 2850.935 1969.195 ;
        RECT 2849.845 1790.525 2850.015 1841.695 ;
        RECT 2849.845 1768.085 2850.015 1769.955 ;
        RECT 2851.225 1577.345 2851.395 1603.695 ;
        RECT 2851.685 1501.865 2851.855 1519.375 ;
        RECT 2849.845 1441.345 2850.015 1462.935 ;
        RECT 2850.305 1217.625 2850.475 1233.435 ;
        RECT 2850.305 1135.005 2850.475 1180.395 ;
        RECT 2850.305 1015.665 2850.475 1018.555 ;
        RECT 2850.305 941.885 2850.475 961.095 ;
        RECT 2850.305 884.085 2850.475 902.275 ;
        RECT 2851.225 809.965 2851.395 876.095 ;
        RECT 2851.685 769.505 2851.855 778.175 ;
        RECT 2852.605 734.825 2852.775 747.915 ;
        RECT 2852.145 293.505 2852.315 324.955 ;
        RECT 2851.685 39.185 2851.855 155.295 ;
        RECT 889.785 15.385 895.935 15.555 ;
        RECT 629.885 6.035 630.055 8.075 ;
        RECT 795.025 7.565 795.195 8.415 ;
        RECT 801.925 7.565 802.095 8.415 ;
        RECT 895.765 7.225 895.935 15.385 ;
        RECT 920.145 7.905 947.915 8.075 ;
        RECT 947.745 7.565 947.915 7.905 ;
        RECT 1254.105 7.225 1254.275 8.755 ;
        RECT 644.605 6.035 644.775 6.715 ;
        RECT 629.885 5.865 644.775 6.035 ;
      LAYER mcon ;
        RECT 2850.765 1969.025 2850.935 1969.195 ;
        RECT 2849.845 1841.525 2850.015 1841.695 ;
        RECT 2849.845 1769.785 2850.015 1769.955 ;
        RECT 2851.225 1603.525 2851.395 1603.695 ;
        RECT 2851.685 1519.205 2851.855 1519.375 ;
        RECT 2849.845 1462.765 2850.015 1462.935 ;
        RECT 2850.305 1233.265 2850.475 1233.435 ;
        RECT 2850.305 1180.225 2850.475 1180.395 ;
        RECT 2850.305 1018.385 2850.475 1018.555 ;
        RECT 2850.305 960.925 2850.475 961.095 ;
        RECT 2850.305 902.105 2850.475 902.275 ;
        RECT 2851.225 875.925 2851.395 876.095 ;
        RECT 2851.685 778.005 2851.855 778.175 ;
        RECT 2852.605 747.745 2852.775 747.915 ;
        RECT 2852.145 324.785 2852.315 324.955 ;
        RECT 2851.685 155.125 2851.855 155.295 ;
        RECT 795.025 8.245 795.195 8.415 ;
        RECT 629.885 7.905 630.055 8.075 ;
        RECT 801.925 8.245 802.095 8.415 ;
        RECT 1254.105 8.585 1254.275 8.755 ;
        RECT 644.605 6.545 644.775 6.715 ;
      LAYER met1 ;
        RECT 2850.690 2325.980 2851.010 2326.240 ;
        RECT 2850.780 2325.560 2850.920 2325.980 ;
        RECT 2850.690 2325.300 2851.010 2325.560 ;
        RECT 2849.770 1969.180 2850.090 1969.240 ;
        RECT 2850.705 1969.180 2850.995 1969.225 ;
        RECT 2849.770 1969.040 2850.995 1969.180 ;
        RECT 2849.770 1968.980 2850.090 1969.040 ;
        RECT 2850.705 1968.995 2850.995 1969.040 ;
        RECT 2849.770 1945.380 2850.090 1945.440 ;
        RECT 2850.705 1945.380 2850.995 1945.425 ;
        RECT 2849.770 1945.240 2850.995 1945.380 ;
        RECT 2849.770 1945.180 2850.090 1945.240 ;
        RECT 2850.705 1945.195 2850.995 1945.240 ;
        RECT 2849.770 1841.680 2850.090 1841.740 ;
        RECT 2849.575 1841.540 2850.090 1841.680 ;
        RECT 2849.770 1841.480 2850.090 1841.540 ;
        RECT 2849.785 1790.680 2850.075 1790.725 ;
        RECT 2849.400 1790.540 2850.075 1790.680 ;
        RECT 2849.400 1789.320 2849.540 1790.540 ;
        RECT 2849.785 1790.495 2850.075 1790.540 ;
        RECT 2849.770 1789.320 2850.090 1789.380 ;
        RECT 2849.400 1789.180 2850.090 1789.320 ;
        RECT 2849.770 1789.120 2850.090 1789.180 ;
        RECT 2849.770 1769.940 2850.090 1770.000 ;
        RECT 2849.770 1769.800 2850.285 1769.940 ;
        RECT 2849.770 1769.740 2850.090 1769.800 ;
        RECT 2849.770 1768.240 2850.090 1768.300 ;
        RECT 2849.770 1768.100 2850.285 1768.240 ;
        RECT 2849.770 1768.040 2850.090 1768.100 ;
        RECT 2849.770 1604.840 2850.090 1605.100 ;
        RECT 2849.860 1604.700 2850.000 1604.840 ;
        RECT 2849.860 1604.560 2851.380 1604.700 ;
        RECT 2851.240 1603.725 2851.380 1604.560 ;
        RECT 2851.165 1603.495 2851.455 1603.725 ;
        RECT 2851.150 1577.500 2851.470 1577.560 ;
        RECT 2850.955 1577.360 2851.470 1577.500 ;
        RECT 2851.150 1577.300 2851.470 1577.360 ;
        RECT 2851.150 1519.360 2851.470 1519.420 ;
        RECT 2851.625 1519.360 2851.915 1519.405 ;
        RECT 2851.150 1519.220 2851.915 1519.360 ;
        RECT 2851.150 1519.160 2851.470 1519.220 ;
        RECT 2851.625 1519.175 2851.915 1519.220 ;
        RECT 2851.625 1502.020 2851.915 1502.065 ;
        RECT 2852.070 1502.020 2852.390 1502.080 ;
        RECT 2851.625 1501.880 2852.390 1502.020 ;
        RECT 2851.625 1501.835 2851.915 1501.880 ;
        RECT 2852.070 1501.820 2852.390 1501.880 ;
        RECT 2849.785 1462.920 2850.075 1462.965 ;
        RECT 2852.070 1462.920 2852.390 1462.980 ;
        RECT 2849.785 1462.780 2852.390 1462.920 ;
        RECT 2849.785 1462.735 2850.075 1462.780 ;
        RECT 2852.070 1462.720 2852.390 1462.780 ;
        RECT 2849.785 1441.500 2850.075 1441.545 ;
        RECT 2851.610 1441.500 2851.930 1441.560 ;
        RECT 2849.785 1441.360 2851.930 1441.500 ;
        RECT 2849.785 1441.315 2850.075 1441.360 ;
        RECT 2851.610 1441.300 2851.930 1441.360 ;
        RECT 2849.770 1351.060 2850.090 1351.120 ;
        RECT 2851.150 1351.060 2851.470 1351.120 ;
        RECT 2849.770 1350.920 2851.470 1351.060 ;
        RECT 2849.770 1350.860 2850.090 1350.920 ;
        RECT 2851.150 1350.860 2851.470 1350.920 ;
        RECT 2850.230 1233.420 2850.550 1233.480 ;
        RECT 2850.035 1233.280 2850.550 1233.420 ;
        RECT 2850.230 1233.220 2850.550 1233.280 ;
        RECT 2849.770 1217.780 2850.090 1217.840 ;
        RECT 2850.245 1217.780 2850.535 1217.825 ;
        RECT 2849.770 1217.640 2850.535 1217.780 ;
        RECT 2849.770 1217.580 2850.090 1217.640 ;
        RECT 2850.245 1217.595 2850.535 1217.640 ;
        RECT 2849.770 1180.380 2850.090 1180.440 ;
        RECT 2850.245 1180.380 2850.535 1180.425 ;
        RECT 2849.770 1180.240 2850.535 1180.380 ;
        RECT 2849.770 1180.180 2850.090 1180.240 ;
        RECT 2850.245 1180.195 2850.535 1180.240 ;
        RECT 2850.230 1135.160 2850.550 1135.220 ;
        RECT 2850.035 1135.020 2850.550 1135.160 ;
        RECT 2850.230 1134.960 2850.550 1135.020 ;
        RECT 2849.770 1018.540 2850.090 1018.600 ;
        RECT 2850.245 1018.540 2850.535 1018.585 ;
        RECT 2849.770 1018.400 2850.535 1018.540 ;
        RECT 2849.770 1018.340 2850.090 1018.400 ;
        RECT 2850.245 1018.355 2850.535 1018.400 ;
        RECT 2849.770 1015.820 2850.090 1015.880 ;
        RECT 2850.245 1015.820 2850.535 1015.865 ;
        RECT 2849.770 1015.680 2850.535 1015.820 ;
        RECT 2849.770 1015.620 2850.090 1015.680 ;
        RECT 2850.245 1015.635 2850.535 1015.680 ;
        RECT 2849.770 961.080 2850.090 961.140 ;
        RECT 2850.245 961.080 2850.535 961.125 ;
        RECT 2849.770 960.940 2850.535 961.080 ;
        RECT 2849.770 960.880 2850.090 960.940 ;
        RECT 2850.245 960.895 2850.535 960.940 ;
        RECT 2849.770 942.040 2850.090 942.100 ;
        RECT 2850.245 942.040 2850.535 942.085 ;
        RECT 2849.770 941.900 2850.535 942.040 ;
        RECT 2849.770 941.840 2850.090 941.900 ;
        RECT 2850.245 941.855 2850.535 941.900 ;
        RECT 2849.770 902.260 2850.090 902.320 ;
        RECT 2850.245 902.260 2850.535 902.305 ;
        RECT 2849.770 902.120 2850.535 902.260 ;
        RECT 2849.770 902.060 2850.090 902.120 ;
        RECT 2850.245 902.075 2850.535 902.120 ;
        RECT 2849.770 884.240 2850.090 884.300 ;
        RECT 2850.245 884.240 2850.535 884.285 ;
        RECT 2849.770 884.100 2850.535 884.240 ;
        RECT 2849.770 884.040 2850.090 884.100 ;
        RECT 2850.245 884.055 2850.535 884.100 ;
        RECT 2849.770 876.080 2850.090 876.140 ;
        RECT 2851.165 876.080 2851.455 876.125 ;
        RECT 2849.770 875.940 2851.455 876.080 ;
        RECT 2849.770 875.880 2850.090 875.940 ;
        RECT 2851.165 875.895 2851.455 875.940 ;
        RECT 2850.230 810.120 2850.550 810.180 ;
        RECT 2851.165 810.120 2851.455 810.165 ;
        RECT 2850.230 809.980 2851.455 810.120 ;
        RECT 2850.230 809.920 2850.550 809.980 ;
        RECT 2851.165 809.935 2851.455 809.980 ;
        RECT 2850.230 778.160 2850.550 778.220 ;
        RECT 2851.625 778.160 2851.915 778.205 ;
        RECT 2850.230 778.020 2851.915 778.160 ;
        RECT 2850.230 777.960 2850.550 778.020 ;
        RECT 2851.625 777.975 2851.915 778.020 ;
        RECT 2850.230 769.660 2850.550 769.720 ;
        RECT 2851.625 769.660 2851.915 769.705 ;
        RECT 2850.230 769.520 2851.915 769.660 ;
        RECT 2850.230 769.460 2850.550 769.520 ;
        RECT 2851.625 769.475 2851.915 769.520 ;
        RECT 2850.230 747.900 2850.550 747.960 ;
        RECT 2852.545 747.900 2852.835 747.945 ;
        RECT 2850.230 747.760 2852.835 747.900 ;
        RECT 2850.230 747.700 2850.550 747.760 ;
        RECT 2852.545 747.715 2852.835 747.760 ;
        RECT 2849.770 734.980 2850.090 735.040 ;
        RECT 2852.545 734.980 2852.835 735.025 ;
        RECT 2849.770 734.840 2852.835 734.980 ;
        RECT 2849.770 734.780 2850.090 734.840 ;
        RECT 2852.545 734.795 2852.835 734.840 ;
        RECT 2849.770 674.600 2850.090 674.860 ;
        RECT 2849.860 673.840 2850.000 674.600 ;
        RECT 2849.770 673.580 2850.090 673.840 ;
        RECT 2849.770 382.400 2850.090 382.460 ;
        RECT 2850.690 382.400 2851.010 382.460 ;
        RECT 2849.770 382.260 2851.010 382.400 ;
        RECT 2849.770 382.200 2850.090 382.260 ;
        RECT 2850.690 382.200 2851.010 382.260 ;
        RECT 2849.770 339.560 2850.090 339.620 ;
        RECT 2850.690 339.560 2851.010 339.620 ;
        RECT 2849.770 339.420 2851.010 339.560 ;
        RECT 2849.770 339.360 2850.090 339.420 ;
        RECT 2850.690 339.360 2851.010 339.420 ;
        RECT 2849.770 324.940 2850.090 325.000 ;
        RECT 2852.085 324.940 2852.375 324.985 ;
        RECT 2849.770 324.800 2852.375 324.940 ;
        RECT 2849.770 324.740 2850.090 324.800 ;
        RECT 2852.085 324.755 2852.375 324.800 ;
        RECT 2849.770 293.660 2850.090 293.720 ;
        RECT 2852.085 293.660 2852.375 293.705 ;
        RECT 2849.770 293.520 2852.375 293.660 ;
        RECT 2849.770 293.460 2850.090 293.520 ;
        RECT 2852.085 293.475 2852.375 293.520 ;
        RECT 2850.690 155.280 2851.010 155.340 ;
        RECT 2851.625 155.280 2851.915 155.325 ;
        RECT 2850.690 155.140 2851.915 155.280 ;
        RECT 2850.690 155.080 2851.010 155.140 ;
        RECT 2851.625 155.095 2851.915 155.140 ;
        RECT 2849.770 39.340 2850.090 39.400 ;
        RECT 2851.625 39.340 2851.915 39.385 ;
        RECT 2849.770 39.200 2851.915 39.340 ;
        RECT 2849.770 39.140 2850.090 39.200 ;
        RECT 2851.625 39.155 2851.915 39.200 ;
        RECT 1250.810 8.740 1251.130 8.800 ;
        RECT 1254.045 8.740 1254.335 8.785 ;
        RECT 1250.810 8.600 1254.335 8.740 ;
        RECT 1250.810 8.540 1251.130 8.600 ;
        RECT 1254.045 8.555 1254.335 8.600 ;
        RECT 675.810 8.400 676.130 8.460 ;
        RECT 685.930 8.400 686.250 8.460 ;
        RECT 675.810 8.260 686.250 8.400 ;
        RECT 675.810 8.200 676.130 8.260 ;
        RECT 685.930 8.200 686.250 8.260 ;
        RECT 794.965 8.400 795.255 8.445 ;
        RECT 801.865 8.400 802.155 8.445 ;
        RECT 794.965 8.260 802.155 8.400 ;
        RECT 794.965 8.215 795.255 8.260 ;
        RECT 801.865 8.215 802.155 8.260 ;
        RECT 2789.970 8.400 2790.290 8.460 ;
        RECT 2848.850 8.400 2849.170 8.460 ;
        RECT 2789.970 8.260 2849.170 8.400 ;
        RECT 2789.970 8.200 2790.290 8.260 ;
        RECT 2848.850 8.200 2849.170 8.260 ;
        RECT 628.890 8.060 629.210 8.120 ;
        RECT 629.825 8.060 630.115 8.105 ;
        RECT 628.890 7.920 630.115 8.060 ;
        RECT 628.890 7.860 629.210 7.920 ;
        RECT 629.825 7.875 630.115 7.920 ;
        RECT 920.085 7.875 920.375 8.105 ;
        RECT 1170.310 8.060 1170.630 8.120 ;
        RECT 1189.630 8.060 1189.950 8.120 ;
        RECT 1170.310 7.920 1189.950 8.060 ;
        RECT 789.890 7.720 790.210 7.780 ;
        RECT 794.965 7.720 795.255 7.765 ;
        RECT 789.890 7.580 795.255 7.720 ;
        RECT 789.890 7.520 790.210 7.580 ;
        RECT 794.965 7.535 795.255 7.580 ;
        RECT 801.865 7.720 802.155 7.765 ;
        RECT 804.610 7.720 804.930 7.780 ;
        RECT 920.160 7.720 920.300 7.875 ;
        RECT 1170.310 7.860 1170.630 7.920 ;
        RECT 1189.630 7.860 1189.950 7.920 ;
        RECT 2577.910 8.060 2578.230 8.120 ;
        RECT 2644.150 8.060 2644.470 8.120 ;
        RECT 2577.910 7.920 2644.470 8.060 ;
        RECT 2577.910 7.860 2578.230 7.920 ;
        RECT 2644.150 7.860 2644.470 7.920 ;
        RECT 801.865 7.580 804.930 7.720 ;
        RECT 801.865 7.535 802.155 7.580 ;
        RECT 804.610 7.520 804.930 7.580 ;
        RECT 899.920 7.580 920.300 7.720 ;
        RECT 947.685 7.720 947.975 7.765 ;
        RECT 949.510 7.720 949.830 7.780 ;
        RECT 947.685 7.580 949.830 7.720 ;
        RECT 895.705 7.380 895.995 7.425 ;
        RECT 899.920 7.380 900.060 7.580 ;
        RECT 947.685 7.535 947.975 7.580 ;
        RECT 949.510 7.520 949.830 7.580 ;
        RECT 950.430 7.720 950.750 7.780 ;
        RECT 952.730 7.720 953.050 7.780 ;
        RECT 950.430 7.580 953.050 7.720 ;
        RECT 950.430 7.520 950.750 7.580 ;
        RECT 952.730 7.520 953.050 7.580 ;
        RECT 1302.420 7.580 1303.480 7.720 ;
        RECT 895.705 7.240 900.060 7.380 ;
        RECT 1254.045 7.380 1254.335 7.425 ;
        RECT 1302.420 7.380 1302.560 7.580 ;
        RECT 1254.045 7.240 1302.560 7.380 ;
        RECT 1303.340 7.380 1303.480 7.580 ;
        RECT 1315.210 7.380 1315.530 7.440 ;
        RECT 1303.340 7.240 1315.530 7.380 ;
        RECT 895.705 7.195 895.995 7.240 ;
        RECT 1254.045 7.195 1254.335 7.240 ;
        RECT 1315.210 7.180 1315.530 7.240 ;
        RECT 644.530 6.700 644.850 6.760 ;
        RECT 644.335 6.560 644.850 6.700 ;
        RECT 644.530 6.500 644.850 6.560 ;
        RECT 440.750 6.020 441.070 6.080 ;
        RECT 442.590 6.020 442.910 6.080 ;
        RECT 440.750 5.880 442.910 6.020 ;
        RECT 440.750 5.820 441.070 5.880 ;
        RECT 442.590 5.820 442.910 5.880 ;
        RECT 460.990 6.020 461.310 6.080 ;
        RECT 465.590 6.020 465.910 6.080 ;
        RECT 460.990 5.880 465.910 6.020 ;
        RECT 460.990 5.820 461.310 5.880 ;
        RECT 465.590 5.820 465.910 5.880 ;
        RECT 2506.610 5.340 2506.930 5.400 ;
        RECT 2563.190 5.340 2563.510 5.400 ;
        RECT 2506.610 5.200 2563.510 5.340 ;
        RECT 2506.610 5.140 2506.930 5.200 ;
        RECT 2563.190 5.140 2563.510 5.200 ;
      LAYER via ;
        RECT 2850.720 2325.980 2850.980 2326.240 ;
        RECT 2850.720 2325.300 2850.980 2325.560 ;
        RECT 2849.800 1968.980 2850.060 1969.240 ;
        RECT 2849.800 1945.180 2850.060 1945.440 ;
        RECT 2849.800 1841.480 2850.060 1841.740 ;
        RECT 2849.800 1789.120 2850.060 1789.380 ;
        RECT 2849.800 1769.740 2850.060 1770.000 ;
        RECT 2849.800 1768.040 2850.060 1768.300 ;
        RECT 2849.800 1604.840 2850.060 1605.100 ;
        RECT 2851.180 1577.300 2851.440 1577.560 ;
        RECT 2851.180 1519.160 2851.440 1519.420 ;
        RECT 2852.100 1501.820 2852.360 1502.080 ;
        RECT 2852.100 1462.720 2852.360 1462.980 ;
        RECT 2851.640 1441.300 2851.900 1441.560 ;
        RECT 2849.800 1350.860 2850.060 1351.120 ;
        RECT 2851.180 1350.860 2851.440 1351.120 ;
        RECT 2850.260 1233.220 2850.520 1233.480 ;
        RECT 2849.800 1217.580 2850.060 1217.840 ;
        RECT 2849.800 1180.180 2850.060 1180.440 ;
        RECT 2850.260 1134.960 2850.520 1135.220 ;
        RECT 2849.800 1018.340 2850.060 1018.600 ;
        RECT 2849.800 1015.620 2850.060 1015.880 ;
        RECT 2849.800 960.880 2850.060 961.140 ;
        RECT 2849.800 941.840 2850.060 942.100 ;
        RECT 2849.800 902.060 2850.060 902.320 ;
        RECT 2849.800 884.040 2850.060 884.300 ;
        RECT 2849.800 875.880 2850.060 876.140 ;
        RECT 2850.260 809.920 2850.520 810.180 ;
        RECT 2850.260 777.960 2850.520 778.220 ;
        RECT 2850.260 769.460 2850.520 769.720 ;
        RECT 2850.260 747.700 2850.520 747.960 ;
        RECT 2849.800 734.780 2850.060 735.040 ;
        RECT 2849.800 674.600 2850.060 674.860 ;
        RECT 2849.800 673.580 2850.060 673.840 ;
        RECT 2849.800 382.200 2850.060 382.460 ;
        RECT 2850.720 382.200 2850.980 382.460 ;
        RECT 2849.800 339.360 2850.060 339.620 ;
        RECT 2850.720 339.360 2850.980 339.620 ;
        RECT 2849.800 324.740 2850.060 325.000 ;
        RECT 2849.800 293.460 2850.060 293.720 ;
        RECT 2850.720 155.080 2850.980 155.340 ;
        RECT 2849.800 39.140 2850.060 39.400 ;
        RECT 1250.840 8.540 1251.100 8.800 ;
        RECT 675.840 8.200 676.100 8.460 ;
        RECT 685.960 8.200 686.220 8.460 ;
        RECT 2790.000 8.200 2790.260 8.460 ;
        RECT 2848.880 8.200 2849.140 8.460 ;
        RECT 628.920 7.860 629.180 8.120 ;
        RECT 789.920 7.520 790.180 7.780 ;
        RECT 804.640 7.520 804.900 7.780 ;
        RECT 1170.340 7.860 1170.600 8.120 ;
        RECT 1189.660 7.860 1189.920 8.120 ;
        RECT 2577.940 7.860 2578.200 8.120 ;
        RECT 2644.180 7.860 2644.440 8.120 ;
        RECT 949.540 7.520 949.800 7.780 ;
        RECT 950.460 7.520 950.720 7.780 ;
        RECT 952.760 7.520 953.020 7.780 ;
        RECT 1315.240 7.180 1315.500 7.440 ;
        RECT 644.560 6.500 644.820 6.760 ;
        RECT 440.780 5.820 441.040 6.080 ;
        RECT 442.620 5.820 442.880 6.080 ;
        RECT 461.020 5.820 461.280 6.080 ;
        RECT 465.620 5.820 465.880 6.080 ;
        RECT 2506.640 5.140 2506.900 5.400 ;
        RECT 2563.220 5.140 2563.480 5.400 ;
      LAYER met2 ;
        RECT 2851.630 2654.450 2851.910 2654.565 ;
        RECT 2850.320 2654.310 2851.910 2654.450 ;
        RECT 2850.320 2650.200 2850.460 2654.310 ;
        RECT 2851.630 2654.195 2851.910 2654.310 ;
        RECT 2848.020 2650.060 2850.460 2650.200 ;
        RECT 2848.020 2622.490 2848.160 2650.060 ;
        RECT 2848.020 2622.350 2848.620 2622.490 ;
        RECT 2848.480 2618.410 2848.620 2622.350 ;
        RECT 2847.560 2618.270 2848.620 2618.410 ;
        RECT 2847.560 2334.340 2847.700 2618.270 ;
        RECT 2849.860 2334.710 2850.920 2334.850 ;
        RECT 2849.860 2334.340 2850.000 2334.710 ;
        RECT 2847.560 2334.200 2850.000 2334.340 ;
        RECT 2850.780 2326.270 2850.920 2334.710 ;
        RECT 2850.720 2325.950 2850.980 2326.270 ;
        RECT 2850.720 2325.270 2850.980 2325.590 ;
        RECT 2850.780 2315.130 2850.920 2325.270 ;
        RECT 2850.320 2314.990 2850.920 2315.130 ;
        RECT 2850.320 2314.450 2850.460 2314.990 ;
        RECT 2847.560 2314.310 2850.460 2314.450 ;
        RECT 2847.560 1974.450 2847.700 2314.310 ;
        RECT 2847.560 1974.310 2850.000 1974.450 ;
        RECT 2849.860 1969.270 2850.000 1974.310 ;
        RECT 2849.800 1968.950 2850.060 1969.270 ;
        RECT 2849.800 1945.210 2850.060 1945.470 ;
        RECT 2847.560 1945.150 2850.060 1945.210 ;
        RECT 2847.560 1945.070 2850.000 1945.150 ;
        RECT 2847.560 1891.490 2847.700 1945.070 ;
        RECT 2847.560 1891.350 2849.080 1891.490 ;
        RECT 2848.940 1886.050 2849.080 1891.350 ;
        RECT 2847.560 1885.910 2849.080 1886.050 ;
        RECT 2847.560 1841.680 2847.700 1885.910 ;
        RECT 2849.800 1841.680 2850.060 1841.770 ;
        RECT 2847.560 1841.540 2850.060 1841.680 ;
        RECT 2849.800 1841.450 2850.060 1841.540 ;
        RECT 2849.800 1789.090 2850.060 1789.410 ;
        RECT 2849.860 1770.030 2850.000 1789.090 ;
        RECT 2849.800 1769.710 2850.060 1770.030 ;
        RECT 2849.800 1768.010 2850.060 1768.330 ;
        RECT 2849.860 1762.290 2850.000 1768.010 ;
        RECT 2849.860 1762.150 2850.460 1762.290 ;
        RECT 2850.320 1740.700 2850.460 1762.150 ;
        RECT 2847.560 1740.560 2850.460 1740.700 ;
        RECT 2847.560 1700.410 2847.700 1740.560 ;
        RECT 2847.560 1700.270 2848.620 1700.410 ;
        RECT 2848.480 1685.450 2848.620 1700.270 ;
        RECT 2847.560 1685.310 2848.620 1685.450 ;
        RECT 2847.560 1651.450 2847.700 1685.310 ;
        RECT 2847.560 1651.310 2850.460 1651.450 ;
        RECT 2850.320 1625.610 2850.460 1651.310 ;
        RECT 2849.860 1625.470 2850.460 1625.610 ;
        RECT 2849.860 1605.130 2850.000 1625.470 ;
        RECT 2849.800 1604.810 2850.060 1605.130 ;
        RECT 2851.180 1577.270 2851.440 1577.590 ;
        RECT 2851.240 1519.450 2851.380 1577.270 ;
        RECT 2851.180 1519.130 2851.440 1519.450 ;
        RECT 2852.100 1501.790 2852.360 1502.110 ;
        RECT 2852.160 1463.010 2852.300 1501.790 ;
        RECT 2852.100 1462.690 2852.360 1463.010 ;
        RECT 2851.640 1441.270 2851.900 1441.590 ;
        RECT 2851.700 1416.850 2851.840 1441.270 ;
        RECT 2850.780 1416.710 2851.840 1416.850 ;
        RECT 2850.780 1388.290 2850.920 1416.710 ;
        RECT 2850.780 1388.150 2851.380 1388.290 ;
        RECT 2851.240 1351.150 2851.380 1388.150 ;
        RECT 2849.800 1350.890 2850.060 1351.150 ;
        RECT 2847.560 1350.830 2850.060 1350.890 ;
        RECT 2851.180 1350.830 2851.440 1351.150 ;
        RECT 2847.560 1350.750 2850.000 1350.830 ;
        RECT 2847.560 1320.970 2847.700 1350.750 ;
        RECT 2847.560 1320.830 2850.460 1320.970 ;
        RECT 2850.320 1300.060 2850.460 1320.830 ;
        RECT 2848.940 1299.920 2850.460 1300.060 ;
        RECT 2848.940 1282.210 2849.080 1299.920 ;
        RECT 2848.940 1282.070 2850.000 1282.210 ;
        RECT 2849.860 1273.370 2850.000 1282.070 ;
        RECT 2849.860 1273.230 2850.460 1273.370 ;
        RECT 2850.320 1233.510 2850.460 1273.230 ;
        RECT 2850.260 1233.190 2850.520 1233.510 ;
        RECT 2849.800 1217.550 2850.060 1217.870 ;
        RECT 2849.860 1180.470 2850.000 1217.550 ;
        RECT 2849.800 1180.150 2850.060 1180.470 ;
        RECT 2850.260 1134.930 2850.520 1135.250 ;
        RECT 2850.320 1023.130 2850.460 1134.930 ;
        RECT 2849.860 1022.990 2850.460 1023.130 ;
        RECT 2849.860 1018.630 2850.000 1022.990 ;
        RECT 2849.800 1018.310 2850.060 1018.630 ;
        RECT 2849.800 1015.650 2850.060 1015.910 ;
        RECT 2847.560 1015.590 2850.060 1015.650 ;
        RECT 2847.560 1015.510 2850.000 1015.590 ;
        RECT 2847.560 961.930 2847.700 1015.510 ;
        RECT 2847.560 961.790 2848.160 961.930 ;
        RECT 2848.020 961.080 2848.160 961.790 ;
        RECT 2849.800 961.080 2850.060 961.170 ;
        RECT 2848.020 960.940 2850.060 961.080 ;
        RECT 2849.800 960.850 2850.060 960.940 ;
        RECT 2849.800 941.810 2850.060 942.130 ;
        RECT 2849.860 902.350 2850.000 941.810 ;
        RECT 2849.800 902.030 2850.060 902.350 ;
        RECT 2849.800 884.010 2850.060 884.330 ;
        RECT 2849.860 876.170 2850.000 884.010 ;
        RECT 2849.800 875.850 2850.060 876.170 ;
        RECT 2850.260 809.890 2850.520 810.210 ;
        RECT 2850.320 778.250 2850.460 809.890 ;
        RECT 2850.260 777.930 2850.520 778.250 ;
        RECT 2850.260 769.430 2850.520 769.750 ;
        RECT 2850.320 747.990 2850.460 769.430 ;
        RECT 2850.260 747.670 2850.520 747.990 ;
        RECT 2849.800 734.980 2850.060 735.070 ;
        RECT 2848.940 734.840 2850.060 734.980 ;
        RECT 2848.940 697.410 2849.080 734.840 ;
        RECT 2849.800 734.750 2850.060 734.840 ;
        RECT 2848.480 697.270 2849.080 697.410 ;
        RECT 2848.480 678.200 2848.620 697.270 ;
        RECT 2848.480 678.060 2849.540 678.200 ;
        RECT 2849.400 674.970 2849.540 678.060 ;
        RECT 2849.400 674.890 2850.000 674.970 ;
        RECT 2849.400 674.830 2850.060 674.890 ;
        RECT 2849.800 674.570 2850.060 674.830 ;
        RECT 2849.800 673.550 2850.060 673.870 ;
        RECT 2849.860 672.250 2850.000 673.550 ;
        RECT 2847.560 672.110 2850.000 672.250 ;
        RECT 2847.560 383.080 2847.700 672.110 ;
        RECT 2847.560 382.940 2848.160 383.080 ;
        RECT 2848.020 382.570 2848.160 382.940 ;
        RECT 2848.020 382.490 2850.000 382.570 ;
        RECT 2848.020 382.430 2850.060 382.490 ;
        RECT 2849.800 382.170 2850.060 382.430 ;
        RECT 2850.720 382.170 2850.980 382.490 ;
        RECT 2850.780 339.650 2850.920 382.170 ;
        RECT 2849.800 339.330 2850.060 339.650 ;
        RECT 2850.720 339.330 2850.980 339.650 ;
        RECT 2849.860 325.030 2850.000 339.330 ;
        RECT 2849.800 324.710 2850.060 325.030 ;
        RECT 2849.800 293.490 2850.060 293.750 ;
        RECT 2847.560 293.430 2850.060 293.490 ;
        RECT 2847.560 293.350 2850.000 293.430 ;
        RECT 2847.560 213.930 2847.700 293.350 ;
        RECT 2847.560 213.790 2848.620 213.930 ;
        RECT 2848.480 210.530 2848.620 213.790 ;
        RECT 2848.480 210.390 2851.380 210.530 ;
        RECT 2851.240 196.930 2851.380 210.390 ;
        RECT 2850.780 196.790 2851.380 196.930 ;
        RECT 2850.780 155.370 2850.920 196.790 ;
        RECT 2850.720 155.050 2850.980 155.370 ;
        RECT 2849.800 39.340 2850.060 39.430 ;
        RECT 2848.940 39.200 2850.060 39.340 ;
        RECT 889.740 15.340 890.000 15.600 ;
        RECT 628.910 8.315 629.190 8.685 ;
        RECT 645.010 8.570 645.290 8.685 ;
        RECT 644.620 8.430 645.290 8.570 ;
        RECT 628.980 8.150 629.120 8.315 ;
        RECT 628.920 7.830 629.180 8.150 ;
        RECT 505.630 6.955 505.910 7.325 ;
        RECT 505.700 6.700 505.840 6.955 ;
        RECT 644.620 6.790 644.760 8.430 ;
        RECT 645.010 8.315 645.290 8.430 ;
        RECT 675.830 8.315 676.110 8.685 ;
        RECT 744.830 8.570 745.110 8.685 ;
        RECT 675.840 8.170 676.100 8.315 ;
        RECT 685.960 8.170 686.220 8.490 ;
        RECT 744.830 8.430 745.500 8.570 ;
        RECT 744.830 8.315 745.110 8.430 ;
        RECT 505.700 6.645 507.220 6.700 ;
        RECT 483.090 6.530 483.370 6.645 ;
        RECT 505.700 6.560 507.290 6.645 ;
        RECT 442.680 6.390 443.740 6.530 ;
        RECT 442.680 6.110 442.820 6.390 ;
        RECT 440.780 6.020 441.040 6.110 ;
        RECT 440.380 5.880 441.040 6.020 ;
        RECT 440.380 5.170 440.520 5.880 ;
        RECT 440.780 5.790 441.040 5.880 ;
        RECT 442.620 5.790 442.880 6.110 ;
        RECT 443.600 5.850 443.740 6.390 ;
        RECT 465.680 6.390 483.370 6.530 ;
        RECT 465.680 6.110 465.820 6.390 ;
        RECT 483.090 6.275 483.370 6.390 ;
        RECT 507.010 6.275 507.290 6.560 ;
        RECT 644.560 6.470 644.820 6.790 ;
        RECT 686.020 6.645 686.160 8.170 ;
        RECT 745.360 6.645 745.500 8.430 ;
        RECT 1160.670 8.315 1160.950 8.685 ;
        RECT 1170.330 8.315 1170.610 8.685 ;
        RECT 1250.840 8.510 1251.100 8.830 ;
        RECT 806.010 7.890 806.290 8.005 ;
        RECT 804.700 7.810 806.290 7.890 ;
        RECT 789.920 7.720 790.180 7.810 ;
        RECT 789.520 7.580 790.180 7.720 ;
        RECT 685.950 6.275 686.230 6.645 ;
        RECT 745.290 6.275 745.570 6.645 ;
        RECT 461.020 5.965 461.280 6.110 ;
        RECT 453.650 5.850 453.930 5.965 ;
        RECT 443.600 5.710 453.930 5.850 ;
        RECT 453.650 5.595 453.930 5.710 ;
        RECT 461.010 5.595 461.290 5.965 ;
        RECT 465.620 5.790 465.880 6.110 ;
        RECT 789.520 5.965 789.660 7.580 ;
        RECT 789.920 7.490 790.180 7.580 ;
        RECT 804.640 7.750 806.290 7.810 ;
        RECT 804.640 7.490 804.900 7.750 ;
        RECT 806.010 7.635 806.290 7.750 ;
        RECT 857.990 7.635 858.270 8.005 ;
        RECT 953.210 7.890 953.490 8.005 ;
        RECT 952.820 7.810 953.490 7.890 ;
        RECT 858.060 7.210 858.200 7.635 ;
        RECT 949.540 7.490 949.800 7.810 ;
        RECT 950.460 7.490 950.720 7.810 ;
        RECT 952.760 7.750 953.490 7.810 ;
        RECT 952.760 7.490 953.020 7.750 ;
        RECT 953.210 7.635 953.490 7.750 ;
        RECT 866.730 7.210 867.010 7.325 ;
        RECT 858.060 7.070 867.010 7.210 ;
        RECT 949.600 7.210 949.740 7.490 ;
        RECT 950.520 7.210 950.660 7.490 ;
        RECT 949.600 7.070 950.660 7.210 ;
        RECT 866.730 6.955 867.010 7.070 ;
        RECT 1160.740 6.645 1160.880 8.315 ;
        RECT 1170.400 8.150 1170.540 8.315 ;
        RECT 1170.340 7.830 1170.600 8.150 ;
        RECT 1189.660 7.830 1189.920 8.150 ;
        RECT 1250.900 7.890 1251.040 8.510 ;
        RECT 1160.670 6.275 1160.950 6.645 ;
        RECT 551.630 5.595 551.910 5.965 ;
        RECT 558.070 5.595 558.350 5.965 ;
        RECT 789.450 5.595 789.730 5.965 ;
        RECT 439.000 5.030 440.520 5.170 ;
        RECT 430.720 3.670 437.760 3.810 ;
        RECT 430.720 2.400 430.860 3.670 ;
        RECT 437.620 3.640 437.760 3.670 ;
        RECT 439.000 3.640 439.140 5.030 ;
        RECT 551.700 5.000 551.840 5.595 ;
        RECT 558.140 5.000 558.280 5.595 ;
        RECT 1189.720 5.340 1189.860 7.830 ;
        RECT 1245.380 7.750 1251.040 7.890 ;
        RECT 1191.030 6.275 1191.310 6.645 ;
        RECT 1191.100 5.340 1191.240 6.275 ;
        RECT 1245.380 5.850 1245.520 7.750 ;
        RECT 1315.240 7.210 1315.500 7.470 ;
        RECT 1315.240 7.150 1325.100 7.210 ;
        RECT 1315.300 7.070 1325.100 7.150 ;
        RECT 1324.960 6.530 1325.100 7.070 ;
        RECT 1326.730 6.530 1327.010 6.645 ;
        RECT 1324.960 6.390 1327.010 6.530 ;
        RECT 1326.730 6.275 1327.010 6.390 ;
        RECT 1357.090 6.530 1357.370 6.645 ;
        RECT 1358.410 6.530 1358.690 9.000 ;
        RECT 1473.010 8.315 1473.290 8.685 ;
        RECT 2848.940 8.490 2849.080 39.200 ;
        RECT 2849.800 39.110 2850.060 39.200 ;
        RECT 1357.090 6.390 1358.690 6.530 ;
        RECT 1357.090 6.275 1357.370 6.390 ;
        RECT 1189.720 5.200 1191.240 5.340 ;
        RECT 1239.400 5.710 1245.520 5.850 ;
        RECT 551.700 4.860 558.280 5.000 ;
        RECT 1238.870 5.170 1239.150 5.285 ;
        RECT 1239.400 5.170 1239.540 5.710 ;
        RECT 1238.870 5.030 1239.540 5.170 ;
        RECT 1238.870 4.915 1239.150 5.030 ;
        RECT 1358.410 5.000 1358.690 6.390 ;
        RECT 1473.080 6.020 1473.220 8.315 ;
        RECT 2790.000 8.170 2790.260 8.490 ;
        RECT 2848.880 8.170 2849.140 8.490 ;
        RECT 1830.890 7.635 1831.170 8.005 ;
        RECT 2034.210 7.635 2034.490 8.005 ;
        RECT 2094.010 7.635 2094.290 8.005 ;
        RECT 2203.490 7.635 2203.770 8.005 ;
        RECT 2577.940 7.830 2578.200 8.150 ;
        RECT 2644.180 7.830 2644.440 8.150 ;
        RECT 1473.080 5.880 1474.140 6.020 ;
        RECT 1830.960 5.965 1831.100 7.635 ;
        RECT 2034.280 6.645 2034.420 7.635 ;
        RECT 2094.080 6.645 2094.220 7.635 ;
        RECT 2034.210 6.275 2034.490 6.645 ;
        RECT 2094.010 6.275 2094.290 6.645 ;
        RECT 2203.560 5.965 2203.700 7.635 ;
        RECT 2506.630 6.275 2506.910 6.645 ;
        RECT 1474.000 3.925 1474.140 5.880 ;
        RECT 1830.890 5.595 1831.170 5.965 ;
        RECT 2203.490 5.595 2203.770 5.965 ;
        RECT 2506.700 5.430 2506.840 6.275 ;
        RECT 2506.640 5.110 2506.900 5.430 ;
        RECT 2563.220 5.110 2563.480 5.430 ;
        RECT 2563.280 3.925 2563.420 5.110 ;
        RECT 2578.000 3.925 2578.140 7.830 ;
        RECT 437.620 3.500 439.140 3.640 ;
        RECT 1473.930 3.555 1474.210 3.925 ;
        RECT 2563.210 3.555 2563.490 3.925 ;
        RECT 2577.930 3.555 2578.210 3.925 ;
        RECT 430.510 -4.800 431.070 2.400 ;
        RECT 2644.240 1.885 2644.380 7.830 ;
        RECT 2693.850 6.275 2694.130 6.645 ;
        RECT 2762.390 6.275 2762.670 6.645 ;
        RECT 2693.920 1.885 2694.060 6.275 ;
        RECT 2762.460 5.850 2762.600 6.275 ;
        RECT 2790.060 5.965 2790.200 8.170 ;
        RECT 2763.770 5.850 2764.050 5.965 ;
        RECT 2762.460 5.710 2764.050 5.850 ;
        RECT 2763.770 5.595 2764.050 5.710 ;
        RECT 2789.990 5.595 2790.270 5.965 ;
        RECT 2644.170 1.515 2644.450 1.885 ;
        RECT 2693.850 1.515 2694.130 1.885 ;
      LAYER via2 ;
        RECT 2851.630 2654.240 2851.910 2654.520 ;
        RECT 628.910 8.360 629.190 8.640 ;
        RECT 505.630 7.000 505.910 7.280 ;
        RECT 645.010 8.360 645.290 8.640 ;
        RECT 675.830 8.360 676.110 8.640 ;
        RECT 744.830 8.360 745.110 8.640 ;
        RECT 483.090 6.320 483.370 6.600 ;
        RECT 507.010 6.320 507.290 6.600 ;
        RECT 1160.670 8.360 1160.950 8.640 ;
        RECT 1170.330 8.360 1170.610 8.640 ;
        RECT 685.950 6.320 686.230 6.600 ;
        RECT 745.290 6.320 745.570 6.600 ;
        RECT 453.650 5.640 453.930 5.920 ;
        RECT 461.010 5.640 461.290 5.920 ;
        RECT 806.010 7.680 806.290 7.960 ;
        RECT 857.990 7.680 858.270 7.960 ;
        RECT 953.210 7.680 953.490 7.960 ;
        RECT 866.730 7.000 867.010 7.280 ;
        RECT 1160.670 6.320 1160.950 6.600 ;
        RECT 551.630 5.640 551.910 5.920 ;
        RECT 558.070 5.640 558.350 5.920 ;
        RECT 789.450 5.640 789.730 5.920 ;
        RECT 1191.030 6.320 1191.310 6.600 ;
        RECT 1326.730 6.320 1327.010 6.600 ;
        RECT 1357.090 6.320 1357.370 6.600 ;
        RECT 1473.010 8.360 1473.290 8.640 ;
        RECT 1238.870 4.960 1239.150 5.240 ;
        RECT 1830.890 7.680 1831.170 7.960 ;
        RECT 2034.210 7.680 2034.490 7.960 ;
        RECT 2094.010 7.680 2094.290 7.960 ;
        RECT 2203.490 7.680 2203.770 7.960 ;
        RECT 2034.210 6.320 2034.490 6.600 ;
        RECT 2094.010 6.320 2094.290 6.600 ;
        RECT 2506.630 6.320 2506.910 6.600 ;
        RECT 1830.890 5.640 1831.170 5.920 ;
        RECT 2203.490 5.640 2203.770 5.920 ;
        RECT 1473.930 3.600 1474.210 3.880 ;
        RECT 2563.210 3.600 2563.490 3.880 ;
        RECT 2577.930 3.600 2578.210 3.880 ;
        RECT 2693.850 6.320 2694.130 6.600 ;
        RECT 2762.390 6.320 2762.670 6.600 ;
        RECT 2763.770 5.640 2764.050 5.920 ;
        RECT 2789.990 5.640 2790.270 5.920 ;
        RECT 2644.170 1.560 2644.450 1.840 ;
        RECT 2693.850 1.560 2694.130 1.840 ;
      LAYER met3 ;
        RECT 2851.000 2657.040 2855.000 2657.640 ;
        RECT 2851.390 2654.545 2851.690 2657.040 ;
        RECT 2851.390 2654.230 2851.935 2654.545 ;
        RECT 2851.605 2654.215 2851.935 2654.230 ;
        RECT 622.190 8.650 622.570 8.660 ;
        RECT 628.885 8.650 629.215 8.665 ;
        RECT 622.190 8.350 629.215 8.650 ;
        RECT 622.190 8.340 622.570 8.350 ;
        RECT 628.885 8.335 629.215 8.350 ;
        RECT 644.985 8.650 645.315 8.665 ;
        RECT 675.805 8.650 676.135 8.665 ;
        RECT 644.985 8.350 676.135 8.650 ;
        RECT 644.985 8.335 645.315 8.350 ;
        RECT 675.805 8.335 676.135 8.350 ;
        RECT 740.870 8.650 741.250 8.660 ;
        RECT 744.805 8.650 745.135 8.665 ;
        RECT 740.870 8.350 745.135 8.650 ;
        RECT 740.870 8.340 741.250 8.350 ;
        RECT 744.805 8.335 745.135 8.350 ;
        RECT 961.670 8.650 962.050 8.660 ;
        RECT 973.630 8.650 974.010 8.660 ;
        RECT 961.670 8.350 974.010 8.650 ;
        RECT 961.670 8.340 962.050 8.350 ;
        RECT 973.630 8.340 974.010 8.350 ;
        RECT 1160.645 8.650 1160.975 8.665 ;
        RECT 1170.305 8.650 1170.635 8.665 ;
        RECT 1160.645 8.350 1170.635 8.650 ;
        RECT 1160.645 8.335 1160.975 8.350 ;
        RECT 1170.305 8.335 1170.635 8.350 ;
        RECT 1472.270 8.650 1472.650 8.660 ;
        RECT 1472.985 8.650 1473.315 8.665 ;
        RECT 1472.270 8.350 1473.315 8.650 ;
        RECT 1472.270 8.340 1472.650 8.350 ;
        RECT 1472.985 8.335 1473.315 8.350 ;
        RECT 729.830 7.970 730.210 7.980 ;
        RECT 736.270 7.970 736.650 7.980 ;
        RECT 729.830 7.670 736.650 7.970 ;
        RECT 729.830 7.660 730.210 7.670 ;
        RECT 736.270 7.660 736.650 7.670 ;
        RECT 805.985 7.970 806.315 7.985 ;
        RECT 846.670 7.970 847.050 7.980 ;
        RECT 805.985 7.670 847.050 7.970 ;
        RECT 805.985 7.655 806.315 7.670 ;
        RECT 846.670 7.660 847.050 7.670 ;
        RECT 855.870 7.970 856.250 7.980 ;
        RECT 857.965 7.970 858.295 7.985 ;
        RECT 855.870 7.670 858.295 7.970 ;
        RECT 855.870 7.660 856.250 7.670 ;
        RECT 857.965 7.655 858.295 7.670 ;
        RECT 953.185 7.970 953.515 7.985 ;
        RECT 979.150 7.970 979.530 7.980 ;
        RECT 953.185 7.670 979.530 7.970 ;
        RECT 953.185 7.655 953.515 7.670 ;
        RECT 979.150 7.660 979.530 7.670 ;
        RECT 1830.865 7.970 1831.195 7.985 ;
        RECT 2034.185 7.970 2034.515 7.985 ;
        RECT 1830.865 7.670 2034.515 7.970 ;
        RECT 1830.865 7.655 1831.195 7.670 ;
        RECT 2034.185 7.655 2034.515 7.670 ;
        RECT 2093.985 7.970 2094.315 7.985 ;
        RECT 2203.465 7.970 2203.795 7.985 ;
        RECT 2093.985 7.670 2203.795 7.970 ;
        RECT 2093.985 7.655 2094.315 7.670 ;
        RECT 2203.465 7.655 2203.795 7.670 ;
        RECT 505.605 7.300 505.935 7.305 ;
        RECT 505.350 7.290 505.935 7.300 ;
        RECT 866.705 7.290 867.035 7.305 ;
        RECT 884.390 7.290 884.770 7.300 ;
        RECT 505.350 6.990 506.160 7.290 ;
        RECT 866.705 6.990 884.770 7.290 ;
        RECT 505.350 6.980 505.935 6.990 ;
        RECT 505.605 6.975 505.935 6.980 ;
        RECT 866.705 6.975 867.035 6.990 ;
        RECT 884.390 6.980 884.770 6.990 ;
        RECT 987.430 7.290 987.810 7.300 ;
        RECT 993.870 7.290 994.250 7.300 ;
        RECT 987.430 6.990 994.250 7.290 ;
        RECT 987.430 6.980 987.810 6.990 ;
        RECT 993.870 6.980 994.250 6.990 ;
        RECT 483.065 6.610 483.395 6.625 ;
        RECT 488.790 6.610 489.170 6.620 ;
        RECT 483.065 6.310 489.170 6.610 ;
        RECT 483.065 6.295 483.395 6.310 ;
        RECT 488.790 6.300 489.170 6.310 ;
        RECT 506.985 6.610 507.315 6.625 ;
        RECT 510.870 6.610 511.250 6.620 ;
        RECT 506.985 6.310 511.250 6.610 ;
        RECT 506.985 6.295 507.315 6.310 ;
        RECT 510.870 6.300 511.250 6.310 ;
        RECT 685.925 6.610 686.255 6.625 ;
        RECT 705.910 6.610 706.290 6.620 ;
        RECT 685.925 6.310 706.290 6.610 ;
        RECT 685.925 6.295 686.255 6.310 ;
        RECT 705.910 6.300 706.290 6.310 ;
        RECT 745.265 6.610 745.595 6.625 ;
        RECT 918.430 6.610 918.810 6.620 ;
        RECT 745.265 6.310 757.540 6.610 ;
        RECT 745.265 6.295 745.595 6.310 ;
        RECT 453.625 5.930 453.955 5.945 ;
        RECT 460.985 5.930 461.315 5.945 ;
        RECT 453.625 5.630 461.315 5.930 ;
        RECT 453.625 5.615 453.955 5.630 ;
        RECT 460.985 5.615 461.315 5.630 ;
        RECT 537.550 5.930 537.930 5.940 ;
        RECT 551.605 5.930 551.935 5.945 ;
        RECT 558.045 5.940 558.375 5.945 ;
        RECT 537.550 5.630 551.935 5.930 ;
        RECT 537.550 5.620 537.930 5.630 ;
        RECT 551.605 5.615 551.935 5.630 ;
        RECT 557.790 5.930 558.375 5.940 ;
        RECT 757.240 5.930 757.540 6.310 ;
        RECT 913.870 6.310 918.810 6.610 ;
        RECT 789.425 5.930 789.755 5.945 ;
        RECT 557.790 5.630 558.600 5.930 ;
        RECT 757.240 5.630 789.755 5.930 ;
        RECT 557.790 5.620 558.375 5.630 ;
        RECT 558.045 5.615 558.375 5.620 ;
        RECT 789.425 5.615 789.755 5.630 ;
        RECT 904.630 5.930 905.010 5.940 ;
        RECT 913.870 5.930 914.170 6.310 ;
        RECT 918.430 6.300 918.810 6.310 ;
        RECT 1146.590 6.610 1146.970 6.620 ;
        RECT 1160.645 6.610 1160.975 6.625 ;
        RECT 1146.590 6.310 1160.975 6.610 ;
        RECT 1146.590 6.300 1146.970 6.310 ;
        RECT 1160.645 6.295 1160.975 6.310 ;
        RECT 1191.005 6.610 1191.335 6.625 ;
        RECT 1227.550 6.610 1227.930 6.620 ;
        RECT 1191.005 6.310 1227.930 6.610 ;
        RECT 1191.005 6.295 1191.335 6.310 ;
        RECT 1227.550 6.300 1227.930 6.310 ;
        RECT 1326.705 6.610 1327.035 6.625 ;
        RECT 1357.065 6.610 1357.395 6.625 ;
        RECT 1326.705 6.310 1357.395 6.610 ;
        RECT 1326.705 6.295 1327.035 6.310 ;
        RECT 1357.065 6.295 1357.395 6.310 ;
        RECT 2034.185 6.610 2034.515 6.625 ;
        RECT 2093.985 6.610 2094.315 6.625 ;
        RECT 2506.605 6.610 2506.935 6.625 ;
        RECT 2034.185 6.310 2094.315 6.610 ;
        RECT 2034.185 6.295 2034.515 6.310 ;
        RECT 2093.985 6.295 2094.315 6.310 ;
        RECT 2411.630 6.310 2506.935 6.610 ;
        RECT 904.630 5.630 914.170 5.930 ;
        RECT 1744.590 5.930 1744.970 5.940 ;
        RECT 1830.865 5.930 1831.195 5.945 ;
        RECT 1744.590 5.630 1831.195 5.930 ;
        RECT 904.630 5.620 905.010 5.630 ;
        RECT 1744.590 5.620 1744.970 5.630 ;
        RECT 1830.865 5.615 1831.195 5.630 ;
        RECT 2203.465 5.930 2203.795 5.945 ;
        RECT 2411.630 5.930 2411.930 6.310 ;
        RECT 2506.605 6.295 2506.935 6.310 ;
        RECT 2693.825 6.610 2694.155 6.625 ;
        RECT 2762.365 6.610 2762.695 6.625 ;
        RECT 2693.825 6.310 2762.695 6.610 ;
        RECT 2693.825 6.295 2694.155 6.310 ;
        RECT 2762.365 6.295 2762.695 6.310 ;
        RECT 2203.465 5.630 2411.930 5.930 ;
        RECT 2763.745 5.930 2764.075 5.945 ;
        RECT 2789.965 5.930 2790.295 5.945 ;
        RECT 2763.745 5.630 2790.295 5.930 ;
        RECT 2203.465 5.615 2203.795 5.630 ;
        RECT 2763.745 5.615 2764.075 5.630 ;
        RECT 2789.965 5.615 2790.295 5.630 ;
        RECT 1237.670 5.250 1238.050 5.260 ;
        RECT 1238.845 5.250 1239.175 5.265 ;
        RECT 1237.670 4.950 1239.175 5.250 ;
        RECT 1237.670 4.940 1238.050 4.950 ;
        RECT 1238.845 4.935 1239.175 4.950 ;
        RECT 1473.905 3.900 1474.235 3.905 ;
        RECT 1473.905 3.890 1474.490 3.900 ;
        RECT 1473.680 3.590 1474.490 3.890 ;
        RECT 1473.905 3.580 1474.490 3.590 ;
        RECT 2563.185 3.890 2563.515 3.905 ;
        RECT 2577.905 3.890 2578.235 3.905 ;
        RECT 2563.185 3.590 2578.235 3.890 ;
        RECT 1473.905 3.575 1474.235 3.580 ;
        RECT 2563.185 3.575 2563.515 3.590 ;
        RECT 2577.905 3.575 2578.235 3.590 ;
        RECT 1052.750 3.210 1053.130 3.220 ;
        RECT 1056.430 3.210 1056.810 3.220 ;
        RECT 1052.750 2.910 1056.810 3.210 ;
        RECT 1052.750 2.900 1053.130 2.910 ;
        RECT 1056.430 2.900 1056.810 2.910 ;
        RECT 2644.145 1.850 2644.475 1.865 ;
        RECT 2693.825 1.850 2694.155 1.865 ;
        RECT 2644.145 1.550 2694.155 1.850 ;
        RECT 2644.145 1.535 2644.475 1.550 ;
        RECT 2693.825 1.535 2694.155 1.550 ;
      LAYER via3 ;
        RECT 622.220 8.340 622.540 8.660 ;
        RECT 740.900 8.340 741.220 8.660 ;
        RECT 961.700 8.340 962.020 8.660 ;
        RECT 973.660 8.340 973.980 8.660 ;
        RECT 1472.300 8.340 1472.620 8.660 ;
        RECT 729.860 7.660 730.180 7.980 ;
        RECT 736.300 7.660 736.620 7.980 ;
        RECT 846.700 7.660 847.020 7.980 ;
        RECT 855.900 7.660 856.220 7.980 ;
        RECT 979.180 7.660 979.500 7.980 ;
        RECT 505.380 6.980 505.700 7.300 ;
        RECT 884.420 6.980 884.740 7.300 ;
        RECT 987.460 6.980 987.780 7.300 ;
        RECT 993.900 6.980 994.220 7.300 ;
        RECT 488.820 6.300 489.140 6.620 ;
        RECT 510.900 6.300 511.220 6.620 ;
        RECT 705.940 6.300 706.260 6.620 ;
        RECT 537.580 5.620 537.900 5.940 ;
        RECT 557.820 5.620 558.140 5.940 ;
        RECT 904.660 5.620 904.980 5.940 ;
        RECT 918.460 6.300 918.780 6.620 ;
        RECT 1146.620 6.300 1146.940 6.620 ;
        RECT 1227.580 6.300 1227.900 6.620 ;
        RECT 1744.620 5.620 1744.940 5.940 ;
        RECT 1237.700 4.940 1238.020 5.260 ;
        RECT 1474.140 3.580 1474.460 3.900 ;
        RECT 1052.780 2.900 1053.100 3.220 ;
        RECT 1056.460 2.900 1056.780 3.220 ;
      LAYER met4 ;
        RECT 977.830 14.710 979.010 15.890 ;
        RECT 1125.030 14.710 1126.210 15.890 ;
        RECT 1134.230 14.710 1135.410 15.890 ;
        RECT 1471.870 14.710 1473.050 15.890 ;
        RECT 1683.470 14.710 1684.650 15.890 ;
        RECT 1744.190 14.710 1745.370 15.890 ;
        RECT 846.710 9.030 850.690 9.330 ;
        RECT 622.215 8.650 622.545 8.665 ;
        RECT 740.895 8.650 741.225 8.665 ;
        RECT 614.870 8.350 622.545 8.650 ;
        RECT 614.870 7.970 615.170 8.350 ;
        RECT 622.215 8.335 622.545 8.350 ;
        RECT 712.390 8.350 725.570 8.650 ;
        RECT 557.830 7.670 615.170 7.970 ;
        RECT 505.375 7.290 505.705 7.305 ;
        RECT 488.830 6.990 505.705 7.290 ;
        RECT 488.830 6.625 489.130 6.990 ;
        RECT 505.375 6.975 505.705 6.990 ;
        RECT 488.815 6.295 489.145 6.625 ;
        RECT 510.895 6.295 511.225 6.625 ;
        RECT 510.910 5.930 511.210 6.295 ;
        RECT 557.830 5.945 558.130 7.670 ;
        RECT 712.390 7.290 712.690 8.350 ;
        RECT 725.270 7.970 725.570 8.350 ;
        RECT 736.310 8.350 741.225 8.650 ;
        RECT 736.310 7.985 736.610 8.350 ;
        RECT 740.895 8.335 741.225 8.350 ;
        RECT 846.710 7.985 847.010 9.030 ;
        RECT 729.855 7.970 730.185 7.985 ;
        RECT 725.270 7.670 730.185 7.970 ;
        RECT 729.855 7.655 730.185 7.670 ;
        RECT 736.295 7.655 736.625 7.985 ;
        RECT 846.695 7.655 847.025 7.985 ;
        RECT 850.390 7.970 850.690 9.030 ;
        RECT 925.830 9.030 939.010 9.330 ;
        RECT 855.895 7.970 856.225 7.985 ;
        RECT 850.390 7.670 856.225 7.970 ;
        RECT 855.895 7.655 856.225 7.670 ;
        RECT 705.950 6.990 712.690 7.290 ;
        RECT 705.950 6.625 706.250 6.990 ;
        RECT 884.415 6.975 884.745 7.305 ;
        RECT 925.830 7.290 926.130 9.030 ;
        RECT 938.710 8.650 939.010 9.030 ;
        RECT 961.695 8.650 962.025 8.665 ;
        RECT 938.710 8.350 962.025 8.650 ;
        RECT 961.695 8.335 962.025 8.350 ;
        RECT 973.655 8.335 973.985 8.665 ;
        RECT 978.270 8.650 978.570 14.710 ;
        RECT 1125.470 12.050 1125.770 14.710 ;
        RECT 1134.670 12.050 1134.970 14.710 ;
        RECT 1125.470 11.750 1128.530 12.050 ;
        RECT 975.510 8.350 978.570 8.650 ;
        RECT 973.670 7.970 973.970 8.335 ;
        RECT 975.510 7.970 975.810 8.350 ;
        RECT 973.670 7.670 975.810 7.970 ;
        RECT 979.175 7.655 979.505 7.985 ;
        RECT 1090.510 7.670 1092.650 7.970 ;
        RECT 918.470 6.990 926.130 7.290 ;
        RECT 979.190 7.290 979.490 7.655 ;
        RECT 987.455 7.290 987.785 7.305 ;
        RECT 979.190 6.990 987.785 7.290 ;
        RECT 705.935 6.295 706.265 6.625 ;
        RECT 537.575 5.930 537.905 5.945 ;
        RECT 510.910 5.630 523.170 5.930 ;
        RECT 522.870 2.290 523.170 5.630 ;
        RECT 536.670 5.630 537.905 5.930 ;
        RECT 536.670 5.250 536.970 5.630 ;
        RECT 537.575 5.615 537.905 5.630 ;
        RECT 557.815 5.615 558.145 5.945 ;
        RECT 884.430 5.930 884.730 6.975 ;
        RECT 918.470 6.625 918.770 6.990 ;
        RECT 987.455 6.975 987.785 6.990 ;
        RECT 993.895 6.975 994.225 7.305 ;
        RECT 1090.510 7.290 1090.810 7.670 ;
        RECT 1086.830 6.990 1090.810 7.290 ;
        RECT 918.455 6.295 918.785 6.625 ;
        RECT 993.910 6.610 994.210 6.975 ;
        RECT 993.910 6.310 1047.570 6.610 ;
        RECT 904.655 5.930 904.985 5.945 ;
        RECT 884.430 5.630 904.985 5.930 ;
        RECT 904.655 5.615 904.985 5.630 ;
        RECT 533.910 4.950 536.970 5.250 ;
        RECT 533.910 2.290 534.210 4.950 ;
        RECT 1047.270 2.530 1047.570 6.310 ;
        RECT 1052.775 2.895 1053.105 3.225 ;
        RECT 1056.455 2.895 1056.785 3.225 ;
        RECT 1052.790 2.530 1053.090 2.895 ;
        RECT 522.430 1.110 523.610 2.290 ;
        RECT 533.470 1.110 534.650 2.290 ;
        RECT 1047.270 2.230 1053.090 2.530 ;
        RECT 1056.470 2.530 1056.770 2.895 ;
        RECT 1086.830 2.530 1087.130 6.990 ;
        RECT 1092.350 3.890 1092.650 7.670 ;
        RECT 1105.230 6.310 1126.690 6.610 ;
        RECT 1105.230 3.890 1105.530 6.310 ;
        RECT 1126.390 5.250 1126.690 6.310 ;
        RECT 1128.230 5.250 1128.530 11.750 ;
        RECT 1130.990 11.750 1134.970 12.050 ;
        RECT 1130.990 6.610 1131.290 11.750 ;
        RECT 1472.310 8.665 1472.610 14.710 ;
        RECT 1472.295 8.335 1472.625 8.665 ;
        RECT 1227.590 6.990 1231.570 7.290 ;
        RECT 1227.590 6.625 1227.890 6.990 ;
        RECT 1130.990 6.310 1134.970 6.610 ;
        RECT 1134.670 5.250 1134.970 6.310 ;
        RECT 1146.615 6.295 1146.945 6.625 ;
        RECT 1227.575 6.295 1227.905 6.625 ;
        RECT 1126.390 4.950 1134.970 5.250 ;
        RECT 1092.350 3.590 1105.530 3.890 ;
        RECT 1128.230 3.890 1128.530 4.950 ;
        RECT 1146.630 3.890 1146.930 6.295 ;
        RECT 1128.230 3.590 1146.930 3.890 ;
        RECT 1056.470 2.230 1057.460 2.530 ;
        RECT 1057.160 1.850 1057.460 2.230 ;
        RECT 1070.270 2.230 1087.130 2.530 ;
        RECT 1070.270 1.850 1070.570 2.230 ;
        RECT 1057.160 1.550 1070.570 1.850 ;
        RECT 1231.270 1.850 1231.570 6.990 ;
        RECT 1237.695 5.250 1238.025 5.265 ;
        RECT 1234.950 4.950 1238.025 5.250 ;
        RECT 1234.950 1.850 1235.250 4.950 ;
        RECT 1237.695 4.935 1238.025 4.950 ;
        RECT 1474.135 3.575 1474.465 3.905 ;
        RECT 1474.150 2.290 1474.450 3.575 ;
        RECT 1683.910 2.290 1684.210 14.710 ;
        RECT 1744.630 5.945 1744.930 14.710 ;
        RECT 1744.615 5.615 1744.945 5.945 ;
        RECT 1231.270 1.550 1235.250 1.850 ;
        RECT 1473.710 1.110 1474.890 2.290 ;
        RECT 1683.470 1.110 1684.650 2.290 ;
      LAYER met5 ;
        RECT 1014.420 21.300 1106.180 22.900 ;
        RECT 1014.420 19.500 1016.020 21.300 ;
        RECT 978.540 17.900 1016.020 19.500 ;
        RECT 1104.580 19.500 1106.180 21.300 ;
        RECT 1134.940 21.300 1297.540 22.900 ;
        RECT 1134.940 19.500 1136.540 21.300 ;
        RECT 1104.580 17.900 1126.420 19.500 ;
        RECT 978.540 16.100 980.140 17.900 ;
        RECT 977.620 14.500 980.140 16.100 ;
        RECT 1124.820 14.500 1126.420 17.900 ;
        RECT 1134.020 17.900 1136.540 19.500 ;
        RECT 1295.940 19.500 1297.540 21.300 ;
        RECT 1295.940 17.900 1308.810 19.500 ;
        RECT 1134.020 14.500 1135.620 17.900 ;
        RECT 1307.210 16.100 1308.810 17.900 ;
        RECT 1683.260 17.900 1745.580 19.500 ;
        RECT 1307.210 14.500 1473.260 16.100 ;
        RECT 1683.260 14.500 1684.860 17.900 ;
        RECT 1743.980 14.500 1745.580 17.900 ;
        RECT 522.220 0.900 534.860 2.500 ;
        RECT 1473.500 0.900 1684.860 2.500 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 957.405 9.265 986.555 9.435 ;
        RECT 918.305 3.825 921.235 3.995 ;
        RECT 921.065 3.315 921.235 3.825 ;
        RECT 957.405 3.655 957.575 9.265 ;
        RECT 986.385 7.735 986.555 9.265 ;
        RECT 986.385 7.565 989.775 7.735 ;
        RECT 953.265 3.485 957.575 3.655 ;
        RECT 953.265 3.315 953.435 3.485 ;
        RECT 921.065 3.145 953.435 3.315 ;
      LAYER mcon ;
        RECT 989.605 7.565 989.775 7.735 ;
      LAYER met1 ;
        RECT 1200.670 8.740 1200.990 8.800 ;
        RECT 1207.570 8.740 1207.890 8.800 ;
        RECT 1200.670 8.600 1207.890 8.740 ;
        RECT 1200.670 8.540 1200.990 8.600 ;
        RECT 1207.570 8.540 1207.890 8.600 ;
        RECT 1268.290 8.740 1268.610 8.800 ;
        RECT 1285.310 8.740 1285.630 8.800 ;
        RECT 1268.290 8.600 1285.630 8.740 ;
        RECT 1268.290 8.540 1268.610 8.600 ;
        RECT 1285.310 8.540 1285.630 8.600 ;
        RECT 1083.830 8.400 1084.150 8.460 ;
        RECT 1100.850 8.400 1101.170 8.460 ;
        RECT 1083.830 8.260 1101.170 8.400 ;
        RECT 1083.830 8.200 1084.150 8.260 ;
        RECT 1100.850 8.200 1101.170 8.260 ;
        RECT 1303.710 8.400 1304.030 8.460 ;
        RECT 1306.470 8.400 1306.790 8.460 ;
        RECT 1303.710 8.260 1306.790 8.400 ;
        RECT 1303.710 8.200 1304.030 8.260 ;
        RECT 1306.470 8.200 1306.790 8.260 ;
        RECT 989.545 7.720 989.835 7.765 ;
        RECT 992.750 7.720 993.070 7.780 ;
        RECT 989.545 7.580 993.070 7.720 ;
        RECT 989.545 7.535 989.835 7.580 ;
        RECT 992.750 7.520 993.070 7.580 ;
        RECT 918.245 3.980 918.535 4.025 ;
        RECT 882.440 3.840 918.535 3.980 ;
        RECT 816.110 3.640 816.430 3.700 ;
        RECT 819.330 3.640 819.650 3.700 ;
        RECT 816.110 3.500 819.650 3.640 ;
        RECT 816.110 3.440 816.430 3.500 ;
        RECT 819.330 3.440 819.650 3.500 ;
        RECT 880.050 3.640 880.370 3.700 ;
        RECT 882.440 3.640 882.580 3.840 ;
        RECT 918.245 3.795 918.535 3.840 ;
        RECT 880.050 3.500 882.580 3.640 ;
        RECT 880.050 3.440 880.370 3.500 ;
      LAYER via ;
        RECT 1200.700 8.540 1200.960 8.800 ;
        RECT 1207.600 8.540 1207.860 8.800 ;
        RECT 1268.320 8.540 1268.580 8.800 ;
        RECT 1285.340 8.540 1285.600 8.800 ;
        RECT 1083.860 8.200 1084.120 8.460 ;
        RECT 1100.880 8.200 1101.140 8.460 ;
        RECT 1303.740 8.200 1304.000 8.460 ;
        RECT 1306.500 8.200 1306.760 8.460 ;
        RECT 992.780 7.520 993.040 7.780 ;
        RECT 816.140 3.440 816.400 3.700 ;
        RECT 819.360 3.440 819.620 3.700 ;
        RECT 880.080 3.440 880.340 3.700 ;
      LAYER met2 ;
        RECT 1000.130 8.570 1000.410 8.685 ;
        RECT 994.220 8.430 1000.410 8.570 ;
        RECT 992.780 7.720 993.040 7.810 ;
        RECT 994.220 7.720 994.360 8.430 ;
        RECT 1000.130 8.315 1000.410 8.430 ;
        RECT 1036.470 8.570 1036.750 8.685 ;
        RECT 1040.610 8.570 1040.890 8.685 ;
        RECT 1036.470 8.430 1040.890 8.570 ;
        RECT 1036.470 8.315 1036.750 8.430 ;
        RECT 1040.610 8.315 1040.890 8.430 ;
        RECT 1083.390 8.570 1083.670 8.685 ;
        RECT 1102.250 8.570 1102.530 8.685 ;
        RECT 1083.390 8.490 1084.060 8.570 ;
        RECT 1100.940 8.490 1102.530 8.570 ;
        RECT 1083.390 8.430 1084.120 8.490 ;
        RECT 1083.390 8.315 1083.670 8.430 ;
        RECT 1083.860 8.170 1084.120 8.430 ;
        RECT 1100.880 8.430 1102.530 8.490 ;
        RECT 1100.880 8.170 1101.140 8.430 ;
        RECT 1102.250 8.315 1102.530 8.430 ;
        RECT 1191.950 8.570 1192.230 8.685 ;
        RECT 1200.700 8.570 1200.960 8.830 ;
        RECT 1191.950 8.510 1200.960 8.570 ;
        RECT 1207.600 8.570 1207.860 8.830 ;
        RECT 1207.600 8.510 1212.400 8.570 ;
        RECT 1268.320 8.510 1268.580 8.830 ;
        RECT 1285.340 8.510 1285.600 8.830 ;
        RECT 1191.950 8.430 1200.900 8.510 ;
        RECT 1207.660 8.430 1212.400 8.510 ;
        RECT 1191.950 8.315 1192.230 8.430 ;
        RECT 992.780 7.580 994.360 7.720 ;
        RECT 992.780 7.490 993.040 7.580 ;
        RECT 1212.260 4.660 1212.400 8.430 ;
        RECT 1226.450 7.210 1226.730 7.325 ;
        RECT 1216.400 7.070 1226.730 7.210 ;
        RECT 1216.400 4.660 1216.540 7.070 ;
        RECT 1226.450 6.955 1226.730 7.070 ;
        RECT 457.330 4.235 457.610 4.605 ;
        RECT 1212.260 4.520 1216.540 4.660 ;
        RECT 1268.380 4.605 1268.520 8.510 ;
        RECT 1285.400 7.325 1285.540 8.510 ;
        RECT 1293.680 8.490 1303.940 8.570 ;
        RECT 1293.680 8.430 1304.000 8.490 ;
        RECT 1293.680 7.890 1293.820 8.430 ;
        RECT 1303.740 8.170 1304.000 8.430 ;
        RECT 1306.500 8.170 1306.760 8.490 ;
        RECT 1290.460 7.750 1293.820 7.890 ;
        RECT 1306.560 7.890 1306.700 8.170 ;
        RECT 1310.170 7.890 1310.450 8.005 ;
        RECT 1306.560 7.750 1310.450 7.890 ;
        RECT 1290.460 7.325 1290.600 7.750 ;
        RECT 1310.170 7.635 1310.450 7.750 ;
        RECT 1354.790 7.635 1355.070 8.005 ;
        RECT 1285.330 6.955 1285.610 7.325 ;
        RECT 1290.390 6.955 1290.670 7.325 ;
        RECT 1354.860 7.210 1355.000 7.635 ;
        RECT 1356.170 7.210 1356.450 7.325 ;
        RECT 1354.860 7.070 1356.450 7.210 ;
        RECT 1356.170 6.955 1356.450 7.070 ;
        RECT 1402.700 7.070 1404.680 7.210 ;
        RECT 1402.700 6.645 1402.840 7.070 ;
        RECT 1402.630 6.275 1402.910 6.645 ;
        RECT 1404.540 5.850 1404.680 7.070 ;
        RECT 1405.790 5.850 1406.070 9.000 ;
        RECT 1404.540 5.710 1406.070 5.850 ;
        RECT 1405.790 5.000 1406.070 5.710 ;
        RECT 1262.330 4.235 1262.610 4.605 ;
        RECT 1264.630 4.490 1264.910 4.605 ;
        RECT 1263.780 4.350 1264.910 4.490 ;
        RECT 457.400 3.640 457.540 4.235 ;
        RECT 448.660 3.500 457.540 3.640 ;
        RECT 807.390 3.810 807.670 3.925 ;
        RECT 808.770 3.810 809.050 3.925 ;
        RECT 807.390 3.670 809.050 3.810 ;
        RECT 807.390 3.555 807.670 3.670 ;
        RECT 808.770 3.555 809.050 3.670 ;
        RECT 815.670 3.810 815.950 3.925 ;
        RECT 815.670 3.730 816.340 3.810 ;
        RECT 815.670 3.670 816.400 3.730 ;
        RECT 815.670 3.555 815.950 3.670 ;
        RECT 448.660 2.400 448.800 3.500 ;
        RECT 816.140 3.410 816.400 3.670 ;
        RECT 819.350 3.555 819.630 3.925 ;
        RECT 880.070 3.555 880.350 3.925 ;
        RECT 1262.400 3.810 1262.540 4.235 ;
        RECT 1263.780 3.810 1263.920 4.350 ;
        RECT 1264.630 4.235 1264.910 4.350 ;
        RECT 1268.310 4.235 1268.590 4.605 ;
        RECT 1262.400 3.670 1263.920 3.810 ;
        RECT 819.360 3.410 819.620 3.555 ;
        RECT 880.080 3.410 880.340 3.555 ;
        RECT 448.450 -4.800 449.010 2.400 ;
      LAYER via2 ;
        RECT 1000.130 8.360 1000.410 8.640 ;
        RECT 1036.470 8.360 1036.750 8.640 ;
        RECT 1040.610 8.360 1040.890 8.640 ;
        RECT 1083.390 8.360 1083.670 8.640 ;
        RECT 1102.250 8.360 1102.530 8.640 ;
        RECT 1191.950 8.360 1192.230 8.640 ;
        RECT 1226.450 7.000 1226.730 7.280 ;
        RECT 457.330 4.280 457.610 4.560 ;
        RECT 1310.170 7.680 1310.450 7.960 ;
        RECT 1354.790 7.680 1355.070 7.960 ;
        RECT 1285.330 7.000 1285.610 7.280 ;
        RECT 1290.390 7.000 1290.670 7.280 ;
        RECT 1356.170 7.000 1356.450 7.280 ;
        RECT 1402.630 6.320 1402.910 6.600 ;
        RECT 1262.330 4.280 1262.610 4.560 ;
        RECT 807.390 3.600 807.670 3.880 ;
        RECT 808.770 3.600 809.050 3.880 ;
        RECT 815.670 3.600 815.950 3.880 ;
        RECT 819.350 3.600 819.630 3.880 ;
        RECT 880.070 3.600 880.350 3.880 ;
        RECT 1264.630 4.280 1264.910 4.560 ;
        RECT 1268.310 4.280 1268.590 4.560 ;
      LAYER met3 ;
        RECT 1000.105 8.650 1000.435 8.665 ;
        RECT 1036.445 8.650 1036.775 8.665 ;
        RECT 1000.105 8.350 1036.775 8.650 ;
        RECT 1000.105 8.335 1000.435 8.350 ;
        RECT 1036.445 8.335 1036.775 8.350 ;
        RECT 1040.585 8.650 1040.915 8.665 ;
        RECT 1083.365 8.650 1083.695 8.665 ;
        RECT 1040.585 8.350 1083.695 8.650 ;
        RECT 1040.585 8.335 1040.915 8.350 ;
        RECT 1083.365 8.335 1083.695 8.350 ;
        RECT 1102.225 8.650 1102.555 8.665 ;
        RECT 1191.925 8.650 1192.255 8.665 ;
        RECT 1102.225 8.350 1159.810 8.650 ;
        RECT 1102.225 8.335 1102.555 8.350 ;
        RECT 1159.510 7.970 1159.810 8.350 ;
        RECT 1190.790 8.350 1192.255 8.650 ;
        RECT 1190.790 7.970 1191.090 8.350 ;
        RECT 1191.925 8.335 1192.255 8.350 ;
        RECT 1159.510 7.670 1191.090 7.970 ;
        RECT 1310.145 7.970 1310.475 7.985 ;
        RECT 1354.765 7.970 1355.095 7.985 ;
        RECT 1310.145 7.670 1341.050 7.970 ;
        RECT 1310.145 7.655 1310.475 7.670 ;
        RECT 1226.425 7.290 1226.755 7.305 ;
        RECT 1233.070 7.290 1233.450 7.300 ;
        RECT 1226.425 6.990 1233.450 7.290 ;
        RECT 1226.425 6.975 1226.755 6.990 ;
        RECT 1233.070 6.980 1233.450 6.990 ;
        RECT 1285.305 7.290 1285.635 7.305 ;
        RECT 1290.365 7.290 1290.695 7.305 ;
        RECT 1285.305 6.990 1290.695 7.290 ;
        RECT 1340.750 7.290 1341.050 7.670 ;
        RECT 1342.590 7.670 1355.095 7.970 ;
        RECT 1342.590 7.290 1342.890 7.670 ;
        RECT 1354.765 7.655 1355.095 7.670 ;
        RECT 1340.750 6.990 1342.890 7.290 ;
        RECT 1356.145 7.290 1356.475 7.305 ;
        RECT 1356.145 6.990 1358.530 7.290 ;
        RECT 1285.305 6.975 1285.635 6.990 ;
        RECT 1290.365 6.975 1290.695 6.990 ;
        RECT 1356.145 6.975 1356.475 6.990 ;
        RECT 1358.230 6.610 1358.530 6.990 ;
        RECT 1402.605 6.610 1402.935 6.625 ;
        RECT 1358.230 6.310 1402.935 6.610 ;
        RECT 1402.605 6.295 1402.935 6.310 ;
        RECT 457.305 4.570 457.635 4.585 ;
        RECT 458.430 4.570 458.810 4.580 ;
        RECT 457.305 4.270 458.810 4.570 ;
        RECT 457.305 4.255 457.635 4.270 ;
        RECT 458.430 4.260 458.810 4.270 ;
        RECT 1259.750 4.570 1260.130 4.580 ;
        RECT 1262.305 4.570 1262.635 4.585 ;
        RECT 1259.750 4.270 1262.635 4.570 ;
        RECT 1259.750 4.260 1260.130 4.270 ;
        RECT 1262.305 4.255 1262.635 4.270 ;
        RECT 1264.605 4.570 1264.935 4.585 ;
        RECT 1268.285 4.570 1268.615 4.585 ;
        RECT 1264.605 4.270 1268.615 4.570 ;
        RECT 1264.605 4.255 1264.935 4.270 ;
        RECT 1268.285 4.255 1268.615 4.270 ;
        RECT 735.350 3.890 735.730 3.900 ;
        RECT 807.365 3.890 807.695 3.905 ;
        RECT 735.350 3.590 782.610 3.890 ;
        RECT 735.350 3.580 735.730 3.590 ;
        RECT 782.310 3.210 782.610 3.590 ;
        RECT 785.070 3.590 807.695 3.890 ;
        RECT 785.070 3.210 785.370 3.590 ;
        RECT 807.365 3.575 807.695 3.590 ;
        RECT 808.745 3.890 809.075 3.905 ;
        RECT 815.645 3.890 815.975 3.905 ;
        RECT 808.745 3.590 815.975 3.890 ;
        RECT 808.745 3.575 809.075 3.590 ;
        RECT 815.645 3.575 815.975 3.590 ;
        RECT 819.325 3.890 819.655 3.905 ;
        RECT 880.045 3.890 880.375 3.905 ;
        RECT 819.325 3.590 880.375 3.890 ;
        RECT 819.325 3.575 819.655 3.590 ;
        RECT 880.045 3.575 880.375 3.590 ;
        RECT 1233.070 3.890 1233.450 3.900 ;
        RECT 1233.070 3.590 1238.930 3.890 ;
        RECT 1233.070 3.580 1233.450 3.590 ;
        RECT 782.310 2.910 785.370 3.210 ;
        RECT 1238.630 3.210 1238.930 3.590 ;
        RECT 1241.350 3.210 1241.730 3.220 ;
        RECT 1238.630 2.910 1241.730 3.210 ;
        RECT 1241.350 2.900 1241.730 2.910 ;
      LAYER via3 ;
        RECT 1233.100 6.980 1233.420 7.300 ;
        RECT 458.460 4.260 458.780 4.580 ;
        RECT 1259.780 4.260 1260.100 4.580 ;
        RECT 735.380 3.580 735.700 3.900 ;
        RECT 1233.100 3.580 1233.420 3.900 ;
        RECT 1241.380 2.900 1241.700 3.220 ;
      LAYER met4 ;
        RECT 1241.390 7.670 1245.370 7.970 ;
        RECT 1233.095 6.975 1233.425 7.305 ;
        RECT 458.030 4.510 459.210 5.690 ;
        RECT 731.270 4.510 732.450 5.690 ;
        RECT 458.455 4.255 458.785 4.510 ;
        RECT 731.710 3.890 732.010 4.510 ;
        RECT 1233.110 3.905 1233.410 6.975 ;
        RECT 735.375 3.890 735.705 3.905 ;
        RECT 731.710 3.590 735.705 3.890 ;
        RECT 735.375 3.575 735.705 3.590 ;
        RECT 1233.095 3.575 1233.425 3.905 ;
        RECT 1241.390 3.225 1241.690 7.670 ;
        RECT 1245.070 3.890 1245.370 7.670 ;
        RECT 1259.775 4.255 1260.105 4.585 ;
        RECT 1259.790 3.890 1260.090 4.255 ;
        RECT 1245.070 3.590 1260.090 3.890 ;
        RECT 1241.375 2.895 1241.705 3.225 ;
      LAYER via4 ;
        RECT 458.030 4.510 459.210 5.690 ;
      LAYER met5 ;
        RECT 457.820 4.300 732.660 5.900 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1157.505 11.305 1162.735 11.475 ;
        RECT 896.225 10.285 959.415 10.455 ;
        RECT 534.205 8.585 535.295 8.755 ;
        RECT 508.445 7.905 510.915 8.075 ;
        RECT 467.045 7.565 483.775 7.735 ;
        RECT 467.045 5.695 467.215 7.565 ;
        RECT 483.605 7.055 483.775 7.565 ;
        RECT 508.445 7.055 508.615 7.905 ;
        RECT 483.605 6.885 508.615 7.055 ;
        RECT 510.745 7.055 510.915 7.905 ;
        RECT 511.665 7.055 511.835 7.395 ;
        RECT 534.205 7.225 534.375 8.585 ;
        RECT 558.125 7.395 558.295 8.755 ;
        RECT 896.225 8.245 896.395 10.285 ;
        RECT 959.245 10.115 959.415 10.285 ;
        RECT 959.245 9.945 987.015 10.115 ;
        RECT 986.845 8.585 987.015 9.945 ;
        RECT 1157.505 8.585 1157.675 11.305 ;
        RECT 1162.565 10.115 1162.735 11.305 ;
        RECT 1162.565 9.945 1196.775 10.115 ;
        RECT 1196.605 8.585 1196.775 9.945 ;
        RECT 1250.425 9.605 1256.115 9.775 ;
        RECT 1200.285 8.585 1208.275 8.755 ;
        RECT 1250.425 8.585 1250.595 9.605 ;
        RECT 1255.945 9.435 1256.115 9.605 ;
        RECT 1255.945 9.265 1257.955 9.435 ;
        RECT 1257.785 8.585 1257.955 9.265 ;
        RECT 1262.845 8.925 1263.935 9.095 ;
        RECT 1262.845 8.585 1263.015 8.925 ;
        RECT 559.965 7.565 561.515 7.735 ;
        RECT 559.965 7.395 560.135 7.565 ;
        RECT 558.125 7.225 560.135 7.395 ;
        RECT 510.745 6.885 511.835 7.055 ;
        RECT 466.585 5.525 467.215 5.695 ;
        RECT 466.585 2.975 466.755 5.525 ;
        RECT 561.345 4.335 561.515 7.565 ;
        RECT 561.345 4.165 562.895 4.335 ;
        RECT 573.765 3.995 573.935 4.335 ;
        RECT 575.145 3.995 575.315 6.375 ;
        RECT 583.425 6.035 583.595 6.375 ;
        RECT 583.425 5.865 584.515 6.035 ;
        RECT 596.305 5.695 596.475 6.035 ;
        RECT 597.685 5.695 597.855 6.035 ;
        RECT 596.305 5.525 597.855 5.695 ;
        RECT 696.585 5.695 696.755 6.035 ;
        RECT 697.505 5.865 698.135 6.035 ;
        RECT 747.645 5.865 749.655 6.035 ;
        RECT 697.505 5.695 697.675 5.865 ;
        RECT 696.585 5.525 697.675 5.695 ;
        RECT 573.765 3.825 575.315 3.995 ;
        RECT 1263.765 3.315 1263.935 8.925 ;
        RECT 1403.145 4.335 1403.315 8.075 ;
        RECT 1401.305 4.165 1403.315 4.335 ;
        RECT 1401.305 3.655 1401.475 4.165 ;
        RECT 1399.925 3.485 1401.475 3.655 ;
        RECT 1263.765 3.145 1297.055 3.315 ;
        RECT 1399.925 3.145 1400.095 3.485 ;
        RECT 466.585 2.805 467.215 2.975 ;
      LAYER mcon ;
        RECT 535.125 8.585 535.295 8.755 ;
        RECT 558.125 8.585 558.295 8.755 ;
        RECT 511.665 7.225 511.835 7.395 ;
        RECT 1208.105 8.585 1208.275 8.755 ;
        RECT 575.145 6.205 575.315 6.375 ;
        RECT 562.725 4.165 562.895 4.335 ;
        RECT 573.765 4.165 573.935 4.335 ;
        RECT 583.425 6.205 583.595 6.375 ;
        RECT 584.345 5.865 584.515 6.035 ;
        RECT 596.305 5.865 596.475 6.035 ;
        RECT 597.685 5.865 597.855 6.035 ;
        RECT 696.585 5.865 696.755 6.035 ;
        RECT 697.965 5.865 698.135 6.035 ;
        RECT 749.485 5.865 749.655 6.035 ;
        RECT 1403.145 7.905 1403.315 8.075 ;
        RECT 1296.885 3.145 1297.055 3.315 ;
        RECT 467.045 2.805 467.215 2.975 ;
      LAYER met1 ;
        RECT 535.065 8.740 535.355 8.785 ;
        RECT 558.065 8.740 558.355 8.785 ;
        RECT 535.065 8.600 558.355 8.740 ;
        RECT 535.065 8.555 535.355 8.600 ;
        RECT 558.065 8.555 558.355 8.600 ;
        RECT 986.785 8.740 987.075 8.785 ;
        RECT 1157.445 8.740 1157.735 8.785 ;
        RECT 986.785 8.600 1157.735 8.740 ;
        RECT 986.785 8.555 987.075 8.600 ;
        RECT 1157.445 8.555 1157.735 8.600 ;
        RECT 1196.545 8.740 1196.835 8.785 ;
        RECT 1200.225 8.740 1200.515 8.785 ;
        RECT 1196.545 8.600 1200.515 8.740 ;
        RECT 1196.545 8.555 1196.835 8.600 ;
        RECT 1200.225 8.555 1200.515 8.600 ;
        RECT 1208.045 8.740 1208.335 8.785 ;
        RECT 1250.365 8.740 1250.655 8.785 ;
        RECT 1208.045 8.600 1250.655 8.740 ;
        RECT 1208.045 8.555 1208.335 8.600 ;
        RECT 1250.365 8.555 1250.655 8.600 ;
        RECT 1257.725 8.740 1258.015 8.785 ;
        RECT 1262.785 8.740 1263.075 8.785 ;
        RECT 1257.725 8.600 1263.075 8.740 ;
        RECT 1257.725 8.555 1258.015 8.600 ;
        RECT 1262.785 8.555 1263.075 8.600 ;
        RECT 895.690 8.400 896.010 8.460 ;
        RECT 896.165 8.400 896.455 8.445 ;
        RECT 895.690 8.260 896.455 8.400 ;
        RECT 895.690 8.200 896.010 8.260 ;
        RECT 896.165 8.215 896.455 8.260 ;
        RECT 1403.085 8.060 1403.375 8.105 ;
        RECT 1451.830 8.060 1452.150 8.120 ;
        RECT 1403.085 7.920 1452.150 8.060 ;
        RECT 1403.085 7.875 1403.375 7.920 ;
        RECT 1451.830 7.860 1452.150 7.920 ;
        RECT 511.605 7.380 511.895 7.425 ;
        RECT 534.145 7.380 534.435 7.425 ;
        RECT 511.605 7.240 534.435 7.380 ;
        RECT 511.605 7.195 511.895 7.240 ;
        RECT 534.145 7.195 534.435 7.240 ;
        RECT 575.085 6.360 575.375 6.405 ;
        RECT 582.430 6.360 582.750 6.420 ;
        RECT 583.350 6.360 583.670 6.420 ;
        RECT 575.085 6.220 582.750 6.360 ;
        RECT 583.155 6.220 583.670 6.360 ;
        RECT 575.085 6.175 575.375 6.220 ;
        RECT 582.430 6.160 582.750 6.220 ;
        RECT 583.350 6.160 583.670 6.220 ;
        RECT 584.285 6.020 584.575 6.065 ;
        RECT 596.245 6.020 596.535 6.065 ;
        RECT 584.285 5.880 596.535 6.020 ;
        RECT 584.285 5.835 584.575 5.880 ;
        RECT 596.245 5.835 596.535 5.880 ;
        RECT 597.625 6.020 597.915 6.065 ;
        RECT 696.525 6.020 696.815 6.065 ;
        RECT 597.625 5.880 696.815 6.020 ;
        RECT 597.625 5.835 597.915 5.880 ;
        RECT 696.525 5.835 696.815 5.880 ;
        RECT 697.905 6.020 698.195 6.065 ;
        RECT 724.110 6.020 724.430 6.080 ;
        RECT 697.905 5.880 724.430 6.020 ;
        RECT 697.905 5.835 698.195 5.880 ;
        RECT 724.110 5.820 724.430 5.880 ;
        RECT 724.570 6.020 724.890 6.080 ;
        RECT 747.585 6.020 747.875 6.065 ;
        RECT 724.570 5.880 747.875 6.020 ;
        RECT 724.570 5.820 724.890 5.880 ;
        RECT 747.585 5.835 747.875 5.880 ;
        RECT 749.425 6.020 749.715 6.065 ;
        RECT 762.290 6.020 762.610 6.080 ;
        RECT 749.425 5.880 762.610 6.020 ;
        RECT 749.425 5.835 749.715 5.880 ;
        RECT 762.290 5.820 762.610 5.880 ;
        RECT 769.190 6.020 769.510 6.080 ;
        RECT 805.530 6.020 805.850 6.080 ;
        RECT 769.190 5.880 803.460 6.020 ;
        RECT 769.190 5.820 769.510 5.880 ;
        RECT 803.320 5.680 803.460 5.880 ;
        RECT 804.700 5.880 805.850 6.020 ;
        RECT 804.700 5.680 804.840 5.880 ;
        RECT 805.530 5.820 805.850 5.880 ;
        RECT 806.450 6.020 806.770 6.080 ;
        RECT 894.770 6.020 895.090 6.080 ;
        RECT 806.450 5.880 895.090 6.020 ;
        RECT 806.450 5.820 806.770 5.880 ;
        RECT 894.770 5.820 895.090 5.880 ;
        RECT 803.320 5.540 804.840 5.680 ;
        RECT 562.665 4.320 562.955 4.365 ;
        RECT 573.705 4.320 573.995 4.365 ;
        RECT 562.665 4.180 573.995 4.320 ;
        RECT 562.665 4.135 562.955 4.180 ;
        RECT 573.705 4.135 573.995 4.180 ;
        RECT 1307.480 3.500 1355.460 3.640 ;
        RECT 1296.825 3.300 1297.115 3.345 ;
        RECT 1307.480 3.300 1307.620 3.500 ;
        RECT 1296.825 3.160 1307.620 3.300 ;
        RECT 1355.320 3.300 1355.460 3.500 ;
        RECT 1399.865 3.300 1400.155 3.345 ;
        RECT 1355.320 3.160 1400.155 3.300 ;
        RECT 1296.825 3.115 1297.115 3.160 ;
        RECT 1399.865 3.115 1400.155 3.160 ;
        RECT 466.970 2.960 467.290 3.020 ;
        RECT 466.970 2.820 467.485 2.960 ;
        RECT 466.970 2.760 467.290 2.820 ;
      LAYER via ;
        RECT 895.720 8.200 895.980 8.460 ;
        RECT 1451.860 7.860 1452.120 8.120 ;
        RECT 582.460 6.160 582.720 6.420 ;
        RECT 583.380 6.160 583.640 6.420 ;
        RECT 724.140 5.820 724.400 6.080 ;
        RECT 724.600 5.820 724.860 6.080 ;
        RECT 762.320 5.820 762.580 6.080 ;
        RECT 769.220 5.820 769.480 6.080 ;
        RECT 805.560 5.820 805.820 6.080 ;
        RECT 806.480 5.820 806.740 6.080 ;
        RECT 894.800 5.820 895.060 6.080 ;
        RECT 467.000 2.760 467.260 3.020 ;
      LAYER met2 ;
        RECT 895.720 8.170 895.980 8.490 ;
        RECT 895.780 6.530 895.920 8.170 ;
        RECT 1451.860 7.890 1452.120 8.150 ;
        RECT 1453.630 7.890 1453.910 9.000 ;
        RECT 1451.860 7.830 1453.910 7.890 ;
        RECT 1451.920 7.750 1453.910 7.830 ;
        RECT 582.520 6.450 583.580 6.530 ;
        RECT 582.460 6.390 583.640 6.450 ;
        RECT 582.460 6.130 582.720 6.390 ;
        RECT 583.380 6.130 583.640 6.390 ;
        RECT 763.760 6.390 768.960 6.530 ;
        RECT 724.140 5.790 724.400 6.110 ;
        RECT 724.600 5.790 724.860 6.110 ;
        RECT 762.320 5.850 762.580 6.110 ;
        RECT 763.760 5.850 763.900 6.390 ;
        RECT 768.820 6.020 768.960 6.390 ;
        RECT 894.860 6.390 895.920 6.530 ;
        RECT 894.860 6.110 895.000 6.390 ;
        RECT 769.220 6.020 769.480 6.110 ;
        RECT 768.820 5.880 769.480 6.020 ;
        RECT 762.320 5.790 763.900 5.850 ;
        RECT 769.220 5.790 769.480 5.880 ;
        RECT 805.560 5.850 805.820 6.110 ;
        RECT 806.480 5.850 806.740 6.110 ;
        RECT 805.560 5.790 806.740 5.850 ;
        RECT 894.800 5.790 895.060 6.110 ;
        RECT 724.200 5.340 724.340 5.790 ;
        RECT 724.660 5.340 724.800 5.790 ;
        RECT 762.380 5.710 763.900 5.790 ;
        RECT 805.620 5.710 806.680 5.790 ;
        RECT 724.200 5.200 724.800 5.340 ;
        RECT 1453.630 5.000 1453.910 7.750 ;
        RECT 467.000 2.960 467.260 3.050 ;
        RECT 466.600 2.820 467.260 2.960 ;
        RECT 466.600 2.400 466.740 2.820 ;
        RECT 467.000 2.730 467.260 2.820 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 739.825 10.285 771.735 10.455 ;
        RECT 531.445 9.945 564.275 10.115 ;
        RECT 531.445 5.865 531.615 9.945 ;
        RECT 564.105 7.735 564.275 9.945 ;
        RECT 579.745 9.265 581.295 9.435 ;
        RECT 564.105 7.565 576.235 7.735 ;
        RECT 576.065 5.355 576.235 7.565 ;
        RECT 579.745 5.355 579.915 9.265 ;
        RECT 581.125 8.925 581.295 9.265 ;
        RECT 628.045 8.245 628.215 9.095 ;
        RECT 672.205 8.925 673.295 9.095 ;
        RECT 734.305 8.925 735.855 9.095 ;
        RECT 739.825 8.925 739.995 10.285 ;
        RECT 672.205 8.585 672.375 8.925 ;
        RECT 771.565 8.755 771.735 10.285 ;
        RECT 781.225 9.605 807.155 9.775 ;
        RECT 771.565 8.585 776.795 8.755 ;
        RECT 576.065 5.185 579.915 5.355 ;
        RECT 776.625 3.995 776.795 8.585 ;
        RECT 781.225 3.995 781.395 9.605 ;
        RECT 806.985 5.355 807.155 9.605 ;
        RECT 1103.685 7.905 1104.315 8.075 ;
        RECT 994.205 7.565 996.215 7.735 ;
        RECT 810.205 7.225 815.435 7.395 ;
        RECT 810.205 5.355 810.375 7.225 ;
        RECT 815.265 7.055 815.435 7.225 ;
        RECT 820.785 7.055 820.955 7.395 ;
        RECT 815.265 6.885 820.955 7.055 ;
        RECT 822.625 7.055 822.795 7.395 ;
        RECT 823.545 7.225 824.635 7.395 ;
        RECT 823.545 7.055 823.715 7.225 ;
        RECT 822.625 6.885 823.715 7.055 ;
        RECT 824.465 6.885 824.635 7.225 ;
        RECT 833.665 6.885 836.135 7.055 ;
        RECT 806.985 5.185 810.375 5.355 ;
        RECT 776.625 3.825 781.395 3.995 ;
        RECT 835.965 3.145 836.135 6.885 ;
        RECT 885.185 3.825 890.415 3.995 ;
        RECT 844.705 3.485 845.795 3.655 ;
        RECT 844.705 3.145 844.875 3.485 ;
        RECT 885.185 3.145 885.355 3.825 ;
        RECT 890.245 3.145 890.415 3.825 ;
        RECT 994.205 3.655 994.375 7.565 ;
        RECT 1014.445 7.395 1014.615 7.735 ;
        RECT 1055.845 7.395 1056.015 7.735 ;
        RECT 1104.145 7.565 1104.315 7.905 ;
        RECT 1122.085 7.735 1122.255 8.075 ;
        RECT 1121.625 7.565 1122.255 7.735 ;
        RECT 1492.385 7.565 1492.555 8.415 ;
        RECT 1014.445 7.225 1056.015 7.395 ;
        RECT 985.005 3.485 994.375 3.655 ;
        RECT 917.385 3.145 918.015 3.315 ;
        RECT 985.005 3.145 985.175 3.485 ;
        RECT 917.845 2.975 918.015 3.145 ;
        RECT 917.845 2.805 919.395 2.975 ;
      LAYER mcon ;
        RECT 628.045 8.925 628.215 9.095 ;
        RECT 673.125 8.925 673.295 9.095 ;
        RECT 735.685 8.925 735.855 9.095 ;
        RECT 1492.385 8.245 1492.555 8.415 ;
        RECT 1122.085 7.905 1122.255 8.075 ;
        RECT 996.045 7.565 996.215 7.735 ;
        RECT 1014.445 7.565 1014.615 7.735 ;
        RECT 820.785 7.225 820.955 7.395 ;
        RECT 822.625 7.225 822.795 7.395 ;
        RECT 845.625 3.485 845.795 3.655 ;
        RECT 1055.845 7.565 1056.015 7.735 ;
        RECT 919.225 2.805 919.395 2.975 ;
      LAYER met1 ;
        RECT 581.065 9.080 581.355 9.125 ;
        RECT 627.985 9.080 628.275 9.125 ;
        RECT 673.065 9.080 673.355 9.125 ;
        RECT 734.245 9.080 734.535 9.125 ;
        RECT 581.065 8.940 628.275 9.080 ;
        RECT 581.065 8.895 581.355 8.940 ;
        RECT 627.985 8.895 628.275 8.940 ;
        RECT 642.780 8.940 652.120 9.080 ;
        RECT 627.985 8.400 628.275 8.445 ;
        RECT 642.780 8.400 642.920 8.940 ;
        RECT 651.980 8.740 652.120 8.940 ;
        RECT 673.065 8.940 734.535 9.080 ;
        RECT 673.065 8.895 673.355 8.940 ;
        RECT 734.245 8.895 734.535 8.940 ;
        RECT 735.625 8.895 735.915 9.125 ;
        RECT 739.765 8.895 740.055 9.125 ;
        RECT 672.145 8.740 672.435 8.785 ;
        RECT 651.980 8.600 672.435 8.740 ;
        RECT 735.700 8.740 735.840 8.895 ;
        RECT 739.840 8.740 739.980 8.895 ;
        RECT 735.700 8.600 739.980 8.740 ;
        RECT 672.145 8.555 672.435 8.600 ;
        RECT 627.985 8.260 642.920 8.400 ;
        RECT 1492.325 8.400 1492.615 8.445 ;
        RECT 1499.670 8.400 1499.990 8.460 ;
        RECT 1492.325 8.260 1499.990 8.400 ;
        RECT 627.985 8.215 628.275 8.260 ;
        RECT 1492.325 8.215 1492.615 8.260 ;
        RECT 1499.670 8.200 1499.990 8.260 ;
        RECT 1103.625 7.875 1103.915 8.105 ;
        RECT 1122.025 8.060 1122.315 8.105 ;
        RECT 1122.025 7.920 1123.620 8.060 ;
        RECT 1122.025 7.875 1122.315 7.920 ;
        RECT 995.985 7.720 996.275 7.765 ;
        RECT 1014.385 7.720 1014.675 7.765 ;
        RECT 995.985 7.580 1014.675 7.720 ;
        RECT 995.985 7.535 996.275 7.580 ;
        RECT 1014.385 7.535 1014.675 7.580 ;
        RECT 1055.785 7.720 1056.075 7.765 ;
        RECT 1103.700 7.720 1103.840 7.875 ;
        RECT 1055.785 7.580 1103.840 7.720 ;
        RECT 1104.085 7.720 1104.375 7.765 ;
        RECT 1121.565 7.720 1121.855 7.765 ;
        RECT 1104.085 7.580 1121.855 7.720 ;
        RECT 1123.480 7.720 1123.620 7.920 ;
        RECT 1301.960 7.920 1303.940 8.060 ;
        RECT 1301.960 7.720 1302.100 7.920 ;
        RECT 1123.480 7.580 1160.420 7.720 ;
        RECT 1055.785 7.535 1056.075 7.580 ;
        RECT 1104.085 7.535 1104.375 7.580 ;
        RECT 1121.565 7.535 1121.855 7.580 ;
        RECT 820.725 7.380 821.015 7.425 ;
        RECT 822.565 7.380 822.855 7.425 ;
        RECT 820.725 7.240 822.855 7.380 ;
        RECT 1160.280 7.380 1160.420 7.580 ;
        RECT 1162.580 7.580 1302.100 7.720 ;
        RECT 1303.800 7.720 1303.940 7.920 ;
        RECT 1428.830 7.720 1429.150 7.780 ;
        RECT 1303.800 7.580 1429.150 7.720 ;
        RECT 1162.580 7.380 1162.720 7.580 ;
        RECT 1428.830 7.520 1429.150 7.580 ;
        RECT 1448.610 7.720 1448.930 7.780 ;
        RECT 1492.325 7.720 1492.615 7.765 ;
        RECT 1448.610 7.580 1492.615 7.720 ;
        RECT 1448.610 7.520 1448.930 7.580 ;
        RECT 1492.325 7.535 1492.615 7.580 ;
        RECT 1160.280 7.240 1162.720 7.380 ;
        RECT 820.725 7.195 821.015 7.240 ;
        RECT 822.565 7.195 822.855 7.240 ;
        RECT 824.405 7.040 824.695 7.085 ;
        RECT 833.605 7.040 833.895 7.085 ;
        RECT 824.405 6.900 833.895 7.040 ;
        RECT 824.405 6.855 824.695 6.900 ;
        RECT 833.605 6.855 833.895 6.900 ;
        RECT 523.090 6.020 523.410 6.080 ;
        RECT 531.385 6.020 531.675 6.065 ;
        RECT 523.090 5.880 531.675 6.020 ;
        RECT 523.090 5.820 523.410 5.880 ;
        RECT 531.385 5.835 531.675 5.880 ;
        RECT 878.210 3.980 878.530 4.040 ;
        RECT 847.940 3.840 878.530 3.980 ;
        RECT 845.565 3.640 845.855 3.685 ;
        RECT 847.940 3.640 848.080 3.840 ;
        RECT 878.210 3.780 878.530 3.840 ;
        RECT 845.565 3.500 848.080 3.640 ;
        RECT 845.565 3.455 845.855 3.500 ;
        RECT 835.905 3.300 836.195 3.345 ;
        RECT 844.645 3.300 844.935 3.345 ;
        RECT 835.905 3.160 844.935 3.300 ;
        RECT 835.905 3.115 836.195 3.160 ;
        RECT 844.645 3.115 844.935 3.160 ;
        RECT 883.270 3.300 883.590 3.360 ;
        RECT 885.125 3.300 885.415 3.345 ;
        RECT 883.270 3.160 885.415 3.300 ;
        RECT 883.270 3.100 883.590 3.160 ;
        RECT 885.125 3.115 885.415 3.160 ;
        RECT 890.185 3.300 890.475 3.345 ;
        RECT 917.325 3.300 917.615 3.345 ;
        RECT 984.945 3.300 985.235 3.345 ;
        RECT 890.185 3.160 917.615 3.300 ;
        RECT 890.185 3.115 890.475 3.160 ;
        RECT 917.325 3.115 917.615 3.160 ;
        RECT 919.240 3.160 985.235 3.300 ;
        RECT 919.240 3.005 919.380 3.160 ;
        RECT 984.945 3.115 985.235 3.160 ;
        RECT 919.165 2.775 919.455 3.005 ;
      LAYER via ;
        RECT 1499.700 8.200 1499.960 8.460 ;
        RECT 1428.860 7.520 1429.120 7.780 ;
        RECT 1448.640 7.520 1448.900 7.780 ;
        RECT 523.120 5.820 523.380 6.080 ;
        RECT 878.240 3.780 878.500 4.040 ;
        RECT 883.300 3.100 883.560 3.360 ;
      LAYER met2 ;
        RECT 1499.760 8.490 1500.820 8.570 ;
        RECT 1499.700 8.430 1500.820 8.490 ;
        RECT 1499.700 8.170 1499.960 8.430 ;
        RECT 1500.680 8.400 1500.820 8.430 ;
        RECT 1501.010 8.400 1501.290 9.000 ;
        RECT 1500.680 8.260 1501.290 8.400 ;
        RECT 1428.920 7.810 1448.840 7.890 ;
        RECT 1428.860 7.750 1448.900 7.810 ;
        RECT 1428.860 7.490 1429.120 7.750 ;
        RECT 1448.640 7.490 1448.900 7.750 ;
        RECT 523.120 5.965 523.380 6.110 ;
        RECT 507.010 5.680 507.290 5.965 ;
        RECT 504.320 5.595 507.290 5.680 ;
        RECT 523.110 5.595 523.390 5.965 ;
        RECT 504.320 5.540 507.220 5.595 ;
        RECT 504.320 5.340 504.460 5.540 ;
        RECT 503.860 5.200 504.460 5.340 ;
        RECT 503.860 4.660 504.000 5.200 ;
        RECT 1501.010 5.000 1501.290 8.260 ;
        RECT 489.600 4.520 504.000 4.660 ;
        RECT 484.540 2.820 485.600 2.960 ;
        RECT 484.540 2.400 484.680 2.820 ;
        RECT 484.330 -4.800 484.890 2.400 ;
        RECT 485.460 0.410 485.600 2.820 ;
        RECT 489.600 0.410 489.740 4.520 ;
        RECT 878.240 3.750 878.500 4.070 ;
        RECT 878.300 1.090 878.440 3.750 ;
        RECT 883.300 3.300 883.560 3.390 ;
        RECT 881.980 3.160 883.560 3.300 ;
        RECT 881.980 1.090 882.120 3.160 ;
        RECT 883.300 3.070 883.560 3.160 ;
        RECT 878.300 0.950 882.120 1.090 ;
        RECT 485.460 0.270 489.740 0.410 ;
      LAYER via2 ;
        RECT 507.010 5.640 507.290 5.920 ;
        RECT 523.110 5.640 523.390 5.920 ;
      LAYER met3 ;
        RECT 506.985 5.930 507.315 5.945 ;
        RECT 523.085 5.930 523.415 5.945 ;
        RECT 506.985 5.630 523.415 5.930 ;
        RECT 506.985 5.615 507.315 5.630 ;
        RECT 523.085 5.615 523.415 5.630 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 809.745 9.605 810.835 9.775 ;
        RECT 550.765 8.925 558.755 9.095 ;
        RECT 513.965 6.545 517.355 6.715 ;
        RECT 513.965 4.675 514.135 6.545 ;
        RECT 511.665 4.505 514.135 4.675 ;
        RECT 511.665 3.485 511.835 4.505 ;
        RECT 517.185 3.995 517.355 6.545 ;
        RECT 537.885 4.165 545.875 4.335 ;
        RECT 537.885 3.995 538.055 4.165 ;
        RECT 517.185 3.825 538.055 3.995 ;
        RECT 545.705 3.995 545.875 4.165 ;
        RECT 550.765 3.995 550.935 8.925 ;
        RECT 558.585 7.735 558.755 8.925 ;
        RECT 581.585 8.925 611.655 9.095 ;
        RECT 559.505 7.905 561.975 8.075 ;
        RECT 575.605 7.905 576.695 8.075 ;
        RECT 559.505 7.735 559.675 7.905 ;
        RECT 558.585 7.565 559.675 7.735 ;
        RECT 576.525 6.885 576.695 7.905 ;
        RECT 581.585 7.395 581.755 8.925 ;
        RECT 581.125 7.225 581.755 7.395 ;
        RECT 581.125 6.885 581.295 7.225 ;
        RECT 611.485 6.885 611.655 8.925 ;
        RECT 664.385 7.565 671.455 7.735 ;
        RECT 658.865 7.225 663.635 7.395 ;
        RECT 658.865 6.885 659.035 7.225 ;
        RECT 663.465 6.715 663.635 7.225 ;
        RECT 664.385 6.715 664.555 7.565 ;
        RECT 671.285 7.395 671.455 7.565 ;
        RECT 674.045 7.565 675.135 7.735 ;
        RECT 671.285 7.225 672.835 7.395 ;
        RECT 663.465 6.545 664.555 6.715 ;
        RECT 672.665 6.715 672.835 7.225 ;
        RECT 674.045 6.715 674.215 7.565 ;
        RECT 674.965 7.395 675.135 7.565 ;
        RECT 674.965 7.225 705.495 7.395 ;
        RECT 672.665 6.545 674.215 6.715 ;
        RECT 705.325 4.335 705.495 7.225 ;
        RECT 715.445 7.225 718.835 7.395 ;
        RECT 706.245 4.335 706.415 7.055 ;
        RECT 715.445 6.885 715.615 7.225 ;
        RECT 718.665 5.355 718.835 7.225 ;
        RECT 718.665 5.185 731.715 5.355 ;
        RECT 731.545 4.505 731.715 5.185 ;
        RECT 705.325 4.165 706.415 4.335 ;
        RECT 736.605 4.335 736.775 4.675 ;
        RECT 750.865 4.335 751.035 4.675 ;
        RECT 736.605 4.165 751.035 4.335 ;
        RECT 545.705 3.825 550.935 3.995 ;
        RECT 783.065 3.485 783.235 7.055 ;
        RECT 809.745 6.885 809.915 9.605 ;
        RECT 810.665 9.435 810.835 9.605 ;
        RECT 810.665 9.265 851.315 9.435 ;
        RECT 851.145 8.585 851.315 9.265 ;
        RECT 1292.745 7.565 1304.875 7.735 ;
        RECT 1292.745 7.395 1292.915 7.565 ;
        RECT 883.805 7.225 888.575 7.395 ;
        RECT 882.425 6.715 882.595 7.055 ;
        RECT 883.805 6.715 883.975 7.225 ;
        RECT 882.425 6.545 883.975 6.715 ;
        RECT 888.405 6.205 888.575 7.225 ;
        RECT 1291.825 7.225 1292.915 7.395 ;
        RECT 900.365 5.865 900.535 7.055 ;
        RECT 949.125 6.375 949.295 7.055 ;
        RECT 952.805 6.715 952.975 7.055 ;
        RECT 1122.545 6.885 1125.475 7.055 ;
        RECT 1291.825 6.885 1291.995 7.225 ;
        RECT 1304.705 7.055 1304.875 7.565 ;
        RECT 1304.705 6.885 1305.335 7.055 ;
        RECT 951.425 6.545 952.975 6.715 ;
        RECT 949.125 6.205 950.675 6.375 ;
        RECT 950.505 6.035 950.675 6.205 ;
        RECT 951.425 6.035 951.595 6.545 ;
        RECT 950.505 5.865 951.595 6.035 ;
        RECT 1425.685 0.935 1425.855 7.055 ;
        RECT 1436.725 1.955 1436.895 7.055 ;
        RECT 1436.725 1.785 1446.555 1.955 ;
        RECT 1446.385 1.275 1446.555 1.785 ;
        RECT 1430.285 1.105 1446.555 1.275 ;
        RECT 1430.285 0.935 1430.455 1.105 ;
        RECT 1425.685 0.765 1430.455 0.935 ;
      LAYER mcon ;
        RECT 561.805 7.905 561.975 8.075 ;
        RECT 706.245 6.885 706.415 7.055 ;
        RECT 783.065 6.885 783.235 7.055 ;
        RECT 882.425 6.885 882.595 7.055 ;
        RECT 736.605 4.505 736.775 4.675 ;
        RECT 750.865 4.505 751.035 4.675 ;
        RECT 900.365 6.885 900.535 7.055 ;
        RECT 949.125 6.885 949.295 7.055 ;
        RECT 952.805 6.885 952.975 7.055 ;
        RECT 1125.305 6.885 1125.475 7.055 ;
        RECT 1305.165 6.885 1305.335 7.055 ;
        RECT 1425.685 6.885 1425.855 7.055 ;
        RECT 1436.725 6.885 1436.895 7.055 ;
      LAYER met1 ;
        RECT 851.085 8.740 851.375 8.785 ;
        RECT 854.750 8.740 855.070 8.800 ;
        RECT 851.085 8.600 855.070 8.740 ;
        RECT 851.085 8.555 851.375 8.600 ;
        RECT 854.750 8.540 855.070 8.600 ;
        RECT 561.745 8.060 562.035 8.105 ;
        RECT 575.545 8.060 575.835 8.105 ;
        RECT 561.745 7.920 575.835 8.060 ;
        RECT 561.745 7.875 562.035 7.920 ;
        RECT 575.545 7.875 575.835 7.920 ;
        RECT 576.465 7.040 576.755 7.085 ;
        RECT 581.065 7.040 581.355 7.085 ;
        RECT 576.465 6.900 581.355 7.040 ;
        RECT 576.465 6.855 576.755 6.900 ;
        RECT 581.065 6.855 581.355 6.900 ;
        RECT 611.425 7.040 611.715 7.085 ;
        RECT 658.805 7.040 659.095 7.085 ;
        RECT 611.425 6.900 659.095 7.040 ;
        RECT 611.425 6.855 611.715 6.900 ;
        RECT 658.805 6.855 659.095 6.900 ;
        RECT 706.185 7.040 706.475 7.085 ;
        RECT 715.385 7.040 715.675 7.085 ;
        RECT 706.185 6.900 715.675 7.040 ;
        RECT 706.185 6.855 706.475 6.900 ;
        RECT 715.385 6.855 715.675 6.900 ;
        RECT 783.005 7.040 783.295 7.085 ;
        RECT 809.685 7.040 809.975 7.085 ;
        RECT 783.005 6.900 809.975 7.040 ;
        RECT 783.005 6.855 783.295 6.900 ;
        RECT 809.685 6.855 809.975 6.900 ;
        RECT 868.090 7.040 868.410 7.100 ;
        RECT 882.365 7.040 882.655 7.085 ;
        RECT 868.090 6.900 882.655 7.040 ;
        RECT 868.090 6.840 868.410 6.900 ;
        RECT 882.365 6.855 882.655 6.900 ;
        RECT 900.305 7.040 900.595 7.085 ;
        RECT 949.065 7.040 949.355 7.085 ;
        RECT 900.305 6.900 949.355 7.040 ;
        RECT 900.305 6.855 900.595 6.900 ;
        RECT 949.065 6.855 949.355 6.900 ;
        RECT 952.745 7.040 953.035 7.085 ;
        RECT 1088.430 7.040 1088.750 7.100 ;
        RECT 952.745 6.900 1088.750 7.040 ;
        RECT 952.745 6.855 953.035 6.900 ;
        RECT 1088.430 6.840 1088.750 6.900 ;
        RECT 1093.950 7.040 1094.270 7.100 ;
        RECT 1122.485 7.040 1122.775 7.085 ;
        RECT 1093.950 6.900 1122.775 7.040 ;
        RECT 1093.950 6.840 1094.270 6.900 ;
        RECT 1122.485 6.855 1122.775 6.900 ;
        RECT 1125.245 7.040 1125.535 7.085 ;
        RECT 1291.765 7.040 1292.055 7.085 ;
        RECT 1125.245 6.900 1292.055 7.040 ;
        RECT 1125.245 6.855 1125.535 6.900 ;
        RECT 1291.765 6.855 1292.055 6.900 ;
        RECT 1305.105 7.040 1305.395 7.085 ;
        RECT 1425.625 7.040 1425.915 7.085 ;
        RECT 1305.105 6.900 1425.915 7.040 ;
        RECT 1305.105 6.855 1305.395 6.900 ;
        RECT 1425.625 6.855 1425.915 6.900 ;
        RECT 1436.665 7.040 1436.955 7.085 ;
        RECT 1546.590 7.040 1546.910 7.100 ;
        RECT 1436.665 6.900 1546.910 7.040 ;
        RECT 1436.665 6.855 1436.955 6.900 ;
        RECT 1546.590 6.840 1546.910 6.900 ;
        RECT 888.330 6.360 888.650 6.420 ;
        RECT 888.330 6.220 888.845 6.360 ;
        RECT 888.330 6.160 888.650 6.220 ;
        RECT 896.150 6.020 896.470 6.080 ;
        RECT 900.305 6.020 900.595 6.065 ;
        RECT 896.150 5.880 900.595 6.020 ;
        RECT 896.150 5.820 896.470 5.880 ;
        RECT 900.305 5.835 900.595 5.880 ;
        RECT 731.485 4.660 731.775 4.705 ;
        RECT 736.545 4.660 736.835 4.705 ;
        RECT 731.485 4.520 736.835 4.660 ;
        RECT 731.485 4.475 731.775 4.520 ;
        RECT 736.545 4.475 736.835 4.520 ;
        RECT 750.805 4.660 751.095 4.705 ;
        RECT 761.830 4.660 762.150 4.720 ;
        RECT 750.805 4.520 762.150 4.660 ;
        RECT 750.805 4.475 751.095 4.520 ;
        RECT 761.830 4.460 762.150 4.520 ;
        RECT 503.770 3.640 504.090 3.700 ;
        RECT 511.605 3.640 511.895 3.685 ;
        RECT 782.990 3.640 783.310 3.700 ;
        RECT 503.770 3.500 511.895 3.640 ;
        RECT 782.795 3.500 783.310 3.640 ;
        RECT 503.770 3.440 504.090 3.500 ;
        RECT 511.605 3.455 511.895 3.500 ;
        RECT 782.990 3.440 783.310 3.500 ;
      LAYER via ;
        RECT 854.780 8.540 855.040 8.800 ;
        RECT 868.120 6.840 868.380 7.100 ;
        RECT 1088.460 6.840 1088.720 7.100 ;
        RECT 1093.980 6.840 1094.240 7.100 ;
        RECT 1546.620 6.840 1546.880 7.100 ;
        RECT 888.360 6.160 888.620 6.420 ;
        RECT 896.180 5.820 896.440 6.080 ;
        RECT 761.860 4.460 762.120 4.720 ;
        RECT 503.800 3.440 504.060 3.700 ;
        RECT 783.020 3.440 783.280 3.700 ;
      LAYER met2 ;
        RECT 854.780 8.510 855.040 8.830 ;
        RECT 854.840 6.530 854.980 8.510 ;
        RECT 1088.520 7.920 1092.800 8.060 ;
        RECT 1088.520 7.130 1088.660 7.920 ;
        RECT 868.120 6.810 868.380 7.130 ;
        RECT 1088.460 6.810 1088.720 7.130 ;
        RECT 1092.660 7.040 1092.800 7.920 ;
        RECT 1548.390 7.210 1548.670 9.000 ;
        RECT 1546.680 7.130 1548.670 7.210 ;
        RECT 1093.980 7.040 1094.240 7.130 ;
        RECT 1092.660 6.900 1094.240 7.040 ;
        RECT 1093.980 6.810 1094.240 6.900 ;
        RECT 1546.620 7.070 1548.670 7.130 ;
        RECT 1546.620 6.810 1546.880 7.070 ;
        RECT 868.180 6.530 868.320 6.810 ;
        RECT 854.840 6.390 868.320 6.530 ;
        RECT 888.360 6.130 888.620 6.450 ;
        RECT 764.220 5.880 768.500 6.020 ;
        RECT 888.420 5.965 888.560 6.130 ;
        RECT 896.180 6.020 896.440 6.110 ;
        RECT 895.780 5.965 896.440 6.020 ;
        RECT 761.860 4.660 762.120 4.750 ;
        RECT 764.220 4.660 764.360 5.880 ;
        RECT 761.860 4.520 764.360 4.660 ;
        RECT 761.860 4.430 762.120 4.520 ;
        RECT 768.360 3.980 768.500 5.880 ;
        RECT 888.350 5.595 888.630 5.965 ;
        RECT 895.710 5.880 896.440 5.965 ;
        RECT 895.710 5.595 895.990 5.880 ;
        RECT 896.180 5.790 896.440 5.880 ;
        RECT 771.580 5.030 776.320 5.170 ;
        RECT 771.580 3.980 771.720 5.030 ;
        RECT 768.360 3.840 771.720 3.980 ;
        RECT 503.800 3.640 504.060 3.730 ;
        RECT 502.480 3.500 504.060 3.640 ;
        RECT 776.180 3.640 776.320 5.030 ;
        RECT 1548.390 5.000 1548.670 7.070 ;
        RECT 783.020 3.640 783.280 3.730 ;
        RECT 776.180 3.500 783.280 3.640 ;
        RECT 502.480 2.400 502.620 3.500 ;
        RECT 503.800 3.410 504.060 3.500 ;
        RECT 783.020 3.410 783.280 3.500 ;
        RECT 502.270 -4.800 502.830 2.400 ;
      LAYER via2 ;
        RECT 888.350 5.640 888.630 5.920 ;
        RECT 895.710 5.640 895.990 5.920 ;
      LAYER met3 ;
        RECT 888.325 5.930 888.655 5.945 ;
        RECT 895.685 5.930 896.015 5.945 ;
        RECT 888.325 5.630 896.015 5.930 ;
        RECT 888.325 5.615 888.655 5.630 ;
        RECT 895.685 5.615 896.015 5.630 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1083.905 9.605 1105.235 9.775 ;
        RECT 1083.905 9.095 1084.075 9.605 ;
        RECT 1075.625 8.925 1084.075 9.095 ;
        RECT 996.965 7.565 1004.035 7.735 ;
        RECT 996.965 7.395 997.135 7.565 ;
        RECT 994.665 7.225 997.135 7.395 ;
        RECT 883.345 4.165 890.875 4.335 ;
        RECT 773.405 1.275 773.575 3.655 ;
        RECT 798.705 1.275 798.875 3.315 ;
        RECT 831.365 2.295 831.535 3.315 ;
        RECT 883.345 2.975 883.515 4.165 ;
        RECT 890.705 3.655 890.875 4.165 ;
        RECT 899.445 3.655 899.615 7.055 ;
        RECT 890.705 3.485 899.615 3.655 ;
        RECT 881.965 2.805 883.515 2.975 ;
        RECT 852.065 2.465 879.375 2.635 ;
        RECT 852.065 2.295 852.235 2.465 ;
        RECT 831.365 2.125 852.235 2.295 ;
        RECT 994.665 2.125 994.835 7.225 ;
        RECT 1003.865 5.695 1004.035 7.565 ;
        RECT 1071.025 6.885 1072.115 7.055 ;
        RECT 1056.305 5.695 1056.475 6.715 ;
        RECT 1071.025 6.545 1071.195 6.885 ;
        RECT 1071.945 6.375 1072.115 6.885 ;
        RECT 1075.625 6.375 1075.795 8.925 ;
        RECT 1071.945 6.205 1075.795 6.375 ;
        RECT 1105.065 6.375 1105.235 9.605 ;
        RECT 1372.785 7.905 1401.935 8.075 ;
        RECT 1366.345 7.565 1370.195 7.735 ;
        RECT 1105.065 6.205 1121.335 6.375 ;
        RECT 1121.165 5.865 1121.335 6.205 ;
        RECT 1003.865 5.525 1056.475 5.695 ;
        RECT 1366.345 3.485 1366.515 7.565 ;
        RECT 1370.025 7.225 1370.195 7.565 ;
        RECT 1372.785 7.225 1372.955 7.905 ;
        RECT 773.405 1.105 798.875 1.275 ;
      LAYER mcon ;
        RECT 899.445 6.885 899.615 7.055 ;
        RECT 773.405 3.485 773.575 3.655 ;
        RECT 798.705 3.145 798.875 3.315 ;
        RECT 831.365 3.145 831.535 3.315 ;
        RECT 879.205 2.465 879.375 2.635 ;
        RECT 1056.305 6.545 1056.475 6.715 ;
        RECT 1401.765 7.905 1401.935 8.075 ;
      LAYER met1 ;
        RECT 920.990 8.060 921.310 8.120 ;
        RECT 1401.705 8.060 1401.995 8.105 ;
        RECT 1402.610 8.060 1402.930 8.120 ;
        RECT 920.990 7.920 953.880 8.060 ;
        RECT 920.990 7.860 921.310 7.920 ;
        RECT 953.740 7.720 953.880 7.920 ;
        RECT 1401.705 7.920 1402.930 8.060 ;
        RECT 1401.705 7.875 1401.995 7.920 ;
        RECT 1402.610 7.860 1402.930 7.920 ;
        RECT 989.070 7.720 989.390 7.780 ;
        RECT 953.740 7.580 989.390 7.720 ;
        RECT 989.070 7.520 989.390 7.580 ;
        RECT 1528.190 7.720 1528.510 7.780 ;
        RECT 1594.430 7.720 1594.750 7.780 ;
        RECT 1528.190 7.580 1594.750 7.720 ;
        RECT 1528.190 7.520 1528.510 7.580 ;
        RECT 1594.430 7.520 1594.750 7.580 ;
        RECT 1369.965 7.380 1370.255 7.425 ;
        RECT 1372.725 7.380 1373.015 7.425 ;
        RECT 1369.965 7.240 1373.015 7.380 ;
        RECT 1369.965 7.195 1370.255 7.240 ;
        RECT 1372.725 7.195 1373.015 7.240 ;
        RECT 899.370 7.040 899.690 7.100 ;
        RECT 899.370 6.900 899.885 7.040 ;
        RECT 899.370 6.840 899.690 6.900 ;
        RECT 1056.245 6.700 1056.535 6.745 ;
        RECT 1070.965 6.700 1071.255 6.745 ;
        RECT 1056.245 6.560 1071.255 6.700 ;
        RECT 1056.245 6.515 1056.535 6.560 ;
        RECT 1070.965 6.515 1071.255 6.560 ;
        RECT 1121.105 6.020 1121.395 6.065 ;
        RECT 1123.850 6.020 1124.170 6.080 ;
        RECT 1121.105 5.880 1124.170 6.020 ;
        RECT 1121.105 5.835 1121.395 5.880 ;
        RECT 1123.850 5.820 1124.170 5.880 ;
        RECT 767.810 3.640 768.130 3.700 ;
        RECT 773.345 3.640 773.635 3.685 ;
        RECT 767.810 3.500 773.635 3.640 ;
        RECT 767.810 3.440 768.130 3.500 ;
        RECT 773.345 3.455 773.635 3.500 ;
        RECT 1355.690 3.640 1356.010 3.700 ;
        RECT 1366.285 3.640 1366.575 3.685 ;
        RECT 1355.690 3.500 1366.575 3.640 ;
        RECT 1355.690 3.440 1356.010 3.500 ;
        RECT 1366.285 3.455 1366.575 3.500 ;
        RECT 798.645 3.300 798.935 3.345 ;
        RECT 804.610 3.300 804.930 3.360 ;
        RECT 798.645 3.160 804.930 3.300 ;
        RECT 798.645 3.115 798.935 3.160 ;
        RECT 804.610 3.100 804.930 3.160 ;
        RECT 830.830 3.300 831.150 3.360 ;
        RECT 831.305 3.300 831.595 3.345 ;
        RECT 830.830 3.160 831.595 3.300 ;
        RECT 830.830 3.100 831.150 3.160 ;
        RECT 831.305 3.115 831.595 3.160 ;
        RECT 1264.150 3.300 1264.470 3.360 ;
        RECT 1296.350 3.300 1296.670 3.360 ;
        RECT 1264.150 3.160 1296.670 3.300 ;
        RECT 1264.150 3.100 1264.470 3.160 ;
        RECT 1296.350 3.100 1296.670 3.160 ;
        RECT 881.905 2.960 882.195 3.005 ;
        RECT 880.140 2.820 882.195 2.960 ;
        RECT 879.145 2.620 879.435 2.665 ;
        RECT 880.140 2.620 880.280 2.820 ;
        RECT 881.905 2.775 882.195 2.820 ;
        RECT 879.145 2.480 880.280 2.620 ;
        RECT 879.145 2.435 879.435 2.480 ;
        RECT 993.670 2.280 993.990 2.340 ;
        RECT 994.605 2.280 994.895 2.325 ;
        RECT 993.670 2.140 994.895 2.280 ;
        RECT 993.670 2.080 993.990 2.140 ;
        RECT 994.605 2.095 994.895 2.140 ;
        RECT 1258.630 2.280 1258.950 2.340 ;
        RECT 1264.150 2.280 1264.470 2.340 ;
        RECT 1258.630 2.140 1264.470 2.280 ;
        RECT 1258.630 2.080 1258.950 2.140 ;
        RECT 1264.150 2.080 1264.470 2.140 ;
        RECT 1300.030 2.280 1300.350 2.340 ;
        RECT 1302.790 2.280 1303.110 2.340 ;
        RECT 1300.030 2.140 1303.110 2.280 ;
        RECT 1300.030 2.080 1300.350 2.140 ;
        RECT 1302.790 2.080 1303.110 2.140 ;
        RECT 1306.010 2.280 1306.330 2.340 ;
        RECT 1314.290 2.280 1314.610 2.340 ;
        RECT 1306.010 2.140 1314.610 2.280 ;
        RECT 1306.010 2.080 1306.330 2.140 ;
        RECT 1314.290 2.080 1314.610 2.140 ;
      LAYER via ;
        RECT 921.020 7.860 921.280 8.120 ;
        RECT 1402.640 7.860 1402.900 8.120 ;
        RECT 989.100 7.520 989.360 7.780 ;
        RECT 1528.220 7.520 1528.480 7.780 ;
        RECT 1594.460 7.520 1594.720 7.780 ;
        RECT 899.400 6.840 899.660 7.100 ;
        RECT 1123.880 5.820 1124.140 6.080 ;
        RECT 767.840 3.440 768.100 3.700 ;
        RECT 1355.720 3.440 1355.980 3.700 ;
        RECT 804.640 3.100 804.900 3.360 ;
        RECT 830.860 3.100 831.120 3.360 ;
        RECT 1264.180 3.100 1264.440 3.360 ;
        RECT 1296.380 3.100 1296.640 3.360 ;
        RECT 993.700 2.080 993.960 2.340 ;
        RECT 1258.660 2.080 1258.920 2.340 ;
        RECT 1264.180 2.080 1264.440 2.340 ;
        RECT 1300.060 2.080 1300.320 2.340 ;
        RECT 1302.820 2.080 1303.080 2.340 ;
        RECT 1306.040 2.080 1306.300 2.340 ;
        RECT 1314.320 2.080 1314.580 2.340 ;
      LAYER met2 ;
        RECT 919.240 8.430 921.220 8.570 ;
        RECT 899.390 7.635 899.670 8.005 ;
        RECT 908.590 7.890 908.870 8.005 ;
        RECT 919.240 7.890 919.380 8.430 ;
        RECT 921.080 8.150 921.220 8.430 ;
        RECT 908.590 7.750 919.380 7.890 ;
        RECT 921.020 7.830 921.280 8.150 ;
        RECT 1402.640 8.005 1402.900 8.150 ;
        RECT 908.590 7.635 908.870 7.750 ;
        RECT 989.100 7.720 989.360 7.810 ;
        RECT 899.460 7.130 899.600 7.635 ;
        RECT 989.100 7.580 991.600 7.720 ;
        RECT 1402.630 7.635 1402.910 8.005 ;
        RECT 1478.070 7.635 1478.350 8.005 ;
        RECT 1481.290 7.890 1481.570 8.005 ;
        RECT 1480.900 7.750 1481.570 7.890 ;
        RECT 989.100 7.490 989.360 7.580 ;
        RECT 899.400 6.810 899.660 7.130 ;
        RECT 991.460 5.850 991.600 7.580 ;
        RECT 1478.140 7.210 1478.280 7.635 ;
        RECT 1480.900 7.210 1481.040 7.750 ;
        RECT 1481.290 7.635 1481.570 7.750 ;
        RECT 1528.210 7.635 1528.490 8.005 ;
        RECT 1595.770 7.890 1596.050 9.000 ;
        RECT 1594.520 7.810 1596.050 7.890 ;
        RECT 1594.460 7.750 1596.050 7.810 ;
        RECT 1528.220 7.490 1528.480 7.635 ;
        RECT 1594.460 7.490 1594.720 7.750 ;
        RECT 1478.140 7.070 1481.040 7.210 ;
        RECT 1236.570 6.275 1236.850 6.645 ;
        RECT 991.460 5.710 992.520 5.850 ;
        RECT 1123.880 5.790 1124.140 6.110 ;
        RECT 992.380 5.170 992.520 5.710 ;
        RECT 992.380 5.030 993.900 5.170 ;
        RECT 519.890 3.555 520.170 3.925 ;
        RECT 519.960 2.400 520.100 3.555 ;
        RECT 755.940 3.500 759.300 3.640 ;
        RECT 754.030 2.450 754.310 2.565 ;
        RECT 755.940 2.450 756.080 3.500 ;
        RECT 759.160 3.130 759.300 3.500 ;
        RECT 767.840 3.410 768.100 3.730 ;
        RECT 767.900 3.130 768.040 3.410 ;
        RECT 759.160 2.990 768.040 3.130 ;
        RECT 804.640 3.130 804.900 3.390 ;
        RECT 830.860 3.300 831.120 3.390 ;
        RECT 808.770 3.130 809.050 3.245 ;
        RECT 804.640 3.070 806.680 3.130 ;
        RECT 804.700 2.990 806.680 3.070 ;
        RECT 519.750 -4.800 520.310 2.400 ;
        RECT 754.030 2.310 756.080 2.450 ;
        RECT 754.030 2.195 754.310 2.310 ;
        RECT 806.540 1.090 806.680 2.990 ;
        RECT 807.460 2.990 809.050 3.130 ;
        RECT 807.460 1.090 807.600 2.990 ;
        RECT 808.770 2.875 809.050 2.990 ;
        RECT 817.510 3.130 817.790 3.245 ;
        RECT 820.340 3.160 831.120 3.300 ;
        RECT 820.340 3.130 820.480 3.160 ;
        RECT 817.510 2.990 820.480 3.130 ;
        RECT 830.860 3.070 831.120 3.160 ;
        RECT 817.510 2.875 817.790 2.990 ;
        RECT 993.760 2.370 993.900 5.030 ;
        RECT 1123.940 4.490 1124.080 5.790 ;
        RECT 1157.450 4.490 1157.730 4.605 ;
        RECT 1123.940 4.350 1157.730 4.490 ;
        RECT 1236.640 4.490 1236.780 6.275 ;
        RECT 1595.770 5.000 1596.050 7.750 ;
        RECT 1236.640 4.350 1240.000 4.490 ;
        RECT 1157.450 4.235 1157.730 4.350 ;
        RECT 1239.860 3.810 1240.000 4.350 ;
        RECT 1239.860 3.670 1256.100 3.810 ;
        RECT 1255.960 3.300 1256.100 3.670 ;
        RECT 1314.310 3.555 1314.590 3.925 ;
        RECT 1329.950 3.810 1330.230 3.925 ;
        RECT 1331.330 3.810 1331.610 3.925 ;
        RECT 1329.950 3.670 1331.610 3.810 ;
        RECT 1329.950 3.555 1330.230 3.670 ;
        RECT 1331.330 3.555 1331.610 3.670 ;
        RECT 1355.250 3.810 1355.530 3.925 ;
        RECT 1355.250 3.730 1355.920 3.810 ;
        RECT 1355.250 3.670 1355.980 3.730 ;
        RECT 1355.250 3.555 1355.530 3.670 ;
        RECT 1255.960 3.160 1258.860 3.300 ;
        RECT 1258.720 2.370 1258.860 3.160 ;
        RECT 1264.180 3.070 1264.440 3.390 ;
        RECT 1296.380 3.130 1296.640 3.390 ;
        RECT 1296.380 3.070 1300.260 3.130 ;
        RECT 1264.240 2.370 1264.380 3.070 ;
        RECT 1296.440 2.990 1300.260 3.070 ;
        RECT 1300.120 2.370 1300.260 2.990 ;
        RECT 1302.880 2.990 1306.240 3.130 ;
        RECT 1302.880 2.370 1303.020 2.990 ;
        RECT 1306.100 2.370 1306.240 2.990 ;
        RECT 1314.380 2.370 1314.520 3.555 ;
        RECT 1355.720 3.410 1355.980 3.670 ;
        RECT 993.700 2.050 993.960 2.370 ;
        RECT 1258.660 2.050 1258.920 2.370 ;
        RECT 1264.180 2.050 1264.440 2.370 ;
        RECT 1300.060 2.050 1300.320 2.370 ;
        RECT 1302.820 2.050 1303.080 2.370 ;
        RECT 1306.040 2.050 1306.300 2.370 ;
        RECT 1314.320 2.050 1314.580 2.370 ;
        RECT 806.540 0.950 807.600 1.090 ;
      LAYER via2 ;
        RECT 899.390 7.680 899.670 7.960 ;
        RECT 908.590 7.680 908.870 7.960 ;
        RECT 1402.630 7.680 1402.910 7.960 ;
        RECT 1478.070 7.680 1478.350 7.960 ;
        RECT 1481.290 7.680 1481.570 7.960 ;
        RECT 1528.210 7.680 1528.490 7.960 ;
        RECT 1236.570 6.320 1236.850 6.600 ;
        RECT 519.890 3.600 520.170 3.880 ;
        RECT 754.030 2.240 754.310 2.520 ;
        RECT 808.770 2.920 809.050 3.200 ;
        RECT 817.510 2.920 817.790 3.200 ;
        RECT 1157.450 4.280 1157.730 4.560 ;
        RECT 1314.310 3.600 1314.590 3.880 ;
        RECT 1329.950 3.600 1330.230 3.880 ;
        RECT 1331.330 3.600 1331.610 3.880 ;
        RECT 1355.250 3.600 1355.530 3.880 ;
      LAYER met3 ;
        RECT 899.365 7.970 899.695 7.985 ;
        RECT 908.565 7.970 908.895 7.985 ;
        RECT 899.365 7.670 908.895 7.970 ;
        RECT 899.365 7.655 899.695 7.670 ;
        RECT 908.565 7.655 908.895 7.670 ;
        RECT 1402.605 7.970 1402.935 7.985 ;
        RECT 1478.045 7.970 1478.375 7.985 ;
        RECT 1402.605 7.670 1427.530 7.970 ;
        RECT 1402.605 7.655 1402.935 7.670 ;
        RECT 1427.230 7.290 1427.530 7.670 ;
        RECT 1429.070 7.670 1478.375 7.970 ;
        RECT 1429.070 7.290 1429.370 7.670 ;
        RECT 1478.045 7.655 1478.375 7.670 ;
        RECT 1481.265 7.970 1481.595 7.985 ;
        RECT 1528.185 7.970 1528.515 7.985 ;
        RECT 1481.265 7.670 1528.515 7.970 ;
        RECT 1481.265 7.655 1481.595 7.670 ;
        RECT 1528.185 7.655 1528.515 7.670 ;
        RECT 1427.230 6.990 1429.370 7.290 ;
        RECT 1228.470 6.610 1228.850 6.620 ;
        RECT 1236.545 6.610 1236.875 6.625 ;
        RECT 1228.470 6.310 1236.875 6.610 ;
        RECT 1228.470 6.300 1228.850 6.310 ;
        RECT 1236.545 6.295 1236.875 6.310 ;
        RECT 1157.425 4.570 1157.755 4.585 ;
        RECT 1163.150 4.570 1163.530 4.580 ;
        RECT 1157.425 4.270 1163.530 4.570 ;
        RECT 1157.425 4.255 1157.755 4.270 ;
        RECT 1163.150 4.260 1163.530 4.270 ;
        RECT 519.865 3.890 520.195 3.905 ;
        RECT 534.790 3.890 535.170 3.900 ;
        RECT 519.865 3.590 535.170 3.890 ;
        RECT 519.865 3.575 520.195 3.590 ;
        RECT 534.790 3.580 535.170 3.590 ;
        RECT 1314.285 3.890 1314.615 3.905 ;
        RECT 1329.925 3.890 1330.255 3.905 ;
        RECT 1314.285 3.590 1330.255 3.890 ;
        RECT 1314.285 3.575 1314.615 3.590 ;
        RECT 1329.925 3.575 1330.255 3.590 ;
        RECT 1331.305 3.890 1331.635 3.905 ;
        RECT 1355.225 3.890 1355.555 3.905 ;
        RECT 1331.305 3.590 1355.555 3.890 ;
        RECT 1331.305 3.575 1331.635 3.590 ;
        RECT 1355.225 3.575 1355.555 3.590 ;
        RECT 808.745 3.210 809.075 3.225 ;
        RECT 817.485 3.210 817.815 3.225 ;
        RECT 808.745 2.910 817.815 3.210 ;
        RECT 808.745 2.895 809.075 2.910 ;
        RECT 817.485 2.895 817.815 2.910 ;
        RECT 754.005 2.540 754.335 2.545 ;
        RECT 753.750 2.530 754.335 2.540 ;
        RECT 753.550 2.230 754.335 2.530 ;
        RECT 753.750 2.220 754.335 2.230 ;
        RECT 754.005 2.215 754.335 2.220 ;
      LAYER via3 ;
        RECT 1228.500 6.300 1228.820 6.620 ;
        RECT 1163.180 4.260 1163.500 4.580 ;
        RECT 534.820 3.580 535.140 3.900 ;
        RECT 753.780 2.220 754.100 2.540 ;
      LAYER met4 ;
        RECT 1228.495 6.295 1228.825 6.625 ;
        RECT 1163.175 4.255 1163.505 4.585 ;
        RECT 534.815 3.890 535.145 3.905 ;
        RECT 1163.190 3.890 1163.490 4.255 ;
        RECT 534.815 3.590 536.050 3.890 ;
        RECT 1163.190 3.590 1166.250 3.890 ;
        RECT 534.815 3.575 535.145 3.590 ;
        RECT 535.750 1.850 536.050 3.590 ;
        RECT 653.510 2.910 672.210 3.210 ;
        RECT 537.150 1.850 538.330 2.290 ;
        RECT 535.750 1.550 538.330 1.850 ;
        RECT 537.150 1.110 538.330 1.550 ;
        RECT 617.190 1.850 618.370 2.290 ;
        RECT 653.510 1.850 653.810 2.910 ;
        RECT 617.190 1.550 653.810 1.850 ;
        RECT 671.910 1.850 672.210 2.910 ;
        RECT 753.775 2.290 754.105 2.545 ;
        RECT 1165.950 2.290 1166.250 3.590 ;
        RECT 1228.510 2.290 1228.810 6.295 ;
        RECT 673.310 1.850 674.490 2.290 ;
        RECT 671.910 1.550 674.490 1.850 ;
        RECT 617.190 1.110 618.370 1.550 ;
        RECT 673.310 1.110 674.490 1.550 ;
        RECT 753.350 1.110 754.530 2.290 ;
        RECT 1165.510 1.110 1166.690 2.290 ;
        RECT 1228.070 1.110 1229.250 2.290 ;
      LAYER met5 ;
        RECT 536.940 0.900 618.580 2.500 ;
        RECT 673.100 0.900 754.740 2.500 ;
        RECT 1165.300 0.900 1229.460 2.500 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 741.665 9.945 758.395 10.115 ;
        RECT 550.305 9.265 559.675 9.435 ;
        RECT 550.305 4.335 550.475 9.265 ;
        RECT 559.505 9.095 559.675 9.265 ;
        RECT 559.045 8.925 559.675 9.095 ;
        RECT 725.105 8.925 733.555 9.095 ;
        RECT 559.045 7.905 559.215 8.925 ;
        RECT 641.845 8.585 646.155 8.755 ;
        RECT 627.585 6.205 627.755 7.395 ;
        RECT 630.345 6.205 630.515 8.075 ;
        RECT 636.785 7.395 636.955 8.075 ;
        RECT 636.785 7.225 640.635 7.395 ;
        RECT 641.845 7.225 642.015 8.585 ;
        RECT 645.985 7.735 646.155 8.585 ;
        RECT 645.985 7.565 664.095 7.735 ;
        RECT 663.925 6.885 664.095 7.565 ;
        RECT 720.045 7.225 721.595 7.395 ;
        RECT 725.105 7.225 725.275 8.925 ;
        RECT 733.385 8.075 733.555 8.925 ;
        RECT 741.665 8.075 741.835 9.945 ;
        RECT 758.225 8.925 758.395 9.945 ;
        RECT 1163.945 9.605 1196.315 9.775 ;
        RECT 1159.805 9.265 1161.355 9.435 ;
        RECT 733.385 7.905 741.835 8.075 ;
        RECT 761.445 7.905 761.615 9.095 ;
        RECT 820.325 8.925 849.015 9.095 ;
        RECT 763.285 7.225 763.455 8.075 ;
        RECT 820.325 7.225 820.495 8.925 ;
        RECT 848.845 7.735 849.015 8.925 ;
        RECT 879.665 8.925 890.875 9.095 ;
        RECT 846.085 7.565 849.015 7.735 ;
        RECT 867.705 7.905 871.095 8.075 ;
        RECT 846.085 7.055 846.255 7.565 ;
        RECT 867.705 7.225 867.875 7.905 ;
        RECT 870.925 7.395 871.095 7.905 ;
        RECT 879.665 7.395 879.835 8.925 ;
        RECT 890.705 7.735 890.875 8.925 ;
        RECT 1055.385 7.905 1056.475 8.075 ;
        RECT 890.705 7.565 893.635 7.735 ;
        RECT 870.925 7.225 879.835 7.395 ;
        RECT 846.085 6.885 847.635 7.055 ;
        RECT 893.465 6.885 893.635 7.565 ;
        RECT 959.705 7.225 983.335 7.395 ;
        RECT 984.545 7.055 984.715 7.395 ;
        RECT 993.745 7.055 993.915 7.735 ;
        RECT 1055.385 7.565 1055.555 7.905 ;
        RECT 1056.305 7.395 1056.475 7.905 ;
        RECT 1056.305 7.225 1057.395 7.395 ;
        RECT 1100.925 7.225 1102.015 7.395 ;
        RECT 1159.805 7.225 1159.975 9.265 ;
        RECT 1161.185 9.095 1161.355 9.265 ;
        RECT 1161.185 8.925 1161.815 9.095 ;
        RECT 1161.645 7.735 1161.815 8.925 ;
        RECT 1163.945 7.735 1164.115 9.605 ;
        RECT 1161.645 7.565 1164.115 7.735 ;
        RECT 1196.145 7.395 1196.315 9.605 ;
        RECT 1196.145 7.225 1207.355 7.395 ;
        RECT 984.545 6.885 993.915 7.055 ;
        RECT 1249.045 7.055 1249.215 7.395 ;
        RECT 1254.565 7.055 1254.735 8.755 ;
        RECT 1249.045 6.885 1254.735 7.055 ;
        RECT 1257.325 7.055 1257.495 8.755 ;
        RECT 1402.225 8.245 1403.775 8.415 ;
        RECT 1402.225 7.735 1402.395 8.245 ;
        RECT 1400.845 7.565 1402.395 7.735 ;
        RECT 1400.845 7.395 1401.015 7.565 ;
        RECT 1302.865 7.225 1304.415 7.395 ;
        RECT 1257.325 6.885 1257.955 7.055 ;
        RECT 1257.785 6.205 1257.955 6.885 ;
        RECT 1304.245 6.715 1304.415 7.225 ;
        RECT 1305.625 7.225 1315.915 7.395 ;
        RECT 1305.625 6.715 1305.795 7.225 ;
        RECT 1304.245 6.545 1305.795 6.715 ;
        RECT 546.625 4.165 550.475 4.335 ;
        RECT 1325.405 3.315 1325.575 7.395 ;
        RECT 1397.625 7.225 1401.015 7.395 ;
        RECT 1325.405 3.145 1335.695 3.315 ;
        RECT 1403.605 2.975 1403.775 8.245 ;
        RECT 1600.945 7.565 1602.495 7.735 ;
        RECT 1447.765 7.225 1451.615 7.395 ;
        RECT 1451.445 5.865 1451.615 7.225 ;
        RECT 1486.405 7.225 1500.375 7.395 ;
        RECT 1408.665 2.975 1408.835 3.655 ;
        RECT 1427.525 3.315 1427.695 3.655 ;
        RECT 1427.525 3.145 1428.155 3.315 ;
        RECT 1403.605 2.805 1408.835 2.975 ;
        RECT 1427.985 2.975 1428.155 3.145 ;
        RECT 1427.985 2.805 1428.615 2.975 ;
        RECT 1428.445 2.635 1428.615 2.805 ;
        RECT 1428.445 2.465 1429.535 2.635 ;
        RECT 1469.845 2.465 1470.015 6.035 ;
        RECT 1486.405 2.975 1486.575 7.225 ;
        RECT 1545.745 6.035 1545.915 7.395 ;
        RECT 1592.205 7.225 1593.295 7.395 ;
        RECT 1600.945 7.225 1601.115 7.565 ;
        RECT 1602.325 7.395 1602.495 7.565 ;
        RECT 1602.325 7.225 1602.955 7.395 ;
        RECT 1602.785 7.055 1602.955 7.225 ;
        RECT 1602.785 6.885 1609.395 7.055 ;
        RECT 1545.745 5.865 1547.295 6.035 ;
        RECT 1485.945 2.805 1486.575 2.975 ;
        RECT 1485.945 2.635 1486.115 2.805 ;
        RECT 1483.645 2.465 1486.115 2.635 ;
        RECT 1609.225 2.465 1609.395 6.885 ;
        RECT 1614.745 4.845 1617.675 5.015 ;
        RECT 1614.745 2.465 1614.915 4.845 ;
        RECT 1617.505 4.505 1617.675 4.845 ;
        RECT 1429.365 1.445 1429.535 2.465 ;
      LAYER mcon ;
        RECT 630.345 7.905 630.515 8.075 ;
        RECT 627.585 7.225 627.755 7.395 ;
        RECT 636.785 7.905 636.955 8.075 ;
        RECT 640.465 7.225 640.635 7.395 ;
        RECT 761.445 8.925 761.615 9.095 ;
        RECT 763.285 7.905 763.455 8.075 ;
        RECT 721.425 7.225 721.595 7.395 ;
        RECT 993.745 7.565 993.915 7.735 ;
        RECT 983.165 7.225 983.335 7.395 ;
        RECT 984.545 7.225 984.715 7.395 ;
        RECT 847.465 6.885 847.635 7.055 ;
        RECT 1057.225 7.225 1057.395 7.395 ;
        RECT 1101.845 7.225 1102.015 7.395 ;
        RECT 1254.565 8.585 1254.735 8.755 ;
        RECT 1207.185 7.225 1207.355 7.395 ;
        RECT 1249.045 7.225 1249.215 7.395 ;
        RECT 1257.325 8.585 1257.495 8.755 ;
        RECT 1315.745 7.225 1315.915 7.395 ;
        RECT 1325.405 7.225 1325.575 7.395 ;
        RECT 1335.525 3.145 1335.695 3.315 ;
        RECT 1500.205 7.225 1500.375 7.395 ;
        RECT 1545.745 7.225 1545.915 7.395 ;
        RECT 1593.125 7.225 1593.295 7.395 ;
        RECT 1469.845 5.865 1470.015 6.035 ;
        RECT 1408.665 3.485 1408.835 3.655 ;
        RECT 1427.525 3.485 1427.695 3.655 ;
        RECT 1547.125 5.865 1547.295 6.035 ;
      LAYER met1 ;
        RECT 758.165 9.080 758.455 9.125 ;
        RECT 761.385 9.080 761.675 9.125 ;
        RECT 758.165 8.940 761.675 9.080 ;
        RECT 758.165 8.895 758.455 8.940 ;
        RECT 761.385 8.895 761.675 8.940 ;
        RECT 951.810 8.740 952.130 8.800 ;
        RECT 955.030 8.740 955.350 8.800 ;
        RECT 951.810 8.600 955.350 8.740 ;
        RECT 951.810 8.540 952.130 8.600 ;
        RECT 955.030 8.540 955.350 8.600 ;
        RECT 1254.505 8.740 1254.795 8.785 ;
        RECT 1257.265 8.740 1257.555 8.785 ;
        RECT 1254.505 8.600 1257.555 8.740 ;
        RECT 1254.505 8.555 1254.795 8.600 ;
        RECT 1257.265 8.555 1257.555 8.600 ;
        RECT 558.985 8.060 559.275 8.105 ;
        RECT 560.810 8.060 561.130 8.120 ;
        RECT 558.985 7.920 561.130 8.060 ;
        RECT 558.985 7.875 559.275 7.920 ;
        RECT 560.810 7.860 561.130 7.920 ;
        RECT 630.285 8.060 630.575 8.105 ;
        RECT 636.725 8.060 637.015 8.105 ;
        RECT 630.285 7.920 637.015 8.060 ;
        RECT 630.285 7.875 630.575 7.920 ;
        RECT 636.725 7.875 637.015 7.920 ;
        RECT 761.385 8.060 761.675 8.105 ;
        RECT 763.225 8.060 763.515 8.105 ;
        RECT 761.385 7.920 763.515 8.060 ;
        RECT 761.385 7.875 761.675 7.920 ;
        RECT 763.225 7.875 763.515 7.920 ;
        RECT 1360.750 8.060 1361.070 8.120 ;
        RECT 1369.490 8.060 1369.810 8.120 ;
        RECT 1360.750 7.920 1369.810 8.060 ;
        RECT 1360.750 7.860 1361.070 7.920 ;
        RECT 1369.490 7.860 1369.810 7.920 ;
        RECT 949.970 7.520 950.290 7.780 ;
        RECT 993.685 7.720 993.975 7.765 ;
        RECT 995.510 7.720 995.830 7.780 ;
        RECT 1055.325 7.720 1055.615 7.765 ;
        RECT 993.685 7.580 995.830 7.720 ;
        RECT 993.685 7.535 993.975 7.580 ;
        RECT 995.510 7.520 995.830 7.580 ;
        RECT 1023.660 7.580 1055.615 7.720 ;
        RECT 613.710 7.380 614.030 7.440 ;
        RECT 627.525 7.380 627.815 7.425 ;
        RECT 613.710 7.240 627.815 7.380 ;
        RECT 613.710 7.180 614.030 7.240 ;
        RECT 627.525 7.195 627.815 7.240 ;
        RECT 640.405 7.380 640.695 7.425 ;
        RECT 641.785 7.380 642.075 7.425 ;
        RECT 719.985 7.380 720.275 7.425 ;
        RECT 640.405 7.240 642.075 7.380 ;
        RECT 640.405 7.195 640.695 7.240 ;
        RECT 641.785 7.195 642.075 7.240 ;
        RECT 671.760 7.240 720.275 7.380 ;
        RECT 663.865 7.040 664.155 7.085 ;
        RECT 671.760 7.040 671.900 7.240 ;
        RECT 719.985 7.195 720.275 7.240 ;
        RECT 721.365 7.380 721.655 7.425 ;
        RECT 725.045 7.380 725.335 7.425 ;
        RECT 721.365 7.240 725.335 7.380 ;
        RECT 721.365 7.195 721.655 7.240 ;
        RECT 725.045 7.195 725.335 7.240 ;
        RECT 763.225 7.380 763.515 7.425 ;
        RECT 820.265 7.380 820.555 7.425 ;
        RECT 763.225 7.240 820.555 7.380 ;
        RECT 763.225 7.195 763.515 7.240 ;
        RECT 820.265 7.195 820.555 7.240 ;
        RECT 867.645 7.195 867.935 7.425 ;
        RECT 913.170 7.380 913.490 7.440 ;
        RECT 950.060 7.380 950.200 7.520 ;
        RECT 913.170 7.240 950.200 7.380 ;
        RECT 959.170 7.380 959.490 7.440 ;
        RECT 959.645 7.380 959.935 7.425 ;
        RECT 959.170 7.240 959.935 7.380 ;
        RECT 663.865 6.900 671.900 7.040 ;
        RECT 847.405 7.040 847.695 7.085 ;
        RECT 867.720 7.040 867.860 7.195 ;
        RECT 913.170 7.180 913.490 7.240 ;
        RECT 959.170 7.180 959.490 7.240 ;
        RECT 959.645 7.195 959.935 7.240 ;
        RECT 983.105 7.380 983.395 7.425 ;
        RECT 984.485 7.380 984.775 7.425 ;
        RECT 983.105 7.240 984.775 7.380 ;
        RECT 983.105 7.195 983.395 7.240 ;
        RECT 984.485 7.195 984.775 7.240 ;
        RECT 1022.650 7.380 1022.970 7.440 ;
        RECT 1023.660 7.380 1023.800 7.580 ;
        RECT 1055.325 7.535 1055.615 7.580 ;
        RECT 1122.100 7.580 1123.160 7.720 ;
        RECT 1022.650 7.240 1023.800 7.380 ;
        RECT 1057.165 7.380 1057.455 7.425 ;
        RECT 1100.865 7.380 1101.155 7.425 ;
        RECT 1057.165 7.240 1101.155 7.380 ;
        RECT 1022.650 7.180 1022.970 7.240 ;
        RECT 1057.165 7.195 1057.455 7.240 ;
        RECT 1100.865 7.195 1101.155 7.240 ;
        RECT 1101.785 7.380 1102.075 7.425 ;
        RECT 1122.100 7.380 1122.240 7.580 ;
        RECT 1101.785 7.240 1122.240 7.380 ;
        RECT 1101.785 7.195 1102.075 7.240 ;
        RECT 847.405 6.900 867.860 7.040 ;
        RECT 893.405 7.040 893.695 7.085 ;
        RECT 898.910 7.040 899.230 7.100 ;
        RECT 893.405 6.900 899.230 7.040 ;
        RECT 1123.020 7.040 1123.160 7.580 ;
        RECT 1159.745 7.380 1160.035 7.425 ;
        RECT 1124.860 7.240 1160.035 7.380 ;
        RECT 1124.860 7.040 1125.000 7.240 ;
        RECT 1159.745 7.195 1160.035 7.240 ;
        RECT 1207.125 7.380 1207.415 7.425 ;
        RECT 1248.985 7.380 1249.275 7.425 ;
        RECT 1207.125 7.240 1249.275 7.380 ;
        RECT 1207.125 7.195 1207.415 7.240 ;
        RECT 1248.985 7.195 1249.275 7.240 ;
        RECT 1302.805 7.195 1303.095 7.425 ;
        RECT 1315.685 7.380 1315.975 7.425 ;
        RECT 1325.345 7.380 1325.635 7.425 ;
        RECT 1315.685 7.240 1325.635 7.380 ;
        RECT 1315.685 7.195 1315.975 7.240 ;
        RECT 1325.345 7.195 1325.635 7.240 ;
        RECT 1347.410 7.380 1347.730 7.440 ;
        RECT 1356.610 7.380 1356.930 7.440 ;
        RECT 1397.550 7.380 1397.870 7.440 ;
        RECT 1347.410 7.240 1356.930 7.380 ;
        RECT 1397.355 7.240 1397.870 7.380 ;
        RECT 1123.020 6.900 1125.000 7.040 ;
        RECT 1295.890 7.040 1296.210 7.100 ;
        RECT 1302.880 7.040 1303.020 7.195 ;
        RECT 1347.410 7.180 1347.730 7.240 ;
        RECT 1356.610 7.180 1356.930 7.240 ;
        RECT 1397.550 7.180 1397.870 7.240 ;
        RECT 1446.770 7.380 1447.090 7.440 ;
        RECT 1447.705 7.380 1447.995 7.425 ;
        RECT 1446.770 7.240 1447.995 7.380 ;
        RECT 1446.770 7.180 1447.090 7.240 ;
        RECT 1447.705 7.195 1447.995 7.240 ;
        RECT 1500.145 7.380 1500.435 7.425 ;
        RECT 1545.685 7.380 1545.975 7.425 ;
        RECT 1500.145 7.240 1545.975 7.380 ;
        RECT 1500.145 7.195 1500.435 7.240 ;
        RECT 1545.685 7.195 1545.975 7.240 ;
        RECT 1592.130 7.380 1592.450 7.440 ;
        RECT 1593.065 7.380 1593.355 7.425 ;
        RECT 1600.885 7.380 1601.175 7.425 ;
        RECT 1592.130 7.240 1592.645 7.380 ;
        RECT 1593.065 7.240 1601.175 7.380 ;
        RECT 1592.130 7.180 1592.450 7.240 ;
        RECT 1593.065 7.195 1593.355 7.240 ;
        RECT 1600.885 7.195 1601.175 7.240 ;
        RECT 1295.890 6.900 1303.020 7.040 ;
        RECT 663.865 6.855 664.155 6.900 ;
        RECT 847.405 6.855 847.695 6.900 ;
        RECT 893.405 6.855 893.695 6.900 ;
        RECT 898.910 6.840 899.230 6.900 ;
        RECT 1295.890 6.840 1296.210 6.900 ;
        RECT 627.525 6.360 627.815 6.405 ;
        RECT 630.285 6.360 630.575 6.405 ;
        RECT 627.525 6.220 630.575 6.360 ;
        RECT 627.525 6.175 627.815 6.220 ;
        RECT 630.285 6.175 630.575 6.220 ;
        RECT 1257.725 6.360 1258.015 6.405 ;
        RECT 1265.530 6.360 1265.850 6.420 ;
        RECT 1257.725 6.220 1265.850 6.360 ;
        RECT 1257.725 6.175 1258.015 6.220 ;
        RECT 1265.530 6.160 1265.850 6.220 ;
        RECT 1356.610 6.360 1356.930 6.420 ;
        RECT 1360.750 6.360 1361.070 6.420 ;
        RECT 1356.610 6.220 1361.070 6.360 ;
        RECT 1356.610 6.160 1356.930 6.220 ;
        RECT 1360.750 6.160 1361.070 6.220 ;
        RECT 1369.490 6.360 1369.810 6.420 ;
        RECT 1397.550 6.360 1397.870 6.420 ;
        RECT 1369.490 6.220 1397.870 6.360 ;
        RECT 1369.490 6.160 1369.810 6.220 ;
        RECT 1397.550 6.160 1397.870 6.220 ;
        RECT 1451.385 6.020 1451.675 6.065 ;
        RECT 1452.750 6.020 1453.070 6.080 ;
        RECT 1451.385 5.880 1453.070 6.020 ;
        RECT 1451.385 5.835 1451.675 5.880 ;
        RECT 1452.750 5.820 1453.070 5.880 ;
        RECT 1455.050 6.020 1455.370 6.080 ;
        RECT 1469.785 6.020 1470.075 6.065 ;
        RECT 1455.050 5.880 1470.075 6.020 ;
        RECT 1455.050 5.820 1455.370 5.880 ;
        RECT 1469.785 5.835 1470.075 5.880 ;
        RECT 1547.065 6.020 1547.355 6.065 ;
        RECT 1592.130 6.020 1592.450 6.080 ;
        RECT 1547.065 5.880 1592.450 6.020 ;
        RECT 1547.065 5.835 1547.355 5.880 ;
        RECT 1592.130 5.820 1592.450 5.880 ;
        RECT 1617.445 4.660 1617.735 4.705 ;
        RECT 1643.650 4.660 1643.970 4.720 ;
        RECT 1617.445 4.520 1643.970 4.660 ;
        RECT 1617.445 4.475 1617.735 4.520 ;
        RECT 1643.650 4.460 1643.970 4.520 ;
        RECT 546.565 4.320 546.855 4.365 ;
        RECT 544.800 4.180 546.855 4.320 ;
        RECT 540.110 3.980 540.430 4.040 ;
        RECT 544.800 3.980 544.940 4.180 ;
        RECT 546.565 4.135 546.855 4.180 ;
        RECT 540.110 3.840 544.940 3.980 ;
        RECT 540.110 3.780 540.430 3.840 ;
        RECT 1408.605 3.640 1408.895 3.685 ;
        RECT 1427.465 3.640 1427.755 3.685 ;
        RECT 1408.605 3.500 1427.755 3.640 ;
        RECT 1408.605 3.455 1408.895 3.500 ;
        RECT 1427.465 3.455 1427.755 3.500 ;
        RECT 1335.465 3.300 1335.755 3.345 ;
        RECT 1335.910 3.300 1336.230 3.360 ;
        RECT 1335.465 3.160 1336.230 3.300 ;
        RECT 1335.465 3.115 1335.755 3.160 ;
        RECT 1335.910 3.100 1336.230 3.160 ;
        RECT 1469.785 2.620 1470.075 2.665 ;
        RECT 1483.585 2.620 1483.875 2.665 ;
        RECT 1469.785 2.480 1483.875 2.620 ;
        RECT 1469.785 2.435 1470.075 2.480 ;
        RECT 1483.585 2.435 1483.875 2.480 ;
        RECT 1609.165 2.620 1609.455 2.665 ;
        RECT 1614.685 2.620 1614.975 2.665 ;
        RECT 1609.165 2.480 1614.975 2.620 ;
        RECT 1609.165 2.435 1609.455 2.480 ;
        RECT 1614.685 2.435 1614.975 2.480 ;
        RECT 1265.530 2.280 1265.850 2.340 ;
        RECT 1295.890 2.280 1296.210 2.340 ;
        RECT 1265.530 2.140 1296.210 2.280 ;
        RECT 1265.530 2.080 1265.850 2.140 ;
        RECT 1295.890 2.080 1296.210 2.140 ;
        RECT 1345.110 2.280 1345.430 2.340 ;
        RECT 1347.410 2.280 1347.730 2.340 ;
        RECT 1345.110 2.140 1347.730 2.280 ;
        RECT 1345.110 2.080 1345.430 2.140 ;
        RECT 1347.410 2.080 1347.730 2.140 ;
        RECT 1429.305 1.600 1429.595 1.645 ;
        RECT 1444.470 1.600 1444.790 1.660 ;
        RECT 1429.305 1.460 1444.790 1.600 ;
        RECT 1429.305 1.415 1429.595 1.460 ;
        RECT 1444.470 1.400 1444.790 1.460 ;
      LAYER via ;
        RECT 951.840 8.540 952.100 8.800 ;
        RECT 955.060 8.540 955.320 8.800 ;
        RECT 560.840 7.860 561.100 8.120 ;
        RECT 1360.780 7.860 1361.040 8.120 ;
        RECT 1369.520 7.860 1369.780 8.120 ;
        RECT 950.000 7.520 950.260 7.780 ;
        RECT 995.540 7.520 995.800 7.780 ;
        RECT 613.740 7.180 614.000 7.440 ;
        RECT 913.200 7.180 913.460 7.440 ;
        RECT 959.200 7.180 959.460 7.440 ;
        RECT 1022.680 7.180 1022.940 7.440 ;
        RECT 898.940 6.840 899.200 7.100 ;
        RECT 1295.920 6.840 1296.180 7.100 ;
        RECT 1347.440 7.180 1347.700 7.440 ;
        RECT 1356.640 7.180 1356.900 7.440 ;
        RECT 1397.580 7.180 1397.840 7.440 ;
        RECT 1446.800 7.180 1447.060 7.440 ;
        RECT 1592.160 7.180 1592.420 7.440 ;
        RECT 1265.560 6.160 1265.820 6.420 ;
        RECT 1356.640 6.160 1356.900 6.420 ;
        RECT 1360.780 6.160 1361.040 6.420 ;
        RECT 1369.520 6.160 1369.780 6.420 ;
        RECT 1397.580 6.160 1397.840 6.420 ;
        RECT 1452.780 5.820 1453.040 6.080 ;
        RECT 1455.080 5.820 1455.340 6.080 ;
        RECT 1592.160 5.820 1592.420 6.080 ;
        RECT 1643.680 4.460 1643.940 4.720 ;
        RECT 540.140 3.780 540.400 4.040 ;
        RECT 1335.940 3.100 1336.200 3.360 ;
        RECT 1265.560 2.080 1265.820 2.340 ;
        RECT 1295.920 2.080 1296.180 2.340 ;
        RECT 1345.140 2.080 1345.400 2.340 ;
        RECT 1347.440 2.080 1347.700 2.340 ;
        RECT 1444.500 1.400 1444.760 1.660 ;
      LAYER met2 ;
        RECT 951.840 8.740 952.100 8.830 ;
        RECT 950.060 8.600 952.100 8.740 ;
        RECT 560.840 8.005 561.100 8.150 ;
        RECT 560.830 7.635 561.110 8.005 ;
        RECT 600.850 7.635 601.130 8.005 ;
        RECT 900.380 7.750 905.580 7.890 ;
        RECT 950.060 7.810 950.200 8.600 ;
        RECT 951.840 8.510 952.100 8.600 ;
        RECT 955.060 8.510 955.320 8.830 ;
        RECT 955.120 7.890 955.260 8.510 ;
        RECT 1000.660 8.260 1022.880 8.400 ;
        RECT 600.920 5.340 601.060 7.635 ;
        RECT 613.740 7.380 614.000 7.470 ;
        RECT 610.580 7.240 614.000 7.380 ;
        RECT 600.920 5.200 604.280 5.340 ;
        RECT 540.140 3.980 540.400 4.070 ;
        RECT 539.740 3.840 540.400 3.980 ;
        RECT 539.740 3.130 539.880 3.840 ;
        RECT 540.140 3.750 540.400 3.840 ;
        RECT 537.900 2.990 539.880 3.130 ;
        RECT 537.900 2.400 538.040 2.990 ;
        RECT 604.140 2.450 604.280 5.200 ;
        RECT 610.580 4.320 610.720 7.240 ;
        RECT 613.740 7.150 614.000 7.240 ;
        RECT 898.940 6.810 899.200 7.130 ;
        RECT 899.000 6.530 899.140 6.810 ;
        RECT 900.380 6.530 900.520 7.750 ;
        RECT 905.440 7.380 905.580 7.750 ;
        RECT 950.000 7.490 950.260 7.810 ;
        RECT 955.120 7.750 958.940 7.890 ;
        RECT 913.200 7.380 913.460 7.470 ;
        RECT 905.440 7.240 913.460 7.380 ;
        RECT 958.800 7.380 958.940 7.750 ;
        RECT 995.530 7.635 995.810 8.005 ;
        RECT 998.750 7.890 999.030 8.005 ;
        RECT 1000.660 7.890 1000.800 8.260 ;
        RECT 998.750 7.750 1000.800 7.890 ;
        RECT 998.750 7.635 999.030 7.750 ;
        RECT 995.540 7.490 995.800 7.635 ;
        RECT 1022.740 7.470 1022.880 8.260 ;
        RECT 1360.780 7.830 1361.040 8.150 ;
        RECT 1369.520 7.830 1369.780 8.150 ;
        RECT 959.200 7.380 959.460 7.470 ;
        RECT 958.800 7.240 959.460 7.380 ;
        RECT 913.200 7.150 913.460 7.240 ;
        RECT 959.200 7.150 959.460 7.240 ;
        RECT 1022.680 7.150 1022.940 7.470 ;
        RECT 1347.440 7.150 1347.700 7.470 ;
        RECT 1356.640 7.150 1356.900 7.470 ;
        RECT 1295.920 6.810 1296.180 7.130 ;
        RECT 899.000 6.390 900.520 6.530 ;
        RECT 1265.560 6.130 1265.820 6.450 ;
        RECT 606.440 4.180 610.720 4.320 ;
        RECT 606.440 2.450 606.580 4.180 ;
        RECT 537.690 -4.800 538.250 2.400 ;
        RECT 604.140 2.310 606.580 2.450 ;
        RECT 1265.620 2.370 1265.760 6.130 ;
        RECT 1295.980 2.370 1296.120 6.810 ;
        RECT 1335.940 3.070 1336.200 3.390 ;
        RECT 1336.000 2.450 1336.140 3.070 ;
        RECT 1336.920 2.990 1345.340 3.130 ;
        RECT 1336.920 2.450 1337.060 2.990 ;
        RECT 1265.560 2.050 1265.820 2.370 ;
        RECT 1295.920 2.050 1296.180 2.370 ;
        RECT 1336.000 2.310 1337.060 2.450 ;
        RECT 1345.200 2.370 1345.340 2.990 ;
        RECT 1347.500 2.370 1347.640 7.150 ;
        RECT 1356.700 6.450 1356.840 7.150 ;
        RECT 1360.840 6.450 1360.980 7.830 ;
        RECT 1369.580 6.450 1369.720 7.830 ;
        RECT 1397.580 7.150 1397.840 7.470 ;
        RECT 1446.800 7.210 1447.060 7.470 ;
        RECT 1444.560 7.150 1447.060 7.210 ;
        RECT 1592.160 7.150 1592.420 7.470 ;
        RECT 1397.640 6.450 1397.780 7.150 ;
        RECT 1444.560 7.070 1447.000 7.150 ;
        RECT 1356.640 6.130 1356.900 6.450 ;
        RECT 1360.780 6.130 1361.040 6.450 ;
        RECT 1369.520 6.130 1369.780 6.450 ;
        RECT 1397.580 6.130 1397.840 6.450 ;
        RECT 1345.140 2.050 1345.400 2.370 ;
        RECT 1347.440 2.050 1347.700 2.370 ;
        RECT 1444.560 1.690 1444.700 7.070 ;
        RECT 1592.220 6.110 1592.360 7.150 ;
        RECT 1452.780 5.790 1453.040 6.110 ;
        RECT 1455.080 5.790 1455.340 6.110 ;
        RECT 1592.160 5.790 1592.420 6.110 ;
        RECT 1452.840 4.490 1452.980 5.790 ;
        RECT 1455.140 4.490 1455.280 5.790 ;
        RECT 1643.610 5.000 1643.890 9.000 ;
        RECT 1643.740 4.750 1643.880 5.000 ;
        RECT 1452.840 4.350 1455.280 4.490 ;
        RECT 1643.680 4.430 1643.940 4.750 ;
        RECT 1444.500 1.370 1444.760 1.690 ;
      LAYER via2 ;
        RECT 560.830 7.680 561.110 7.960 ;
        RECT 600.850 7.680 601.130 7.960 ;
        RECT 995.530 7.680 995.810 7.960 ;
        RECT 998.750 7.680 999.030 7.960 ;
      LAYER met3 ;
        RECT 560.805 7.970 561.135 7.985 ;
        RECT 600.825 7.970 601.155 7.985 ;
        RECT 560.805 7.670 601.155 7.970 ;
        RECT 560.805 7.655 561.135 7.670 ;
        RECT 600.825 7.655 601.155 7.670 ;
        RECT 995.505 7.970 995.835 7.985 ;
        RECT 998.725 7.970 999.055 7.985 ;
        RECT 995.505 7.670 999.055 7.970 ;
        RECT 995.505 7.655 995.835 7.670 ;
        RECT 998.725 7.655 999.055 7.670 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 640.925 9.605 672.375 9.775 ;
        RECT 627.125 9.265 631.435 9.435 ;
        RECT 574.685 6.205 574.855 7.395 ;
        RECT 610.565 6.205 610.735 7.395 ;
        RECT 627.125 6.205 627.295 9.265 ;
        RECT 631.265 8.415 631.435 9.265 ;
        RECT 640.925 8.415 641.095 9.605 ;
        RECT 672.205 9.435 672.375 9.605 ;
        RECT 1452.365 9.605 1470.935 9.775 ;
        RECT 672.205 9.265 693.995 9.435 ;
        RECT 693.825 8.755 693.995 9.265 ;
        RECT 693.825 8.585 702.735 8.755 ;
        RECT 631.265 8.245 637.415 8.415 ;
        RECT 637.245 7.905 637.415 8.245 ;
        RECT 640.465 8.245 641.095 8.415 ;
        RECT 708.085 8.415 708.255 8.755 ;
        RECT 748.565 8.585 750.575 8.755 ;
        RECT 1452.365 8.585 1452.535 9.605 ;
        RECT 1470.765 9.095 1470.935 9.605 ;
        RECT 1470.765 8.925 1476.455 9.095 ;
        RECT 1476.285 8.585 1476.455 8.925 ;
        RECT 708.085 8.245 716.075 8.415 ;
        RECT 640.465 7.905 640.635 8.245 ;
        RECT 715.905 8.075 716.075 8.245 ;
        RECT 726.485 8.245 733.095 8.415 ;
        RECT 715.905 7.905 722.515 8.075 ;
        RECT 722.345 7.055 722.515 7.905 ;
        RECT 726.485 7.055 726.655 8.245 ;
        RECT 732.925 7.735 733.095 8.245 ;
        RECT 732.925 7.565 742.295 7.735 ;
        RECT 722.345 6.885 726.655 7.055 ;
        RECT 742.125 6.715 742.295 7.565 ;
        RECT 748.565 6.715 748.735 8.585 ;
        RECT 742.125 6.545 748.735 6.715 ;
        RECT 755.925 5.015 756.095 8.075 ;
        RECT 787.205 6.375 787.375 8.075 ;
        RECT 1327.245 7.225 1327.875 7.395 ;
        RECT 759.145 6.205 762.995 6.375 ;
        RECT 787.205 6.205 791.515 6.375 ;
        RECT 759.145 5.015 759.315 6.205 ;
        RECT 1327.705 5.695 1327.875 7.225 ;
        RECT 755.925 4.845 759.315 5.015 ;
        RECT 847.925 2.975 848.095 5.695 ;
        RECT 1327.705 5.525 1336.155 5.695 ;
        RECT 851.145 2.975 851.315 3.315 ;
        RECT 847.925 2.805 851.315 2.975 ;
        RECT 879.665 2.295 879.835 2.975 ;
        RECT 879.205 2.125 879.835 2.295 ;
        RECT 879.205 1.275 879.375 2.125 ;
        RECT 901.285 1.275 901.455 4.335 ;
        RECT 1335.985 3.315 1336.155 5.525 ;
        RECT 1428.905 3.485 1429.075 7.055 ;
        RECT 1335.985 3.145 1336.615 3.315 ;
        RECT 879.205 1.105 901.455 1.275 ;
      LAYER mcon ;
        RECT 574.685 7.225 574.855 7.395 ;
        RECT 610.565 7.225 610.735 7.395 ;
        RECT 702.565 8.585 702.735 8.755 ;
        RECT 708.085 8.585 708.255 8.755 ;
        RECT 750.405 8.585 750.575 8.755 ;
        RECT 755.925 7.905 756.095 8.075 ;
        RECT 787.205 7.905 787.375 8.075 ;
        RECT 762.825 6.205 762.995 6.375 ;
        RECT 791.345 6.205 791.515 6.375 ;
        RECT 1428.905 6.885 1429.075 7.055 ;
        RECT 847.925 5.525 848.095 5.695 ;
        RECT 901.285 4.165 901.455 4.335 ;
        RECT 851.145 3.145 851.315 3.315 ;
        RECT 879.665 2.805 879.835 2.975 ;
        RECT 1336.445 3.145 1336.615 3.315 ;
      LAYER met1 ;
        RECT 702.505 8.740 702.795 8.785 ;
        RECT 708.025 8.740 708.315 8.785 ;
        RECT 702.505 8.600 708.315 8.740 ;
        RECT 702.505 8.555 702.795 8.600 ;
        RECT 708.025 8.555 708.315 8.600 ;
        RECT 750.345 8.740 750.635 8.785 ;
        RECT 1451.370 8.740 1451.690 8.800 ;
        RECT 1452.305 8.740 1452.595 8.785 ;
        RECT 750.345 8.600 751.480 8.740 ;
        RECT 750.345 8.555 750.635 8.600 ;
        RECT 751.340 8.400 751.480 8.600 ;
        RECT 1451.370 8.600 1452.595 8.740 ;
        RECT 1451.370 8.540 1451.690 8.600 ;
        RECT 1452.305 8.555 1452.595 8.600 ;
        RECT 1476.225 8.740 1476.515 8.785 ;
        RECT 1689.190 8.740 1689.510 8.800 ;
        RECT 1476.225 8.600 1689.510 8.740 ;
        RECT 1476.225 8.555 1476.515 8.600 ;
        RECT 1689.190 8.540 1689.510 8.600 ;
        RECT 751.340 8.260 752.860 8.400 ;
        RECT 637.185 8.060 637.475 8.105 ;
        RECT 640.405 8.060 640.695 8.105 ;
        RECT 637.185 7.920 640.695 8.060 ;
        RECT 752.720 8.060 752.860 8.260 ;
        RECT 755.865 8.060 756.155 8.105 ;
        RECT 752.720 7.920 756.155 8.060 ;
        RECT 637.185 7.875 637.475 7.920 ;
        RECT 640.405 7.875 640.695 7.920 ;
        RECT 755.865 7.875 756.155 7.920 ;
        RECT 785.290 8.060 785.610 8.120 ;
        RECT 787.145 8.060 787.435 8.105 ;
        RECT 785.290 7.920 787.435 8.060 ;
        RECT 785.290 7.860 785.610 7.920 ;
        RECT 787.145 7.875 787.435 7.920 ;
        RECT 1160.190 8.060 1160.510 8.120 ;
        RECT 1162.490 8.060 1162.810 8.120 ;
        RECT 1160.190 7.920 1162.810 8.060 ;
        RECT 1160.190 7.860 1160.510 7.920 ;
        RECT 1162.490 7.860 1162.810 7.920 ;
        RECT 574.625 7.380 574.915 7.425 ;
        RECT 610.505 7.380 610.795 7.425 ;
        RECT 574.625 7.240 610.795 7.380 ;
        RECT 574.625 7.195 574.915 7.240 ;
        RECT 610.505 7.195 610.795 7.240 ;
        RECT 960.550 7.380 960.870 7.440 ;
        RECT 982.630 7.380 982.950 7.440 ;
        RECT 960.550 7.240 982.950 7.380 ;
        RECT 960.550 7.180 960.870 7.240 ;
        RECT 982.630 7.180 982.950 7.240 ;
        RECT 984.930 7.380 985.250 7.440 ;
        RECT 1001.030 7.380 1001.350 7.440 ;
        RECT 984.930 7.240 1001.350 7.380 ;
        RECT 984.930 7.180 985.250 7.240 ;
        RECT 1001.030 7.180 1001.350 7.240 ;
        RECT 1162.950 7.380 1163.270 7.440 ;
        RECT 1165.710 7.380 1166.030 7.440 ;
        RECT 1327.170 7.380 1327.490 7.440 ;
        RECT 1162.950 7.240 1166.030 7.380 ;
        RECT 1326.975 7.240 1327.490 7.380 ;
        RECT 1162.950 7.180 1163.270 7.240 ;
        RECT 1165.710 7.180 1166.030 7.240 ;
        RECT 1327.170 7.180 1327.490 7.240 ;
        RECT 1410.890 7.380 1411.210 7.440 ;
        RECT 1410.890 7.240 1426.300 7.380 ;
        RECT 1410.890 7.180 1411.210 7.240 ;
        RECT 1426.160 7.040 1426.300 7.240 ;
        RECT 1428.845 7.040 1429.135 7.085 ;
        RECT 1426.160 6.900 1429.135 7.040 ;
        RECT 1428.845 6.855 1429.135 6.900 ;
        RECT 559.430 6.360 559.750 6.420 ;
        RECT 574.625 6.360 574.915 6.405 ;
        RECT 559.430 6.220 574.915 6.360 ;
        RECT 559.430 6.160 559.750 6.220 ;
        RECT 574.625 6.175 574.915 6.220 ;
        RECT 610.505 6.360 610.795 6.405 ;
        RECT 627.065 6.360 627.355 6.405 ;
        RECT 610.505 6.220 627.355 6.360 ;
        RECT 610.505 6.175 610.795 6.220 ;
        RECT 627.065 6.175 627.355 6.220 ;
        RECT 762.765 6.360 763.055 6.405 ;
        RECT 763.210 6.360 763.530 6.420 ;
        RECT 762.765 6.220 763.530 6.360 ;
        RECT 762.765 6.175 763.055 6.220 ;
        RECT 763.210 6.160 763.530 6.220 ;
        RECT 791.285 6.360 791.575 6.405 ;
        RECT 793.110 6.360 793.430 6.420 ;
        RECT 791.285 6.220 793.430 6.360 ;
        RECT 791.285 6.175 791.575 6.220 ;
        RECT 793.110 6.160 793.430 6.220 ;
        RECT 1256.790 6.020 1257.110 6.080 ;
        RECT 1302.790 6.020 1303.110 6.080 ;
        RECT 1256.790 5.880 1303.110 6.020 ;
        RECT 1256.790 5.820 1257.110 5.880 ;
        RECT 1302.790 5.820 1303.110 5.880 ;
        RECT 845.090 5.680 845.410 5.740 ;
        RECT 847.865 5.680 848.155 5.725 ;
        RECT 845.090 5.540 848.155 5.680 ;
        RECT 845.090 5.480 845.410 5.540 ;
        RECT 847.865 5.495 848.155 5.540 ;
        RECT 901.225 4.320 901.515 4.365 ;
        RECT 903.050 4.320 903.370 4.380 ;
        RECT 901.225 4.180 903.370 4.320 ;
        RECT 901.225 4.135 901.515 4.180 ;
        RECT 903.050 4.120 903.370 4.180 ;
        RECT 879.590 3.640 879.910 3.700 ;
        RECT 851.160 3.500 879.910 3.640 ;
        RECT 851.160 3.345 851.300 3.500 ;
        RECT 879.590 3.440 879.910 3.500 ;
        RECT 1428.845 3.640 1429.135 3.685 ;
        RECT 1451.370 3.640 1451.690 3.700 ;
        RECT 1428.845 3.500 1451.690 3.640 ;
        RECT 1428.845 3.455 1429.135 3.500 ;
        RECT 1451.370 3.440 1451.690 3.500 ;
        RECT 851.085 3.115 851.375 3.345 ;
        RECT 1336.385 3.300 1336.675 3.345 ;
        RECT 1354.770 3.300 1355.090 3.360 ;
        RECT 1336.385 3.160 1355.090 3.300 ;
        RECT 1336.385 3.115 1336.675 3.160 ;
        RECT 1354.770 3.100 1355.090 3.160 ;
        RECT 1400.310 3.300 1400.630 3.360 ;
        RECT 1407.670 3.300 1407.990 3.360 ;
        RECT 1400.310 3.160 1407.990 3.300 ;
        RECT 1400.310 3.100 1400.630 3.160 ;
        RECT 1407.670 3.100 1407.990 3.160 ;
        RECT 879.590 2.960 879.910 3.020 ;
        RECT 879.395 2.820 879.910 2.960 ;
        RECT 879.590 2.760 879.910 2.820 ;
      LAYER via ;
        RECT 1451.400 8.540 1451.660 8.800 ;
        RECT 1689.220 8.540 1689.480 8.800 ;
        RECT 785.320 7.860 785.580 8.120 ;
        RECT 1160.220 7.860 1160.480 8.120 ;
        RECT 1162.520 7.860 1162.780 8.120 ;
        RECT 960.580 7.180 960.840 7.440 ;
        RECT 982.660 7.180 982.920 7.440 ;
        RECT 984.960 7.180 985.220 7.440 ;
        RECT 1001.060 7.180 1001.320 7.440 ;
        RECT 1162.980 7.180 1163.240 7.440 ;
        RECT 1165.740 7.180 1166.000 7.440 ;
        RECT 1327.200 7.180 1327.460 7.440 ;
        RECT 1410.920 7.180 1411.180 7.440 ;
        RECT 559.460 6.160 559.720 6.420 ;
        RECT 763.240 6.160 763.500 6.420 ;
        RECT 793.140 6.160 793.400 6.420 ;
        RECT 1256.820 5.820 1257.080 6.080 ;
        RECT 1302.820 5.820 1303.080 6.080 ;
        RECT 845.120 5.480 845.380 5.740 ;
        RECT 903.080 4.120 903.340 4.380 ;
        RECT 879.620 3.440 879.880 3.700 ;
        RECT 1451.400 3.440 1451.660 3.700 ;
        RECT 1354.800 3.100 1355.060 3.360 ;
        RECT 1400.340 3.100 1400.600 3.360 ;
        RECT 1407.700 3.100 1407.960 3.360 ;
        RECT 879.620 2.760 879.880 3.020 ;
      LAYER met2 ;
        RECT 1451.400 8.510 1451.660 8.830 ;
        RECT 1689.220 8.570 1689.480 8.830 ;
        RECT 1690.990 8.570 1691.270 9.000 ;
        RECT 1689.220 8.510 1691.270 8.570 ;
        RECT 1123.940 8.260 1129.140 8.400 ;
        RECT 785.320 7.830 785.580 8.150 ;
        RECT 810.220 7.920 820.020 8.060 ;
        RECT 763.300 7.580 765.280 7.720 ;
        RECT 763.300 6.450 763.440 7.580 ;
        RECT 765.140 7.380 765.280 7.580 ;
        RECT 770.200 7.580 784.140 7.720 ;
        RECT 770.200 7.380 770.340 7.580 ;
        RECT 765.140 7.240 770.340 7.380 ;
        RECT 784.000 7.380 784.140 7.580 ;
        RECT 785.380 7.380 785.520 7.830 ;
        RECT 784.000 7.240 785.520 7.380 ;
        RECT 559.460 6.130 559.720 6.450 ;
        RECT 763.240 6.130 763.500 6.450 ;
        RECT 793.140 6.130 793.400 6.450 ;
        RECT 797.730 6.275 798.010 6.645 ;
        RECT 809.230 6.530 809.510 6.645 ;
        RECT 810.220 6.530 810.360 7.920 ;
        RECT 819.880 7.210 820.020 7.920 ;
        RECT 1001.120 7.750 1001.720 7.890 ;
        RECT 1001.120 7.470 1001.260 7.750 ;
        RECT 1001.580 7.720 1001.720 7.750 ;
        RECT 1022.210 7.720 1022.490 8.005 ;
        RECT 1001.580 7.635 1022.490 7.720 ;
        RECT 1001.580 7.580 1022.420 7.635 ;
        RECT 821.190 7.210 821.470 7.325 ;
        RECT 819.880 7.070 821.470 7.210 ;
        RECT 821.190 6.955 821.470 7.070 ;
        RECT 845.110 6.955 845.390 7.325 ;
        RECT 960.580 7.150 960.840 7.470 ;
        RECT 982.660 7.150 982.920 7.470 ;
        RECT 984.960 7.380 985.220 7.470 ;
        RECT 984.100 7.240 985.220 7.380 ;
        RECT 809.230 6.390 810.360 6.530 ;
        RECT 809.230 6.275 809.510 6.390 ;
        RECT 559.520 4.660 559.660 6.130 ;
        RECT 793.200 5.965 793.340 6.130 ;
        RECT 793.130 5.595 793.410 5.965 ;
        RECT 796.350 5.595 796.630 5.965 ;
        RECT 796.420 5.340 796.560 5.595 ;
        RECT 797.800 5.340 797.940 6.275 ;
        RECT 845.180 5.770 845.320 6.955 ;
        RECT 903.140 6.220 904.660 6.360 ;
        RECT 845.120 5.450 845.380 5.770 ;
        RECT 796.420 5.200 797.940 5.340 ;
        RECT 555.840 4.520 559.660 4.660 ;
        RECT 555.840 2.400 555.980 4.520 ;
        RECT 903.140 4.410 903.280 6.220 ;
        RECT 903.080 4.090 903.340 4.410 ;
        RECT 904.520 4.320 904.660 6.220 ;
        RECT 917.860 4.350 921.680 4.490 ;
        RECT 917.860 4.320 918.000 4.350 ;
        RECT 904.520 4.180 918.000 4.320 ;
        RECT 921.540 3.810 921.680 4.350 ;
        RECT 960.640 3.980 960.780 7.150 ;
        RECT 982.720 5.170 982.860 7.150 ;
        RECT 984.100 5.170 984.240 7.240 ;
        RECT 984.960 7.150 985.220 7.240 ;
        RECT 1001.060 7.150 1001.320 7.470 ;
        RECT 1083.850 7.210 1084.130 7.325 ;
        RECT 1084.770 7.210 1085.050 7.325 ;
        RECT 1083.850 7.070 1085.050 7.210 ;
        RECT 1083.850 6.955 1084.130 7.070 ;
        RECT 1084.770 6.955 1085.050 7.070 ;
        RECT 1090.750 7.210 1091.030 7.325 ;
        RECT 1090.750 7.070 1091.880 7.210 ;
        RECT 1090.750 6.955 1091.030 7.070 ;
        RECT 1091.740 6.530 1091.880 7.070 ;
        RECT 1123.940 6.530 1124.080 8.260 ;
        RECT 1129.000 7.890 1129.140 8.260 ;
        RECT 1160.220 8.060 1160.480 8.150 ;
        RECT 1129.390 7.890 1129.670 8.005 ;
        RECT 1129.000 7.750 1129.670 7.890 ;
        RECT 1129.390 7.635 1129.670 7.750 ;
        RECT 1158.830 7.635 1159.110 8.005 ;
        RECT 1159.820 7.920 1160.480 8.060 ;
        RECT 1158.900 7.380 1159.040 7.635 ;
        RECT 1159.820 7.380 1159.960 7.920 ;
        RECT 1160.220 7.830 1160.480 7.920 ;
        RECT 1162.520 8.060 1162.780 8.150 ;
        RECT 1162.520 7.920 1163.180 8.060 ;
        RECT 1162.520 7.830 1162.780 7.920 ;
        RECT 1163.040 7.470 1163.180 7.920 ;
        RECT 1408.220 7.750 1411.120 7.890 ;
        RECT 1158.900 7.240 1159.960 7.380 ;
        RECT 1162.980 7.150 1163.240 7.470 ;
        RECT 1165.740 7.380 1166.000 7.470 ;
        RECT 1165.740 7.240 1166.400 7.380 ;
        RECT 1165.740 7.150 1166.000 7.240 ;
        RECT 1091.740 6.390 1107.980 6.530 ;
        RECT 982.720 5.030 984.240 5.170 ;
        RECT 921.930 3.810 922.210 3.925 ;
        RECT 879.620 3.410 879.880 3.730 ;
        RECT 921.540 3.670 922.210 3.810 ;
        RECT 921.930 3.555 922.210 3.670 ;
        RECT 957.880 3.840 960.780 3.980 ;
        RECT 1107.840 3.980 1107.980 6.390 ;
        RECT 1123.480 6.390 1124.080 6.530 ;
        RECT 1107.840 3.840 1121.780 3.980 ;
        RECT 957.880 3.640 958.020 3.840 ;
        RECT 956.500 3.500 958.020 3.640 ;
        RECT 879.680 3.050 879.820 3.410 ;
        RECT 879.620 2.730 879.880 3.050 ;
        RECT 956.500 2.565 956.640 3.500 ;
        RECT 1121.640 2.620 1121.780 3.840 ;
        RECT 1123.480 2.620 1123.620 6.390 ;
        RECT 1166.260 4.490 1166.400 7.240 ;
        RECT 1304.260 7.070 1307.160 7.210 ;
        RECT 1327.200 7.150 1327.460 7.470 ;
        RECT 1254.120 6.390 1257.020 6.530 ;
        RECT 1252.670 4.915 1252.950 5.285 ;
        RECT 1166.650 4.490 1166.930 4.605 ;
        RECT 1166.260 4.350 1166.930 4.490 ;
        RECT 1252.740 4.490 1252.880 4.915 ;
        RECT 1254.120 4.490 1254.260 6.390 ;
        RECT 1256.880 6.110 1257.020 6.390 ;
        RECT 1256.820 5.790 1257.080 6.110 ;
        RECT 1302.820 5.790 1303.080 6.110 ;
        RECT 1252.740 4.350 1254.260 4.490 ;
        RECT 1302.880 4.490 1303.020 5.790 ;
        RECT 1304.260 4.490 1304.400 7.070 ;
        RECT 1307.020 6.645 1307.160 7.070 ;
        RECT 1306.950 6.275 1307.230 6.645 ;
        RECT 1313.390 6.530 1313.670 6.645 ;
        RECT 1313.390 6.390 1314.060 6.530 ;
        RECT 1313.390 6.275 1313.670 6.390 ;
        RECT 1313.920 5.850 1314.060 6.390 ;
        RECT 1327.260 5.850 1327.400 7.150 ;
        RECT 1313.920 5.710 1325.560 5.850 ;
        RECT 1325.420 5.170 1325.560 5.710 ;
        RECT 1326.800 5.710 1327.400 5.850 ;
        RECT 1326.800 5.170 1326.940 5.710 ;
        RECT 1325.420 5.030 1326.940 5.170 ;
        RECT 1302.880 4.350 1304.400 4.490 ;
        RECT 1166.650 4.235 1166.930 4.350 ;
        RECT 1356.170 3.555 1356.450 3.925 ;
        RECT 1399.410 3.555 1399.690 3.925 ;
        RECT 1354.800 3.130 1355.060 3.390 ;
        RECT 1356.240 3.130 1356.380 3.555 ;
        RECT 1354.800 3.070 1356.380 3.130 ;
        RECT 1354.860 2.990 1356.380 3.070 ;
        RECT 1399.480 3.130 1399.620 3.555 ;
        RECT 1400.340 3.130 1400.600 3.390 ;
        RECT 1399.480 3.070 1400.600 3.130 ;
        RECT 1407.700 3.300 1407.960 3.390 ;
        RECT 1408.220 3.300 1408.360 7.750 ;
        RECT 1410.980 7.470 1411.120 7.750 ;
        RECT 1410.920 7.150 1411.180 7.470 ;
        RECT 1451.460 3.730 1451.600 8.510 ;
        RECT 1689.280 8.430 1691.270 8.510 ;
        RECT 1690.990 5.000 1691.270 8.430 ;
        RECT 1451.400 3.410 1451.660 3.730 ;
        RECT 1407.700 3.160 1408.360 3.300 ;
        RECT 1407.700 3.070 1407.960 3.160 ;
        RECT 1399.480 2.990 1400.540 3.070 ;
        RECT 555.630 -4.800 556.190 2.400 ;
        RECT 956.430 2.195 956.710 2.565 ;
        RECT 1121.640 2.480 1123.620 2.620 ;
      LAYER via2 ;
        RECT 797.730 6.320 798.010 6.600 ;
        RECT 809.230 6.320 809.510 6.600 ;
        RECT 1022.210 7.680 1022.490 7.960 ;
        RECT 821.190 7.000 821.470 7.280 ;
        RECT 845.110 7.000 845.390 7.280 ;
        RECT 793.130 5.640 793.410 5.920 ;
        RECT 796.350 5.640 796.630 5.920 ;
        RECT 1083.850 7.000 1084.130 7.280 ;
        RECT 1084.770 7.000 1085.050 7.280 ;
        RECT 1090.750 7.000 1091.030 7.280 ;
        RECT 1129.390 7.680 1129.670 7.960 ;
        RECT 1158.830 7.680 1159.110 7.960 ;
        RECT 921.930 3.600 922.210 3.880 ;
        RECT 1252.670 4.960 1252.950 5.240 ;
        RECT 1166.650 4.280 1166.930 4.560 ;
        RECT 1306.950 6.320 1307.230 6.600 ;
        RECT 1313.390 6.320 1313.670 6.600 ;
        RECT 1356.170 3.600 1356.450 3.880 ;
        RECT 1399.410 3.600 1399.690 3.880 ;
        RECT 956.430 2.240 956.710 2.520 ;
      LAYER met3 ;
        RECT 1022.185 7.970 1022.515 7.985 ;
        RECT 1023.310 7.970 1023.690 7.980 ;
        RECT 1022.185 7.670 1023.690 7.970 ;
        RECT 1022.185 7.655 1022.515 7.670 ;
        RECT 1023.310 7.660 1023.690 7.670 ;
        RECT 1129.365 7.970 1129.695 7.985 ;
        RECT 1158.805 7.970 1159.135 7.985 ;
        RECT 1129.365 7.670 1159.135 7.970 ;
        RECT 1129.365 7.655 1129.695 7.670 ;
        RECT 1158.805 7.655 1159.135 7.670 ;
        RECT 821.165 7.290 821.495 7.305 ;
        RECT 845.085 7.290 845.415 7.305 ;
        RECT 821.165 6.990 845.415 7.290 ;
        RECT 821.165 6.975 821.495 6.990 ;
        RECT 845.085 6.975 845.415 6.990 ;
        RECT 1041.710 7.290 1042.090 7.300 ;
        RECT 1049.070 7.290 1049.450 7.300 ;
        RECT 1083.825 7.290 1084.155 7.305 ;
        RECT 1041.710 6.990 1049.450 7.290 ;
        RECT 1041.710 6.980 1042.090 6.990 ;
        RECT 1049.070 6.980 1049.450 6.990 ;
        RECT 1073.030 6.990 1084.155 7.290 ;
        RECT 797.705 6.610 798.035 6.625 ;
        RECT 809.205 6.610 809.535 6.625 ;
        RECT 797.705 6.310 809.535 6.610 ;
        RECT 797.705 6.295 798.035 6.310 ;
        RECT 809.205 6.295 809.535 6.310 ;
        RECT 1049.990 6.610 1050.370 6.620 ;
        RECT 1073.030 6.610 1073.330 6.990 ;
        RECT 1083.825 6.975 1084.155 6.990 ;
        RECT 1084.745 7.290 1085.075 7.305 ;
        RECT 1090.725 7.290 1091.055 7.305 ;
        RECT 1084.745 6.990 1091.055 7.290 ;
        RECT 1084.745 6.975 1085.075 6.990 ;
        RECT 1090.725 6.975 1091.055 6.990 ;
        RECT 1049.990 6.310 1073.330 6.610 ;
        RECT 1306.925 6.610 1307.255 6.625 ;
        RECT 1313.365 6.610 1313.695 6.625 ;
        RECT 1306.925 6.310 1313.695 6.610 ;
        RECT 1049.990 6.300 1050.370 6.310 ;
        RECT 1306.925 6.295 1307.255 6.310 ;
        RECT 1313.365 6.295 1313.695 6.310 ;
        RECT 793.105 5.930 793.435 5.945 ;
        RECT 796.325 5.930 796.655 5.945 ;
        RECT 793.105 5.630 796.655 5.930 ;
        RECT 793.105 5.615 793.435 5.630 ;
        RECT 796.325 5.615 796.655 5.630 ;
        RECT 1239.510 5.250 1239.890 5.260 ;
        RECT 1252.645 5.250 1252.975 5.265 ;
        RECT 1239.510 4.950 1252.975 5.250 ;
        RECT 1239.510 4.940 1239.890 4.950 ;
        RECT 1252.645 4.935 1252.975 4.950 ;
        RECT 1166.625 4.580 1166.955 4.585 ;
        RECT 1166.625 4.570 1167.210 4.580 ;
        RECT 1166.400 4.270 1167.210 4.570 ;
        RECT 1166.625 4.260 1167.210 4.270 ;
        RECT 1166.625 4.255 1166.955 4.260 ;
        RECT 921.905 3.890 922.235 3.905 ;
        RECT 951.550 3.890 951.930 3.900 ;
        RECT 921.905 3.590 951.930 3.890 ;
        RECT 921.905 3.575 922.235 3.590 ;
        RECT 951.550 3.580 951.930 3.590 ;
        RECT 1225.710 3.890 1226.090 3.900 ;
        RECT 1232.150 3.890 1232.530 3.900 ;
        RECT 1225.710 3.590 1232.530 3.890 ;
        RECT 1225.710 3.580 1226.090 3.590 ;
        RECT 1232.150 3.580 1232.530 3.590 ;
        RECT 1356.145 3.890 1356.475 3.905 ;
        RECT 1399.385 3.890 1399.715 3.905 ;
        RECT 1356.145 3.590 1399.715 3.890 ;
        RECT 1356.145 3.575 1356.475 3.590 ;
        RECT 1399.385 3.575 1399.715 3.590 ;
        RECT 954.310 2.530 954.690 2.540 ;
        RECT 956.405 2.530 956.735 2.545 ;
        RECT 954.310 2.230 956.735 2.530 ;
        RECT 954.310 2.220 954.690 2.230 ;
        RECT 956.405 2.215 956.735 2.230 ;
      LAYER via3 ;
        RECT 1023.340 7.660 1023.660 7.980 ;
        RECT 1041.740 6.980 1042.060 7.300 ;
        RECT 1049.100 6.980 1049.420 7.300 ;
        RECT 1050.020 6.300 1050.340 6.620 ;
        RECT 1239.540 4.940 1239.860 5.260 ;
        RECT 1166.860 4.260 1167.180 4.580 ;
        RECT 951.580 3.580 951.900 3.900 ;
        RECT 1225.740 3.580 1226.060 3.900 ;
        RECT 1232.180 3.580 1232.500 3.900 ;
        RECT 954.340 2.220 954.660 2.540 ;
      LAYER met4 ;
        RECT 1023.350 8.350 1025.490 8.650 ;
        RECT 1023.350 7.985 1023.650 8.350 ;
        RECT 1023.335 7.655 1023.665 7.985 ;
        RECT 1025.190 7.290 1025.490 8.350 ;
        RECT 1041.735 7.290 1042.065 7.305 ;
        RECT 1025.190 6.990 1042.065 7.290 ;
        RECT 1041.735 6.975 1042.065 6.990 ;
        RECT 1049.095 7.290 1049.425 7.305 ;
        RECT 1049.095 6.990 1050.330 7.290 ;
        RECT 1049.095 6.975 1049.425 6.990 ;
        RECT 1050.030 6.625 1050.330 6.990 ;
        RECT 1050.015 6.295 1050.345 6.625 ;
        RECT 1234.030 5.630 1238.930 5.930 ;
        RECT 1166.855 4.255 1167.185 4.585 ;
        RECT 951.575 3.575 951.905 3.905 ;
        RECT 951.590 2.530 951.890 3.575 ;
        RECT 1166.870 3.210 1167.170 4.255 ;
        RECT 1225.735 3.575 1226.065 3.905 ;
        RECT 1232.175 3.575 1232.505 3.905 ;
        RECT 1166.870 2.910 1168.090 3.210 ;
        RECT 954.335 2.530 954.665 2.545 ;
        RECT 951.590 2.230 954.665 2.530 ;
        RECT 954.335 2.215 954.665 2.230 ;
        RECT 1167.790 1.850 1168.090 2.910 ;
        RECT 1225.750 1.850 1226.050 3.575 ;
        RECT 1232.190 3.210 1232.490 3.575 ;
        RECT 1234.030 3.210 1234.330 5.630 ;
        RECT 1238.630 5.250 1238.930 5.630 ;
        RECT 1239.535 5.250 1239.865 5.265 ;
        RECT 1238.630 4.950 1239.865 5.250 ;
        RECT 1239.535 4.935 1239.865 4.950 ;
        RECT 1232.190 2.910 1234.330 3.210 ;
        RECT 1167.790 1.550 1226.050 1.850 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1303.325 8.245 1307.175 8.415 ;
        RECT 1448.685 8.075 1448.855 8.755 ;
        RECT 682.785 7.905 685.255 8.075 ;
        RECT 1448.685 7.905 1452.535 8.075 ;
        RECT 789.505 7.565 792.435 7.735 ;
        RECT 640.005 6.545 641.095 6.715 ;
        RECT 640.005 6.205 640.175 6.545 ;
        RECT 792.265 6.375 792.435 7.565 ;
        RECT 792.265 6.205 793.815 6.375 ;
        RECT 1190.165 6.205 1191.255 6.375 ;
        RECT 1193.385 6.205 1194.935 6.375 ;
        RECT 844.705 5.865 848.555 6.035 ;
        RECT 829.525 5.525 835.215 5.695 ;
        RECT 844.705 5.525 844.875 5.865 ;
        RECT 848.385 5.525 848.555 5.865 ;
        RECT 1089.425 5.525 1090.975 5.695 ;
        RECT 815.725 3.995 815.895 4.675 ;
        RECT 821.705 4.505 822.795 4.675 ;
        RECT 822.625 4.165 822.795 4.505 ;
        RECT 829.525 4.165 829.695 5.525 ;
        RECT 1090.805 5.355 1090.975 5.525 ;
        RECT 1090.805 5.185 1108.455 5.355 ;
        RECT 805.605 3.825 806.235 3.995 ;
        RECT 815.265 3.825 815.895 3.995 ;
        RECT 1108.285 3.655 1108.455 5.185 ;
        RECT 1190.165 4.335 1190.335 6.205 ;
        RECT 1194.765 6.035 1194.935 6.205 ;
        RECT 1196.605 6.035 1196.775 6.375 ;
        RECT 1194.765 5.865 1196.775 6.035 ;
        RECT 1159.805 4.165 1190.335 4.335 ;
        RECT 1534.245 4.165 1534.415 5.015 ;
        RECT 1120.705 3.825 1121.335 3.995 ;
        RECT 1159.805 3.825 1159.975 4.165 ;
        RECT 1120.705 3.655 1120.875 3.825 ;
        RECT 1108.285 3.485 1120.875 3.655 ;
      LAYER mcon ;
        RECT 1448.685 8.585 1448.855 8.755 ;
        RECT 1307.005 8.245 1307.175 8.415 ;
        RECT 685.085 7.905 685.255 8.075 ;
        RECT 1452.365 7.905 1452.535 8.075 ;
        RECT 640.925 6.545 641.095 6.715 ;
        RECT 793.645 6.205 793.815 6.375 ;
        RECT 1191.085 6.205 1191.255 6.375 ;
        RECT 835.045 5.525 835.215 5.695 ;
        RECT 815.725 4.505 815.895 4.675 ;
        RECT 806.065 3.825 806.235 3.995 ;
        RECT 1196.605 6.205 1196.775 6.375 ;
        RECT 1534.245 4.845 1534.415 5.015 ;
        RECT 1121.165 3.825 1121.335 3.995 ;
      LAYER met1 ;
        RECT 1401.230 8.740 1401.550 8.800 ;
        RECT 1448.625 8.740 1448.915 8.785 ;
        RECT 1401.230 8.600 1448.915 8.740 ;
        RECT 1401.230 8.540 1401.550 8.600 ;
        RECT 1448.625 8.555 1448.915 8.600 ;
        RECT 750.790 8.400 751.110 8.460 ;
        RECT 704.880 8.260 751.110 8.400 ;
        RECT 644.070 8.060 644.390 8.120 ;
        RECT 682.725 8.060 683.015 8.105 ;
        RECT 644.070 7.920 683.015 8.060 ;
        RECT 644.070 7.860 644.390 7.920 ;
        RECT 682.725 7.875 683.015 7.920 ;
        RECT 685.025 8.060 685.315 8.105 ;
        RECT 704.880 8.060 705.020 8.260 ;
        RECT 750.790 8.200 751.110 8.260 ;
        RECT 753.090 8.400 753.410 8.460 ;
        RECT 1292.210 8.400 1292.530 8.460 ;
        RECT 1303.265 8.400 1303.555 8.445 ;
        RECT 753.090 8.260 787.820 8.400 ;
        RECT 753.090 8.200 753.410 8.260 ;
        RECT 685.025 7.920 705.020 8.060 ;
        RECT 685.025 7.875 685.315 7.920 ;
        RECT 787.680 7.720 787.820 8.260 ;
        RECT 1292.210 8.260 1303.555 8.400 ;
        RECT 1292.210 8.200 1292.530 8.260 ;
        RECT 1303.265 8.215 1303.555 8.260 ;
        RECT 1306.945 8.400 1307.235 8.445 ;
        RECT 1308.770 8.400 1309.090 8.460 ;
        RECT 1306.945 8.260 1309.090 8.400 ;
        RECT 1306.945 8.215 1307.235 8.260 ;
        RECT 1308.770 8.200 1309.090 8.260 ;
        RECT 1452.305 8.060 1452.595 8.105 ;
        RECT 1454.590 8.060 1454.910 8.120 ;
        RECT 1452.305 7.920 1454.910 8.060 ;
        RECT 1452.305 7.875 1452.595 7.920 ;
        RECT 1454.590 7.860 1454.910 7.920 ;
        RECT 789.445 7.720 789.735 7.765 ;
        RECT 787.680 7.580 789.735 7.720 ;
        RECT 789.445 7.535 789.735 7.580 ;
        RECT 640.865 6.700 641.155 6.745 ;
        RECT 643.150 6.700 643.470 6.760 ;
        RECT 640.865 6.560 643.470 6.700 ;
        RECT 640.865 6.515 641.155 6.560 ;
        RECT 643.150 6.500 643.470 6.560 ;
        RECT 630.730 6.360 631.050 6.420 ;
        RECT 639.945 6.360 640.235 6.405 ;
        RECT 630.730 6.220 640.235 6.360 ;
        RECT 630.730 6.160 631.050 6.220 ;
        RECT 639.945 6.175 640.235 6.220 ;
        RECT 793.585 6.360 793.875 6.405 ;
        RECT 794.030 6.360 794.350 6.420 ;
        RECT 793.585 6.220 794.350 6.360 ;
        RECT 793.585 6.175 793.875 6.220 ;
        RECT 794.030 6.160 794.350 6.220 ;
        RECT 1191.025 6.360 1191.315 6.405 ;
        RECT 1193.325 6.360 1193.615 6.405 ;
        RECT 1196.530 6.360 1196.850 6.420 ;
        RECT 1191.025 6.220 1193.615 6.360 ;
        RECT 1196.335 6.220 1196.850 6.360 ;
        RECT 1191.025 6.175 1191.315 6.220 ;
        RECT 1193.325 6.175 1193.615 6.220 ;
        RECT 1196.530 6.160 1196.850 6.220 ;
        RECT 579.670 5.680 579.990 5.740 ;
        RECT 614.170 5.680 614.490 5.740 ;
        RECT 579.670 5.540 614.490 5.680 ;
        RECT 579.670 5.480 579.990 5.540 ;
        RECT 614.170 5.480 614.490 5.540 ;
        RECT 834.985 5.680 835.275 5.725 ;
        RECT 844.645 5.680 844.935 5.725 ;
        RECT 834.985 5.540 844.935 5.680 ;
        RECT 834.985 5.495 835.275 5.540 ;
        RECT 844.645 5.495 844.935 5.540 ;
        RECT 848.325 5.680 848.615 5.725 ;
        RECT 1089.365 5.680 1089.655 5.725 ;
        RECT 848.325 5.540 1089.655 5.680 ;
        RECT 848.325 5.495 848.615 5.540 ;
        RECT 1089.365 5.495 1089.655 5.540 ;
        RECT 1227.810 5.340 1228.130 5.400 ;
        RECT 1235.630 5.340 1235.950 5.400 ;
        RECT 1227.810 5.200 1235.950 5.340 ;
        RECT 1227.810 5.140 1228.130 5.200 ;
        RECT 1235.630 5.140 1235.950 5.200 ;
        RECT 1484.490 5.000 1484.810 5.060 ;
        RECT 1534.185 5.000 1534.475 5.045 ;
        RECT 1484.490 4.860 1534.475 5.000 ;
        RECT 1484.490 4.800 1484.810 4.860 ;
        RECT 1534.185 4.815 1534.475 4.860 ;
        RECT 815.665 4.660 815.955 4.705 ;
        RECT 821.645 4.660 821.935 4.705 ;
        RECT 815.665 4.520 821.935 4.660 ;
        RECT 815.665 4.475 815.955 4.520 ;
        RECT 821.645 4.475 821.935 4.520 ;
        RECT 822.565 4.320 822.855 4.365 ;
        RECT 829.465 4.320 829.755 4.365 ;
        RECT 822.565 4.180 829.755 4.320 ;
        RECT 822.565 4.135 822.855 4.180 ;
        RECT 829.465 4.135 829.755 4.180 ;
        RECT 1534.185 4.320 1534.475 4.365 ;
        RECT 1549.810 4.320 1550.130 4.380 ;
        RECT 1534.185 4.180 1550.130 4.320 ;
        RECT 1534.185 4.135 1534.475 4.180 ;
        RECT 1549.810 4.120 1550.130 4.180 ;
        RECT 804.150 3.980 804.470 4.040 ;
        RECT 805.545 3.980 805.835 4.025 ;
        RECT 804.150 3.840 805.835 3.980 ;
        RECT 804.150 3.780 804.470 3.840 ;
        RECT 805.545 3.795 805.835 3.840 ;
        RECT 806.005 3.980 806.295 4.025 ;
        RECT 815.205 3.980 815.495 4.025 ;
        RECT 806.005 3.840 815.495 3.980 ;
        RECT 806.005 3.795 806.295 3.840 ;
        RECT 815.205 3.795 815.495 3.840 ;
        RECT 1121.105 3.980 1121.395 4.025 ;
        RECT 1159.745 3.980 1160.035 4.025 ;
        RECT 1121.105 3.840 1160.035 3.980 ;
        RECT 1121.105 3.795 1121.395 3.840 ;
        RECT 1159.745 3.795 1160.035 3.840 ;
      LAYER via ;
        RECT 1401.260 8.540 1401.520 8.800 ;
        RECT 644.100 7.860 644.360 8.120 ;
        RECT 750.820 8.200 751.080 8.460 ;
        RECT 753.120 8.200 753.380 8.460 ;
        RECT 1292.240 8.200 1292.500 8.460 ;
        RECT 1308.800 8.200 1309.060 8.460 ;
        RECT 1454.620 7.860 1454.880 8.120 ;
        RECT 643.180 6.500 643.440 6.760 ;
        RECT 630.760 6.160 631.020 6.420 ;
        RECT 794.060 6.160 794.320 6.420 ;
        RECT 1196.560 6.160 1196.820 6.420 ;
        RECT 579.700 5.480 579.960 5.740 ;
        RECT 614.200 5.480 614.460 5.740 ;
        RECT 1227.840 5.140 1228.100 5.400 ;
        RECT 1235.660 5.140 1235.920 5.400 ;
        RECT 1484.520 4.800 1484.780 5.060 ;
        RECT 1549.840 4.120 1550.100 4.380 ;
        RECT 804.180 3.780 804.440 4.040 ;
      LAYER met2 ;
        RECT 1401.260 8.740 1401.520 8.830 ;
        RECT 1238.940 8.685 1250.580 8.740 ;
        RECT 1238.940 8.600 1250.650 8.685 ;
        RECT 750.820 8.400 751.080 8.490 ;
        RECT 753.120 8.400 753.380 8.490 ;
        RECT 750.820 8.260 753.380 8.400 ;
        RECT 750.820 8.170 751.080 8.260 ;
        RECT 753.120 8.170 753.380 8.260 ;
        RECT 644.100 8.060 644.360 8.150 ;
        RECT 643.240 7.920 644.360 8.060 ;
        RECT 577.920 7.070 579.900 7.210 ;
        RECT 577.920 3.130 578.060 7.070 ;
        RECT 579.760 5.770 579.900 7.070 ;
        RECT 643.240 6.790 643.380 7.920 ;
        RECT 644.100 7.830 644.360 7.920 ;
        RECT 1238.940 7.890 1239.080 8.600 ;
        RECT 1250.370 8.315 1250.650 8.600 ;
        RECT 1290.390 8.400 1290.670 8.685 ;
        RECT 1292.240 8.400 1292.500 8.490 ;
        RECT 1290.390 8.315 1292.500 8.400 ;
        RECT 1290.460 8.260 1292.500 8.315 ;
        RECT 1292.240 8.170 1292.500 8.260 ;
        RECT 1308.800 8.400 1309.060 8.490 ;
        RECT 1310.170 8.400 1310.450 8.685 ;
        RECT 1344.210 8.570 1344.490 8.685 ;
        RECT 1308.800 8.315 1310.450 8.400 ;
        RECT 1343.360 8.430 1344.490 8.570 ;
        RECT 1308.800 8.260 1310.380 8.315 ;
        RECT 1308.800 8.170 1309.060 8.260 ;
        RECT 1235.720 7.750 1239.080 7.890 ;
        RECT 1341.910 7.890 1342.190 8.005 ;
        RECT 1343.360 7.890 1343.500 8.430 ;
        RECT 1344.210 8.315 1344.490 8.430 ;
        RECT 1400.860 8.600 1401.520 8.740 ;
        RECT 1400.860 8.005 1401.000 8.600 ;
        RECT 1401.260 8.510 1401.520 8.600 ;
        RECT 1454.680 8.430 1455.740 8.570 ;
        RECT 1454.680 8.150 1454.820 8.430 ;
        RECT 1341.910 7.750 1343.500 7.890 ;
        RECT 1398.950 7.890 1399.230 8.005 ;
        RECT 1399.870 7.890 1400.150 8.005 ;
        RECT 1398.950 7.750 1400.150 7.890 ;
        RECT 643.180 6.470 643.440 6.790 ;
        RECT 630.760 6.360 631.020 6.450 ;
        RECT 614.260 6.220 631.020 6.360 ;
        RECT 614.260 5.770 614.400 6.220 ;
        RECT 630.760 6.130 631.020 6.220 ;
        RECT 794.060 6.130 794.320 6.450 ;
        RECT 1196.560 6.130 1196.820 6.450 ;
        RECT 579.700 5.450 579.960 5.770 ;
        RECT 614.200 5.450 614.460 5.770 ;
        RECT 794.120 3.640 794.260 6.130 ;
        RECT 796.880 4.350 804.380 4.490 ;
        RECT 796.880 3.640 797.020 4.350 ;
        RECT 804.240 4.070 804.380 4.350 ;
        RECT 804.180 3.750 804.440 4.070 ;
        RECT 1196.620 3.925 1196.760 6.130 ;
        RECT 1235.720 5.430 1235.860 7.750 ;
        RECT 1341.910 7.635 1342.190 7.750 ;
        RECT 1398.950 7.635 1399.230 7.750 ;
        RECT 1399.870 7.635 1400.150 7.750 ;
        RECT 1400.790 7.635 1401.070 8.005 ;
        RECT 1454.620 7.830 1454.880 8.150 ;
        RECT 1227.840 5.340 1228.100 5.430 ;
        RECT 1227.440 5.200 1228.100 5.340 ;
        RECT 1227.440 3.980 1227.580 5.200 ;
        RECT 1227.840 5.110 1228.100 5.200 ;
        RECT 1235.660 5.110 1235.920 5.430 ;
        RECT 1455.600 5.170 1455.740 8.430 ;
        RECT 1609.630 8.315 1609.910 8.685 ;
        RECT 1737.050 8.570 1737.330 8.685 ;
        RECT 1738.370 8.570 1738.650 9.000 ;
        RECT 1737.050 8.430 1738.650 8.570 ;
        RECT 1737.050 8.315 1737.330 8.430 ;
        RECT 1609.700 5.965 1609.840 8.315 ;
        RECT 1549.830 5.595 1550.110 5.965 ;
        RECT 1609.630 5.595 1609.910 5.965 ;
        RECT 1469.330 5.170 1469.610 5.285 ;
        RECT 1455.600 5.030 1469.610 5.170 ;
        RECT 1469.330 4.915 1469.610 5.030 ;
        RECT 1484.510 4.915 1484.790 5.285 ;
        RECT 1484.520 4.770 1484.780 4.915 ;
        RECT 1549.900 4.410 1550.040 5.595 ;
        RECT 1738.370 5.000 1738.650 8.430 ;
        RECT 1549.840 4.090 1550.100 4.410 ;
        RECT 1225.140 3.925 1227.580 3.980 ;
        RECT 794.120 3.500 797.020 3.640 ;
        RECT 1196.550 3.555 1196.830 3.925 ;
        RECT 1225.070 3.840 1227.580 3.925 ;
        RECT 1225.070 3.555 1225.350 3.840 ;
        RECT 573.780 2.990 578.060 3.130 ;
        RECT 573.780 2.400 573.920 2.990 ;
        RECT 573.570 -4.800 574.130 2.400 ;
      LAYER via2 ;
        RECT 1250.370 8.360 1250.650 8.640 ;
        RECT 1290.390 8.360 1290.670 8.640 ;
        RECT 1310.170 8.360 1310.450 8.640 ;
        RECT 1341.910 7.680 1342.190 7.960 ;
        RECT 1344.210 8.360 1344.490 8.640 ;
        RECT 1398.950 7.680 1399.230 7.960 ;
        RECT 1399.870 7.680 1400.150 7.960 ;
        RECT 1400.790 7.680 1401.070 7.960 ;
        RECT 1609.630 8.360 1609.910 8.640 ;
        RECT 1737.050 8.360 1737.330 8.640 ;
        RECT 1549.830 5.640 1550.110 5.920 ;
        RECT 1609.630 5.640 1609.910 5.920 ;
        RECT 1469.330 4.960 1469.610 5.240 ;
        RECT 1484.510 4.960 1484.790 5.240 ;
        RECT 1196.550 3.600 1196.830 3.880 ;
        RECT 1225.070 3.600 1225.350 3.880 ;
      LAYER met3 ;
        RECT 1250.345 8.650 1250.675 8.665 ;
        RECT 1290.365 8.650 1290.695 8.665 ;
        RECT 1250.345 8.350 1290.695 8.650 ;
        RECT 1250.345 8.335 1250.675 8.350 ;
        RECT 1290.365 8.335 1290.695 8.350 ;
        RECT 1310.145 8.650 1310.475 8.665 ;
        RECT 1344.185 8.650 1344.515 8.665 ;
        RECT 1609.605 8.650 1609.935 8.665 ;
        RECT 1737.025 8.650 1737.355 8.665 ;
        RECT 1310.145 8.350 1341.970 8.650 ;
        RECT 1310.145 8.335 1310.475 8.350 ;
        RECT 1341.670 7.985 1341.970 8.350 ;
        RECT 1344.185 8.350 1360.370 8.650 ;
        RECT 1344.185 8.335 1344.515 8.350 ;
        RECT 1341.670 7.670 1342.215 7.985 ;
        RECT 1360.070 7.970 1360.370 8.350 ;
        RECT 1609.605 8.350 1737.355 8.650 ;
        RECT 1609.605 8.335 1609.935 8.350 ;
        RECT 1737.025 8.335 1737.355 8.350 ;
        RECT 1398.925 7.970 1399.255 7.985 ;
        RECT 1360.070 7.670 1399.255 7.970 ;
        RECT 1341.885 7.655 1342.215 7.670 ;
        RECT 1398.925 7.655 1399.255 7.670 ;
        RECT 1399.845 7.970 1400.175 7.985 ;
        RECT 1400.765 7.970 1401.095 7.985 ;
        RECT 1399.845 7.670 1401.095 7.970 ;
        RECT 1399.845 7.655 1400.175 7.670 ;
        RECT 1400.765 7.655 1401.095 7.670 ;
        RECT 1549.805 5.930 1550.135 5.945 ;
        RECT 1609.605 5.930 1609.935 5.945 ;
        RECT 1549.805 5.630 1609.935 5.930 ;
        RECT 1549.805 5.615 1550.135 5.630 ;
        RECT 1609.605 5.615 1609.935 5.630 ;
        RECT 1469.305 5.250 1469.635 5.265 ;
        RECT 1484.485 5.250 1484.815 5.265 ;
        RECT 1469.305 4.950 1484.815 5.250 ;
        RECT 1469.305 4.935 1469.635 4.950 ;
        RECT 1484.485 4.935 1484.815 4.950 ;
        RECT 1196.525 3.890 1196.855 3.905 ;
        RECT 1225.045 3.890 1225.375 3.905 ;
        RECT 1196.525 3.590 1225.375 3.890 ;
        RECT 1196.525 3.575 1196.855 3.590 ;
        RECT 1225.045 3.575 1225.375 3.590 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 793.645 8.925 805.775 9.095 ;
        RECT 786.285 8.245 787.835 8.415 ;
        RECT 712.225 6.205 714.695 6.375 ;
        RECT 766.965 6.205 768.055 6.375 ;
        RECT 772.945 6.205 774.495 6.375 ;
        RECT 698.425 5.525 703.655 5.695 ;
        RECT 603.665 0.935 603.835 3.995 ;
        RECT 698.425 2.975 698.595 5.525 ;
        RECT 711.305 5.355 711.475 5.695 ;
        RECT 712.225 5.355 712.395 6.205 ;
        RECT 766.965 6.035 767.135 6.205 ;
        RECT 711.305 5.185 712.395 5.355 ;
        RECT 766.045 5.865 767.135 6.035 ;
        RECT 766.045 3.825 766.215 5.865 ;
        RECT 648.285 2.805 698.595 2.975 ;
        RECT 774.325 2.975 774.495 6.205 ;
        RECT 786.285 2.975 786.455 8.245 ;
        RECT 787.665 8.075 787.835 8.245 ;
        RECT 787.665 7.905 788.295 8.075 ;
        RECT 793.645 7.905 793.815 8.925 ;
        RECT 805.605 7.905 805.775 8.925 ;
        RECT 983.165 8.925 985.175 9.095 ;
        RECT 893.005 8.585 894.555 8.755 ;
        RECT 893.005 8.245 893.175 8.585 ;
        RECT 983.165 8.245 983.335 8.925 ;
        RECT 985.005 8.245 985.175 8.925 ;
        RECT 1120.245 8.585 1123.635 8.755 ;
        RECT 1120.245 8.245 1120.415 8.585 ;
        RECT 1123.465 8.245 1123.635 8.585 ;
        RECT 1158.885 8.245 1159.515 8.415 ;
        RECT 1159.345 5.355 1159.515 8.245 ;
        RECT 1166.705 5.355 1166.875 8.415 ;
        RECT 1291.365 8.075 1291.535 8.415 ;
        RECT 1292.745 8.075 1292.915 9.095 ;
        RECT 1312.525 8.585 1313.155 8.755 ;
        RECT 1312.985 8.415 1313.155 8.585 ;
        RECT 1312.985 8.245 1314.535 8.415 ;
        RECT 1291.365 7.905 1292.915 8.075 ;
        RECT 1159.345 5.185 1166.875 5.355 ;
        RECT 1598.645 3.655 1598.815 7.055 ;
        RECT 1596.805 3.485 1598.815 3.655 ;
        RECT 1596.805 3.145 1596.975 3.485 ;
        RECT 774.325 2.805 786.455 2.975 ;
        RECT 648.285 0.935 648.455 2.805 ;
        RECT 603.665 0.765 648.455 0.935 ;
      LAYER mcon ;
        RECT 714.525 6.205 714.695 6.375 ;
        RECT 767.885 6.205 768.055 6.375 ;
        RECT 703.485 5.525 703.655 5.695 ;
        RECT 711.305 5.525 711.475 5.695 ;
        RECT 603.665 3.825 603.835 3.995 ;
        RECT 788.125 7.905 788.295 8.075 ;
        RECT 894.385 8.585 894.555 8.755 ;
        RECT 1292.745 8.925 1292.915 9.095 ;
        RECT 1166.705 8.245 1166.875 8.415 ;
        RECT 1291.365 8.245 1291.535 8.415 ;
        RECT 1314.365 8.245 1314.535 8.415 ;
        RECT 1598.645 6.885 1598.815 7.055 ;
      LAYER met1 ;
        RECT 1292.685 9.080 1292.975 9.125 ;
        RECT 1292.685 8.940 1309.920 9.080 ;
        RECT 1292.685 8.895 1292.975 8.940 ;
        RECT 894.325 8.740 894.615 8.785 ;
        RECT 894.325 8.600 896.840 8.740 ;
        RECT 894.325 8.555 894.615 8.600 ;
        RECT 896.700 8.460 896.840 8.600 ;
        RECT 892.945 8.400 893.235 8.445 ;
        RECT 848.400 8.260 893.235 8.400 ;
        RECT 788.065 8.060 788.355 8.105 ;
        RECT 793.585 8.060 793.875 8.105 ;
        RECT 788.065 7.920 793.875 8.060 ;
        RECT 788.065 7.875 788.355 7.920 ;
        RECT 793.585 7.875 793.875 7.920 ;
        RECT 805.545 8.060 805.835 8.105 ;
        RECT 848.400 8.060 848.540 8.260 ;
        RECT 892.945 8.215 893.235 8.260 ;
        RECT 896.610 8.200 896.930 8.460 ;
        RECT 897.530 8.400 897.850 8.460 ;
        RECT 983.105 8.400 983.395 8.445 ;
        RECT 897.530 8.260 983.395 8.400 ;
        RECT 897.530 8.200 897.850 8.260 ;
        RECT 983.105 8.215 983.395 8.260 ;
        RECT 984.945 8.400 985.235 8.445 ;
        RECT 1120.185 8.400 1120.475 8.445 ;
        RECT 984.945 8.260 1083.600 8.400 ;
        RECT 984.945 8.215 985.235 8.260 ;
        RECT 805.545 7.920 848.540 8.060 ;
        RECT 1083.460 8.060 1083.600 8.260 ;
        RECT 1101.400 8.260 1120.475 8.400 ;
        RECT 1101.400 8.060 1101.540 8.260 ;
        RECT 1120.185 8.215 1120.475 8.260 ;
        RECT 1123.405 8.400 1123.695 8.445 ;
        RECT 1158.825 8.400 1159.115 8.445 ;
        RECT 1123.405 8.260 1159.115 8.400 ;
        RECT 1123.405 8.215 1123.695 8.260 ;
        RECT 1158.825 8.215 1159.115 8.260 ;
        RECT 1166.645 8.400 1166.935 8.445 ;
        RECT 1291.305 8.400 1291.595 8.445 ;
        RECT 1166.645 8.260 1291.595 8.400 ;
        RECT 1309.780 8.400 1309.920 8.940 ;
        RECT 1312.465 8.555 1312.755 8.785 ;
        RECT 1312.540 8.400 1312.680 8.555 ;
        RECT 1309.780 8.260 1312.680 8.400 ;
        RECT 1314.305 8.400 1314.595 8.445 ;
        RECT 1484.030 8.400 1484.350 8.460 ;
        RECT 1314.305 8.260 1484.350 8.400 ;
        RECT 1166.645 8.215 1166.935 8.260 ;
        RECT 1291.305 8.215 1291.595 8.260 ;
        RECT 1314.305 8.215 1314.595 8.260 ;
        RECT 1484.030 8.200 1484.350 8.260 ;
        RECT 1083.460 7.920 1101.540 8.060 ;
        RECT 805.545 7.875 805.835 7.920 ;
        RECT 1598.585 7.040 1598.875 7.085 ;
        RECT 1783.950 7.040 1784.270 7.100 ;
        RECT 1598.585 6.900 1784.270 7.040 ;
        RECT 1598.585 6.855 1598.875 6.900 ;
        RECT 1783.950 6.840 1784.270 6.900 ;
        RECT 751.800 6.560 759.300 6.700 ;
        RECT 714.465 6.360 714.755 6.405 ;
        RECT 751.800 6.360 751.940 6.560 ;
        RECT 714.465 6.220 751.940 6.360 ;
        RECT 759.160 6.360 759.300 6.560 ;
        RECT 760.450 6.360 760.770 6.420 ;
        RECT 759.160 6.220 760.770 6.360 ;
        RECT 714.465 6.175 714.755 6.220 ;
        RECT 760.450 6.160 760.770 6.220 ;
        RECT 767.825 6.360 768.115 6.405 ;
        RECT 772.885 6.360 773.175 6.405 ;
        RECT 767.825 6.220 773.175 6.360 ;
        RECT 767.825 6.175 768.115 6.220 ;
        RECT 772.885 6.175 773.175 6.220 ;
        RECT 703.425 5.680 703.715 5.725 ;
        RECT 711.245 5.680 711.535 5.725 ;
        RECT 703.425 5.540 711.535 5.680 ;
        RECT 703.425 5.495 703.715 5.540 ;
        RECT 711.245 5.495 711.535 5.540 ;
        RECT 603.590 3.980 603.910 4.040 ;
        RECT 603.395 3.840 603.910 3.980 ;
        RECT 603.590 3.780 603.910 3.840 ;
        RECT 760.450 3.980 760.770 4.040 ;
        RECT 765.985 3.980 766.275 4.025 ;
        RECT 760.450 3.840 766.275 3.980 ;
        RECT 760.450 3.780 760.770 3.840 ;
        RECT 765.985 3.795 766.275 3.840 ;
        RECT 1503.810 3.300 1504.130 3.360 ;
        RECT 1596.745 3.300 1597.035 3.345 ;
        RECT 1503.810 3.160 1597.035 3.300 ;
        RECT 1503.810 3.100 1504.130 3.160 ;
        RECT 1596.745 3.115 1597.035 3.160 ;
      LAYER via ;
        RECT 896.640 8.200 896.900 8.460 ;
        RECT 897.560 8.200 897.820 8.460 ;
        RECT 1484.060 8.200 1484.320 8.460 ;
        RECT 1783.980 6.840 1784.240 7.100 ;
        RECT 760.480 6.160 760.740 6.420 ;
        RECT 603.620 3.780 603.880 4.040 ;
        RECT 760.480 3.780 760.740 4.040 ;
        RECT 1503.840 3.100 1504.100 3.360 ;
      LAYER met2 ;
        RECT 1484.120 8.490 1493.460 8.570 ;
        RECT 896.640 8.400 896.900 8.490 ;
        RECT 897.560 8.400 897.820 8.490 ;
        RECT 896.640 8.260 897.820 8.400 ;
        RECT 896.640 8.170 896.900 8.260 ;
        RECT 897.560 8.170 897.820 8.260 ;
        RECT 1484.060 8.430 1493.460 8.490 ;
        RECT 1484.060 8.170 1484.320 8.430 ;
        RECT 760.480 6.130 760.740 6.450 ;
        RECT 591.260 4.350 603.820 4.490 ;
        RECT 591.260 2.400 591.400 4.350 ;
        RECT 603.680 4.070 603.820 4.350 ;
        RECT 760.540 4.070 760.680 6.130 ;
        RECT 1493.320 4.490 1493.460 8.430 ;
        RECT 1785.750 7.210 1786.030 9.000 ;
        RECT 1784.040 7.130 1786.030 7.210 ;
        RECT 1783.980 7.070 1786.030 7.130 ;
        RECT 1783.980 6.810 1784.240 7.070 ;
        RECT 1785.750 5.000 1786.030 7.070 ;
        RECT 1493.320 4.350 1502.660 4.490 ;
        RECT 603.620 3.750 603.880 4.070 ;
        RECT 760.480 3.750 760.740 4.070 ;
        RECT 1502.520 2.450 1502.660 4.350 ;
        RECT 1503.840 3.070 1504.100 3.390 ;
        RECT 1503.900 2.450 1504.040 3.070 ;
        RECT 591.050 -4.800 591.610 2.400 ;
        RECT 1502.520 2.310 1504.040 2.450 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1304.705 10.285 1307.175 10.455 ;
        RECT 1304.705 9.775 1304.875 10.285 ;
        RECT 1293.205 9.605 1304.875 9.775 ;
        RECT 1293.205 9.435 1293.375 9.605 ;
        RECT 898.985 9.265 904.215 9.435 ;
        RECT 706.705 7.905 715.615 8.075 ;
        RECT 674.505 6.885 679.735 7.055 ;
        RECT 693.365 6.885 705.035 7.055 ;
        RECT 674.505 6.375 674.675 6.885 ;
        RECT 673.585 6.205 674.675 6.375 ;
        RECT 704.865 3.995 705.035 6.885 ;
        RECT 706.705 3.995 706.875 7.905 ;
        RECT 715.445 7.735 715.615 7.905 ;
        RECT 715.445 7.565 719.295 7.735 ;
        RECT 719.125 7.055 719.295 7.565 ;
        RECT 719.125 6.885 720.215 7.055 ;
        RECT 720.045 5.695 720.215 6.885 ;
        RECT 836.425 6.205 850.395 6.375 ;
        RECT 720.045 5.525 739.075 5.695 ;
        RECT 738.905 5.185 739.075 5.525 ;
        RECT 704.865 3.825 706.875 3.995 ;
        RECT 835.505 2.975 835.675 3.315 ;
        RECT 836.425 2.975 836.595 6.205 ;
        RECT 879.205 6.035 879.375 6.375 ;
        RECT 879.205 5.865 891.335 6.035 ;
        RECT 891.165 3.995 891.335 5.865 ;
        RECT 898.985 3.995 899.155 9.265 ;
        RECT 904.045 7.225 904.215 9.265 ;
        RECT 1292.285 9.265 1293.375 9.435 ;
        RECT 1169.465 8.925 1183.895 9.095 ;
        RECT 1292.285 8.925 1292.455 9.265 ;
        RECT 1307.005 9.095 1307.175 10.285 ;
        RECT 1307.005 8.925 1310.395 9.095 ;
        RECT 1343.805 8.925 1344.895 9.095 ;
        RECT 912.785 5.355 912.955 7.395 ;
        RECT 955.105 6.375 955.275 6.715 ;
        RECT 955.105 6.205 955.735 6.375 ;
        RECT 912.785 5.185 945.615 5.355 ;
        RECT 945.445 4.675 945.615 5.185 ;
        RECT 955.565 4.675 955.735 6.205 ;
        RECT 1126.225 5.865 1128.235 6.035 ;
        RECT 945.445 4.505 955.735 4.675 ;
        RECT 1123.005 5.525 1125.475 5.695 ;
        RECT 1123.005 3.995 1123.175 5.525 ;
        RECT 1125.305 5.355 1125.475 5.525 ;
        RECT 1126.225 5.355 1126.395 5.865 ;
        RECT 1128.065 5.525 1128.235 5.865 ;
        RECT 1125.305 5.185 1126.395 5.355 ;
        RECT 891.165 3.825 899.155 3.995 ;
        RECT 1121.625 3.825 1123.175 3.995 ;
        RECT 1158.425 3.995 1158.595 5.695 ;
        RECT 1169.465 4.675 1169.635 8.925 ;
        RECT 1343.805 8.585 1343.975 8.925 ;
        RECT 1159.345 4.505 1169.635 4.675 ;
        RECT 1159.345 3.995 1159.515 4.505 ;
        RECT 1158.425 3.825 1159.515 3.995 ;
        RECT 1121.625 3.145 1121.795 3.825 ;
        RECT 835.505 2.805 836.595 2.975 ;
      LAYER mcon ;
        RECT 679.565 6.885 679.735 7.055 ;
        RECT 850.225 6.205 850.395 6.375 ;
        RECT 879.205 6.205 879.375 6.375 ;
        RECT 835.505 3.145 835.675 3.315 ;
        RECT 1183.725 8.925 1183.895 9.095 ;
        RECT 1310.225 8.925 1310.395 9.095 ;
        RECT 1344.725 8.925 1344.895 9.095 ;
        RECT 912.785 7.225 912.955 7.395 ;
        RECT 955.105 6.545 955.275 6.715 ;
        RECT 1158.425 5.525 1158.595 5.695 ;
      LAYER met1 ;
        RECT 1183.665 9.080 1183.955 9.125 ;
        RECT 1292.225 9.080 1292.515 9.125 ;
        RECT 1183.665 8.940 1292.515 9.080 ;
        RECT 1183.665 8.895 1183.955 8.940 ;
        RECT 1292.225 8.895 1292.515 8.940 ;
        RECT 1310.165 9.080 1310.455 9.125 ;
        RECT 1344.665 9.080 1344.955 9.125 ;
        RECT 1310.165 8.940 1313.140 9.080 ;
        RECT 1310.165 8.895 1310.455 8.940 ;
        RECT 1313.000 8.740 1313.140 8.940 ;
        RECT 1344.665 8.940 1838.920 9.080 ;
        RECT 1344.665 8.895 1344.955 8.940 ;
        RECT 1343.745 8.740 1344.035 8.785 ;
        RECT 1313.000 8.600 1344.035 8.740 ;
        RECT 1838.780 8.740 1838.920 8.940 ;
        RECT 1879.630 8.740 1879.950 8.800 ;
        RECT 1838.780 8.600 1879.950 8.740 ;
        RECT 1343.745 8.555 1344.035 8.600 ;
        RECT 1879.630 8.540 1879.950 8.600 ;
        RECT 903.985 7.380 904.275 7.425 ;
        RECT 912.725 7.380 913.015 7.425 ;
        RECT 903.985 7.240 913.015 7.380 ;
        RECT 903.985 7.195 904.275 7.240 ;
        RECT 912.725 7.195 913.015 7.240 ;
        RECT 679.505 7.040 679.795 7.085 ;
        RECT 693.305 7.040 693.595 7.085 ;
        RECT 679.505 6.900 693.595 7.040 ;
        RECT 679.505 6.855 679.795 6.900 ;
        RECT 693.305 6.855 693.595 6.900 ;
        RECT 954.110 6.700 954.430 6.760 ;
        RECT 955.045 6.700 955.335 6.745 ;
        RECT 954.110 6.560 955.335 6.700 ;
        RECT 954.110 6.500 954.430 6.560 ;
        RECT 955.045 6.515 955.335 6.560 ;
        RECT 673.050 6.360 673.370 6.420 ;
        RECT 673.525 6.360 673.815 6.405 ;
        RECT 673.050 6.220 673.815 6.360 ;
        RECT 673.050 6.160 673.370 6.220 ;
        RECT 673.525 6.175 673.815 6.220 ;
        RECT 850.165 6.360 850.455 6.405 ;
        RECT 879.145 6.360 879.435 6.405 ;
        RECT 850.165 6.220 879.435 6.360 ;
        RECT 850.165 6.175 850.455 6.220 ;
        RECT 879.145 6.175 879.435 6.220 ;
        RECT 748.950 6.020 749.270 6.080 ;
        RECT 748.120 5.880 749.270 6.020 ;
        RECT 748.120 5.680 748.260 5.880 ;
        RECT 748.950 5.820 749.270 5.880 ;
        RECT 740.300 5.540 748.260 5.680 ;
        RECT 1128.005 5.680 1128.295 5.725 ;
        RECT 1158.365 5.680 1158.655 5.725 ;
        RECT 1128.005 5.540 1158.655 5.680 ;
        RECT 738.845 5.340 739.135 5.385 ;
        RECT 740.300 5.340 740.440 5.540 ;
        RECT 1128.005 5.495 1128.295 5.540 ;
        RECT 1158.365 5.495 1158.655 5.540 ;
        RECT 738.845 5.200 740.440 5.340 ;
        RECT 738.845 5.155 739.135 5.200 ;
        RECT 833.130 3.300 833.450 3.360 ;
        RECT 835.445 3.300 835.735 3.345 ;
        RECT 833.130 3.160 835.735 3.300 ;
        RECT 833.130 3.100 833.450 3.160 ;
        RECT 835.445 3.115 835.735 3.160 ;
        RECT 1121.090 3.300 1121.410 3.360 ;
        RECT 1121.565 3.300 1121.855 3.345 ;
        RECT 1121.090 3.160 1121.855 3.300 ;
        RECT 1121.090 3.100 1121.410 3.160 ;
        RECT 1121.565 3.115 1121.855 3.160 ;
      LAYER via ;
        RECT 1879.660 8.540 1879.920 8.800 ;
        RECT 954.140 6.500 954.400 6.760 ;
        RECT 673.080 6.160 673.340 6.420 ;
        RECT 748.980 5.820 749.240 6.080 ;
        RECT 833.160 3.100 833.420 3.360 ;
        RECT 1121.120 3.100 1121.380 3.360 ;
      LAYER met2 ;
        RECT 1879.660 8.570 1879.920 8.830 ;
        RECT 1880.970 8.570 1881.250 9.000 ;
        RECT 1879.660 8.510 1881.250 8.570 ;
        RECT 1879.720 8.430 1881.250 8.510 ;
        RECT 648.760 6.900 659.020 7.040 ;
        RECT 648.760 4.320 648.900 6.900 ;
        RECT 658.880 5.850 659.020 6.900 ;
        RECT 954.140 6.470 954.400 6.790 ;
        RECT 673.080 6.360 673.340 6.450 ;
        RECT 662.560 6.220 673.340 6.360 ;
        RECT 662.560 5.850 662.700 6.220 ;
        RECT 673.080 6.130 673.340 6.220 ;
        RECT 658.880 5.710 662.700 5.850 ;
        RECT 748.980 5.790 749.240 6.110 ;
        RECT 954.200 5.965 954.340 6.470 ;
        RECT 1045.280 6.390 1046.800 6.530 ;
        RECT 1045.280 5.965 1045.420 6.390 ;
        RECT 749.040 4.660 749.180 5.790 ;
        RECT 954.130 5.595 954.410 5.965 ;
        RECT 1045.210 5.595 1045.490 5.965 ;
        RECT 1046.660 5.850 1046.800 6.390 ;
        RECT 1047.510 5.850 1047.790 5.965 ;
        RECT 1046.660 5.710 1047.790 5.850 ;
        RECT 1047.510 5.595 1047.790 5.710 ;
        RECT 1059.470 5.680 1059.750 5.965 ;
        RECT 1059.470 5.595 1069.800 5.680 ;
        RECT 1059.540 5.540 1069.800 5.595 ;
        RECT 833.150 4.915 833.430 5.285 ;
        RECT 749.040 4.520 753.780 4.660 ;
        RECT 647.840 4.180 648.900 4.320 ;
        RECT 647.840 3.130 647.980 4.180 ;
        RECT 627.140 2.990 647.980 3.130 ;
        RECT 753.640 3.130 753.780 4.520 ;
        RECT 833.220 3.390 833.360 4.915 ;
        RECT 1069.660 4.490 1069.800 5.540 ;
        RECT 1074.260 5.030 1104.300 5.170 ;
        RECT 1074.260 4.490 1074.400 5.030 ;
        RECT 1069.660 4.350 1074.400 4.490 ;
        RECT 1104.160 4.490 1104.300 5.030 ;
        RECT 1880.970 5.000 1881.250 8.430 ;
        RECT 1104.160 4.350 1107.520 4.490 ;
        RECT 755.410 3.130 755.690 3.245 ;
        RECT 753.640 2.990 755.690 3.130 ;
        RECT 833.160 3.070 833.420 3.390 ;
        RECT 1107.380 3.300 1107.520 4.350 ;
        RECT 1121.120 3.300 1121.380 3.390 ;
        RECT 1107.380 3.160 1121.380 3.300 ;
        RECT 1121.120 3.070 1121.380 3.160 ;
        RECT 627.140 2.400 627.280 2.990 ;
        RECT 755.410 2.875 755.690 2.990 ;
        RECT 626.930 -4.800 627.490 2.400 ;
      LAYER via2 ;
        RECT 954.130 5.640 954.410 5.920 ;
        RECT 1045.210 5.640 1045.490 5.920 ;
        RECT 1047.510 5.640 1047.790 5.920 ;
        RECT 1059.470 5.640 1059.750 5.920 ;
        RECT 833.150 4.960 833.430 5.240 ;
        RECT 755.410 2.920 755.690 3.200 ;
      LAYER met3 ;
        RECT 954.105 5.930 954.435 5.945 ;
        RECT 955.230 5.930 955.610 5.940 ;
        RECT 1045.185 5.930 1045.515 5.945 ;
        RECT 954.105 5.630 955.610 5.930 ;
        RECT 954.105 5.615 954.435 5.630 ;
        RECT 955.230 5.620 955.610 5.630 ;
        RECT 991.150 5.630 1045.515 5.930 ;
        RECT 819.070 5.250 819.450 5.260 ;
        RECT 833.125 5.250 833.455 5.265 ;
        RECT 819.070 4.950 833.455 5.250 ;
        RECT 819.070 4.940 819.450 4.950 ;
        RECT 833.125 4.935 833.455 4.950 ;
        RECT 986.510 5.250 986.890 5.260 ;
        RECT 991.150 5.250 991.450 5.630 ;
        RECT 1045.185 5.615 1045.515 5.630 ;
        RECT 1047.485 5.930 1047.815 5.945 ;
        RECT 1059.445 5.930 1059.775 5.945 ;
        RECT 1047.485 5.630 1059.775 5.930 ;
        RECT 1047.485 5.615 1047.815 5.630 ;
        RECT 1059.445 5.615 1059.775 5.630 ;
        RECT 986.510 4.950 991.450 5.250 ;
        RECT 986.510 4.940 986.890 4.950 ;
        RECT 755.385 3.210 755.715 3.225 ;
        RECT 756.510 3.210 756.890 3.220 ;
        RECT 755.385 2.910 756.890 3.210 ;
        RECT 755.385 2.895 755.715 2.910 ;
        RECT 756.510 2.900 756.890 2.910 ;
      LAYER via3 ;
        RECT 955.260 5.620 955.580 5.940 ;
        RECT 819.100 4.940 819.420 5.260 ;
        RECT 986.540 4.940 986.860 5.260 ;
        RECT 756.540 2.900 756.860 3.220 ;
      LAYER met4 ;
        RECT 955.255 5.615 955.585 5.945 ;
        RECT 819.095 4.935 819.425 5.265 ;
        RECT 955.270 5.250 955.570 5.615 ;
        RECT 986.535 5.250 986.865 5.265 ;
        RECT 955.270 4.950 986.865 5.250 ;
        RECT 986.535 4.935 986.865 4.950 ;
        RECT 756.535 3.210 756.865 3.225 ;
        RECT 756.535 2.910 757.770 3.210 ;
        RECT 756.535 2.895 756.865 2.910 ;
        RECT 757.470 2.290 757.770 2.910 ;
        RECT 819.110 2.290 819.410 4.935 ;
        RECT 757.030 1.110 758.210 2.290 ;
        RECT 818.670 1.110 819.850 2.290 ;
      LAYER met5 ;
        RECT 756.820 0.900 820.060 2.500 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 358.945 8.245 359.575 8.415 ;
        RECT 606.885 8.245 607.515 8.415 ;
        RECT 245.325 5.865 245.495 7.395 ;
        RECT 358.945 6.885 359.115 8.245 ;
        RECT 316.625 4.505 316.795 6.035 ;
        RECT 607.345 4.845 607.515 8.245 ;
        RECT 609.185 2.635 609.355 5.015 ;
        RECT 626.205 4.505 645.695 4.675 ;
        RECT 626.205 3.655 626.375 4.505 ;
        RECT 622.985 3.485 626.375 3.655 ;
        RECT 622.985 2.635 623.155 3.485 ;
        RECT 609.185 2.465 623.155 2.635 ;
      LAYER mcon ;
        RECT 359.405 8.245 359.575 8.415 ;
        RECT 245.325 7.225 245.495 7.395 ;
        RECT 316.625 5.865 316.795 6.035 ;
        RECT 609.185 4.845 609.355 5.015 ;
        RECT 645.525 4.505 645.695 4.675 ;
      LAYER met1 ;
        RECT 359.345 8.400 359.635 8.445 ;
        RECT 606.825 8.400 607.115 8.445 ;
        RECT 359.345 8.260 607.115 8.400 ;
        RECT 359.345 8.215 359.635 8.260 ;
        RECT 606.825 8.215 607.115 8.260 ;
        RECT 245.265 7.380 245.555 7.425 ;
        RECT 289.870 7.380 290.190 7.440 ;
        RECT 245.265 7.240 290.190 7.380 ;
        RECT 245.265 7.195 245.555 7.240 ;
        RECT 289.870 7.180 290.190 7.240 ;
        RECT 344.610 7.040 344.930 7.100 ;
        RECT 358.885 7.040 359.175 7.085 ;
        RECT 344.610 6.900 359.175 7.040 ;
        RECT 344.610 6.840 344.930 6.900 ;
        RECT 358.885 6.855 359.175 6.900 ;
        RECT 196.950 6.020 197.270 6.080 ;
        RECT 245.265 6.020 245.555 6.065 ;
        RECT 196.950 5.880 245.555 6.020 ;
        RECT 196.950 5.820 197.270 5.880 ;
        RECT 245.265 5.835 245.555 5.880 ;
        RECT 289.870 6.020 290.190 6.080 ;
        RECT 316.565 6.020 316.855 6.065 ;
        RECT 289.870 5.880 316.855 6.020 ;
        RECT 289.870 5.820 290.190 5.880 ;
        RECT 316.565 5.835 316.855 5.880 ;
        RECT 607.285 5.000 607.575 5.045 ;
        RECT 609.125 5.000 609.415 5.045 ;
        RECT 607.285 4.860 609.415 5.000 ;
        RECT 607.285 4.815 607.575 4.860 ;
        RECT 609.125 4.815 609.415 4.860 ;
        RECT 316.565 4.660 316.855 4.705 ;
        RECT 324.370 4.660 324.690 4.720 ;
        RECT 316.565 4.520 324.690 4.660 ;
        RECT 316.565 4.475 316.855 4.520 ;
        RECT 324.370 4.460 324.690 4.520 ;
        RECT 645.450 4.660 645.770 4.720 ;
        RECT 645.450 4.520 645.965 4.660 ;
        RECT 645.450 4.460 645.770 4.520 ;
      LAYER via ;
        RECT 289.900 7.180 290.160 7.440 ;
        RECT 344.640 6.840 344.900 7.100 ;
        RECT 196.980 5.820 197.240 6.080 ;
        RECT 289.900 5.820 290.160 6.080 ;
        RECT 324.400 4.460 324.660 4.720 ;
        RECT 645.480 4.460 645.740 4.720 ;
      LAYER met2 ;
        RECT 163.390 7.635 163.670 8.005 ;
        RECT 196.970 7.635 197.250 8.005 ;
        RECT 163.460 2.400 163.600 7.635 ;
        RECT 197.040 6.110 197.180 7.635 ;
        RECT 289.900 7.150 290.160 7.470 ;
        RECT 289.960 6.110 290.100 7.150 ;
        RECT 344.640 6.810 344.900 7.130 ;
        RECT 196.980 5.790 197.240 6.110 ;
        RECT 289.900 5.790 290.160 6.110 ;
        RECT 344.700 5.850 344.840 6.810 ;
        RECT 340.560 5.710 344.840 5.850 ;
        RECT 324.400 4.490 324.660 4.750 ;
        RECT 324.400 4.430 325.060 4.490 ;
        RECT 324.460 4.350 325.060 4.430 ;
        RECT 324.920 2.450 325.060 4.350 ;
        RECT 340.560 2.565 340.700 5.710 ;
        RECT 645.870 5.170 646.150 9.000 ;
        RECT 645.540 5.030 646.150 5.170 ;
        RECT 645.540 4.750 645.680 5.030 ;
        RECT 645.870 5.000 646.150 5.030 ;
        RECT 645.480 4.430 645.740 4.750 ;
        RECT 326.690 2.450 326.970 2.565 ;
        RECT 163.250 -4.800 163.810 2.400 ;
        RECT 324.920 2.310 326.970 2.450 ;
        RECT 326.690 2.195 326.970 2.310 ;
        RECT 340.490 2.195 340.770 2.565 ;
      LAYER via2 ;
        RECT 163.390 7.680 163.670 7.960 ;
        RECT 196.970 7.680 197.250 7.960 ;
        RECT 326.690 2.240 326.970 2.520 ;
        RECT 340.490 2.240 340.770 2.520 ;
      LAYER met3 ;
        RECT 163.365 7.970 163.695 7.985 ;
        RECT 196.945 7.970 197.275 7.985 ;
        RECT 163.365 7.670 197.275 7.970 ;
        RECT 163.365 7.655 163.695 7.670 ;
        RECT 196.945 7.655 197.275 7.670 ;
        RECT 326.665 2.530 326.995 2.545 ;
        RECT 340.465 2.530 340.795 2.545 ;
        RECT 326.665 2.230 340.795 2.530 ;
        RECT 326.665 2.215 326.995 2.230 ;
        RECT 340.465 2.215 340.795 2.230 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 626.665 9.605 631.895 9.775 ;
        RECT 245.325 7.735 245.495 8.075 ;
        RECT 244.405 7.565 245.495 7.735 ;
        RECT 556.285 6.205 556.455 8.075 ;
        RECT 559.045 6.545 560.595 6.715 ;
        RECT 559.045 6.205 559.215 6.545 ;
        RECT 560.425 5.865 560.595 6.545 ;
        RECT 582.965 5.865 583.135 8.075 ;
        RECT 626.665 7.905 626.835 9.605 ;
        RECT 631.725 9.435 631.895 9.605 ;
        RECT 631.725 9.265 637.875 9.435 ;
        RECT 637.705 7.735 637.875 9.265 ;
        RECT 651.505 8.925 652.595 9.095 ;
        RECT 646.905 8.585 647.995 8.755 ;
        RECT 651.505 8.585 651.675 8.925 ;
        RECT 671.285 8.755 671.455 9.095 ;
        RECT 671.285 8.585 671.915 8.755 ;
        RECT 646.905 8.245 647.075 8.585 ;
        RECT 671.745 8.415 671.915 8.585 ;
        RECT 671.745 8.245 673.295 8.415 ;
        RECT 675.425 8.245 686.635 8.415 ;
        RECT 640.925 7.735 641.095 8.075 ;
        RECT 637.705 7.565 641.095 7.735 ;
      LAYER mcon ;
        RECT 245.325 7.905 245.495 8.075 ;
        RECT 556.285 7.905 556.455 8.075 ;
        RECT 582.965 7.905 583.135 8.075 ;
        RECT 652.425 8.925 652.595 9.095 ;
        RECT 671.285 8.925 671.455 9.095 ;
        RECT 647.825 8.585 647.995 8.755 ;
        RECT 673.125 8.245 673.295 8.415 ;
        RECT 686.465 8.245 686.635 8.415 ;
        RECT 640.925 7.905 641.095 8.075 ;
      LAYER met1 ;
        RECT 652.365 9.080 652.655 9.125 ;
        RECT 671.225 9.080 671.515 9.125 ;
        RECT 652.365 8.940 671.515 9.080 ;
        RECT 652.365 8.895 652.655 8.940 ;
        RECT 671.225 8.895 671.515 8.940 ;
        RECT 647.765 8.740 648.055 8.785 ;
        RECT 651.445 8.740 651.735 8.785 ;
        RECT 647.765 8.600 651.735 8.740 ;
        RECT 647.765 8.555 648.055 8.600 ;
        RECT 651.445 8.555 651.735 8.600 ;
        RECT 646.845 8.400 647.135 8.445 ;
        RECT 643.700 8.260 647.135 8.400 ;
        RECT 245.265 8.060 245.555 8.105 ;
        RECT 556.225 8.060 556.515 8.105 ;
        RECT 245.265 7.920 556.515 8.060 ;
        RECT 245.265 7.875 245.555 7.920 ;
        RECT 556.225 7.875 556.515 7.920 ;
        RECT 582.905 8.060 583.195 8.105 ;
        RECT 626.605 8.060 626.895 8.105 ;
        RECT 582.905 7.920 626.895 8.060 ;
        RECT 582.905 7.875 583.195 7.920 ;
        RECT 626.605 7.875 626.895 7.920 ;
        RECT 640.865 8.060 641.155 8.105 ;
        RECT 643.700 8.060 643.840 8.260 ;
        RECT 646.845 8.215 647.135 8.260 ;
        RECT 673.065 8.400 673.355 8.445 ;
        RECT 675.365 8.400 675.655 8.445 ;
        RECT 673.065 8.260 675.655 8.400 ;
        RECT 673.065 8.215 673.355 8.260 ;
        RECT 675.365 8.215 675.655 8.260 ;
        RECT 686.405 8.400 686.695 8.445 ;
        RECT 691.450 8.400 691.770 8.460 ;
        RECT 686.405 8.260 691.770 8.400 ;
        RECT 686.405 8.215 686.695 8.260 ;
        RECT 691.450 8.200 691.770 8.260 ;
        RECT 640.865 7.920 643.840 8.060 ;
        RECT 640.865 7.875 641.155 7.920 ;
        RECT 180.850 7.720 181.170 7.780 ;
        RECT 180.850 7.580 197.640 7.720 ;
        RECT 180.850 7.520 181.170 7.580 ;
        RECT 197.500 7.380 197.640 7.580 ;
        RECT 244.345 7.535 244.635 7.765 ;
        RECT 244.420 7.380 244.560 7.535 ;
        RECT 197.500 7.240 244.560 7.380 ;
        RECT 556.225 6.360 556.515 6.405 ;
        RECT 558.985 6.360 559.275 6.405 ;
        RECT 556.225 6.220 559.275 6.360 ;
        RECT 556.225 6.175 556.515 6.220 ;
        RECT 558.985 6.175 559.275 6.220 ;
        RECT 560.365 6.020 560.655 6.065 ;
        RECT 582.905 6.020 583.195 6.065 ;
        RECT 560.365 5.880 583.195 6.020 ;
        RECT 560.365 5.835 560.655 5.880 ;
        RECT 582.905 5.835 583.195 5.880 ;
      LAYER via ;
        RECT 691.480 8.200 691.740 8.460 ;
        RECT 180.880 7.520 181.140 7.780 ;
      LAYER met2 ;
        RECT 691.480 8.170 691.740 8.490 ;
        RECT 691.540 7.890 691.680 8.170 ;
        RECT 693.250 7.890 693.530 9.000 ;
        RECT 180.880 7.490 181.140 7.810 ;
        RECT 691.540 7.750 693.530 7.890 ;
        RECT 180.940 2.400 181.080 7.490 ;
        RECT 693.250 5.000 693.530 7.750 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 316.165 6.375 316.335 8.415 ;
        RECT 317.085 6.375 317.255 6.715 ;
        RECT 335.025 6.545 335.195 7.735 ;
        RECT 414.145 7.565 417.535 7.735 ;
        RECT 437.605 6.885 437.775 7.735 ;
        RECT 459.225 6.885 462.155 7.055 ;
        RECT 461.985 6.545 462.155 6.885 ;
        RECT 316.165 6.205 317.255 6.375 ;
      LAYER mcon ;
        RECT 316.165 8.245 316.335 8.415 ;
        RECT 335.025 7.565 335.195 7.735 ;
        RECT 417.365 7.565 417.535 7.735 ;
        RECT 437.605 7.565 437.775 7.735 ;
        RECT 317.085 6.545 317.255 6.715 ;
      LAYER met1 ;
        RECT 559.890 8.740 560.210 8.800 ;
        RECT 559.890 8.600 607.500 8.740 ;
        RECT 559.890 8.540 560.210 8.600 ;
        RECT 227.770 8.400 228.090 8.460 ;
        RECT 214.060 8.260 228.090 8.400 ;
        RECT 212.590 8.060 212.910 8.120 ;
        RECT 214.060 8.060 214.200 8.260 ;
        RECT 227.770 8.200 228.090 8.260 ;
        RECT 289.410 8.400 289.730 8.460 ;
        RECT 316.105 8.400 316.395 8.445 ;
        RECT 289.410 8.260 316.395 8.400 ;
        RECT 607.360 8.400 607.500 8.600 ;
        RECT 622.910 8.400 623.230 8.460 ;
        RECT 607.360 8.260 623.230 8.400 ;
        RECT 289.410 8.200 289.730 8.260 ;
        RECT 316.105 8.215 316.395 8.260 ;
        RECT 622.910 8.200 623.230 8.260 ;
        RECT 212.590 7.920 214.200 8.060 ;
        RECT 212.590 7.860 212.910 7.920 ;
        RECT 334.965 7.720 335.255 7.765 ;
        RECT 414.085 7.720 414.375 7.765 ;
        RECT 334.965 7.580 414.375 7.720 ;
        RECT 334.965 7.535 335.255 7.580 ;
        RECT 414.085 7.535 414.375 7.580 ;
        RECT 417.305 7.720 417.595 7.765 ;
        RECT 437.545 7.720 437.835 7.765 ;
        RECT 417.305 7.580 437.835 7.720 ;
        RECT 417.305 7.535 417.595 7.580 ;
        RECT 437.545 7.535 437.835 7.580 ;
        RECT 437.545 7.040 437.835 7.085 ;
        RECT 459.165 7.040 459.455 7.085 ;
        RECT 437.545 6.900 459.455 7.040 ;
        RECT 437.545 6.855 437.835 6.900 ;
        RECT 459.165 6.855 459.455 6.900 ;
        RECT 317.025 6.700 317.315 6.745 ;
        RECT 334.965 6.700 335.255 6.745 ;
        RECT 317.025 6.560 335.255 6.700 ;
        RECT 317.025 6.515 317.315 6.560 ;
        RECT 334.965 6.515 335.255 6.560 ;
        RECT 461.925 6.700 462.215 6.745 ;
        RECT 461.925 6.560 463.520 6.700 ;
        RECT 461.925 6.515 462.215 6.560 ;
        RECT 463.380 6.420 463.520 6.560 ;
        RECT 463.290 6.160 463.610 6.420 ;
      LAYER via ;
        RECT 559.920 8.540 560.180 8.800 ;
        RECT 212.620 7.860 212.880 8.120 ;
        RECT 227.800 8.200 228.060 8.460 ;
        RECT 289.440 8.200 289.700 8.460 ;
        RECT 622.940 8.200 623.200 8.460 ;
        RECT 463.320 6.160 463.580 6.420 ;
      LAYER met2 ;
        RECT 559.920 8.740 560.180 8.830 ;
        RECT 502.410 8.570 502.690 8.685 ;
        RECT 227.800 8.170 228.060 8.490 ;
        RECT 289.440 8.170 289.700 8.490 ;
        RECT 485.460 8.430 502.690 8.570 ;
        RECT 212.620 8.005 212.880 8.150 ;
        RECT 198.810 7.635 199.090 8.005 ;
        RECT 212.610 7.635 212.890 8.005 ;
        RECT 198.880 2.400 199.020 7.635 ;
        RECT 227.860 7.210 228.000 8.170 ;
        RECT 289.500 8.005 289.640 8.170 ;
        RECT 289.430 7.635 289.710 8.005 ;
        RECT 482.170 7.890 482.450 8.005 ;
        RECT 464.300 7.750 482.450 7.890 ;
        RECT 228.250 7.210 228.530 7.325 ;
        RECT 227.860 7.070 228.530 7.210 ;
        RECT 228.250 6.955 228.530 7.070 ;
        RECT 463.320 6.360 463.580 6.450 ;
        RECT 464.300 6.360 464.440 7.750 ;
        RECT 482.170 7.635 482.450 7.750 ;
        RECT 483.090 7.635 483.370 8.005 ;
        RECT 483.160 7.210 483.300 7.635 ;
        RECT 485.460 7.210 485.600 8.430 ;
        RECT 502.410 8.315 502.690 8.430 ;
        RECT 557.150 8.315 557.430 8.685 ;
        RECT 558.140 8.600 560.180 8.740 ;
        RECT 557.220 7.890 557.360 8.315 ;
        RECT 558.140 7.890 558.280 8.600 ;
        RECT 559.920 8.510 560.180 8.600 ;
        RECT 705.730 8.570 706.010 8.685 ;
        RECT 622.940 8.170 623.200 8.490 ;
        RECT 703.960 8.430 706.010 8.570 ;
        RECT 629.440 8.260 639.700 8.400 ;
        RECT 557.220 7.750 558.280 7.890 ;
        RECT 623.000 7.380 623.140 8.170 ;
        RECT 629.440 7.380 629.580 8.260 ;
        RECT 623.000 7.240 629.580 7.380 ;
        RECT 639.560 7.325 639.700 8.260 ;
        RECT 703.960 8.005 704.100 8.430 ;
        RECT 705.730 8.315 706.010 8.430 ;
        RECT 740.230 8.570 740.510 8.685 ;
        RECT 741.090 8.570 741.370 9.000 ;
        RECT 740.230 8.430 741.370 8.570 ;
        RECT 740.230 8.315 740.510 8.430 ;
        RECT 674.450 7.635 674.730 8.005 ;
        RECT 703.890 7.635 704.170 8.005 ;
        RECT 483.160 7.070 485.600 7.210 ;
        RECT 639.490 6.955 639.770 7.325 ;
        RECT 674.520 6.530 674.660 7.635 ;
        RECT 675.370 6.530 675.650 6.645 ;
        RECT 674.520 6.390 675.650 6.530 ;
        RECT 463.320 6.220 464.440 6.360 ;
        RECT 675.370 6.275 675.650 6.390 ;
        RECT 679.510 6.530 679.790 6.645 ;
        RECT 681.810 6.530 682.090 6.645 ;
        RECT 679.510 6.390 682.090 6.530 ;
        RECT 679.510 6.275 679.790 6.390 ;
        RECT 681.810 6.275 682.090 6.390 ;
        RECT 463.320 6.130 463.580 6.220 ;
        RECT 741.090 5.000 741.370 8.430 ;
        RECT 198.670 -4.800 199.230 2.400 ;
      LAYER via2 ;
        RECT 198.810 7.680 199.090 7.960 ;
        RECT 212.610 7.680 212.890 7.960 ;
        RECT 289.430 7.680 289.710 7.960 ;
        RECT 228.250 7.000 228.530 7.280 ;
        RECT 482.170 7.680 482.450 7.960 ;
        RECT 483.090 7.680 483.370 7.960 ;
        RECT 502.410 8.360 502.690 8.640 ;
        RECT 557.150 8.360 557.430 8.640 ;
        RECT 705.730 8.360 706.010 8.640 ;
        RECT 740.230 8.360 740.510 8.640 ;
        RECT 674.450 7.680 674.730 7.960 ;
        RECT 703.890 7.680 704.170 7.960 ;
        RECT 639.490 7.000 639.770 7.280 ;
        RECT 675.370 6.320 675.650 6.600 ;
        RECT 679.510 6.320 679.790 6.600 ;
        RECT 681.810 6.320 682.090 6.600 ;
      LAYER met3 ;
        RECT 502.385 8.650 502.715 8.665 ;
        RECT 513.670 8.650 515.580 8.820 ;
        RECT 557.125 8.650 557.455 8.665 ;
        RECT 502.385 8.520 557.455 8.650 ;
        RECT 502.385 8.350 513.970 8.520 ;
        RECT 515.280 8.350 557.455 8.520 ;
        RECT 502.385 8.335 502.715 8.350 ;
        RECT 557.125 8.335 557.455 8.350 ;
        RECT 705.705 8.650 706.035 8.665 ;
        RECT 731.670 8.650 732.050 8.660 ;
        RECT 740.205 8.650 740.535 8.665 ;
        RECT 705.705 8.350 707.860 8.650 ;
        RECT 705.705 8.335 706.035 8.350 ;
        RECT 198.785 7.970 199.115 7.985 ;
        RECT 212.585 7.970 212.915 7.985 ;
        RECT 289.405 7.970 289.735 7.985 ;
        RECT 198.785 7.670 212.915 7.970 ;
        RECT 198.785 7.655 199.115 7.670 ;
        RECT 212.585 7.655 212.915 7.670 ;
        RECT 274.470 7.670 289.735 7.970 ;
        RECT 228.225 7.290 228.555 7.305 ;
        RECT 274.470 7.290 274.770 7.670 ;
        RECT 289.405 7.655 289.735 7.670 ;
        RECT 482.145 7.970 482.475 7.985 ;
        RECT 483.065 7.970 483.395 7.985 ;
        RECT 674.425 7.970 674.755 7.985 ;
        RECT 703.865 7.970 704.195 7.985 ;
        RECT 482.145 7.670 483.395 7.970 ;
        RECT 482.145 7.655 482.475 7.670 ;
        RECT 483.065 7.655 483.395 7.670 ;
        RECT 644.080 7.670 674.755 7.970 ;
        RECT 644.080 7.460 644.380 7.670 ;
        RECT 674.425 7.655 674.755 7.670 ;
        RECT 683.640 7.670 704.195 7.970 ;
        RECT 707.560 7.970 707.860 8.350 ;
        RECT 731.670 8.350 740.535 8.650 ;
        RECT 731.670 8.340 732.050 8.350 ;
        RECT 740.205 8.335 740.535 8.350 ;
        RECT 724.310 7.970 724.690 7.980 ;
        RECT 707.560 7.670 724.690 7.970 ;
        RECT 228.225 6.990 274.770 7.290 ;
        RECT 639.465 7.290 639.795 7.305 ;
        RECT 643.390 7.290 644.380 7.460 ;
        RECT 639.465 7.160 644.380 7.290 ;
        RECT 639.465 6.990 643.690 7.160 ;
        RECT 228.225 6.975 228.555 6.990 ;
        RECT 639.465 6.975 639.795 6.990 ;
        RECT 675.345 6.610 675.675 6.625 ;
        RECT 679.485 6.610 679.815 6.625 ;
        RECT 675.345 6.310 679.815 6.610 ;
        RECT 675.345 6.295 675.675 6.310 ;
        RECT 679.485 6.295 679.815 6.310 ;
        RECT 681.785 6.610 682.115 6.625 ;
        RECT 683.640 6.610 683.940 7.670 ;
        RECT 703.865 7.655 704.195 7.670 ;
        RECT 724.310 7.660 724.690 7.670 ;
        RECT 681.785 6.310 683.940 6.610 ;
        RECT 681.785 6.295 682.115 6.310 ;
      LAYER via3 ;
        RECT 731.700 8.340 732.020 8.660 ;
        RECT 724.340 7.660 724.660 7.980 ;
      LAYER met4 ;
        RECT 731.695 8.335 732.025 8.665 ;
        RECT 724.335 7.655 724.665 7.985 ;
        RECT 724.350 7.290 724.650 7.655 ;
        RECT 731.710 7.290 732.010 8.335 ;
        RECT 724.350 6.990 732.010 7.290 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 435.765 9.265 464.915 9.435 ;
        RECT 373.205 8.585 393.615 8.755 ;
        RECT 317.545 4.165 318.175 4.335 ;
        RECT 318.005 1.105 318.175 4.165 ;
        RECT 373.205 2.295 373.375 8.585 ;
        RECT 393.445 7.225 393.615 8.585 ;
        RECT 435.765 8.415 435.935 9.265 ;
        RECT 464.745 8.755 464.915 9.265 ;
        RECT 464.745 8.585 466.755 8.755 ;
        RECT 413.225 8.245 435.935 8.415 ;
        RECT 413.225 7.225 413.395 8.245 ;
        RECT 466.585 5.865 466.755 8.585 ;
        RECT 522.705 5.865 522.875 7.735 ;
        RECT 683.245 7.565 684.335 7.735 ;
        RECT 712.225 7.565 715.155 7.735 ;
        RECT 720.505 7.565 722.055 7.735 ;
        RECT 725.565 7.565 726.195 7.735 ;
        RECT 757.765 5.525 757.935 8.075 ;
        RECT 764.205 5.525 764.375 7.055 ;
        RECT 782.605 6.205 782.775 7.055 ;
        RECT 786.745 6.205 786.915 7.735 ;
        RECT 367.685 2.125 373.375 2.295 ;
        RECT 367.685 1.105 367.855 2.125 ;
      LAYER mcon ;
        RECT 757.765 7.905 757.935 8.075 ;
        RECT 522.705 7.565 522.875 7.735 ;
        RECT 684.165 7.565 684.335 7.735 ;
        RECT 714.985 7.565 715.155 7.735 ;
        RECT 721.885 7.565 722.055 7.735 ;
        RECT 726.025 7.565 726.195 7.735 ;
        RECT 786.745 7.565 786.915 7.735 ;
        RECT 764.205 6.885 764.375 7.055 ;
        RECT 782.605 6.885 782.775 7.055 ;
      LAYER met1 ;
        RECT 757.705 8.060 757.995 8.105 ;
        RECT 756.860 7.920 757.995 8.060 ;
        RECT 522.645 7.720 522.935 7.765 ;
        RECT 683.185 7.720 683.475 7.765 ;
        RECT 522.645 7.580 647.060 7.720 ;
        RECT 522.645 7.535 522.935 7.580 ;
        RECT 393.385 7.380 393.675 7.425 ;
        RECT 413.165 7.380 413.455 7.425 ;
        RECT 393.385 7.240 413.455 7.380 ;
        RECT 646.920 7.380 647.060 7.580 ;
        RECT 648.300 7.580 683.475 7.720 ;
        RECT 648.300 7.380 648.440 7.580 ;
        RECT 683.185 7.535 683.475 7.580 ;
        RECT 684.105 7.720 684.395 7.765 ;
        RECT 712.165 7.720 712.455 7.765 ;
        RECT 684.105 7.580 712.455 7.720 ;
        RECT 684.105 7.535 684.395 7.580 ;
        RECT 712.165 7.535 712.455 7.580 ;
        RECT 714.925 7.720 715.215 7.765 ;
        RECT 720.445 7.720 720.735 7.765 ;
        RECT 714.925 7.580 720.735 7.720 ;
        RECT 714.925 7.535 715.215 7.580 ;
        RECT 720.445 7.535 720.735 7.580 ;
        RECT 721.825 7.720 722.115 7.765 ;
        RECT 725.505 7.720 725.795 7.765 ;
        RECT 721.825 7.580 725.795 7.720 ;
        RECT 721.825 7.535 722.115 7.580 ;
        RECT 725.505 7.535 725.795 7.580 ;
        RECT 725.965 7.720 726.255 7.765 ;
        RECT 756.860 7.720 757.000 7.920 ;
        RECT 757.705 7.875 757.995 7.920 ;
        RECT 786.670 7.720 786.990 7.780 ;
        RECT 725.965 7.580 757.000 7.720 ;
        RECT 786.475 7.580 786.990 7.720 ;
        RECT 725.965 7.535 726.255 7.580 ;
        RECT 786.670 7.520 786.990 7.580 ;
        RECT 646.920 7.240 648.440 7.380 ;
        RECT 393.385 7.195 393.675 7.240 ;
        RECT 413.165 7.195 413.455 7.240 ;
        RECT 764.145 7.040 764.435 7.085 ;
        RECT 782.545 7.040 782.835 7.085 ;
        RECT 764.145 6.900 782.835 7.040 ;
        RECT 764.145 6.855 764.435 6.900 ;
        RECT 782.545 6.855 782.835 6.900 ;
        RECT 782.545 6.360 782.835 6.405 ;
        RECT 786.685 6.360 786.975 6.405 ;
        RECT 782.545 6.220 786.975 6.360 ;
        RECT 782.545 6.175 782.835 6.220 ;
        RECT 786.685 6.175 786.975 6.220 ;
        RECT 466.525 6.020 466.815 6.065 ;
        RECT 522.645 6.020 522.935 6.065 ;
        RECT 466.525 5.880 522.935 6.020 ;
        RECT 466.525 5.835 466.815 5.880 ;
        RECT 522.645 5.835 522.935 5.880 ;
        RECT 757.705 5.680 757.995 5.725 ;
        RECT 764.145 5.680 764.435 5.725 ;
        RECT 757.705 5.540 764.435 5.680 ;
        RECT 757.705 5.495 757.995 5.540 ;
        RECT 764.145 5.495 764.435 5.540 ;
        RECT 317.485 4.320 317.775 4.365 ;
        RECT 234.760 4.180 317.775 4.320 ;
        RECT 216.730 3.980 217.050 4.040 ;
        RECT 234.760 3.980 234.900 4.180 ;
        RECT 317.485 4.135 317.775 4.180 ;
        RECT 216.730 3.840 234.900 3.980 ;
        RECT 216.730 3.780 217.050 3.840 ;
        RECT 317.945 1.260 318.235 1.305 ;
        RECT 334.490 1.260 334.810 1.320 ;
        RECT 317.945 1.120 334.810 1.260 ;
        RECT 317.945 1.075 318.235 1.120 ;
        RECT 334.490 1.060 334.810 1.120 ;
        RECT 367.610 1.260 367.930 1.320 ;
        RECT 367.610 1.120 368.125 1.260 ;
        RECT 367.610 1.060 367.930 1.120 ;
      LAYER via ;
        RECT 786.700 7.520 786.960 7.780 ;
        RECT 216.760 3.780 217.020 4.040 ;
        RECT 334.520 1.060 334.780 1.320 ;
        RECT 367.640 1.060 367.900 1.320 ;
      LAYER met2 ;
        RECT 788.470 7.890 788.750 9.000 ;
        RECT 786.760 7.810 788.750 7.890 ;
        RECT 786.700 7.750 788.750 7.810 ;
        RECT 786.700 7.490 786.960 7.750 ;
        RECT 788.470 5.000 788.750 7.750 ;
        RECT 216.760 3.750 217.020 4.070 ;
        RECT 216.820 2.400 216.960 3.750 ;
        RECT 216.610 -4.800 217.170 2.400 ;
        RECT 334.520 1.205 334.780 1.350 ;
        RECT 367.640 1.205 367.900 1.350 ;
        RECT 334.510 0.835 334.790 1.205 ;
        RECT 367.630 0.835 367.910 1.205 ;
      LAYER via2 ;
        RECT 334.510 0.880 334.790 1.160 ;
        RECT 367.630 0.880 367.910 1.160 ;
      LAYER met3 ;
        RECT 334.485 1.170 334.815 1.185 ;
        RECT 367.605 1.170 367.935 1.185 ;
        RECT 334.485 0.870 367.935 1.170 ;
        RECT 334.485 0.855 334.815 0.870 ;
        RECT 367.605 0.855 367.935 0.870 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 381.025 7.565 382.115 7.735 ;
        RECT 306.505 4.505 306.675 6.715 ;
        RECT 364.925 5.865 366.015 6.035 ;
        RECT 381.025 5.865 381.195 7.565 ;
        RECT 381.945 7.225 382.115 7.565 ;
        RECT 557.205 5.695 557.375 8.075 ;
        RECT 643.685 6.545 643.855 7.395 ;
        RECT 646.445 7.225 648.915 7.395 ;
        RECT 559.965 5.695 560.135 6.035 ;
        RECT 557.205 5.525 560.135 5.695 ;
        RECT 670.825 5.695 670.995 7.395 ;
        RECT 670.825 5.525 674.675 5.695 ;
        RECT 248.545 3.145 248.715 3.995 ;
      LAYER mcon ;
        RECT 557.205 7.905 557.375 8.075 ;
        RECT 306.505 6.545 306.675 6.715 ;
        RECT 365.845 5.865 366.015 6.035 ;
        RECT 643.685 7.225 643.855 7.395 ;
        RECT 648.745 7.225 648.915 7.395 ;
        RECT 670.825 7.225 670.995 7.395 ;
        RECT 559.965 5.865 560.135 6.035 ;
        RECT 674.505 5.525 674.675 5.695 ;
        RECT 248.545 3.825 248.715 3.995 ;
      LAYER met1 ;
        RECT 556.670 8.060 556.990 8.120 ;
        RECT 557.145 8.060 557.435 8.105 ;
        RECT 556.670 7.920 557.435 8.060 ;
        RECT 556.670 7.860 556.990 7.920 ;
        RECT 557.145 7.875 557.435 7.920 ;
        RECT 381.885 7.380 382.175 7.425 ;
        RECT 392.910 7.380 393.230 7.440 ;
        RECT 381.885 7.240 393.230 7.380 ;
        RECT 381.885 7.195 382.175 7.240 ;
        RECT 392.910 7.180 393.230 7.240 ;
        RECT 643.625 7.380 643.915 7.425 ;
        RECT 646.385 7.380 646.675 7.425 ;
        RECT 643.625 7.240 646.675 7.380 ;
        RECT 643.625 7.195 643.915 7.240 ;
        RECT 646.385 7.195 646.675 7.240 ;
        RECT 648.685 7.380 648.975 7.425 ;
        RECT 670.765 7.380 671.055 7.425 ;
        RECT 648.685 7.240 671.055 7.380 ;
        RECT 648.685 7.195 648.975 7.240 ;
        RECT 670.765 7.195 671.055 7.240 ;
        RECT 295.850 6.700 296.170 6.760 ;
        RECT 306.445 6.700 306.735 6.745 ;
        RECT 295.850 6.560 306.735 6.700 ;
        RECT 295.850 6.500 296.170 6.560 ;
        RECT 306.445 6.515 306.735 6.560 ;
        RECT 643.625 6.515 643.915 6.745 ;
        RECT 642.690 6.360 643.010 6.420 ;
        RECT 643.700 6.360 643.840 6.515 ;
        RECT 642.690 6.220 643.840 6.360 ;
        RECT 642.690 6.160 643.010 6.220 ;
        RECT 334.490 6.020 334.810 6.080 ;
        RECT 364.865 6.020 365.155 6.065 ;
        RECT 334.490 5.880 365.155 6.020 ;
        RECT 334.490 5.820 334.810 5.880 ;
        RECT 364.865 5.835 365.155 5.880 ;
        RECT 365.785 6.020 366.075 6.065 ;
        RECT 380.965 6.020 381.255 6.065 ;
        RECT 559.890 6.020 560.210 6.080 ;
        RECT 365.785 5.880 381.255 6.020 ;
        RECT 559.695 5.880 560.210 6.020 ;
        RECT 365.785 5.835 366.075 5.880 ;
        RECT 380.965 5.835 381.255 5.880 ;
        RECT 559.890 5.820 560.210 5.880 ;
        RECT 674.445 5.680 674.735 5.725 ;
        RECT 701.110 5.680 701.430 5.740 ;
        RECT 674.445 5.540 701.430 5.680 ;
        RECT 674.445 5.495 674.735 5.540 ;
        RECT 701.110 5.480 701.430 5.540 ;
        RECT 792.190 5.680 792.510 5.740 ;
        RECT 802.770 5.680 803.090 5.740 ;
        RECT 792.190 5.540 803.090 5.680 ;
        RECT 792.190 5.480 792.510 5.540 ;
        RECT 802.770 5.480 803.090 5.540 ;
        RECT 805.070 5.680 805.390 5.740 ;
        RECT 834.510 5.680 834.830 5.740 ;
        RECT 805.070 5.540 834.830 5.680 ;
        RECT 805.070 5.480 805.390 5.540 ;
        RECT 834.510 5.480 834.830 5.540 ;
        RECT 306.445 4.660 306.735 4.705 ;
        RECT 314.710 4.660 315.030 4.720 ;
        RECT 306.445 4.520 315.030 4.660 ;
        RECT 306.445 4.475 306.735 4.520 ;
        RECT 314.710 4.460 315.030 4.520 ;
        RECT 248.485 3.980 248.775 4.025 ;
        RECT 276.070 3.980 276.390 4.040 ;
        RECT 248.485 3.840 276.390 3.980 ;
        RECT 248.485 3.795 248.775 3.840 ;
        RECT 276.070 3.780 276.390 3.840 ;
        RECT 234.670 3.300 234.990 3.360 ;
        RECT 248.485 3.300 248.775 3.345 ;
        RECT 234.670 3.160 248.775 3.300 ;
        RECT 234.670 3.100 234.990 3.160 ;
        RECT 248.485 3.115 248.775 3.160 ;
      LAYER via ;
        RECT 556.700 7.860 556.960 8.120 ;
        RECT 392.940 7.180 393.200 7.440 ;
        RECT 295.880 6.500 296.140 6.760 ;
        RECT 642.720 6.160 642.980 6.420 ;
        RECT 334.520 5.820 334.780 6.080 ;
        RECT 559.920 5.820 560.180 6.080 ;
        RECT 701.140 5.480 701.400 5.740 ;
        RECT 792.220 5.480 792.480 5.740 ;
        RECT 802.800 5.480 803.060 5.740 ;
        RECT 805.100 5.480 805.360 5.740 ;
        RECT 834.540 5.480 834.800 5.740 ;
        RECT 314.740 4.460 315.000 4.720 ;
        RECT 276.100 3.780 276.360 4.040 ;
        RECT 234.700 3.100 234.960 3.360 ;
      LAYER met2 ;
        RECT 276.090 8.315 276.370 8.685 ;
        RECT 295.410 8.315 295.690 8.685 ;
        RECT 413.700 8.430 417.060 8.570 ;
        RECT 276.160 4.070 276.300 8.315 ;
        RECT 295.480 6.700 295.620 8.315 ;
        RECT 392.930 7.635 393.210 8.005 ;
        RECT 411.330 7.635 411.610 8.005 ;
        RECT 393.000 7.470 393.140 7.635 ;
        RECT 314.730 6.955 315.010 7.325 ;
        RECT 334.510 6.955 334.790 7.325 ;
        RECT 392.940 7.150 393.200 7.470 ;
        RECT 295.880 6.700 296.140 6.790 ;
        RECT 295.480 6.560 296.140 6.700 ;
        RECT 295.880 6.470 296.140 6.560 ;
        RECT 314.800 4.750 314.940 6.955 ;
        RECT 334.580 6.110 334.720 6.955 ;
        RECT 334.520 5.790 334.780 6.110 ;
        RECT 411.400 5.850 411.540 7.635 ;
        RECT 413.700 6.530 413.840 8.430 ;
        RECT 416.920 7.890 417.060 8.430 ;
        RECT 554.000 8.430 556.900 8.570 ;
        RECT 416.920 7.750 417.980 7.890 ;
        RECT 417.840 7.210 417.980 7.750 ;
        RECT 504.780 7.580 506.300 7.720 ;
        RECT 504.780 7.325 504.920 7.580 ;
        RECT 418.230 7.210 418.510 7.325 ;
        RECT 417.840 7.070 418.510 7.210 ;
        RECT 418.230 6.955 418.510 7.070 ;
        RECT 504.710 6.955 504.990 7.325 ;
        RECT 506.160 7.210 506.300 7.580 ;
        RECT 554.000 7.325 554.140 8.430 ;
        RECT 556.760 8.150 556.900 8.430 ;
        RECT 556.700 7.830 556.960 8.150 ;
        RECT 506.550 7.210 506.830 7.325 ;
        RECT 506.160 7.070 506.830 7.210 ;
        RECT 506.550 6.955 506.830 7.070 ;
        RECT 513.910 7.210 514.190 7.325 ;
        RECT 515.290 7.210 515.570 7.325 ;
        RECT 513.910 7.070 515.570 7.210 ;
        RECT 513.910 6.955 514.190 7.070 ;
        RECT 515.290 6.955 515.570 7.070 ;
        RECT 553.930 6.955 554.210 7.325 ;
        RECT 559.910 6.955 560.190 7.325 ;
        RECT 603.150 7.210 603.430 7.325 ;
        RECT 604.530 7.210 604.810 7.325 ;
        RECT 603.150 7.070 604.810 7.210 ;
        RECT 603.150 6.955 603.430 7.070 ;
        RECT 604.530 6.955 604.810 7.070 ;
        RECT 638.570 6.955 638.850 7.325 ;
        RECT 701.130 6.955 701.410 7.325 ;
        RECT 706.190 7.210 706.470 7.325 ;
        RECT 707.570 7.210 707.850 7.325 ;
        RECT 706.190 7.070 707.850 7.210 ;
        RECT 706.190 6.955 706.470 7.070 ;
        RECT 707.570 6.955 707.850 7.070 ;
        RECT 757.710 7.210 757.990 7.325 ;
        RECT 759.090 7.210 759.370 7.325 ;
        RECT 757.710 7.070 759.370 7.210 ;
        RECT 757.710 6.955 757.990 7.070 ;
        RECT 759.090 6.955 759.370 7.070 ;
        RECT 789.910 6.955 790.190 7.325 ;
        RECT 412.320 6.390 413.840 6.530 ;
        RECT 412.320 5.850 412.460 6.390 ;
        RECT 559.980 6.110 560.120 6.955 ;
        RECT 638.640 6.360 638.780 6.955 ;
        RECT 642.720 6.360 642.980 6.450 ;
        RECT 638.640 6.220 642.980 6.360 ;
        RECT 642.720 6.130 642.980 6.220 ;
        RECT 411.400 5.710 412.460 5.850 ;
        RECT 559.920 5.790 560.180 6.110 ;
        RECT 701.200 5.770 701.340 6.955 ;
        RECT 789.980 5.850 790.120 6.955 ;
        RECT 790.370 5.850 790.650 5.965 ;
        RECT 701.140 5.450 701.400 5.770 ;
        RECT 789.980 5.710 790.650 5.850 ;
        RECT 790.370 5.595 790.650 5.710 ;
        RECT 792.210 5.595 792.490 5.965 ;
        RECT 835.850 5.850 836.130 9.000 ;
        RECT 834.600 5.770 836.130 5.850 ;
        RECT 802.800 5.680 803.060 5.770 ;
        RECT 805.100 5.680 805.360 5.770 ;
        RECT 792.220 5.450 792.480 5.595 ;
        RECT 802.800 5.540 805.360 5.680 ;
        RECT 802.800 5.450 803.060 5.540 ;
        RECT 805.100 5.450 805.360 5.540 ;
        RECT 834.540 5.710 836.130 5.770 ;
        RECT 834.540 5.450 834.800 5.710 ;
        RECT 835.850 5.000 836.130 5.710 ;
        RECT 314.740 4.430 315.000 4.750 ;
        RECT 276.100 3.750 276.360 4.070 ;
        RECT 234.700 3.070 234.960 3.390 ;
        RECT 234.760 2.400 234.900 3.070 ;
        RECT 234.550 -4.800 235.110 2.400 ;
      LAYER via2 ;
        RECT 276.090 8.360 276.370 8.640 ;
        RECT 295.410 8.360 295.690 8.640 ;
        RECT 392.930 7.680 393.210 7.960 ;
        RECT 411.330 7.680 411.610 7.960 ;
        RECT 314.730 7.000 315.010 7.280 ;
        RECT 334.510 7.000 334.790 7.280 ;
        RECT 418.230 7.000 418.510 7.280 ;
        RECT 504.710 7.000 504.990 7.280 ;
        RECT 506.550 7.000 506.830 7.280 ;
        RECT 513.910 7.000 514.190 7.280 ;
        RECT 515.290 7.000 515.570 7.280 ;
        RECT 553.930 7.000 554.210 7.280 ;
        RECT 559.910 7.000 560.190 7.280 ;
        RECT 603.150 7.000 603.430 7.280 ;
        RECT 604.530 7.000 604.810 7.280 ;
        RECT 638.570 7.000 638.850 7.280 ;
        RECT 701.130 7.000 701.410 7.280 ;
        RECT 706.190 7.000 706.470 7.280 ;
        RECT 707.570 7.000 707.850 7.280 ;
        RECT 757.710 7.000 757.990 7.280 ;
        RECT 759.090 7.000 759.370 7.280 ;
        RECT 789.910 7.000 790.190 7.280 ;
        RECT 790.370 5.640 790.650 5.920 ;
        RECT 792.210 5.640 792.490 5.920 ;
      LAYER met3 ;
        RECT 276.065 8.650 276.395 8.665 ;
        RECT 295.385 8.650 295.715 8.665 ;
        RECT 276.065 8.350 295.715 8.650 ;
        RECT 276.065 8.335 276.395 8.350 ;
        RECT 295.385 8.335 295.715 8.350 ;
        RECT 392.905 7.970 393.235 7.985 ;
        RECT 411.305 7.970 411.635 7.985 ;
        RECT 392.905 7.670 411.635 7.970 ;
        RECT 392.905 7.655 393.235 7.670 ;
        RECT 411.305 7.655 411.635 7.670 ;
        RECT 314.705 7.290 315.035 7.305 ;
        RECT 334.485 7.290 334.815 7.305 ;
        RECT 314.705 6.990 334.815 7.290 ;
        RECT 314.705 6.975 315.035 6.990 ;
        RECT 334.485 6.975 334.815 6.990 ;
        RECT 418.205 7.290 418.535 7.305 ;
        RECT 504.685 7.290 505.015 7.305 ;
        RECT 418.205 6.990 456.010 7.290 ;
        RECT 418.205 6.975 418.535 6.990 ;
        RECT 455.710 6.610 456.010 6.990 ;
        RECT 460.310 6.990 505.015 7.290 ;
        RECT 460.310 6.610 460.610 6.990 ;
        RECT 504.685 6.975 505.015 6.990 ;
        RECT 506.525 7.290 506.855 7.305 ;
        RECT 513.885 7.290 514.215 7.305 ;
        RECT 506.525 6.990 514.215 7.290 ;
        RECT 506.525 6.975 506.855 6.990 ;
        RECT 513.885 6.975 514.215 6.990 ;
        RECT 515.265 7.290 515.595 7.305 ;
        RECT 553.905 7.290 554.235 7.305 ;
        RECT 515.265 6.990 554.235 7.290 ;
        RECT 515.265 6.975 515.595 6.990 ;
        RECT 553.905 6.975 554.235 6.990 ;
        RECT 559.885 7.290 560.215 7.305 ;
        RECT 603.125 7.290 603.455 7.305 ;
        RECT 559.885 6.990 603.455 7.290 ;
        RECT 559.885 6.975 560.215 6.990 ;
        RECT 603.125 6.975 603.455 6.990 ;
        RECT 604.505 7.290 604.835 7.305 ;
        RECT 638.545 7.290 638.875 7.305 ;
        RECT 604.505 6.990 638.875 7.290 ;
        RECT 604.505 6.975 604.835 6.990 ;
        RECT 638.545 6.975 638.875 6.990 ;
        RECT 701.105 7.290 701.435 7.305 ;
        RECT 706.165 7.290 706.495 7.305 ;
        RECT 701.105 6.990 706.495 7.290 ;
        RECT 701.105 6.975 701.435 6.990 ;
        RECT 706.165 6.975 706.495 6.990 ;
        RECT 707.545 7.290 707.875 7.305 ;
        RECT 757.685 7.290 758.015 7.305 ;
        RECT 707.545 6.990 758.015 7.290 ;
        RECT 707.545 6.975 707.875 6.990 ;
        RECT 757.685 6.975 758.015 6.990 ;
        RECT 759.065 7.290 759.395 7.305 ;
        RECT 789.885 7.300 790.215 7.305 ;
        RECT 787.790 7.290 788.170 7.300 ;
        RECT 789.630 7.290 790.215 7.300 ;
        RECT 759.065 6.990 788.170 7.290 ;
        RECT 789.430 6.990 790.215 7.290 ;
        RECT 759.065 6.975 759.395 6.990 ;
        RECT 787.790 6.980 788.170 6.990 ;
        RECT 789.630 6.980 790.215 6.990 ;
        RECT 789.885 6.975 790.215 6.980 ;
        RECT 455.710 6.310 460.610 6.610 ;
        RECT 790.345 5.930 790.675 5.945 ;
        RECT 792.185 5.930 792.515 5.945 ;
        RECT 790.345 5.630 792.515 5.930 ;
        RECT 790.345 5.615 790.675 5.630 ;
        RECT 792.185 5.615 792.515 5.630 ;
      LAYER via3 ;
        RECT 787.820 6.980 788.140 7.300 ;
        RECT 789.660 6.980 789.980 7.300 ;
      LAYER met4 ;
        RECT 787.815 7.290 788.145 7.305 ;
        RECT 789.655 7.290 789.985 7.305 ;
        RECT 787.815 6.990 789.985 7.290 ;
        RECT 787.815 6.975 788.145 6.990 ;
        RECT 789.655 6.975 789.985 6.990 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2610.645 3396.345 2610.815 3401.955 ;
        RECT 2809.365 3396.345 2809.535 3401.615 ;
        RECT 2.905 77.265 3.075 120.275 ;
        RECT 26.825 7.225 27.455 7.395 ;
      LAYER mcon ;
        RECT 2610.645 3401.785 2610.815 3401.955 ;
        RECT 2809.365 3401.445 2809.535 3401.615 ;
        RECT 2.905 120.105 3.075 120.275 ;
        RECT 27.285 7.225 27.455 7.395 ;
      LAYER met1 ;
        RECT 2610.570 3401.940 2610.890 3402.000 ;
        RECT 2610.375 3401.800 2610.890 3401.940 ;
        RECT 2610.570 3401.740 2610.890 3401.800 ;
        RECT 2809.290 3401.600 2809.610 3401.660 ;
        RECT 2809.290 3401.460 2809.805 3401.600 ;
        RECT 2809.290 3401.400 2809.610 3401.460 ;
        RECT 2610.585 3396.500 2610.875 3396.545 ;
        RECT 2809.305 3396.500 2809.595 3396.545 ;
        RECT 2610.585 3396.360 2809.595 3396.500 ;
        RECT 2610.585 3396.315 2610.875 3396.360 ;
        RECT 2809.305 3396.315 2809.595 3396.360 ;
        RECT 2.845 120.260 3.135 120.305 ;
        RECT 7.430 120.260 7.750 120.320 ;
        RECT 2.845 120.120 7.750 120.260 ;
        RECT 2.845 120.075 3.135 120.120 ;
        RECT 7.430 120.060 7.750 120.120 ;
        RECT 2.845 77.420 3.135 77.465 ;
        RECT 9.730 77.420 10.050 77.480 ;
        RECT 2.845 77.280 10.050 77.420 ;
        RECT 2.845 77.235 3.135 77.280 ;
        RECT 9.730 77.220 10.050 77.280 ;
        RECT 17.550 7.380 17.870 7.440 ;
        RECT 26.765 7.380 27.055 7.425 ;
        RECT 17.550 7.240 27.055 7.380 ;
        RECT 17.550 7.180 17.870 7.240 ;
        RECT 26.765 7.195 27.055 7.240 ;
        RECT 27.225 7.380 27.515 7.425 ;
        RECT 34.110 7.380 34.430 7.440 ;
        RECT 27.225 7.240 34.430 7.380 ;
        RECT 27.225 7.195 27.515 7.240 ;
        RECT 34.110 7.180 34.430 7.240 ;
      LAYER via ;
        RECT 2610.600 3401.740 2610.860 3402.000 ;
        RECT 2809.320 3401.400 2809.580 3401.660 ;
        RECT 7.460 120.060 7.720 120.320 ;
        RECT 9.760 77.220 10.020 77.480 ;
        RECT 17.580 7.180 17.840 7.440 ;
        RECT 34.140 7.180 34.400 7.440 ;
      LAYER met2 ;
        RECT 2609.150 3401.770 2609.430 3405.000 ;
        RECT 2610.600 3401.770 2610.860 3402.030 ;
        RECT 2609.150 3401.710 2610.860 3401.770 ;
        RECT 2609.150 3401.630 2610.800 3401.710 ;
        RECT 2609.150 3401.000 2609.430 3401.630 ;
        RECT 2809.310 3401.515 2809.590 3401.885 ;
        RECT 2809.320 3401.370 2809.580 3401.515 ;
        RECT 7.450 128.675 7.730 129.045 ;
        RECT 7.520 120.350 7.660 128.675 ;
        RECT 7.460 120.030 7.720 120.350 ;
        RECT 9.760 77.420 10.020 77.510 ;
        RECT 9.760 77.280 11.800 77.420 ;
        RECT 9.760 77.190 10.020 77.280 ;
        RECT 11.660 75.720 11.800 77.280 ;
        RECT 11.660 75.580 17.780 75.720 ;
        RECT 17.640 7.470 17.780 75.580 ;
        RECT 34.130 8.315 34.410 8.685 ;
        RECT 56.210 8.315 56.490 8.685 ;
        RECT 34.200 7.470 34.340 8.315 ;
        RECT 17.580 7.150 17.840 7.470 ;
        RECT 34.140 7.150 34.400 7.470 ;
        RECT 56.280 2.400 56.420 8.315 ;
        RECT 56.070 -4.800 56.630 2.400 ;
      LAYER via2 ;
        RECT 2809.310 3401.560 2809.590 3401.840 ;
        RECT 7.450 128.720 7.730 129.000 ;
        RECT 34.130 8.360 34.410 8.640 ;
        RECT 56.210 8.360 56.490 8.640 ;
      LAYER met3 ;
        RECT 2809.285 3401.850 2809.615 3401.865 ;
        RECT 2811.790 3401.850 2812.170 3401.860 ;
        RECT 2809.285 3401.550 2812.170 3401.850 ;
        RECT 2809.285 3401.535 2809.615 3401.550 ;
        RECT 2811.790 3401.540 2812.170 3401.550 ;
        RECT 4.870 129.010 5.250 129.020 ;
        RECT 7.425 129.010 7.755 129.025 ;
        RECT 4.870 128.710 7.755 129.010 ;
        RECT 4.870 128.700 5.250 128.710 ;
        RECT 7.425 128.695 7.755 128.710 ;
        RECT 34.105 8.650 34.435 8.665 ;
        RECT 56.185 8.650 56.515 8.665 ;
        RECT 34.105 8.350 56.515 8.650 ;
        RECT 34.105 8.335 34.435 8.350 ;
        RECT 56.185 8.335 56.515 8.350 ;
      LAYER via3 ;
        RECT 2811.820 3401.540 2812.140 3401.860 ;
        RECT 4.900 128.700 5.220 129.020 ;
      LAYER met4 ;
        RECT 2811.815 3401.535 2812.145 3401.865 ;
        RECT 2811.830 172.290 2812.130 3401.535 ;
        RECT 4.470 171.110 5.650 172.290 ;
        RECT 2811.390 171.110 2812.570 172.290 ;
        RECT 4.910 129.025 5.210 171.110 ;
        RECT 4.895 128.695 5.225 129.025 ;
      LAYER met5 ;
        RECT 4.260 170.900 2812.780 172.500 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 244.865 8.245 245.955 8.415 ;
        RECT 214.505 3.825 214.675 8.075 ;
        RECT 244.865 7.905 245.035 8.245 ;
        RECT 245.785 6.885 245.955 8.245 ;
        RECT 266.485 1.105 266.655 7.055 ;
        RECT 512.125 6.715 512.295 7.735 ;
        RECT 511.205 6.545 512.295 6.715 ;
        RECT 663.005 5.355 663.175 7.055 ;
        RECT 677.265 6.545 697.675 6.715 ;
        RECT 663.005 5.185 674.215 5.355 ;
        RECT 674.045 4.505 674.215 5.185 ;
        RECT 676.345 4.335 676.515 4.675 ;
        RECT 677.265 4.335 677.435 6.545 ;
        RECT 697.505 6.375 697.675 6.545 ;
        RECT 703.945 6.545 704.575 6.715 ;
        RECT 1074.245 6.545 1074.415 8.075 ;
        RECT 1093.565 7.225 1094.655 7.395 ;
        RECT 1093.565 6.885 1093.735 7.225 ;
        RECT 703.945 6.375 704.115 6.545 ;
        RECT 697.505 6.205 704.115 6.375 ;
        RECT 704.405 6.205 704.575 6.545 ;
        RECT 1094.485 6.035 1094.655 7.225 ;
        RECT 1094.485 5.865 1119.955 6.035 ;
        RECT 1119.785 5.355 1119.955 5.865 ;
        RECT 1122.085 5.865 1125.935 6.035 ;
        RECT 1122.085 5.355 1122.255 5.865 ;
        RECT 1125.765 5.525 1125.935 5.865 ;
        RECT 1119.785 5.185 1122.255 5.355 ;
        RECT 676.345 4.165 677.435 4.335 ;
        RECT 1469.385 4.165 1469.555 7.395 ;
        RECT 2641.005 4.505 2641.175 8.415 ;
      LAYER mcon ;
        RECT 214.505 7.905 214.675 8.075 ;
        RECT 2641.005 8.245 2641.175 8.415 ;
        RECT 1074.245 7.905 1074.415 8.075 ;
        RECT 512.125 7.565 512.295 7.735 ;
        RECT 266.485 6.885 266.655 7.055 ;
        RECT 663.005 6.885 663.175 7.055 ;
        RECT 676.345 4.505 676.515 4.675 ;
        RECT 1469.385 7.225 1469.555 7.395 ;
      LAYER met1 ;
        RECT 2545.250 8.400 2545.570 8.460 ;
        RECT 2640.945 8.400 2641.235 8.445 ;
        RECT 2545.250 8.260 2641.235 8.400 ;
        RECT 2545.250 8.200 2545.570 8.260 ;
        RECT 2640.945 8.215 2641.235 8.260 ;
        RECT 214.445 8.060 214.735 8.105 ;
        RECT 244.805 8.060 245.095 8.105 ;
        RECT 214.445 7.920 245.095 8.060 ;
        RECT 214.445 7.875 214.735 7.920 ;
        RECT 244.805 7.875 245.095 7.920 ;
        RECT 1072.330 8.060 1072.650 8.120 ;
        RECT 1074.185 8.060 1074.475 8.105 ;
        RECT 1072.330 7.920 1074.475 8.060 ;
        RECT 1072.330 7.860 1072.650 7.920 ;
        RECT 1074.185 7.875 1074.475 7.920 ;
        RECT 1369.950 8.060 1370.270 8.120 ;
        RECT 1401.230 8.060 1401.550 8.120 ;
        RECT 1369.950 7.920 1401.550 8.060 ;
        RECT 1369.950 7.860 1370.270 7.920 ;
        RECT 1401.230 7.860 1401.550 7.920 ;
        RECT 2217.270 8.060 2217.590 8.120 ;
        RECT 2266.030 8.060 2266.350 8.120 ;
        RECT 2217.270 7.920 2266.350 8.060 ;
        RECT 2217.270 7.860 2217.590 7.920 ;
        RECT 2266.030 7.860 2266.350 7.920 ;
        RECT 512.065 7.720 512.355 7.765 ;
        RECT 516.650 7.720 516.970 7.780 ;
        RECT 512.065 7.580 516.970 7.720 ;
        RECT 512.065 7.535 512.355 7.580 ;
        RECT 516.650 7.520 516.970 7.580 ;
        RECT 1451.830 7.380 1452.150 7.440 ;
        RECT 1469.325 7.380 1469.615 7.425 ;
        RECT 1451.830 7.240 1469.615 7.380 ;
        RECT 1451.830 7.180 1452.150 7.240 ;
        RECT 1469.325 7.195 1469.615 7.240 ;
        RECT 1546.130 7.380 1546.450 7.440 ;
        RECT 1549.810 7.380 1550.130 7.440 ;
        RECT 1546.130 7.240 1550.130 7.380 ;
        RECT 1546.130 7.180 1546.450 7.240 ;
        RECT 1549.810 7.180 1550.130 7.240 ;
        RECT 245.725 7.040 246.015 7.085 ;
        RECT 266.425 7.040 266.715 7.085 ;
        RECT 662.945 7.040 663.235 7.085 ;
        RECT 1093.505 7.040 1093.795 7.085 ;
        RECT 245.725 6.900 266.715 7.040 ;
        RECT 245.725 6.855 246.015 6.900 ;
        RECT 266.425 6.855 266.715 6.900 ;
        RECT 659.340 6.900 663.235 7.040 ;
        RECT 511.130 6.700 511.450 6.760 ;
        RECT 510.935 6.560 511.450 6.700 ;
        RECT 511.130 6.500 511.450 6.560 ;
        RECT 646.370 6.700 646.690 6.760 ;
        RECT 659.340 6.700 659.480 6.900 ;
        RECT 662.945 6.855 663.235 6.900 ;
        RECT 1092.660 6.900 1093.795 7.040 ;
        RECT 646.370 6.560 659.480 6.700 ;
        RECT 1074.185 6.700 1074.475 6.745 ;
        RECT 1092.660 6.700 1092.800 6.900 ;
        RECT 1093.505 6.855 1093.795 6.900 ;
        RECT 1074.185 6.560 1092.800 6.700 ;
        RECT 646.370 6.500 646.690 6.560 ;
        RECT 1074.185 6.515 1074.475 6.560 ;
        RECT 516.650 6.360 516.970 6.420 ;
        RECT 533.210 6.360 533.530 6.420 ;
        RECT 516.650 6.220 533.530 6.360 ;
        RECT 516.650 6.160 516.970 6.220 ;
        RECT 533.210 6.160 533.530 6.220 ;
        RECT 704.345 6.360 704.635 6.405 ;
        RECT 713.990 6.360 714.310 6.420 ;
        RECT 704.345 6.220 714.310 6.360 ;
        RECT 704.345 6.175 704.635 6.220 ;
        RECT 713.990 6.160 714.310 6.220 ;
        RECT 1125.705 5.680 1125.995 5.725 ;
        RECT 1126.150 5.680 1126.470 5.740 ;
        RECT 1125.705 5.540 1126.470 5.680 ;
        RECT 1125.705 5.495 1125.995 5.540 ;
        RECT 1126.150 5.480 1126.470 5.540 ;
        RECT 673.985 4.660 674.275 4.705 ;
        RECT 676.285 4.660 676.575 4.705 ;
        RECT 673.985 4.520 676.575 4.660 ;
        RECT 673.985 4.475 674.275 4.520 ;
        RECT 676.285 4.475 676.575 4.520 ;
        RECT 2640.945 4.660 2641.235 4.705 ;
        RECT 2694.750 4.660 2695.070 4.720 ;
        RECT 2640.945 4.520 2695.070 4.660 ;
        RECT 2640.945 4.475 2641.235 4.520 ;
        RECT 2694.750 4.460 2695.070 4.520 ;
        RECT 1469.325 4.320 1469.615 4.365 ;
        RECT 1533.710 4.320 1534.030 4.380 ;
        RECT 1469.325 4.180 1534.030 4.320 ;
        RECT 1469.325 4.135 1469.615 4.180 ;
        RECT 1533.710 4.120 1534.030 4.180 ;
        RECT 210.290 3.980 210.610 4.040 ;
        RECT 214.445 3.980 214.735 4.025 ;
        RECT 210.290 3.840 214.735 3.980 ;
        RECT 210.290 3.780 210.610 3.840 ;
        RECT 214.445 3.795 214.735 3.840 ;
        RECT 2381.950 3.640 2382.270 3.700 ;
        RECT 2450.950 3.640 2451.270 3.700 ;
        RECT 2381.950 3.500 2451.270 3.640 ;
        RECT 2381.950 3.440 2382.270 3.500 ;
        RECT 2450.950 3.440 2451.270 3.500 ;
        RECT 1308.770 2.620 1309.090 2.680 ;
        RECT 1327.170 2.620 1327.490 2.680 ;
        RECT 1308.770 2.480 1327.490 2.620 ;
        RECT 1308.770 2.420 1309.090 2.480 ;
        RECT 1327.170 2.420 1327.490 2.480 ;
        RECT 266.425 1.260 266.715 1.305 ;
        RECT 277.910 1.260 278.230 1.320 ;
        RECT 266.425 1.120 278.230 1.260 ;
        RECT 266.425 1.075 266.715 1.120 ;
        RECT 277.910 1.060 278.230 1.120 ;
      LAYER via ;
        RECT 2545.280 8.200 2545.540 8.460 ;
        RECT 1072.360 7.860 1072.620 8.120 ;
        RECT 1369.980 7.860 1370.240 8.120 ;
        RECT 1401.260 7.860 1401.520 8.120 ;
        RECT 2217.300 7.860 2217.560 8.120 ;
        RECT 2266.060 7.860 2266.320 8.120 ;
        RECT 516.680 7.520 516.940 7.780 ;
        RECT 1451.860 7.180 1452.120 7.440 ;
        RECT 1546.160 7.180 1546.420 7.440 ;
        RECT 1549.840 7.180 1550.100 7.440 ;
        RECT 511.160 6.500 511.420 6.760 ;
        RECT 646.400 6.500 646.660 6.760 ;
        RECT 516.680 6.160 516.940 6.420 ;
        RECT 533.240 6.160 533.500 6.420 ;
        RECT 714.020 6.160 714.280 6.420 ;
        RECT 1126.180 5.480 1126.440 5.740 ;
        RECT 2694.780 4.460 2695.040 4.720 ;
        RECT 1533.740 4.120 1534.000 4.380 ;
        RECT 210.320 3.780 210.580 4.040 ;
        RECT 2381.980 3.440 2382.240 3.700 ;
        RECT 2450.980 3.440 2451.240 3.700 ;
        RECT 1308.800 2.420 1309.060 2.680 ;
        RECT 1327.200 2.420 1327.460 2.680 ;
        RECT 277.940 1.060 278.200 1.320 ;
      LAYER met2 ;
        RECT 1342.370 8.570 1342.650 8.685 ;
        RECT 1327.720 8.430 1342.650 8.570 ;
        RECT 1044.820 8.260 1057.380 8.400 ;
        RECT 516.680 7.490 516.940 7.810 ;
        RECT 459.630 7.210 459.910 7.325 ;
        RECT 459.630 7.070 460.300 7.210 ;
        RECT 459.630 6.955 459.910 7.070 ;
        RECT 460.160 6.530 460.300 7.070 ;
        RECT 461.010 6.530 461.290 6.645 ;
        RECT 460.160 6.390 461.290 6.530 ;
        RECT 511.160 6.530 511.420 6.790 ;
        RECT 511.610 6.530 511.890 6.645 ;
        RECT 511.160 6.470 511.890 6.530 ;
        RECT 511.220 6.390 511.890 6.470 ;
        RECT 516.740 6.450 516.880 7.490 ;
        RECT 646.400 6.470 646.660 6.790 ;
        RECT 461.010 6.275 461.290 6.390 ;
        RECT 511.610 6.275 511.890 6.390 ;
        RECT 516.680 6.130 516.940 6.450 ;
        RECT 533.240 6.130 533.500 6.450 ;
        RECT 210.310 5.595 210.590 5.965 ;
        RECT 291.730 5.595 292.010 5.965 ;
        RECT 210.380 4.070 210.520 5.595 ;
        RECT 210.320 3.750 210.580 4.070 ;
        RECT 291.800 3.980 291.940 5.595 ;
        RECT 533.300 5.000 533.440 6.130 ;
        RECT 533.300 4.860 533.900 5.000 ;
        RECT 287.200 3.840 291.940 3.980 ;
        RECT 79.280 2.820 80.340 2.960 ;
        RECT 79.280 1.885 79.420 2.820 ;
        RECT 80.200 2.400 80.340 2.820 ;
        RECT 79.210 1.515 79.490 1.885 ;
        RECT 79.990 -4.800 80.550 2.400 ;
        RECT 277.940 1.030 278.200 1.350 ;
        RECT 287.200 1.205 287.340 3.840 ;
        RECT 533.760 2.450 533.900 4.860 ;
        RECT 536.910 3.555 537.190 3.925 ;
        RECT 645.470 3.810 645.750 3.925 ;
        RECT 646.460 3.810 646.600 6.470 ;
        RECT 714.020 6.130 714.280 6.450 ;
        RECT 645.470 3.670 646.600 3.810 ;
        RECT 645.470 3.555 645.750 3.670 ;
        RECT 536.980 2.450 537.120 3.555 ;
        RECT 714.080 3.300 714.220 6.130 ;
        RECT 1044.820 5.340 1044.960 8.260 ;
        RECT 1057.240 7.210 1057.380 8.260 ;
        RECT 1072.360 7.830 1072.620 8.150 ;
        RECT 1060.850 7.210 1061.130 7.325 ;
        RECT 1057.240 7.070 1061.130 7.210 ;
        RECT 1060.850 6.955 1061.130 7.070 ;
        RECT 1071.890 7.210 1072.170 7.325 ;
        RECT 1072.420 7.210 1072.560 7.830 ;
        RECT 1071.890 7.070 1072.560 7.210 ;
        RECT 1071.890 6.955 1072.170 7.070 ;
        RECT 1126.170 6.275 1126.450 6.645 ;
        RECT 1046.130 5.595 1046.410 5.965 ;
        RECT 1126.240 5.770 1126.380 6.275 ;
        RECT 1046.200 5.340 1046.340 5.595 ;
        RECT 1126.180 5.450 1126.440 5.770 ;
        RECT 1044.820 5.200 1046.340 5.340 ;
        RECT 1279.350 4.915 1279.630 5.285 ;
        RECT 1279.420 3.810 1279.560 4.915 ;
        RECT 1279.810 3.810 1280.090 3.925 ;
        RECT 748.120 3.670 753.320 3.810 ;
        RECT 1279.420 3.670 1280.090 3.810 ;
        RECT 714.080 3.160 718.360 3.300 ;
        RECT 718.220 3.130 718.360 3.160 ;
        RECT 718.220 2.990 723.420 3.130 ;
        RECT 533.760 2.310 537.120 2.450 ;
        RECT 723.280 1.770 723.420 2.990 ;
        RECT 748.120 2.960 748.260 3.670 ;
        RECT 724.200 2.820 748.260 2.960 ;
        RECT 724.200 1.770 724.340 2.820 ;
        RECT 723.280 1.630 724.340 1.770 ;
        RECT 753.180 1.770 753.320 3.670 ;
        RECT 1279.810 3.555 1280.090 3.670 ;
        RECT 1304.190 3.810 1304.470 3.925 ;
        RECT 1304.190 3.670 1309.000 3.810 ;
        RECT 1304.190 3.555 1304.470 3.670 ;
        RECT 757.250 3.130 757.530 3.245 ;
        RECT 756.400 2.990 757.530 3.130 ;
        RECT 756.400 1.770 756.540 2.990 ;
        RECT 757.250 2.875 757.530 2.990 ;
        RECT 1308.860 2.710 1309.000 3.670 ;
        RECT 1327.720 3.130 1327.860 8.430 ;
        RECT 1342.370 8.315 1342.650 8.430 ;
        RECT 1401.780 8.430 1405.600 8.570 ;
        RECT 1369.980 7.830 1370.240 8.150 ;
        RECT 1401.260 8.060 1401.520 8.150 ;
        RECT 1401.780 8.060 1401.920 8.430 ;
        RECT 1401.260 7.920 1401.920 8.060 ;
        RECT 1401.260 7.830 1401.520 7.920 ;
        RECT 1367.670 6.955 1367.950 7.325 ;
        RECT 1367.740 5.850 1367.880 6.955 ;
        RECT 1370.040 5.850 1370.180 7.830 ;
        RECT 1404.930 6.530 1405.210 6.645 ;
        RECT 1405.460 6.530 1405.600 8.430 ;
        RECT 1549.830 8.315 1550.110 8.685 ;
        RECT 2180.030 8.315 2180.310 8.685 ;
        RECT 2217.290 8.315 2217.570 8.685 ;
        RECT 1536.030 7.635 1536.310 8.005 ;
        RECT 1546.150 7.635 1546.430 8.005 ;
        RECT 1451.860 7.150 1452.120 7.470 ;
        RECT 1404.930 6.390 1405.600 6.530 ;
        RECT 1404.930 6.275 1405.210 6.390 ;
        RECT 1451.920 5.965 1452.060 7.150 ;
        RECT 1367.740 5.710 1370.180 5.850 ;
        RECT 1451.850 5.595 1452.130 5.965 ;
        RECT 1533.740 4.320 1534.000 4.410 ;
        RECT 1536.100 4.320 1536.240 7.635 ;
        RECT 1546.220 7.470 1546.360 7.635 ;
        RECT 1549.900 7.470 1550.040 8.315 ;
        RECT 1829.970 7.635 1830.250 8.005 ;
        RECT 1546.160 7.150 1546.420 7.470 ;
        RECT 1549.840 7.150 1550.100 7.470 ;
        RECT 1830.040 6.645 1830.180 7.635 ;
        RECT 2180.100 6.645 2180.240 8.315 ;
        RECT 2217.360 8.150 2217.500 8.315 ;
        RECT 2545.280 8.170 2545.540 8.490 ;
        RECT 2217.300 7.830 2217.560 8.150 ;
        RECT 2266.060 8.005 2266.320 8.150 ;
        RECT 2266.050 7.635 2266.330 8.005 ;
        RECT 2312.970 7.635 2313.250 8.005 ;
        RECT 2313.040 6.645 2313.180 7.635 ;
        RECT 1829.970 6.275 1830.250 6.645 ;
        RECT 2180.030 6.275 2180.310 6.645 ;
        RECT 2312.970 6.275 2313.250 6.645 ;
        RECT 2381.970 6.275 2382.250 6.645 ;
        RECT 1533.740 4.180 1536.240 4.320 ;
        RECT 1533.740 4.090 1534.000 4.180 ;
        RECT 2382.040 3.730 2382.180 6.275 ;
        RECT 2381.980 3.410 2382.240 3.730 ;
        RECT 2450.980 3.410 2451.240 3.730 ;
        RECT 2451.040 3.245 2451.180 3.410 ;
        RECT 2545.340 3.245 2545.480 8.170 ;
        RECT 2796.890 7.635 2797.170 8.005 ;
        RECT 2829.090 7.890 2829.370 8.005 ;
        RECT 2830.870 7.890 2831.150 9.000 ;
        RECT 2829.090 7.750 2831.150 7.890 ;
        RECT 2829.090 7.635 2829.370 7.750 ;
        RECT 2694.780 4.430 2695.040 4.750 ;
        RECT 1327.260 2.990 1327.860 3.130 ;
        RECT 1327.260 2.710 1327.400 2.990 ;
        RECT 2450.970 2.875 2451.250 3.245 ;
        RECT 2545.270 2.875 2545.550 3.245 ;
        RECT 1308.800 2.390 1309.060 2.710 ;
        RECT 1327.200 2.390 1327.460 2.710 ;
        RECT 2694.840 1.885 2694.980 4.430 ;
        RECT 2796.960 1.885 2797.100 7.635 ;
        RECT 2830.870 5.000 2831.150 7.750 ;
        RECT 753.180 1.630 756.540 1.770 ;
        RECT 2694.770 1.515 2695.050 1.885 ;
        RECT 2796.890 1.515 2797.170 1.885 ;
        RECT 280.690 1.090 280.970 1.205 ;
        RECT 278.000 0.580 278.140 1.030 ;
        RECT 280.300 0.950 280.970 1.090 ;
        RECT 280.300 0.580 280.440 0.950 ;
        RECT 280.690 0.835 280.970 0.950 ;
        RECT 287.130 0.835 287.410 1.205 ;
        RECT 278.000 0.440 280.440 0.580 ;
      LAYER via2 ;
        RECT 459.630 7.000 459.910 7.280 ;
        RECT 461.010 6.320 461.290 6.600 ;
        RECT 511.610 6.320 511.890 6.600 ;
        RECT 210.310 5.640 210.590 5.920 ;
        RECT 291.730 5.640 292.010 5.920 ;
        RECT 79.210 1.560 79.490 1.840 ;
        RECT 536.910 3.600 537.190 3.880 ;
        RECT 645.470 3.600 645.750 3.880 ;
        RECT 1060.850 7.000 1061.130 7.280 ;
        RECT 1071.890 7.000 1072.170 7.280 ;
        RECT 1126.170 6.320 1126.450 6.600 ;
        RECT 1046.130 5.640 1046.410 5.920 ;
        RECT 1279.350 4.960 1279.630 5.240 ;
        RECT 1279.810 3.600 1280.090 3.880 ;
        RECT 1304.190 3.600 1304.470 3.880 ;
        RECT 757.250 2.920 757.530 3.200 ;
        RECT 1342.370 8.360 1342.650 8.640 ;
        RECT 1367.670 7.000 1367.950 7.280 ;
        RECT 1404.930 6.320 1405.210 6.600 ;
        RECT 1549.830 8.360 1550.110 8.640 ;
        RECT 2180.030 8.360 2180.310 8.640 ;
        RECT 2217.290 8.360 2217.570 8.640 ;
        RECT 1536.030 7.680 1536.310 7.960 ;
        RECT 1546.150 7.680 1546.430 7.960 ;
        RECT 1451.850 5.640 1452.130 5.920 ;
        RECT 1829.970 7.680 1830.250 7.960 ;
        RECT 2266.050 7.680 2266.330 7.960 ;
        RECT 2312.970 7.680 2313.250 7.960 ;
        RECT 1829.970 6.320 1830.250 6.600 ;
        RECT 2180.030 6.320 2180.310 6.600 ;
        RECT 2312.970 6.320 2313.250 6.600 ;
        RECT 2381.970 6.320 2382.250 6.600 ;
        RECT 2796.890 7.680 2797.170 7.960 ;
        RECT 2829.090 7.680 2829.370 7.960 ;
        RECT 2450.970 2.920 2451.250 3.200 ;
        RECT 2545.270 2.920 2545.550 3.200 ;
        RECT 2694.770 1.560 2695.050 1.840 ;
        RECT 2796.890 1.560 2797.170 1.840 ;
        RECT 280.690 0.880 280.970 1.160 ;
        RECT 287.130 0.880 287.410 1.160 ;
      LAYER met3 ;
        RECT 412.430 8.650 412.810 8.660 ;
        RECT 1226.630 8.650 1227.010 8.660 ;
        RECT 384.870 8.350 412.810 8.650 ;
        RECT 382.070 7.970 382.450 7.980 ;
        RECT 384.870 7.970 385.170 8.350 ;
        RECT 412.430 8.340 412.810 8.350 ;
        RECT 1192.630 8.350 1227.010 8.650 ;
        RECT 382.070 7.670 385.170 7.970 ;
        RECT 415.190 7.970 415.570 7.980 ;
        RECT 415.190 7.670 456.930 7.970 ;
        RECT 382.070 7.660 382.450 7.670 ;
        RECT 415.190 7.660 415.570 7.670 ;
        RECT 456.630 7.290 456.930 7.670 ;
        RECT 459.605 7.290 459.935 7.305 ;
        RECT 456.630 6.990 459.935 7.290 ;
        RECT 459.605 6.975 459.935 6.990 ;
        RECT 798.830 7.290 799.210 7.300 ;
        RECT 806.190 7.290 806.570 7.300 ;
        RECT 798.830 6.990 806.570 7.290 ;
        RECT 798.830 6.980 799.210 6.990 ;
        RECT 806.190 6.980 806.570 6.990 ;
        RECT 1060.825 7.290 1061.155 7.305 ;
        RECT 1071.865 7.290 1072.195 7.305 ;
        RECT 1192.630 7.290 1192.930 8.350 ;
        RECT 1226.630 8.340 1227.010 8.350 ;
        RECT 1342.345 8.650 1342.675 8.665 ;
        RECT 1343.470 8.650 1343.850 8.660 ;
        RECT 1342.345 8.350 1343.850 8.650 ;
        RECT 1342.345 8.335 1342.675 8.350 ;
        RECT 1343.470 8.340 1343.850 8.350 ;
        RECT 1549.805 8.650 1550.135 8.665 ;
        RECT 1552.310 8.650 1552.690 8.660 ;
        RECT 1549.805 8.350 1552.690 8.650 ;
        RECT 1549.805 8.335 1550.135 8.350 ;
        RECT 1552.310 8.340 1552.690 8.350 ;
        RECT 2180.005 8.650 2180.335 8.665 ;
        RECT 2217.265 8.650 2217.595 8.665 ;
        RECT 2180.005 8.350 2217.595 8.650 ;
        RECT 2180.005 8.335 2180.335 8.350 ;
        RECT 2217.265 8.335 2217.595 8.350 ;
        RECT 1536.005 7.970 1536.335 7.985 ;
        RECT 1546.125 7.970 1546.455 7.985 ;
        RECT 1536.005 7.670 1546.455 7.970 ;
        RECT 1536.005 7.655 1536.335 7.670 ;
        RECT 1546.125 7.655 1546.455 7.670 ;
        RECT 1771.270 7.970 1771.650 7.980 ;
        RECT 1829.945 7.970 1830.275 7.985 ;
        RECT 1771.270 7.670 1830.275 7.970 ;
        RECT 1771.270 7.660 1771.650 7.670 ;
        RECT 1829.945 7.655 1830.275 7.670 ;
        RECT 2266.025 7.970 2266.355 7.985 ;
        RECT 2312.945 7.970 2313.275 7.985 ;
        RECT 2266.025 7.670 2313.275 7.970 ;
        RECT 2266.025 7.655 2266.355 7.670 ;
        RECT 2312.945 7.655 2313.275 7.670 ;
        RECT 2796.865 7.970 2797.195 7.985 ;
        RECT 2829.065 7.970 2829.395 7.985 ;
        RECT 2796.865 7.670 2829.395 7.970 ;
        RECT 2796.865 7.655 2797.195 7.670 ;
        RECT 2829.065 7.655 2829.395 7.670 ;
        RECT 1367.645 7.300 1367.975 7.305 ;
        RECT 1367.390 7.290 1367.975 7.300 ;
        RECT 1060.825 6.990 1072.195 7.290 ;
        RECT 1060.825 6.975 1061.155 6.990 ;
        RECT 1071.865 6.975 1072.195 6.990 ;
        RECT 1128.230 6.990 1192.930 7.290 ;
        RECT 1367.190 6.990 1367.975 7.290 ;
        RECT 460.985 6.610 461.315 6.625 ;
        RECT 511.585 6.620 511.915 6.625 ;
        RECT 482.350 6.610 482.730 6.620 ;
        RECT 460.985 6.310 482.730 6.610 ;
        RECT 460.985 6.295 461.315 6.310 ;
        RECT 482.350 6.300 482.730 6.310 ;
        RECT 501.670 6.610 502.050 6.620 ;
        RECT 506.270 6.610 506.650 6.620 ;
        RECT 501.670 6.310 506.650 6.610 ;
        RECT 501.670 6.300 502.050 6.310 ;
        RECT 506.270 6.300 506.650 6.310 ;
        RECT 511.585 6.610 512.170 6.620 ;
        RECT 809.870 6.610 810.250 6.620 ;
        RECT 817.230 6.610 817.610 6.620 ;
        RECT 511.585 6.310 512.370 6.610 ;
        RECT 809.870 6.310 817.610 6.610 ;
        RECT 511.585 6.300 512.170 6.310 ;
        RECT 809.870 6.300 810.250 6.310 ;
        RECT 817.230 6.300 817.610 6.310 ;
        RECT 1126.145 6.610 1126.475 6.625 ;
        RECT 1128.230 6.610 1128.530 6.990 ;
        RECT 1367.390 6.980 1367.975 6.990 ;
        RECT 1367.645 6.975 1367.975 6.980 ;
        RECT 1404.905 6.620 1405.235 6.625 ;
        RECT 1126.145 6.310 1128.530 6.610 ;
        RECT 1239.510 6.610 1239.890 6.620 ;
        RECT 1252.390 6.610 1252.770 6.620 ;
        RECT 1404.905 6.610 1405.490 6.620 ;
        RECT 1239.510 6.310 1252.770 6.610 ;
        RECT 1404.680 6.310 1405.490 6.610 ;
        RECT 511.585 6.295 511.915 6.300 ;
        RECT 1126.145 6.295 1126.475 6.310 ;
        RECT 1239.510 6.300 1239.890 6.310 ;
        RECT 1252.390 6.300 1252.770 6.310 ;
        RECT 1404.905 6.300 1405.490 6.310 ;
        RECT 1829.945 6.610 1830.275 6.625 ;
        RECT 1862.350 6.610 1862.730 6.620 ;
        RECT 1829.945 6.310 1862.730 6.610 ;
        RECT 1404.905 6.295 1405.235 6.300 ;
        RECT 1829.945 6.295 1830.275 6.310 ;
        RECT 1862.350 6.300 1862.730 6.310 ;
        RECT 2096.950 6.610 2097.330 6.620 ;
        RECT 2180.005 6.610 2180.335 6.625 ;
        RECT 2096.950 6.310 2180.335 6.610 ;
        RECT 2096.950 6.300 2097.330 6.310 ;
        RECT 2180.005 6.295 2180.335 6.310 ;
        RECT 2312.945 6.610 2313.275 6.625 ;
        RECT 2381.945 6.610 2382.275 6.625 ;
        RECT 2312.945 6.310 2382.275 6.610 ;
        RECT 2312.945 6.295 2313.275 6.310 ;
        RECT 2381.945 6.295 2382.275 6.310 ;
        RECT 197.150 5.930 197.530 5.940 ;
        RECT 210.285 5.930 210.615 5.945 ;
        RECT 197.150 5.630 210.615 5.930 ;
        RECT 197.150 5.620 197.530 5.630 ;
        RECT 210.285 5.615 210.615 5.630 ;
        RECT 291.705 5.930 292.035 5.945 ;
        RECT 1046.105 5.940 1046.435 5.945 ;
        RECT 1451.825 5.940 1452.155 5.945 ;
        RECT 302.950 5.930 303.330 5.940 ;
        RECT 291.705 5.630 303.330 5.930 ;
        RECT 291.705 5.615 292.035 5.630 ;
        RECT 302.950 5.620 303.330 5.630 ;
        RECT 1046.105 5.930 1046.690 5.940 ;
        RECT 1451.825 5.930 1452.410 5.940 ;
        RECT 1046.105 5.630 1046.890 5.930 ;
        RECT 1451.825 5.630 1452.610 5.930 ;
        RECT 1046.105 5.620 1046.690 5.630 ;
        RECT 1451.825 5.620 1452.410 5.630 ;
        RECT 1046.105 5.615 1046.435 5.620 ;
        RECT 1451.825 5.615 1452.155 5.620 ;
        RECT 318.590 5.250 318.970 5.260 ;
        RECT 364.590 5.250 364.970 5.260 ;
        RECT 318.590 4.950 364.970 5.250 ;
        RECT 318.590 4.940 318.970 4.950 ;
        RECT 364.590 4.940 364.970 4.950 ;
        RECT 1267.110 5.250 1267.490 5.260 ;
        RECT 1279.325 5.250 1279.655 5.265 ;
        RECT 1267.110 4.950 1279.655 5.250 ;
        RECT 1267.110 4.940 1267.490 4.950 ;
        RECT 1279.325 4.935 1279.655 4.950 ;
        RECT 536.885 3.890 537.215 3.905 ;
        RECT 538.470 3.890 538.850 3.900 ;
        RECT 536.885 3.590 538.850 3.890 ;
        RECT 536.885 3.575 537.215 3.590 ;
        RECT 538.470 3.580 538.850 3.590 ;
        RECT 614.830 3.890 615.210 3.900 ;
        RECT 645.445 3.890 645.775 3.905 ;
        RECT 614.830 3.590 645.775 3.890 ;
        RECT 614.830 3.580 615.210 3.590 ;
        RECT 645.445 3.575 645.775 3.590 ;
        RECT 1279.785 3.890 1280.115 3.905 ;
        RECT 1304.165 3.900 1304.495 3.905 ;
        RECT 1291.030 3.890 1291.410 3.900 ;
        RECT 1303.910 3.890 1304.495 3.900 ;
        RECT 1279.785 3.590 1291.410 3.890 ;
        RECT 1303.710 3.590 1304.495 3.890 ;
        RECT 1279.785 3.575 1280.115 3.590 ;
        RECT 1291.030 3.580 1291.410 3.590 ;
        RECT 1303.910 3.580 1304.495 3.590 ;
        RECT 1304.165 3.575 1304.495 3.580 ;
        RECT 757.225 3.210 757.555 3.225 ;
        RECT 781.350 3.210 781.730 3.220 ;
        RECT 757.225 2.910 781.730 3.210 ;
        RECT 757.225 2.895 757.555 2.910 ;
        RECT 781.350 2.900 781.730 2.910 ;
        RECT 2450.945 3.210 2451.275 3.225 ;
        RECT 2545.245 3.210 2545.575 3.225 ;
        RECT 2450.945 2.910 2545.575 3.210 ;
        RECT 2450.945 2.895 2451.275 2.910 ;
        RECT 2545.245 2.895 2545.575 2.910 ;
        RECT 74.790 1.850 75.170 1.860 ;
        RECT 79.185 1.850 79.515 1.865 ;
        RECT 74.790 1.550 79.515 1.850 ;
        RECT 74.790 1.540 75.170 1.550 ;
        RECT 79.185 1.535 79.515 1.550 ;
        RECT 2694.745 1.850 2695.075 1.865 ;
        RECT 2796.865 1.850 2797.195 1.865 ;
        RECT 2694.745 1.550 2797.195 1.850 ;
        RECT 2694.745 1.535 2695.075 1.550 ;
        RECT 2796.865 1.535 2797.195 1.550 ;
        RECT 280.665 1.170 280.995 1.185 ;
        RECT 287.105 1.170 287.435 1.185 ;
        RECT 280.665 0.870 287.435 1.170 ;
        RECT 280.665 0.855 280.995 0.870 ;
        RECT 287.105 0.855 287.435 0.870 ;
      LAYER via3 ;
        RECT 382.100 7.660 382.420 7.980 ;
        RECT 412.460 8.340 412.780 8.660 ;
        RECT 415.220 7.660 415.540 7.980 ;
        RECT 798.860 6.980 799.180 7.300 ;
        RECT 806.220 6.980 806.540 7.300 ;
        RECT 1226.660 8.340 1226.980 8.660 ;
        RECT 1343.500 8.340 1343.820 8.660 ;
        RECT 1552.340 8.340 1552.660 8.660 ;
        RECT 1771.300 7.660 1771.620 7.980 ;
        RECT 482.380 6.300 482.700 6.620 ;
        RECT 501.700 6.300 502.020 6.620 ;
        RECT 506.300 6.300 506.620 6.620 ;
        RECT 511.820 6.300 512.140 6.620 ;
        RECT 809.900 6.300 810.220 6.620 ;
        RECT 817.260 6.300 817.580 6.620 ;
        RECT 1367.420 6.980 1367.740 7.300 ;
        RECT 1239.540 6.300 1239.860 6.620 ;
        RECT 1252.420 6.300 1252.740 6.620 ;
        RECT 1405.140 6.300 1405.460 6.620 ;
        RECT 1862.380 6.300 1862.700 6.620 ;
        RECT 2096.980 6.300 2097.300 6.620 ;
        RECT 197.180 5.620 197.500 5.940 ;
        RECT 302.980 5.620 303.300 5.940 ;
        RECT 1046.340 5.620 1046.660 5.940 ;
        RECT 1452.060 5.620 1452.380 5.940 ;
        RECT 318.620 4.940 318.940 5.260 ;
        RECT 364.620 4.940 364.940 5.260 ;
        RECT 1267.140 4.940 1267.460 5.260 ;
        RECT 538.500 3.580 538.820 3.900 ;
        RECT 614.860 3.580 615.180 3.900 ;
        RECT 1291.060 3.580 1291.380 3.900 ;
        RECT 1303.940 3.580 1304.260 3.900 ;
        RECT 781.380 2.900 781.700 3.220 ;
        RECT 74.820 1.540 75.140 1.860 ;
      LAYER met4 ;
        RECT 74.390 14.710 75.570 15.890 ;
        RECT 144.310 14.710 145.490 15.890 ;
        RECT 1555.590 14.710 1556.770 15.890 ;
        RECT 1770.870 14.710 1772.050 15.890 ;
        RECT 1862.180 14.710 1863.360 15.890 ;
        RECT 2096.550 14.710 2097.730 15.890 ;
        RECT 74.830 1.865 75.130 14.710 ;
        RECT 144.750 2.290 145.050 14.710 ;
        RECT 1556.030 12.050 1556.330 14.710 ;
        RECT 1552.350 11.750 1556.330 12.050 ;
        RECT 1552.350 8.665 1552.650 11.750 ;
        RECT 412.455 8.650 412.785 8.665 ;
        RECT 1226.655 8.650 1226.985 8.665 ;
        RECT 1343.495 8.650 1343.825 8.665 ;
        RECT 412.455 8.350 414.610 8.650 ;
        RECT 412.455 8.335 412.785 8.350 ;
        RECT 382.095 7.970 382.425 7.985 ;
        RECT 378.430 7.670 382.425 7.970 ;
        RECT 414.310 7.970 414.610 8.350 ;
        RECT 1226.655 8.350 1237.090 8.650 ;
        RECT 1226.655 8.335 1226.985 8.350 ;
        RECT 415.215 7.970 415.545 7.985 ;
        RECT 414.310 7.670 415.545 7.970 ;
        RECT 1236.790 7.970 1237.090 8.350 ;
        RECT 1343.495 8.350 1360.370 8.650 ;
        RECT 1343.495 8.335 1343.825 8.350 ;
        RECT 1236.790 7.670 1239.850 7.970 ;
        RECT 197.175 5.615 197.505 5.945 ;
        RECT 302.975 5.615 303.305 5.945 ;
        RECT 197.190 2.290 197.490 5.615 ;
        RECT 302.990 5.250 303.290 5.615 ;
        RECT 318.615 5.250 318.945 5.265 ;
        RECT 302.990 4.950 318.945 5.250 ;
        RECT 318.615 4.935 318.945 4.950 ;
        RECT 364.615 4.935 364.945 5.265 ;
        RECT 364.630 4.570 364.930 4.935 ;
        RECT 378.430 4.570 378.730 7.670 ;
        RECT 382.095 7.655 382.425 7.670 ;
        RECT 415.215 7.655 415.545 7.670 ;
        RECT 506.310 6.990 512.130 7.290 ;
        RECT 506.310 6.625 506.610 6.990 ;
        RECT 511.830 6.625 512.130 6.990 ;
        RECT 798.855 6.975 799.185 7.305 ;
        RECT 806.215 6.975 806.545 7.305 ;
        RECT 482.375 6.295 482.705 6.625 ;
        RECT 501.695 6.610 502.025 6.625 ;
        RECT 489.750 6.310 502.025 6.610 ;
        RECT 482.390 5.930 482.690 6.295 ;
        RECT 489.750 5.930 490.050 6.310 ;
        RECT 501.695 6.295 502.025 6.310 ;
        RECT 506.295 6.295 506.625 6.625 ;
        RECT 511.815 6.295 512.145 6.625 ;
        RECT 482.390 5.630 490.050 5.930 ;
        RECT 364.630 4.270 378.730 4.570 ;
        RECT 538.495 3.890 538.825 3.905 ;
        RECT 614.855 3.890 615.185 3.905 ;
        RECT 798.870 3.890 799.170 6.975 ;
        RECT 806.230 5.250 806.530 6.975 ;
        RECT 1239.550 6.625 1239.850 7.670 ;
        RECT 1360.070 7.290 1360.370 8.350 ;
        RECT 1552.335 8.335 1552.665 8.665 ;
        RECT 1771.310 7.985 1771.610 14.710 ;
        RECT 1362.830 7.670 1367.730 7.970 ;
        RECT 1362.830 7.290 1363.130 7.670 ;
        RECT 1367.430 7.305 1367.730 7.670 ;
        RECT 1771.295 7.655 1771.625 7.985 ;
        RECT 1360.070 6.990 1363.130 7.290 ;
        RECT 1367.415 6.975 1367.745 7.305 ;
        RECT 1862.390 6.625 1862.690 14.710 ;
        RECT 2096.990 6.625 2097.290 14.710 ;
        RECT 809.895 6.295 810.225 6.625 ;
        RECT 817.255 6.295 817.585 6.625 ;
        RECT 1239.535 6.295 1239.865 6.625 ;
        RECT 1252.415 6.295 1252.745 6.625 ;
        RECT 1405.135 6.610 1405.465 6.625 ;
        RECT 1405.135 6.310 1408.210 6.610 ;
        RECT 1405.135 6.295 1405.465 6.310 ;
        RECT 809.910 5.250 810.210 6.295 ;
        RECT 817.270 5.930 817.570 6.295 ;
        RECT 1046.335 5.930 1046.665 5.945 ;
        RECT 817.270 5.630 823.090 5.930 ;
        RECT 806.230 4.950 810.210 5.250 ;
        RECT 538.495 3.590 540.650 3.890 ;
        RECT 538.495 3.575 538.825 3.590 ;
        RECT 74.815 1.535 75.145 1.865 ;
        RECT 144.310 1.110 145.490 2.290 ;
        RECT 196.750 1.110 197.930 2.290 ;
        RECT 540.350 1.850 540.650 3.590 ;
        RECT 612.110 3.590 615.185 3.890 ;
        RECT 612.110 1.850 612.410 3.590 ;
        RECT 614.855 3.575 615.185 3.590 ;
        RECT 781.390 3.590 799.170 3.890 ;
        RECT 781.390 3.225 781.690 3.590 ;
        RECT 781.375 2.895 781.705 3.225 ;
        RECT 822.790 2.290 823.090 5.630 ;
        RECT 992.760 5.630 1030.090 5.930 ;
        RECT 992.760 5.250 993.060 5.630 ;
        RECT 991.150 4.950 993.060 5.250 ;
        RECT 991.150 4.570 991.450 4.950 ;
        RECT 990.460 4.270 991.450 4.570 ;
        RECT 990.460 3.890 990.760 4.270 ;
        RECT 845.790 3.590 851.610 3.890 ;
        RECT 845.790 2.290 846.090 3.590 ;
        RECT 540.350 1.550 567.330 1.850 ;
        RECT 567.030 1.170 567.330 1.550 ;
        RECT 576.230 1.550 612.410 1.850 ;
        RECT 576.230 1.170 576.530 1.550 ;
        RECT 567.030 0.870 576.530 1.170 ;
        RECT 822.350 1.110 823.530 2.290 ;
        RECT 845.350 1.110 846.530 2.290 ;
        RECT 851.310 1.850 851.610 3.590 ;
        RECT 983.790 3.590 990.760 3.890 ;
        RECT 1029.790 3.890 1030.090 5.630 ;
        RECT 1043.590 5.630 1046.665 5.930 ;
        RECT 1252.430 5.930 1252.730 6.295 ;
        RECT 1252.430 5.630 1264.690 5.930 ;
        RECT 1043.590 3.890 1043.890 5.630 ;
        RECT 1046.335 5.615 1046.665 5.630 ;
        RECT 1264.390 5.250 1264.690 5.630 ;
        RECT 1267.135 5.250 1267.465 5.265 ;
        RECT 1264.390 4.950 1267.465 5.250 ;
        RECT 1267.135 4.935 1267.465 4.950 ;
        RECT 1302.110 4.270 1304.250 4.570 ;
        RECT 1029.790 3.590 1043.890 3.890 ;
        RECT 1291.055 3.890 1291.385 3.905 ;
        RECT 1291.055 3.590 1296.890 3.890 ;
        RECT 983.790 2.290 984.090 3.590 ;
        RECT 1291.055 3.575 1291.385 3.590 ;
        RECT 1296.590 3.210 1296.890 3.590 ;
        RECT 1302.110 3.210 1302.410 4.270 ;
        RECT 1303.950 3.905 1304.250 4.270 ;
        RECT 1303.935 3.575 1304.265 3.905 ;
        RECT 1296.590 2.910 1302.410 3.210 ;
        RECT 1407.910 2.290 1408.210 6.310 ;
        RECT 1862.375 6.295 1862.705 6.625 ;
        RECT 2096.975 6.295 2097.305 6.625 ;
        RECT 1452.055 5.615 1452.385 5.945 ;
        RECT 1452.070 2.290 1452.370 5.615 ;
        RECT 881.230 1.850 882.410 2.290 ;
        RECT 851.310 1.550 882.410 1.850 ;
        RECT 881.230 1.110 882.410 1.550 ;
        RECT 983.350 1.110 984.530 2.290 ;
        RECT 1407.470 1.110 1408.650 2.290 ;
        RECT 1451.630 1.110 1452.810 2.290 ;
      LAYER met5 ;
        RECT 1665.780 21.300 1772.260 22.900 ;
        RECT 74.180 17.900 145.700 19.500 ;
        RECT 74.180 14.500 75.780 17.900 ;
        RECT 144.100 14.500 145.700 17.900 ;
        RECT 1555.380 17.900 1643.460 19.500 ;
        RECT 1555.380 14.500 1556.980 17.900 ;
        RECT 1641.860 16.100 1643.460 17.900 ;
        RECT 1665.780 16.100 1667.380 21.300 ;
        RECT 1641.860 14.500 1667.380 16.100 ;
        RECT 1770.660 14.500 1772.260 21.300 ;
        RECT 1948.220 21.300 2016.060 22.900 ;
        RECT 1948.220 19.500 1949.820 21.300 ;
        RECT 1861.970 17.900 1943.380 19.500 ;
        RECT 1861.970 14.500 1863.570 17.900 ;
        RECT 1941.780 16.100 1943.380 17.900 ;
        RECT 1947.300 17.900 1949.820 19.500 ;
        RECT 2014.460 19.500 2016.060 21.300 ;
        RECT 2014.460 17.900 2097.940 19.500 ;
        RECT 1947.300 16.100 1948.900 17.900 ;
        RECT 1941.780 14.500 1948.900 16.100 ;
        RECT 2096.340 14.500 2097.940 17.900 ;
        RECT 144.100 0.900 198.140 2.500 ;
        RECT 822.140 0.900 846.740 2.500 ;
        RECT 881.020 0.900 984.740 2.500 ;
        RECT 1407.260 0.900 1453.020 2.500 ;
    END
  END wbs_sel_i[1]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2803.845 3395.665 2804.015 3401.615 ;
      LAYER mcon ;
        RECT 2803.845 3401.445 2804.015 3401.615 ;
      LAYER met1 ;
        RECT 2803.770 3401.600 2804.090 3401.660 ;
        RECT 2803.575 3401.460 2804.090 3401.600 ;
        RECT 2803.770 3401.400 2804.090 3401.460 ;
        RECT 2803.785 3395.820 2804.075 3395.865 ;
        RECT 2863.570 3395.820 2863.890 3395.880 ;
        RECT 2803.785 3395.680 2863.890 3395.820 ;
        RECT 2803.785 3395.635 2804.075 3395.680 ;
        RECT 2863.570 3395.620 2863.890 3395.680 ;
        RECT 5.590 4.320 5.910 4.380 ;
        RECT 24.910 4.320 25.230 4.380 ;
        RECT 5.590 4.180 25.230 4.320 ;
        RECT 5.590 4.120 5.910 4.180 ;
        RECT 24.910 4.120 25.230 4.180 ;
      LAYER via ;
        RECT 2803.800 3401.400 2804.060 3401.660 ;
        RECT 2863.600 3395.620 2863.860 3395.880 ;
        RECT 5.620 4.120 5.880 4.380 ;
        RECT 24.940 4.120 25.200 4.380 ;
      LAYER met2 ;
        RECT 2803.790 3401.515 2804.070 3401.885 ;
        RECT 2803.800 3401.370 2804.060 3401.515 ;
        RECT 2863.600 3395.590 2863.860 3395.910 ;
        RECT 2863.660 3337.285 2863.800 3395.590 ;
        RECT 2863.590 3336.915 2863.870 3337.285 ;
        RECT 6.070 134.115 6.350 134.485 ;
        RECT 6.140 52.090 6.280 134.115 ;
        RECT 5.680 51.950 6.280 52.090 ;
        RECT 5.680 4.410 5.820 51.950 ;
        RECT 5.620 4.090 5.880 4.410 ;
        RECT 24.940 4.090 25.200 4.410 ;
        RECT 25.000 3.810 25.140 4.090 ;
        RECT 25.000 3.670 26.520 3.810 ;
        RECT 26.380 2.400 26.520 3.670 ;
        RECT 26.170 -4.800 26.730 2.400 ;
      LAYER via2 ;
        RECT 2803.790 3401.560 2804.070 3401.840 ;
        RECT 2863.590 3336.960 2863.870 3337.240 ;
        RECT 6.070 134.160 6.350 134.440 ;
      LAYER met3 ;
        RECT 2803.765 3401.860 2804.095 3401.865 ;
        RECT 2803.510 3401.850 2804.095 3401.860 ;
        RECT 2803.310 3401.550 2804.095 3401.850 ;
        RECT 2803.510 3401.540 2804.095 3401.550 ;
        RECT 2803.765 3401.535 2804.095 3401.540 ;
        RECT 2851.000 3337.250 2855.000 3337.640 ;
        RECT 2863.565 3337.250 2863.895 3337.265 ;
        RECT 2851.000 3337.040 2863.895 3337.250 ;
        RECT 2854.300 3336.950 2863.895 3337.040 ;
        RECT 2863.565 3336.935 2863.895 3336.950 ;
        RECT 6.045 134.450 6.375 134.465 ;
        RECT 6.710 134.450 7.090 134.460 ;
        RECT 6.045 134.150 7.090 134.450 ;
        RECT 6.045 134.135 6.375 134.150 ;
        RECT 6.710 134.140 7.090 134.150 ;
      LAYER via3 ;
        RECT 2803.540 3401.540 2803.860 3401.860 ;
        RECT 6.740 134.140 7.060 134.460 ;
      LAYER met4 ;
        RECT 2803.535 3401.535 2803.865 3401.865 ;
        RECT 2803.550 3303.250 2803.850 3401.535 ;
        RECT 2801.710 3302.950 2803.850 3303.250 ;
        RECT 2801.710 3269.250 2802.010 3302.950 ;
        RECT 2801.710 3268.950 2804.770 3269.250 ;
        RECT 2804.470 3106.050 2804.770 3268.950 ;
        RECT 2802.630 3105.750 2804.770 3106.050 ;
        RECT 2802.630 3075.450 2802.930 3105.750 ;
        RECT 2802.630 3075.150 2803.850 3075.450 ;
        RECT 2803.550 3041.450 2803.850 3075.150 ;
        RECT 2801.710 3041.150 2803.850 3041.450 ;
        RECT 2801.710 3024.450 2802.010 3041.150 ;
        RECT 2801.710 3024.150 2802.930 3024.450 ;
        RECT 2802.630 2970.050 2802.930 3024.150 ;
        RECT 2802.630 2969.750 2803.850 2970.050 ;
        RECT 2803.550 2895.250 2803.850 2969.750 ;
        RECT 2802.630 2894.950 2803.850 2895.250 ;
        RECT 2802.630 2813.650 2802.930 2894.950 ;
        RECT 2802.630 2813.350 2803.850 2813.650 ;
        RECT 2803.550 2769.450 2803.850 2813.350 ;
        RECT 2803.550 2769.150 2804.770 2769.450 ;
        RECT 2804.470 2718.450 2804.770 2769.150 ;
        RECT 2801.710 2718.150 2804.770 2718.450 ;
        RECT 2801.710 2674.250 2802.010 2718.150 ;
        RECT 2801.710 2673.950 2803.850 2674.250 ;
        RECT 2803.550 2650.450 2803.850 2673.950 ;
        RECT 2802.630 2650.150 2803.850 2650.450 ;
        RECT 2802.630 2623.250 2802.930 2650.150 ;
        RECT 2801.710 2622.950 2802.930 2623.250 ;
        RECT 2801.710 2599.450 2802.010 2622.950 ;
        RECT 2801.710 2599.150 2802.930 2599.450 ;
        RECT 2802.630 2592.650 2802.930 2599.150 ;
        RECT 2800.790 2592.350 2802.930 2592.650 ;
        RECT 2800.790 2548.450 2801.090 2592.350 ;
        RECT 2800.790 2548.150 2803.850 2548.450 ;
        RECT 2803.550 2524.650 2803.850 2548.150 ;
        RECT 2803.550 2524.350 2804.770 2524.650 ;
        RECT 2804.470 2477.050 2804.770 2524.350 ;
        RECT 2802.630 2476.750 2804.770 2477.050 ;
        RECT 2802.630 2426.050 2802.930 2476.750 ;
        RECT 2802.630 2425.750 2803.850 2426.050 ;
        RECT 2803.550 2402.250 2803.850 2425.750 ;
        RECT 2803.550 2401.950 2804.770 2402.250 ;
        RECT 2804.470 2354.650 2804.770 2401.950 ;
        RECT 2803.550 2354.350 2804.770 2354.650 ;
        RECT 2803.550 2256.050 2803.850 2354.350 ;
        RECT 2801.710 2255.750 2803.850 2256.050 ;
        RECT 2801.710 2228.850 2802.010 2255.750 ;
        RECT 2801.710 2228.550 2803.850 2228.850 ;
        RECT 2803.550 2184.650 2803.850 2228.550 ;
        RECT 2802.630 2184.350 2803.850 2184.650 ;
        RECT 2802.630 2143.850 2802.930 2184.350 ;
        RECT 2800.790 2143.550 2802.930 2143.850 ;
        RECT 2800.790 2092.850 2801.090 2143.550 ;
        RECT 2800.790 2092.550 2803.850 2092.850 ;
        RECT 2803.550 2062.250 2803.850 2092.550 ;
        RECT 2803.550 2061.950 2804.770 2062.250 ;
        RECT 2804.470 2038.450 2804.770 2061.950 ;
        RECT 2801.710 2038.150 2804.770 2038.450 ;
        RECT 2801.710 2014.650 2802.010 2038.150 ;
        RECT 2801.710 2014.350 2802.930 2014.650 ;
        RECT 2802.630 1990.850 2802.930 2014.350 ;
        RECT 2802.630 1990.550 2803.850 1990.850 ;
        RECT 2803.550 1902.450 2803.850 1990.550 ;
        RECT 2798.950 1902.150 2803.850 1902.450 ;
        RECT 2798.950 1895.650 2799.250 1902.150 ;
        RECT 2798.950 1895.350 2801.090 1895.650 ;
        RECT 2800.790 1848.050 2801.090 1895.350 ;
        RECT 2800.790 1847.750 2802.930 1848.050 ;
        RECT 2802.630 1800.450 2802.930 1847.750 ;
        RECT 2802.630 1800.150 2803.850 1800.450 ;
        RECT 2803.550 1725.650 2803.850 1800.150 ;
        RECT 2803.550 1725.350 2804.770 1725.650 ;
        RECT 2804.470 1674.650 2804.770 1725.350 ;
        RECT 2803.550 1674.350 2804.770 1674.650 ;
        RECT 2803.550 1667.850 2803.850 1674.350 ;
        RECT 2800.790 1667.550 2803.850 1667.850 ;
        RECT 2800.790 1627.050 2801.090 1667.550 ;
        RECT 2800.790 1626.750 2802.010 1627.050 ;
        RECT 2801.710 1620.250 2802.010 1626.750 ;
        RECT 2801.710 1619.950 2802.930 1620.250 ;
        RECT 2802.630 1616.850 2802.930 1619.950 ;
        RECT 2802.630 1616.550 2803.850 1616.850 ;
        RECT 2803.550 1531.850 2803.850 1616.550 ;
        RECT 2803.550 1531.550 2804.770 1531.850 ;
        RECT 2804.470 1453.650 2804.770 1531.550 ;
        RECT 2802.630 1453.350 2804.770 1453.650 ;
        RECT 2802.630 1433.250 2802.930 1453.350 ;
        RECT 2802.630 1432.950 2803.850 1433.250 ;
        RECT 2803.550 1416.250 2803.850 1432.950 ;
        RECT 2801.710 1415.950 2803.850 1416.250 ;
        RECT 2801.710 1361.850 2802.010 1415.950 ;
        RECT 2801.710 1361.550 2802.930 1361.850 ;
        RECT 2802.630 1321.050 2802.930 1361.550 ;
        RECT 2801.710 1320.750 2802.930 1321.050 ;
        RECT 2801.710 1314.250 2802.010 1320.750 ;
        RECT 2801.710 1313.950 2803.850 1314.250 ;
        RECT 2803.550 1270.050 2803.850 1313.950 ;
        RECT 2801.710 1269.750 2803.850 1270.050 ;
        RECT 2801.710 1168.050 2802.010 1269.750 ;
        RECT 2801.710 1167.750 2803.850 1168.050 ;
        RECT 2803.550 1140.850 2803.850 1167.750 ;
        RECT 2803.550 1140.550 2804.770 1140.850 ;
        RECT 2804.470 1117.050 2804.770 1140.550 ;
        RECT 2802.630 1116.750 2804.770 1117.050 ;
        RECT 2802.630 1079.650 2802.930 1116.750 ;
        RECT 2802.630 1079.350 2803.850 1079.650 ;
        RECT 2803.550 1072.850 2803.850 1079.350 ;
        RECT 2801.710 1072.550 2803.850 1072.850 ;
        RECT 2801.710 1035.450 2802.010 1072.550 ;
        RECT 2801.710 1035.150 2803.850 1035.450 ;
        RECT 2803.550 1025.250 2803.850 1035.150 ;
        RECT 2802.630 1024.950 2803.850 1025.250 ;
        RECT 2802.630 981.050 2802.930 1024.950 ;
        RECT 2801.710 980.750 2802.930 981.050 ;
        RECT 2801.710 950.450 2802.010 980.750 ;
        RECT 2801.710 950.150 2802.930 950.450 ;
        RECT 2802.630 936.850 2802.930 950.150 ;
        RECT 2801.710 936.550 2802.930 936.850 ;
        RECT 2801.710 930.050 2802.010 936.550 ;
        RECT 2801.710 929.750 2803.850 930.050 ;
        RECT 2803.550 882.450 2803.850 929.750 ;
        RECT 2803.550 882.150 2804.770 882.450 ;
        RECT 2804.470 834.850 2804.770 882.150 ;
        RECT 2802.630 834.550 2804.770 834.850 ;
        RECT 2802.630 783.850 2802.930 834.550 ;
        RECT 2802.630 783.550 2803.850 783.850 ;
        RECT 2803.550 760.050 2803.850 783.550 ;
        RECT 2803.550 759.750 2804.770 760.050 ;
        RECT 2804.470 712.450 2804.770 759.750 ;
        RECT 2803.550 712.150 2804.770 712.450 ;
        RECT 2803.550 658.050 2803.850 712.150 ;
        RECT 2803.550 657.750 2804.770 658.050 ;
        RECT 2804.470 641.050 2804.770 657.750 ;
        RECT 2803.550 640.750 2804.770 641.050 ;
        RECT 2803.550 613.850 2803.850 640.750 ;
        RECT 2803.550 613.550 2804.770 613.850 ;
        RECT 2804.470 566.250 2804.770 613.550 ;
        RECT 2803.550 565.950 2804.770 566.250 ;
        RECT 2803.550 545.850 2803.850 565.950 ;
        RECT 2803.550 545.550 2804.770 545.850 ;
        RECT 2804.470 522.050 2804.770 545.550 ;
        RECT 2803.550 521.750 2804.770 522.050 ;
        RECT 2803.550 518.650 2803.850 521.750 ;
        RECT 2802.630 518.350 2803.850 518.650 ;
        RECT 2802.630 498.250 2802.930 518.350 ;
        RECT 2802.630 497.950 2803.850 498.250 ;
        RECT 2803.550 491.450 2803.850 497.950 ;
        RECT 2800.790 491.150 2803.850 491.450 ;
        RECT 2800.790 454.050 2801.090 491.150 ;
        RECT 2800.790 453.750 2802.010 454.050 ;
        RECT 2801.710 382.650 2802.010 453.750 ;
        RECT 2801.710 382.350 2802.930 382.650 ;
        RECT 2802.630 348.650 2802.930 382.350 ;
        RECT 2802.630 348.350 2803.850 348.650 ;
        RECT 2803.550 273.850 2803.850 348.350 ;
        RECT 2801.710 273.550 2803.850 273.850 ;
        RECT 2801.710 250.050 2802.010 273.550 ;
        RECT 2801.710 249.750 2804.770 250.050 ;
        RECT 2804.470 226.250 2804.770 249.750 ;
        RECT 2802.630 225.950 2804.770 226.250 ;
        RECT 2802.630 202.450 2802.930 225.950 ;
        RECT 2802.630 202.150 2803.850 202.450 ;
        RECT 2803.550 145.090 2803.850 202.150 ;
        RECT 6.310 143.910 7.490 145.090 ;
        RECT 2803.110 143.910 2804.290 145.090 ;
        RECT 6.750 134.465 7.050 143.910 ;
        RECT 6.735 134.135 7.065 134.465 ;
      LAYER met5 ;
        RECT 6.100 143.700 2804.500 145.300 ;
    END
  END wbs_stb_i
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -14.580 -9.220 -11.580 3528.900 ;
        RECT 2931.200 -9.220 2934.200 3528.900 ;
      LAYER via4 ;
        RECT -13.670 3527.610 -12.490 3528.790 ;
        RECT -13.670 3526.010 -12.490 3527.190 ;
        RECT -13.670 3341.090 -12.490 3342.270 ;
        RECT -13.670 3339.490 -12.490 3340.670 ;
        RECT -13.670 3161.090 -12.490 3162.270 ;
        RECT -13.670 3159.490 -12.490 3160.670 ;
        RECT -13.670 2981.090 -12.490 2982.270 ;
        RECT -13.670 2979.490 -12.490 2980.670 ;
        RECT -13.670 2801.090 -12.490 2802.270 ;
        RECT -13.670 2799.490 -12.490 2800.670 ;
        RECT -13.670 2621.090 -12.490 2622.270 ;
        RECT -13.670 2619.490 -12.490 2620.670 ;
        RECT -13.670 2441.090 -12.490 2442.270 ;
        RECT -13.670 2439.490 -12.490 2440.670 ;
        RECT -13.670 2261.090 -12.490 2262.270 ;
        RECT -13.670 2259.490 -12.490 2260.670 ;
        RECT -13.670 2081.090 -12.490 2082.270 ;
        RECT -13.670 2079.490 -12.490 2080.670 ;
        RECT -13.670 1901.090 -12.490 1902.270 ;
        RECT -13.670 1899.490 -12.490 1900.670 ;
        RECT -13.670 1721.090 -12.490 1722.270 ;
        RECT -13.670 1719.490 -12.490 1720.670 ;
        RECT -13.670 1541.090 -12.490 1542.270 ;
        RECT -13.670 1539.490 -12.490 1540.670 ;
        RECT -13.670 1361.090 -12.490 1362.270 ;
        RECT -13.670 1359.490 -12.490 1360.670 ;
        RECT -13.670 1181.090 -12.490 1182.270 ;
        RECT -13.670 1179.490 -12.490 1180.670 ;
        RECT -13.670 1001.090 -12.490 1002.270 ;
        RECT -13.670 999.490 -12.490 1000.670 ;
        RECT -13.670 821.090 -12.490 822.270 ;
        RECT -13.670 819.490 -12.490 820.670 ;
        RECT -13.670 641.090 -12.490 642.270 ;
        RECT -13.670 639.490 -12.490 640.670 ;
        RECT -13.670 461.090 -12.490 462.270 ;
        RECT -13.670 459.490 -12.490 460.670 ;
        RECT -13.670 281.090 -12.490 282.270 ;
        RECT -13.670 279.490 -12.490 280.670 ;
        RECT -13.670 101.090 -12.490 102.270 ;
        RECT -13.670 99.490 -12.490 100.670 ;
        RECT -13.670 -7.510 -12.490 -6.330 ;
        RECT -13.670 -9.110 -12.490 -7.930 ;
        RECT 2932.110 3527.610 2933.290 3528.790 ;
        RECT 2932.110 3526.010 2933.290 3527.190 ;
        RECT 2932.110 3341.090 2933.290 3342.270 ;
        RECT 2932.110 3339.490 2933.290 3340.670 ;
        RECT 2932.110 3161.090 2933.290 3162.270 ;
        RECT 2932.110 3159.490 2933.290 3160.670 ;
        RECT 2932.110 2981.090 2933.290 2982.270 ;
        RECT 2932.110 2979.490 2933.290 2980.670 ;
        RECT 2932.110 2801.090 2933.290 2802.270 ;
        RECT 2932.110 2799.490 2933.290 2800.670 ;
        RECT 2932.110 2621.090 2933.290 2622.270 ;
        RECT 2932.110 2619.490 2933.290 2620.670 ;
        RECT 2932.110 2441.090 2933.290 2442.270 ;
        RECT 2932.110 2439.490 2933.290 2440.670 ;
        RECT 2932.110 2261.090 2933.290 2262.270 ;
        RECT 2932.110 2259.490 2933.290 2260.670 ;
        RECT 2932.110 2081.090 2933.290 2082.270 ;
        RECT 2932.110 2079.490 2933.290 2080.670 ;
        RECT 2932.110 1901.090 2933.290 1902.270 ;
        RECT 2932.110 1899.490 2933.290 1900.670 ;
        RECT 2932.110 1721.090 2933.290 1722.270 ;
        RECT 2932.110 1719.490 2933.290 1720.670 ;
        RECT 2932.110 1541.090 2933.290 1542.270 ;
        RECT 2932.110 1539.490 2933.290 1540.670 ;
        RECT 2932.110 1361.090 2933.290 1362.270 ;
        RECT 2932.110 1359.490 2933.290 1360.670 ;
        RECT 2932.110 1181.090 2933.290 1182.270 ;
        RECT 2932.110 1179.490 2933.290 1180.670 ;
        RECT 2932.110 1001.090 2933.290 1002.270 ;
        RECT 2932.110 999.490 2933.290 1000.670 ;
        RECT 2932.110 821.090 2933.290 822.270 ;
        RECT 2932.110 819.490 2933.290 820.670 ;
        RECT 2932.110 641.090 2933.290 642.270 ;
        RECT 2932.110 639.490 2933.290 640.670 ;
        RECT 2932.110 461.090 2933.290 462.270 ;
        RECT 2932.110 459.490 2933.290 460.670 ;
        RECT 2932.110 281.090 2933.290 282.270 ;
        RECT 2932.110 279.490 2933.290 280.670 ;
        RECT 2932.110 101.090 2933.290 102.270 ;
        RECT 2932.110 99.490 2933.290 100.670 ;
        RECT 2932.110 -7.510 2933.290 -6.330 ;
        RECT 2932.110 -9.110 2933.290 -7.930 ;
      LAYER met5 ;
        RECT -14.580 3528.900 -11.580 3528.910 ;
        RECT 2931.200 3528.900 2934.200 3528.910 ;
        RECT -14.580 3525.900 2934.200 3528.900 ;
        RECT -14.580 3525.890 -11.580 3525.900 ;
        RECT 2931.200 3525.890 2934.200 3525.900 ;
        RECT -14.580 3342.380 -11.580 3342.390 ;
        RECT 2931.200 3342.380 2934.200 3342.390 ;
        RECT -14.580 3339.380 2934.200 3342.380 ;
        RECT -14.580 3339.370 -11.580 3339.380 ;
        RECT 2931.200 3339.370 2934.200 3339.380 ;
        RECT -14.580 3162.380 -11.580 3162.390 ;
        RECT 2931.200 3162.380 2934.200 3162.390 ;
        RECT -14.580 3159.380 2934.200 3162.380 ;
        RECT -14.580 3159.370 -11.580 3159.380 ;
        RECT 2931.200 3159.370 2934.200 3159.380 ;
        RECT -14.580 2982.380 -11.580 2982.390 ;
        RECT 2931.200 2982.380 2934.200 2982.390 ;
        RECT -14.580 2979.380 2934.200 2982.380 ;
        RECT -14.580 2979.370 -11.580 2979.380 ;
        RECT 2931.200 2979.370 2934.200 2979.380 ;
        RECT -14.580 2802.380 -11.580 2802.390 ;
        RECT 2931.200 2802.380 2934.200 2802.390 ;
        RECT -14.580 2799.380 2934.200 2802.380 ;
        RECT -14.580 2799.370 -11.580 2799.380 ;
        RECT 2931.200 2799.370 2934.200 2799.380 ;
        RECT -14.580 2622.380 -11.580 2622.390 ;
        RECT 2931.200 2622.380 2934.200 2622.390 ;
        RECT -14.580 2619.380 2934.200 2622.380 ;
        RECT -14.580 2619.370 -11.580 2619.380 ;
        RECT 2931.200 2619.370 2934.200 2619.380 ;
        RECT -14.580 2442.380 -11.580 2442.390 ;
        RECT 2931.200 2442.380 2934.200 2442.390 ;
        RECT -14.580 2439.380 2934.200 2442.380 ;
        RECT -14.580 2439.370 -11.580 2439.380 ;
        RECT 2931.200 2439.370 2934.200 2439.380 ;
        RECT -14.580 2262.380 -11.580 2262.390 ;
        RECT 2931.200 2262.380 2934.200 2262.390 ;
        RECT -14.580 2259.380 2934.200 2262.380 ;
        RECT -14.580 2259.370 -11.580 2259.380 ;
        RECT 2931.200 2259.370 2934.200 2259.380 ;
        RECT -14.580 2082.380 -11.580 2082.390 ;
        RECT 2931.200 2082.380 2934.200 2082.390 ;
        RECT -14.580 2079.380 2934.200 2082.380 ;
        RECT -14.580 2079.370 -11.580 2079.380 ;
        RECT 2931.200 2079.370 2934.200 2079.380 ;
        RECT -14.580 1902.380 -11.580 1902.390 ;
        RECT 2931.200 1902.380 2934.200 1902.390 ;
        RECT -14.580 1899.380 2934.200 1902.380 ;
        RECT -14.580 1899.370 -11.580 1899.380 ;
        RECT 2931.200 1899.370 2934.200 1899.380 ;
        RECT -14.580 1722.380 -11.580 1722.390 ;
        RECT 2931.200 1722.380 2934.200 1722.390 ;
        RECT -14.580 1719.380 2934.200 1722.380 ;
        RECT -14.580 1719.370 -11.580 1719.380 ;
        RECT 2931.200 1719.370 2934.200 1719.380 ;
        RECT -14.580 1542.380 -11.580 1542.390 ;
        RECT 2931.200 1542.380 2934.200 1542.390 ;
        RECT -14.580 1539.380 2934.200 1542.380 ;
        RECT -14.580 1539.370 -11.580 1539.380 ;
        RECT 2931.200 1539.370 2934.200 1539.380 ;
        RECT -14.580 1362.380 -11.580 1362.390 ;
        RECT 2931.200 1362.380 2934.200 1362.390 ;
        RECT -14.580 1359.380 2934.200 1362.380 ;
        RECT -14.580 1359.370 -11.580 1359.380 ;
        RECT 2931.200 1359.370 2934.200 1359.380 ;
        RECT -14.580 1182.380 -11.580 1182.390 ;
        RECT 2931.200 1182.380 2934.200 1182.390 ;
        RECT -14.580 1179.380 2934.200 1182.380 ;
        RECT -14.580 1179.370 -11.580 1179.380 ;
        RECT 2931.200 1179.370 2934.200 1179.380 ;
        RECT -14.580 1002.380 -11.580 1002.390 ;
        RECT 2931.200 1002.380 2934.200 1002.390 ;
        RECT -14.580 999.380 2934.200 1002.380 ;
        RECT -14.580 999.370 -11.580 999.380 ;
        RECT 2931.200 999.370 2934.200 999.380 ;
        RECT -14.580 822.380 -11.580 822.390 ;
        RECT 2931.200 822.380 2934.200 822.390 ;
        RECT -14.580 819.380 2934.200 822.380 ;
        RECT -14.580 819.370 -11.580 819.380 ;
        RECT 2931.200 819.370 2934.200 819.380 ;
        RECT -14.580 642.380 -11.580 642.390 ;
        RECT 2931.200 642.380 2934.200 642.390 ;
        RECT -14.580 639.380 2934.200 642.380 ;
        RECT -14.580 639.370 -11.580 639.380 ;
        RECT 2931.200 639.370 2934.200 639.380 ;
        RECT -14.580 462.380 -11.580 462.390 ;
        RECT 2931.200 462.380 2934.200 462.390 ;
        RECT -14.580 459.380 2934.200 462.380 ;
        RECT -14.580 459.370 -11.580 459.380 ;
        RECT 2931.200 459.370 2934.200 459.380 ;
        RECT -14.580 282.380 -11.580 282.390 ;
        RECT 2931.200 282.380 2934.200 282.390 ;
        RECT -14.580 279.380 2934.200 282.380 ;
        RECT -14.580 279.370 -11.580 279.380 ;
        RECT 2931.200 279.370 2934.200 279.380 ;
        RECT -14.580 102.380 -11.580 102.390 ;
        RECT 2931.200 102.380 2934.200 102.390 ;
        RECT -14.580 99.380 2934.200 102.380 ;
        RECT -14.580 99.370 -11.580 99.380 ;
        RECT 2931.200 99.370 2934.200 99.380 ;
        RECT -14.580 -6.220 -11.580 -6.210 ;
        RECT 2931.200 -6.220 2934.200 -6.210 ;
        RECT -14.580 -9.220 2934.200 -6.220 ;
        RECT -14.580 -9.230 -11.580 -9.220 ;
        RECT 2931.200 -9.230 2934.200 -9.220 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.180 -13.820 -16.180 3533.500 ;
        RECT 2935.800 -13.820 2938.800 3533.500 ;
      LAYER via4 ;
        RECT -18.270 3532.210 -17.090 3533.390 ;
        RECT -18.270 3530.610 -17.090 3531.790 ;
        RECT -18.270 3449.090 -17.090 3450.270 ;
        RECT -18.270 3447.490 -17.090 3448.670 ;
        RECT -18.270 3269.090 -17.090 3270.270 ;
        RECT -18.270 3267.490 -17.090 3268.670 ;
        RECT -18.270 3089.090 -17.090 3090.270 ;
        RECT -18.270 3087.490 -17.090 3088.670 ;
        RECT -18.270 2909.090 -17.090 2910.270 ;
        RECT -18.270 2907.490 -17.090 2908.670 ;
        RECT -18.270 2729.090 -17.090 2730.270 ;
        RECT -18.270 2727.490 -17.090 2728.670 ;
        RECT -18.270 2549.090 -17.090 2550.270 ;
        RECT -18.270 2547.490 -17.090 2548.670 ;
        RECT -18.270 2369.090 -17.090 2370.270 ;
        RECT -18.270 2367.490 -17.090 2368.670 ;
        RECT -18.270 2189.090 -17.090 2190.270 ;
        RECT -18.270 2187.490 -17.090 2188.670 ;
        RECT -18.270 2009.090 -17.090 2010.270 ;
        RECT -18.270 2007.490 -17.090 2008.670 ;
        RECT -18.270 1829.090 -17.090 1830.270 ;
        RECT -18.270 1827.490 -17.090 1828.670 ;
        RECT -18.270 1649.090 -17.090 1650.270 ;
        RECT -18.270 1647.490 -17.090 1648.670 ;
        RECT -18.270 1469.090 -17.090 1470.270 ;
        RECT -18.270 1467.490 -17.090 1468.670 ;
        RECT -18.270 1289.090 -17.090 1290.270 ;
        RECT -18.270 1287.490 -17.090 1288.670 ;
        RECT -18.270 1109.090 -17.090 1110.270 ;
        RECT -18.270 1107.490 -17.090 1108.670 ;
        RECT -18.270 929.090 -17.090 930.270 ;
        RECT -18.270 927.490 -17.090 928.670 ;
        RECT -18.270 749.090 -17.090 750.270 ;
        RECT -18.270 747.490 -17.090 748.670 ;
        RECT -18.270 569.090 -17.090 570.270 ;
        RECT -18.270 567.490 -17.090 568.670 ;
        RECT -18.270 389.090 -17.090 390.270 ;
        RECT -18.270 387.490 -17.090 388.670 ;
        RECT -18.270 209.090 -17.090 210.270 ;
        RECT -18.270 207.490 -17.090 208.670 ;
        RECT -18.270 29.090 -17.090 30.270 ;
        RECT -18.270 27.490 -17.090 28.670 ;
        RECT -18.270 -12.110 -17.090 -10.930 ;
        RECT -18.270 -13.710 -17.090 -12.530 ;
        RECT 2936.710 3532.210 2937.890 3533.390 ;
        RECT 2936.710 3530.610 2937.890 3531.790 ;
        RECT 2936.710 3449.090 2937.890 3450.270 ;
        RECT 2936.710 3447.490 2937.890 3448.670 ;
        RECT 2936.710 3269.090 2937.890 3270.270 ;
        RECT 2936.710 3267.490 2937.890 3268.670 ;
        RECT 2936.710 3089.090 2937.890 3090.270 ;
        RECT 2936.710 3087.490 2937.890 3088.670 ;
        RECT 2936.710 2909.090 2937.890 2910.270 ;
        RECT 2936.710 2907.490 2937.890 2908.670 ;
        RECT 2936.710 2729.090 2937.890 2730.270 ;
        RECT 2936.710 2727.490 2937.890 2728.670 ;
        RECT 2936.710 2549.090 2937.890 2550.270 ;
        RECT 2936.710 2547.490 2937.890 2548.670 ;
        RECT 2936.710 2369.090 2937.890 2370.270 ;
        RECT 2936.710 2367.490 2937.890 2368.670 ;
        RECT 2936.710 2189.090 2937.890 2190.270 ;
        RECT 2936.710 2187.490 2937.890 2188.670 ;
        RECT 2936.710 2009.090 2937.890 2010.270 ;
        RECT 2936.710 2007.490 2937.890 2008.670 ;
        RECT 2936.710 1829.090 2937.890 1830.270 ;
        RECT 2936.710 1827.490 2937.890 1828.670 ;
        RECT 2936.710 1649.090 2937.890 1650.270 ;
        RECT 2936.710 1647.490 2937.890 1648.670 ;
        RECT 2936.710 1469.090 2937.890 1470.270 ;
        RECT 2936.710 1467.490 2937.890 1468.670 ;
        RECT 2936.710 1289.090 2937.890 1290.270 ;
        RECT 2936.710 1287.490 2937.890 1288.670 ;
        RECT 2936.710 1109.090 2937.890 1110.270 ;
        RECT 2936.710 1107.490 2937.890 1108.670 ;
        RECT 2936.710 929.090 2937.890 930.270 ;
        RECT 2936.710 927.490 2937.890 928.670 ;
        RECT 2936.710 749.090 2937.890 750.270 ;
        RECT 2936.710 747.490 2937.890 748.670 ;
        RECT 2936.710 569.090 2937.890 570.270 ;
        RECT 2936.710 567.490 2937.890 568.670 ;
        RECT 2936.710 389.090 2937.890 390.270 ;
        RECT 2936.710 387.490 2937.890 388.670 ;
        RECT 2936.710 209.090 2937.890 210.270 ;
        RECT 2936.710 207.490 2937.890 208.670 ;
        RECT 2936.710 29.090 2937.890 30.270 ;
        RECT 2936.710 27.490 2937.890 28.670 ;
        RECT 2936.710 -12.110 2937.890 -10.930 ;
        RECT 2936.710 -13.710 2937.890 -12.530 ;
      LAYER met5 ;
        RECT -19.180 3533.500 -16.180 3533.510 ;
        RECT 2935.800 3533.500 2938.800 3533.510 ;
        RECT -19.180 3530.500 2938.800 3533.500 ;
        RECT -19.180 3530.490 -16.180 3530.500 ;
        RECT 2935.800 3530.490 2938.800 3530.500 ;
        RECT -19.180 3450.380 -16.180 3450.390 ;
        RECT 2935.800 3450.380 2938.800 3450.390 ;
        RECT -23.780 3447.380 2943.400 3450.380 ;
        RECT -19.180 3447.370 -16.180 3447.380 ;
        RECT 2935.800 3447.370 2938.800 3447.380 ;
        RECT -19.180 3270.380 -16.180 3270.390 ;
        RECT 2935.800 3270.380 2938.800 3270.390 ;
        RECT -23.780 3267.380 2943.400 3270.380 ;
        RECT -19.180 3267.370 -16.180 3267.380 ;
        RECT 2935.800 3267.370 2938.800 3267.380 ;
        RECT -19.180 3090.380 -16.180 3090.390 ;
        RECT 2935.800 3090.380 2938.800 3090.390 ;
        RECT -23.780 3087.380 2943.400 3090.380 ;
        RECT -19.180 3087.370 -16.180 3087.380 ;
        RECT 2935.800 3087.370 2938.800 3087.380 ;
        RECT -19.180 2910.380 -16.180 2910.390 ;
        RECT 2935.800 2910.380 2938.800 2910.390 ;
        RECT -23.780 2907.380 2943.400 2910.380 ;
        RECT -19.180 2907.370 -16.180 2907.380 ;
        RECT 2935.800 2907.370 2938.800 2907.380 ;
        RECT -19.180 2730.380 -16.180 2730.390 ;
        RECT 2935.800 2730.380 2938.800 2730.390 ;
        RECT -23.780 2727.380 2943.400 2730.380 ;
        RECT -19.180 2727.370 -16.180 2727.380 ;
        RECT 2935.800 2727.370 2938.800 2727.380 ;
        RECT -19.180 2550.380 -16.180 2550.390 ;
        RECT 2935.800 2550.380 2938.800 2550.390 ;
        RECT -23.780 2547.380 2943.400 2550.380 ;
        RECT -19.180 2547.370 -16.180 2547.380 ;
        RECT 2935.800 2547.370 2938.800 2547.380 ;
        RECT -19.180 2370.380 -16.180 2370.390 ;
        RECT 2935.800 2370.380 2938.800 2370.390 ;
        RECT -23.780 2367.380 2943.400 2370.380 ;
        RECT -19.180 2367.370 -16.180 2367.380 ;
        RECT 2935.800 2367.370 2938.800 2367.380 ;
        RECT -19.180 2190.380 -16.180 2190.390 ;
        RECT 2935.800 2190.380 2938.800 2190.390 ;
        RECT -23.780 2187.380 2943.400 2190.380 ;
        RECT -19.180 2187.370 -16.180 2187.380 ;
        RECT 2935.800 2187.370 2938.800 2187.380 ;
        RECT -19.180 2010.380 -16.180 2010.390 ;
        RECT 2935.800 2010.380 2938.800 2010.390 ;
        RECT -23.780 2007.380 2943.400 2010.380 ;
        RECT -19.180 2007.370 -16.180 2007.380 ;
        RECT 2935.800 2007.370 2938.800 2007.380 ;
        RECT -19.180 1830.380 -16.180 1830.390 ;
        RECT 2935.800 1830.380 2938.800 1830.390 ;
        RECT -23.780 1827.380 2943.400 1830.380 ;
        RECT -19.180 1827.370 -16.180 1827.380 ;
        RECT 2935.800 1827.370 2938.800 1827.380 ;
        RECT -19.180 1650.380 -16.180 1650.390 ;
        RECT 2935.800 1650.380 2938.800 1650.390 ;
        RECT -23.780 1647.380 2943.400 1650.380 ;
        RECT -19.180 1647.370 -16.180 1647.380 ;
        RECT 2935.800 1647.370 2938.800 1647.380 ;
        RECT -19.180 1470.380 -16.180 1470.390 ;
        RECT 2935.800 1470.380 2938.800 1470.390 ;
        RECT -23.780 1467.380 2943.400 1470.380 ;
        RECT -19.180 1467.370 -16.180 1467.380 ;
        RECT 2935.800 1467.370 2938.800 1467.380 ;
        RECT -19.180 1290.380 -16.180 1290.390 ;
        RECT 2935.800 1290.380 2938.800 1290.390 ;
        RECT -23.780 1287.380 2943.400 1290.380 ;
        RECT -19.180 1287.370 -16.180 1287.380 ;
        RECT 2935.800 1287.370 2938.800 1287.380 ;
        RECT -19.180 1110.380 -16.180 1110.390 ;
        RECT 2935.800 1110.380 2938.800 1110.390 ;
        RECT -23.780 1107.380 2943.400 1110.380 ;
        RECT -19.180 1107.370 -16.180 1107.380 ;
        RECT 2935.800 1107.370 2938.800 1107.380 ;
        RECT -19.180 930.380 -16.180 930.390 ;
        RECT 2935.800 930.380 2938.800 930.390 ;
        RECT -23.780 927.380 2943.400 930.380 ;
        RECT -19.180 927.370 -16.180 927.380 ;
        RECT 2935.800 927.370 2938.800 927.380 ;
        RECT -19.180 750.380 -16.180 750.390 ;
        RECT 2935.800 750.380 2938.800 750.390 ;
        RECT -23.780 747.380 2943.400 750.380 ;
        RECT -19.180 747.370 -16.180 747.380 ;
        RECT 2935.800 747.370 2938.800 747.380 ;
        RECT -19.180 570.380 -16.180 570.390 ;
        RECT 2935.800 570.380 2938.800 570.390 ;
        RECT -23.780 567.380 2943.400 570.380 ;
        RECT -19.180 567.370 -16.180 567.380 ;
        RECT 2935.800 567.370 2938.800 567.380 ;
        RECT -19.180 390.380 -16.180 390.390 ;
        RECT 2935.800 390.380 2938.800 390.390 ;
        RECT -23.780 387.380 2943.400 390.380 ;
        RECT -19.180 387.370 -16.180 387.380 ;
        RECT 2935.800 387.370 2938.800 387.380 ;
        RECT -19.180 210.380 -16.180 210.390 ;
        RECT 2935.800 210.380 2938.800 210.390 ;
        RECT -23.780 207.380 2943.400 210.380 ;
        RECT -19.180 207.370 -16.180 207.380 ;
        RECT 2935.800 207.370 2938.800 207.380 ;
        RECT -19.180 30.380 -16.180 30.390 ;
        RECT 2935.800 30.380 2938.800 30.390 ;
        RECT -23.780 27.380 2943.400 30.380 ;
        RECT -19.180 27.370 -16.180 27.380 ;
        RECT 2935.800 27.370 2938.800 27.380 ;
        RECT -19.180 -10.820 -16.180 -10.810 ;
        RECT 2935.800 -10.820 2938.800 -10.810 ;
        RECT -19.180 -13.820 2938.800 -10.820 ;
        RECT -19.180 -13.830 -16.180 -13.820 ;
        RECT 2935.800 -13.830 2938.800 -13.820 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -23.780 -18.420 -20.780 3538.100 ;
        RECT 2940.400 -18.420 2943.400 3538.100 ;
      LAYER via4 ;
        RECT -22.870 3536.810 -21.690 3537.990 ;
        RECT -22.870 3535.210 -21.690 3536.390 ;
        RECT -22.870 3359.090 -21.690 3360.270 ;
        RECT -22.870 3357.490 -21.690 3358.670 ;
        RECT -22.870 3179.090 -21.690 3180.270 ;
        RECT -22.870 3177.490 -21.690 3178.670 ;
        RECT -22.870 2999.090 -21.690 3000.270 ;
        RECT -22.870 2997.490 -21.690 2998.670 ;
        RECT -22.870 2819.090 -21.690 2820.270 ;
        RECT -22.870 2817.490 -21.690 2818.670 ;
        RECT -22.870 2639.090 -21.690 2640.270 ;
        RECT -22.870 2637.490 -21.690 2638.670 ;
        RECT -22.870 2459.090 -21.690 2460.270 ;
        RECT -22.870 2457.490 -21.690 2458.670 ;
        RECT -22.870 2279.090 -21.690 2280.270 ;
        RECT -22.870 2277.490 -21.690 2278.670 ;
        RECT -22.870 2099.090 -21.690 2100.270 ;
        RECT -22.870 2097.490 -21.690 2098.670 ;
        RECT -22.870 1919.090 -21.690 1920.270 ;
        RECT -22.870 1917.490 -21.690 1918.670 ;
        RECT -22.870 1739.090 -21.690 1740.270 ;
        RECT -22.870 1737.490 -21.690 1738.670 ;
        RECT -22.870 1559.090 -21.690 1560.270 ;
        RECT -22.870 1557.490 -21.690 1558.670 ;
        RECT -22.870 1379.090 -21.690 1380.270 ;
        RECT -22.870 1377.490 -21.690 1378.670 ;
        RECT -22.870 1199.090 -21.690 1200.270 ;
        RECT -22.870 1197.490 -21.690 1198.670 ;
        RECT -22.870 1019.090 -21.690 1020.270 ;
        RECT -22.870 1017.490 -21.690 1018.670 ;
        RECT -22.870 839.090 -21.690 840.270 ;
        RECT -22.870 837.490 -21.690 838.670 ;
        RECT -22.870 659.090 -21.690 660.270 ;
        RECT -22.870 657.490 -21.690 658.670 ;
        RECT -22.870 479.090 -21.690 480.270 ;
        RECT -22.870 477.490 -21.690 478.670 ;
        RECT -22.870 299.090 -21.690 300.270 ;
        RECT -22.870 297.490 -21.690 298.670 ;
        RECT -22.870 119.090 -21.690 120.270 ;
        RECT -22.870 117.490 -21.690 118.670 ;
        RECT -22.870 -16.710 -21.690 -15.530 ;
        RECT -22.870 -18.310 -21.690 -17.130 ;
        RECT 2941.310 3536.810 2942.490 3537.990 ;
        RECT 2941.310 3535.210 2942.490 3536.390 ;
        RECT 2941.310 3359.090 2942.490 3360.270 ;
        RECT 2941.310 3357.490 2942.490 3358.670 ;
        RECT 2941.310 3179.090 2942.490 3180.270 ;
        RECT 2941.310 3177.490 2942.490 3178.670 ;
        RECT 2941.310 2999.090 2942.490 3000.270 ;
        RECT 2941.310 2997.490 2942.490 2998.670 ;
        RECT 2941.310 2819.090 2942.490 2820.270 ;
        RECT 2941.310 2817.490 2942.490 2818.670 ;
        RECT 2941.310 2639.090 2942.490 2640.270 ;
        RECT 2941.310 2637.490 2942.490 2638.670 ;
        RECT 2941.310 2459.090 2942.490 2460.270 ;
        RECT 2941.310 2457.490 2942.490 2458.670 ;
        RECT 2941.310 2279.090 2942.490 2280.270 ;
        RECT 2941.310 2277.490 2942.490 2278.670 ;
        RECT 2941.310 2099.090 2942.490 2100.270 ;
        RECT 2941.310 2097.490 2942.490 2098.670 ;
        RECT 2941.310 1919.090 2942.490 1920.270 ;
        RECT 2941.310 1917.490 2942.490 1918.670 ;
        RECT 2941.310 1739.090 2942.490 1740.270 ;
        RECT 2941.310 1737.490 2942.490 1738.670 ;
        RECT 2941.310 1559.090 2942.490 1560.270 ;
        RECT 2941.310 1557.490 2942.490 1558.670 ;
        RECT 2941.310 1379.090 2942.490 1380.270 ;
        RECT 2941.310 1377.490 2942.490 1378.670 ;
        RECT 2941.310 1199.090 2942.490 1200.270 ;
        RECT 2941.310 1197.490 2942.490 1198.670 ;
        RECT 2941.310 1019.090 2942.490 1020.270 ;
        RECT 2941.310 1017.490 2942.490 1018.670 ;
        RECT 2941.310 839.090 2942.490 840.270 ;
        RECT 2941.310 837.490 2942.490 838.670 ;
        RECT 2941.310 659.090 2942.490 660.270 ;
        RECT 2941.310 657.490 2942.490 658.670 ;
        RECT 2941.310 479.090 2942.490 480.270 ;
        RECT 2941.310 477.490 2942.490 478.670 ;
        RECT 2941.310 299.090 2942.490 300.270 ;
        RECT 2941.310 297.490 2942.490 298.670 ;
        RECT 2941.310 119.090 2942.490 120.270 ;
        RECT 2941.310 117.490 2942.490 118.670 ;
        RECT 2941.310 -16.710 2942.490 -15.530 ;
        RECT 2941.310 -18.310 2942.490 -17.130 ;
      LAYER met5 ;
        RECT -23.780 3538.100 -20.780 3538.110 ;
        RECT 2940.400 3538.100 2943.400 3538.110 ;
        RECT -23.780 3535.100 2943.400 3538.100 ;
        RECT -23.780 3535.090 -20.780 3535.100 ;
        RECT 2940.400 3535.090 2943.400 3535.100 ;
        RECT -23.780 3360.380 -20.780 3360.390 ;
        RECT 2940.400 3360.380 2943.400 3360.390 ;
        RECT -23.780 3357.380 2943.400 3360.380 ;
        RECT -23.780 3357.370 -20.780 3357.380 ;
        RECT 2940.400 3357.370 2943.400 3357.380 ;
        RECT -23.780 3180.380 -20.780 3180.390 ;
        RECT 2940.400 3180.380 2943.400 3180.390 ;
        RECT -23.780 3177.380 2943.400 3180.380 ;
        RECT -23.780 3177.370 -20.780 3177.380 ;
        RECT 2940.400 3177.370 2943.400 3177.380 ;
        RECT -23.780 3000.380 -20.780 3000.390 ;
        RECT 2940.400 3000.380 2943.400 3000.390 ;
        RECT -23.780 2997.380 2943.400 3000.380 ;
        RECT -23.780 2997.370 -20.780 2997.380 ;
        RECT 2940.400 2997.370 2943.400 2997.380 ;
        RECT -23.780 2820.380 -20.780 2820.390 ;
        RECT 2940.400 2820.380 2943.400 2820.390 ;
        RECT -23.780 2817.380 2943.400 2820.380 ;
        RECT -23.780 2817.370 -20.780 2817.380 ;
        RECT 2940.400 2817.370 2943.400 2817.380 ;
        RECT -23.780 2640.380 -20.780 2640.390 ;
        RECT 2940.400 2640.380 2943.400 2640.390 ;
        RECT -23.780 2637.380 2943.400 2640.380 ;
        RECT -23.780 2637.370 -20.780 2637.380 ;
        RECT 2940.400 2637.370 2943.400 2637.380 ;
        RECT -23.780 2460.380 -20.780 2460.390 ;
        RECT 2940.400 2460.380 2943.400 2460.390 ;
        RECT -23.780 2457.380 2943.400 2460.380 ;
        RECT -23.780 2457.370 -20.780 2457.380 ;
        RECT 2940.400 2457.370 2943.400 2457.380 ;
        RECT -23.780 2280.380 -20.780 2280.390 ;
        RECT 2940.400 2280.380 2943.400 2280.390 ;
        RECT -23.780 2277.380 2943.400 2280.380 ;
        RECT -23.780 2277.370 -20.780 2277.380 ;
        RECT 2940.400 2277.370 2943.400 2277.380 ;
        RECT -23.780 2100.380 -20.780 2100.390 ;
        RECT 2940.400 2100.380 2943.400 2100.390 ;
        RECT -23.780 2097.380 2943.400 2100.380 ;
        RECT -23.780 2097.370 -20.780 2097.380 ;
        RECT 2940.400 2097.370 2943.400 2097.380 ;
        RECT -23.780 1920.380 -20.780 1920.390 ;
        RECT 2940.400 1920.380 2943.400 1920.390 ;
        RECT -23.780 1917.380 2943.400 1920.380 ;
        RECT -23.780 1917.370 -20.780 1917.380 ;
        RECT 2940.400 1917.370 2943.400 1917.380 ;
        RECT -23.780 1740.380 -20.780 1740.390 ;
        RECT 2940.400 1740.380 2943.400 1740.390 ;
        RECT -23.780 1737.380 2943.400 1740.380 ;
        RECT -23.780 1737.370 -20.780 1737.380 ;
        RECT 2940.400 1737.370 2943.400 1737.380 ;
        RECT -23.780 1560.380 -20.780 1560.390 ;
        RECT 2940.400 1560.380 2943.400 1560.390 ;
        RECT -23.780 1557.380 2943.400 1560.380 ;
        RECT -23.780 1557.370 -20.780 1557.380 ;
        RECT 2940.400 1557.370 2943.400 1557.380 ;
        RECT -23.780 1380.380 -20.780 1380.390 ;
        RECT 2940.400 1380.380 2943.400 1380.390 ;
        RECT -23.780 1377.380 2943.400 1380.380 ;
        RECT -23.780 1377.370 -20.780 1377.380 ;
        RECT 2940.400 1377.370 2943.400 1377.380 ;
        RECT -23.780 1200.380 -20.780 1200.390 ;
        RECT 2940.400 1200.380 2943.400 1200.390 ;
        RECT -23.780 1197.380 2943.400 1200.380 ;
        RECT -23.780 1197.370 -20.780 1197.380 ;
        RECT 2940.400 1197.370 2943.400 1197.380 ;
        RECT -23.780 1020.380 -20.780 1020.390 ;
        RECT 2940.400 1020.380 2943.400 1020.390 ;
        RECT -23.780 1017.380 2943.400 1020.380 ;
        RECT -23.780 1017.370 -20.780 1017.380 ;
        RECT 2940.400 1017.370 2943.400 1017.380 ;
        RECT -23.780 840.380 -20.780 840.390 ;
        RECT 2940.400 840.380 2943.400 840.390 ;
        RECT -23.780 837.380 2943.400 840.380 ;
        RECT -23.780 837.370 -20.780 837.380 ;
        RECT 2940.400 837.370 2943.400 837.380 ;
        RECT -23.780 660.380 -20.780 660.390 ;
        RECT 2940.400 660.380 2943.400 660.390 ;
        RECT -23.780 657.380 2943.400 660.380 ;
        RECT -23.780 657.370 -20.780 657.380 ;
        RECT 2940.400 657.370 2943.400 657.380 ;
        RECT -23.780 480.380 -20.780 480.390 ;
        RECT 2940.400 480.380 2943.400 480.390 ;
        RECT -23.780 477.380 2943.400 480.380 ;
        RECT -23.780 477.370 -20.780 477.380 ;
        RECT 2940.400 477.370 2943.400 477.380 ;
        RECT -23.780 300.380 -20.780 300.390 ;
        RECT 2940.400 300.380 2943.400 300.390 ;
        RECT -23.780 297.380 2943.400 300.380 ;
        RECT -23.780 297.370 -20.780 297.380 ;
        RECT 2940.400 297.370 2943.400 297.380 ;
        RECT -23.780 120.380 -20.780 120.390 ;
        RECT 2940.400 120.380 2943.400 120.390 ;
        RECT -23.780 117.380 2943.400 120.380 ;
        RECT -23.780 117.370 -20.780 117.380 ;
        RECT 2940.400 117.370 2943.400 117.380 ;
        RECT -23.780 -15.420 -20.780 -15.410 ;
        RECT 2940.400 -15.420 2943.400 -15.410 ;
        RECT -23.780 -18.420 2943.400 -15.420 ;
        RECT -23.780 -18.430 -20.780 -18.420 ;
        RECT 2940.400 -18.430 2943.400 -18.420 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -28.380 -23.020 -25.380 3542.700 ;
        RECT 2945.000 -23.020 2948.000 3542.700 ;
      LAYER via4 ;
        RECT -27.470 3541.410 -26.290 3542.590 ;
        RECT -27.470 3539.810 -26.290 3540.990 ;
        RECT -27.470 3467.090 -26.290 3468.270 ;
        RECT -27.470 3465.490 -26.290 3466.670 ;
        RECT -27.470 3287.090 -26.290 3288.270 ;
        RECT -27.470 3285.490 -26.290 3286.670 ;
        RECT -27.470 3107.090 -26.290 3108.270 ;
        RECT -27.470 3105.490 -26.290 3106.670 ;
        RECT -27.470 2927.090 -26.290 2928.270 ;
        RECT -27.470 2925.490 -26.290 2926.670 ;
        RECT -27.470 2747.090 -26.290 2748.270 ;
        RECT -27.470 2745.490 -26.290 2746.670 ;
        RECT -27.470 2567.090 -26.290 2568.270 ;
        RECT -27.470 2565.490 -26.290 2566.670 ;
        RECT -27.470 2387.090 -26.290 2388.270 ;
        RECT -27.470 2385.490 -26.290 2386.670 ;
        RECT -27.470 2207.090 -26.290 2208.270 ;
        RECT -27.470 2205.490 -26.290 2206.670 ;
        RECT -27.470 2027.090 -26.290 2028.270 ;
        RECT -27.470 2025.490 -26.290 2026.670 ;
        RECT -27.470 1847.090 -26.290 1848.270 ;
        RECT -27.470 1845.490 -26.290 1846.670 ;
        RECT -27.470 1667.090 -26.290 1668.270 ;
        RECT -27.470 1665.490 -26.290 1666.670 ;
        RECT -27.470 1487.090 -26.290 1488.270 ;
        RECT -27.470 1485.490 -26.290 1486.670 ;
        RECT -27.470 1307.090 -26.290 1308.270 ;
        RECT -27.470 1305.490 -26.290 1306.670 ;
        RECT -27.470 1127.090 -26.290 1128.270 ;
        RECT -27.470 1125.490 -26.290 1126.670 ;
        RECT -27.470 947.090 -26.290 948.270 ;
        RECT -27.470 945.490 -26.290 946.670 ;
        RECT -27.470 767.090 -26.290 768.270 ;
        RECT -27.470 765.490 -26.290 766.670 ;
        RECT -27.470 587.090 -26.290 588.270 ;
        RECT -27.470 585.490 -26.290 586.670 ;
        RECT -27.470 407.090 -26.290 408.270 ;
        RECT -27.470 405.490 -26.290 406.670 ;
        RECT -27.470 227.090 -26.290 228.270 ;
        RECT -27.470 225.490 -26.290 226.670 ;
        RECT -27.470 47.090 -26.290 48.270 ;
        RECT -27.470 45.490 -26.290 46.670 ;
        RECT -27.470 -21.310 -26.290 -20.130 ;
        RECT -27.470 -22.910 -26.290 -21.730 ;
        RECT 2945.910 3541.410 2947.090 3542.590 ;
        RECT 2945.910 3539.810 2947.090 3540.990 ;
        RECT 2945.910 3467.090 2947.090 3468.270 ;
        RECT 2945.910 3465.490 2947.090 3466.670 ;
        RECT 2945.910 3287.090 2947.090 3288.270 ;
        RECT 2945.910 3285.490 2947.090 3286.670 ;
        RECT 2945.910 3107.090 2947.090 3108.270 ;
        RECT 2945.910 3105.490 2947.090 3106.670 ;
        RECT 2945.910 2927.090 2947.090 2928.270 ;
        RECT 2945.910 2925.490 2947.090 2926.670 ;
        RECT 2945.910 2747.090 2947.090 2748.270 ;
        RECT 2945.910 2745.490 2947.090 2746.670 ;
        RECT 2945.910 2567.090 2947.090 2568.270 ;
        RECT 2945.910 2565.490 2947.090 2566.670 ;
        RECT 2945.910 2387.090 2947.090 2388.270 ;
        RECT 2945.910 2385.490 2947.090 2386.670 ;
        RECT 2945.910 2207.090 2947.090 2208.270 ;
        RECT 2945.910 2205.490 2947.090 2206.670 ;
        RECT 2945.910 2027.090 2947.090 2028.270 ;
        RECT 2945.910 2025.490 2947.090 2026.670 ;
        RECT 2945.910 1847.090 2947.090 1848.270 ;
        RECT 2945.910 1845.490 2947.090 1846.670 ;
        RECT 2945.910 1667.090 2947.090 1668.270 ;
        RECT 2945.910 1665.490 2947.090 1666.670 ;
        RECT 2945.910 1487.090 2947.090 1488.270 ;
        RECT 2945.910 1485.490 2947.090 1486.670 ;
        RECT 2945.910 1307.090 2947.090 1308.270 ;
        RECT 2945.910 1305.490 2947.090 1306.670 ;
        RECT 2945.910 1127.090 2947.090 1128.270 ;
        RECT 2945.910 1125.490 2947.090 1126.670 ;
        RECT 2945.910 947.090 2947.090 948.270 ;
        RECT 2945.910 945.490 2947.090 946.670 ;
        RECT 2945.910 767.090 2947.090 768.270 ;
        RECT 2945.910 765.490 2947.090 766.670 ;
        RECT 2945.910 587.090 2947.090 588.270 ;
        RECT 2945.910 585.490 2947.090 586.670 ;
        RECT 2945.910 407.090 2947.090 408.270 ;
        RECT 2945.910 405.490 2947.090 406.670 ;
        RECT 2945.910 227.090 2947.090 228.270 ;
        RECT 2945.910 225.490 2947.090 226.670 ;
        RECT 2945.910 47.090 2947.090 48.270 ;
        RECT 2945.910 45.490 2947.090 46.670 ;
        RECT 2945.910 -21.310 2947.090 -20.130 ;
        RECT 2945.910 -22.910 2947.090 -21.730 ;
      LAYER met5 ;
        RECT -28.380 3542.700 -25.380 3542.710 ;
        RECT 2945.000 3542.700 2948.000 3542.710 ;
        RECT -28.380 3539.700 2948.000 3542.700 ;
        RECT -28.380 3539.690 -25.380 3539.700 ;
        RECT 2945.000 3539.690 2948.000 3539.700 ;
        RECT -28.380 3468.380 -25.380 3468.390 ;
        RECT 2945.000 3468.380 2948.000 3468.390 ;
        RECT -32.980 3465.380 2952.600 3468.380 ;
        RECT -28.380 3465.370 -25.380 3465.380 ;
        RECT 2945.000 3465.370 2948.000 3465.380 ;
        RECT -28.380 3288.380 -25.380 3288.390 ;
        RECT 2945.000 3288.380 2948.000 3288.390 ;
        RECT -32.980 3285.380 2952.600 3288.380 ;
        RECT -28.380 3285.370 -25.380 3285.380 ;
        RECT 2945.000 3285.370 2948.000 3285.380 ;
        RECT -28.380 3108.380 -25.380 3108.390 ;
        RECT 2945.000 3108.380 2948.000 3108.390 ;
        RECT -32.980 3105.380 2952.600 3108.380 ;
        RECT -28.380 3105.370 -25.380 3105.380 ;
        RECT 2945.000 3105.370 2948.000 3105.380 ;
        RECT -28.380 2928.380 -25.380 2928.390 ;
        RECT 2945.000 2928.380 2948.000 2928.390 ;
        RECT -32.980 2925.380 2952.600 2928.380 ;
        RECT -28.380 2925.370 -25.380 2925.380 ;
        RECT 2945.000 2925.370 2948.000 2925.380 ;
        RECT -28.380 2748.380 -25.380 2748.390 ;
        RECT 2945.000 2748.380 2948.000 2748.390 ;
        RECT -32.980 2745.380 2952.600 2748.380 ;
        RECT -28.380 2745.370 -25.380 2745.380 ;
        RECT 2945.000 2745.370 2948.000 2745.380 ;
        RECT -28.380 2568.380 -25.380 2568.390 ;
        RECT 2945.000 2568.380 2948.000 2568.390 ;
        RECT -32.980 2565.380 2952.600 2568.380 ;
        RECT -28.380 2565.370 -25.380 2565.380 ;
        RECT 2945.000 2565.370 2948.000 2565.380 ;
        RECT -28.380 2388.380 -25.380 2388.390 ;
        RECT 2945.000 2388.380 2948.000 2388.390 ;
        RECT -32.980 2385.380 2952.600 2388.380 ;
        RECT -28.380 2385.370 -25.380 2385.380 ;
        RECT 2945.000 2385.370 2948.000 2385.380 ;
        RECT -28.380 2208.380 -25.380 2208.390 ;
        RECT 2945.000 2208.380 2948.000 2208.390 ;
        RECT -32.980 2205.380 2952.600 2208.380 ;
        RECT -28.380 2205.370 -25.380 2205.380 ;
        RECT 2945.000 2205.370 2948.000 2205.380 ;
        RECT -28.380 2028.380 -25.380 2028.390 ;
        RECT 2945.000 2028.380 2948.000 2028.390 ;
        RECT -32.980 2025.380 2952.600 2028.380 ;
        RECT -28.380 2025.370 -25.380 2025.380 ;
        RECT 2945.000 2025.370 2948.000 2025.380 ;
        RECT -28.380 1848.380 -25.380 1848.390 ;
        RECT 2945.000 1848.380 2948.000 1848.390 ;
        RECT -32.980 1845.380 2952.600 1848.380 ;
        RECT -28.380 1845.370 -25.380 1845.380 ;
        RECT 2945.000 1845.370 2948.000 1845.380 ;
        RECT -28.380 1668.380 -25.380 1668.390 ;
        RECT 2945.000 1668.380 2948.000 1668.390 ;
        RECT -32.980 1665.380 2952.600 1668.380 ;
        RECT -28.380 1665.370 -25.380 1665.380 ;
        RECT 2945.000 1665.370 2948.000 1665.380 ;
        RECT -28.380 1488.380 -25.380 1488.390 ;
        RECT 2945.000 1488.380 2948.000 1488.390 ;
        RECT -32.980 1485.380 2952.600 1488.380 ;
        RECT -28.380 1485.370 -25.380 1485.380 ;
        RECT 2945.000 1485.370 2948.000 1485.380 ;
        RECT -28.380 1308.380 -25.380 1308.390 ;
        RECT 2945.000 1308.380 2948.000 1308.390 ;
        RECT -32.980 1305.380 2952.600 1308.380 ;
        RECT -28.380 1305.370 -25.380 1305.380 ;
        RECT 2945.000 1305.370 2948.000 1305.380 ;
        RECT -28.380 1128.380 -25.380 1128.390 ;
        RECT 2945.000 1128.380 2948.000 1128.390 ;
        RECT -32.980 1125.380 2952.600 1128.380 ;
        RECT -28.380 1125.370 -25.380 1125.380 ;
        RECT 2945.000 1125.370 2948.000 1125.380 ;
        RECT -28.380 948.380 -25.380 948.390 ;
        RECT 2945.000 948.380 2948.000 948.390 ;
        RECT -32.980 945.380 2952.600 948.380 ;
        RECT -28.380 945.370 -25.380 945.380 ;
        RECT 2945.000 945.370 2948.000 945.380 ;
        RECT -28.380 768.380 -25.380 768.390 ;
        RECT 2945.000 768.380 2948.000 768.390 ;
        RECT -32.980 765.380 2952.600 768.380 ;
        RECT -28.380 765.370 -25.380 765.380 ;
        RECT 2945.000 765.370 2948.000 765.380 ;
        RECT -28.380 588.380 -25.380 588.390 ;
        RECT 2945.000 588.380 2948.000 588.390 ;
        RECT -32.980 585.380 2952.600 588.380 ;
        RECT -28.380 585.370 -25.380 585.380 ;
        RECT 2945.000 585.370 2948.000 585.380 ;
        RECT -28.380 408.380 -25.380 408.390 ;
        RECT 2945.000 408.380 2948.000 408.390 ;
        RECT -32.980 405.380 2952.600 408.380 ;
        RECT -28.380 405.370 -25.380 405.380 ;
        RECT 2945.000 405.370 2948.000 405.380 ;
        RECT -28.380 228.380 -25.380 228.390 ;
        RECT 2945.000 228.380 2948.000 228.390 ;
        RECT -32.980 225.380 2952.600 228.380 ;
        RECT -28.380 225.370 -25.380 225.380 ;
        RECT 2945.000 225.370 2948.000 225.380 ;
        RECT -28.380 48.380 -25.380 48.390 ;
        RECT 2945.000 48.380 2948.000 48.390 ;
        RECT -32.980 45.380 2952.600 48.380 ;
        RECT -28.380 45.370 -25.380 45.380 ;
        RECT 2945.000 45.370 2948.000 45.380 ;
        RECT -28.380 -20.020 -25.380 -20.010 ;
        RECT 2945.000 -20.020 2948.000 -20.010 ;
        RECT -28.380 -23.020 2948.000 -20.020 ;
        RECT -28.380 -23.030 -25.380 -23.020 ;
        RECT 2945.000 -23.030 2948.000 -23.020 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -32.980 -27.620 -29.980 3547.300 ;
        RECT 2949.600 -27.620 2952.600 3547.300 ;
      LAYER via4 ;
        RECT -32.070 3546.010 -30.890 3547.190 ;
        RECT -32.070 3544.410 -30.890 3545.590 ;
        RECT -32.070 3377.090 -30.890 3378.270 ;
        RECT -32.070 3375.490 -30.890 3376.670 ;
        RECT -32.070 3197.090 -30.890 3198.270 ;
        RECT -32.070 3195.490 -30.890 3196.670 ;
        RECT -32.070 3017.090 -30.890 3018.270 ;
        RECT -32.070 3015.490 -30.890 3016.670 ;
        RECT -32.070 2837.090 -30.890 2838.270 ;
        RECT -32.070 2835.490 -30.890 2836.670 ;
        RECT -32.070 2657.090 -30.890 2658.270 ;
        RECT -32.070 2655.490 -30.890 2656.670 ;
        RECT -32.070 2477.090 -30.890 2478.270 ;
        RECT -32.070 2475.490 -30.890 2476.670 ;
        RECT -32.070 2297.090 -30.890 2298.270 ;
        RECT -32.070 2295.490 -30.890 2296.670 ;
        RECT -32.070 2117.090 -30.890 2118.270 ;
        RECT -32.070 2115.490 -30.890 2116.670 ;
        RECT -32.070 1937.090 -30.890 1938.270 ;
        RECT -32.070 1935.490 -30.890 1936.670 ;
        RECT -32.070 1757.090 -30.890 1758.270 ;
        RECT -32.070 1755.490 -30.890 1756.670 ;
        RECT -32.070 1577.090 -30.890 1578.270 ;
        RECT -32.070 1575.490 -30.890 1576.670 ;
        RECT -32.070 1397.090 -30.890 1398.270 ;
        RECT -32.070 1395.490 -30.890 1396.670 ;
        RECT -32.070 1217.090 -30.890 1218.270 ;
        RECT -32.070 1215.490 -30.890 1216.670 ;
        RECT -32.070 1037.090 -30.890 1038.270 ;
        RECT -32.070 1035.490 -30.890 1036.670 ;
        RECT -32.070 857.090 -30.890 858.270 ;
        RECT -32.070 855.490 -30.890 856.670 ;
        RECT -32.070 677.090 -30.890 678.270 ;
        RECT -32.070 675.490 -30.890 676.670 ;
        RECT -32.070 497.090 -30.890 498.270 ;
        RECT -32.070 495.490 -30.890 496.670 ;
        RECT -32.070 317.090 -30.890 318.270 ;
        RECT -32.070 315.490 -30.890 316.670 ;
        RECT -32.070 137.090 -30.890 138.270 ;
        RECT -32.070 135.490 -30.890 136.670 ;
        RECT -32.070 -25.910 -30.890 -24.730 ;
        RECT -32.070 -27.510 -30.890 -26.330 ;
        RECT 2950.510 3546.010 2951.690 3547.190 ;
        RECT 2950.510 3544.410 2951.690 3545.590 ;
        RECT 2950.510 3377.090 2951.690 3378.270 ;
        RECT 2950.510 3375.490 2951.690 3376.670 ;
        RECT 2950.510 3197.090 2951.690 3198.270 ;
        RECT 2950.510 3195.490 2951.690 3196.670 ;
        RECT 2950.510 3017.090 2951.690 3018.270 ;
        RECT 2950.510 3015.490 2951.690 3016.670 ;
        RECT 2950.510 2837.090 2951.690 2838.270 ;
        RECT 2950.510 2835.490 2951.690 2836.670 ;
        RECT 2950.510 2657.090 2951.690 2658.270 ;
        RECT 2950.510 2655.490 2951.690 2656.670 ;
        RECT 2950.510 2477.090 2951.690 2478.270 ;
        RECT 2950.510 2475.490 2951.690 2476.670 ;
        RECT 2950.510 2297.090 2951.690 2298.270 ;
        RECT 2950.510 2295.490 2951.690 2296.670 ;
        RECT 2950.510 2117.090 2951.690 2118.270 ;
        RECT 2950.510 2115.490 2951.690 2116.670 ;
        RECT 2950.510 1937.090 2951.690 1938.270 ;
        RECT 2950.510 1935.490 2951.690 1936.670 ;
        RECT 2950.510 1757.090 2951.690 1758.270 ;
        RECT 2950.510 1755.490 2951.690 1756.670 ;
        RECT 2950.510 1577.090 2951.690 1578.270 ;
        RECT 2950.510 1575.490 2951.690 1576.670 ;
        RECT 2950.510 1397.090 2951.690 1398.270 ;
        RECT 2950.510 1395.490 2951.690 1396.670 ;
        RECT 2950.510 1217.090 2951.690 1218.270 ;
        RECT 2950.510 1215.490 2951.690 1216.670 ;
        RECT 2950.510 1037.090 2951.690 1038.270 ;
        RECT 2950.510 1035.490 2951.690 1036.670 ;
        RECT 2950.510 857.090 2951.690 858.270 ;
        RECT 2950.510 855.490 2951.690 856.670 ;
        RECT 2950.510 677.090 2951.690 678.270 ;
        RECT 2950.510 675.490 2951.690 676.670 ;
        RECT 2950.510 497.090 2951.690 498.270 ;
        RECT 2950.510 495.490 2951.690 496.670 ;
        RECT 2950.510 317.090 2951.690 318.270 ;
        RECT 2950.510 315.490 2951.690 316.670 ;
        RECT 2950.510 137.090 2951.690 138.270 ;
        RECT 2950.510 135.490 2951.690 136.670 ;
        RECT 2950.510 -25.910 2951.690 -24.730 ;
        RECT 2950.510 -27.510 2951.690 -26.330 ;
      LAYER met5 ;
        RECT -32.980 3547.300 -29.980 3547.310 ;
        RECT 2949.600 3547.300 2952.600 3547.310 ;
        RECT -32.980 3544.300 2952.600 3547.300 ;
        RECT -32.980 3544.290 -29.980 3544.300 ;
        RECT 2949.600 3544.290 2952.600 3544.300 ;
        RECT -32.980 3378.380 -29.980 3378.390 ;
        RECT 2949.600 3378.380 2952.600 3378.390 ;
        RECT -32.980 3375.380 2952.600 3378.380 ;
        RECT -32.980 3375.370 -29.980 3375.380 ;
        RECT 2949.600 3375.370 2952.600 3375.380 ;
        RECT -32.980 3198.380 -29.980 3198.390 ;
        RECT 2949.600 3198.380 2952.600 3198.390 ;
        RECT -32.980 3195.380 2952.600 3198.380 ;
        RECT -32.980 3195.370 -29.980 3195.380 ;
        RECT 2949.600 3195.370 2952.600 3195.380 ;
        RECT -32.980 3018.380 -29.980 3018.390 ;
        RECT 2949.600 3018.380 2952.600 3018.390 ;
        RECT -32.980 3015.380 2952.600 3018.380 ;
        RECT -32.980 3015.370 -29.980 3015.380 ;
        RECT 2949.600 3015.370 2952.600 3015.380 ;
        RECT -32.980 2838.380 -29.980 2838.390 ;
        RECT 2949.600 2838.380 2952.600 2838.390 ;
        RECT -32.980 2835.380 2952.600 2838.380 ;
        RECT -32.980 2835.370 -29.980 2835.380 ;
        RECT 2949.600 2835.370 2952.600 2835.380 ;
        RECT -32.980 2658.380 -29.980 2658.390 ;
        RECT 2949.600 2658.380 2952.600 2658.390 ;
        RECT -32.980 2655.380 2952.600 2658.380 ;
        RECT -32.980 2655.370 -29.980 2655.380 ;
        RECT 2949.600 2655.370 2952.600 2655.380 ;
        RECT -32.980 2478.380 -29.980 2478.390 ;
        RECT 2949.600 2478.380 2952.600 2478.390 ;
        RECT -32.980 2475.380 2952.600 2478.380 ;
        RECT -32.980 2475.370 -29.980 2475.380 ;
        RECT 2949.600 2475.370 2952.600 2475.380 ;
        RECT -32.980 2298.380 -29.980 2298.390 ;
        RECT 2949.600 2298.380 2952.600 2298.390 ;
        RECT -32.980 2295.380 2952.600 2298.380 ;
        RECT -32.980 2295.370 -29.980 2295.380 ;
        RECT 2949.600 2295.370 2952.600 2295.380 ;
        RECT -32.980 2118.380 -29.980 2118.390 ;
        RECT 2949.600 2118.380 2952.600 2118.390 ;
        RECT -32.980 2115.380 2952.600 2118.380 ;
        RECT -32.980 2115.370 -29.980 2115.380 ;
        RECT 2949.600 2115.370 2952.600 2115.380 ;
        RECT -32.980 1938.380 -29.980 1938.390 ;
        RECT 2949.600 1938.380 2952.600 1938.390 ;
        RECT -32.980 1935.380 2952.600 1938.380 ;
        RECT -32.980 1935.370 -29.980 1935.380 ;
        RECT 2949.600 1935.370 2952.600 1935.380 ;
        RECT -32.980 1758.380 -29.980 1758.390 ;
        RECT 2949.600 1758.380 2952.600 1758.390 ;
        RECT -32.980 1755.380 2952.600 1758.380 ;
        RECT -32.980 1755.370 -29.980 1755.380 ;
        RECT 2949.600 1755.370 2952.600 1755.380 ;
        RECT -32.980 1578.380 -29.980 1578.390 ;
        RECT 2949.600 1578.380 2952.600 1578.390 ;
        RECT -32.980 1575.380 2952.600 1578.380 ;
        RECT -32.980 1575.370 -29.980 1575.380 ;
        RECT 2949.600 1575.370 2952.600 1575.380 ;
        RECT -32.980 1398.380 -29.980 1398.390 ;
        RECT 2949.600 1398.380 2952.600 1398.390 ;
        RECT -32.980 1395.380 2952.600 1398.380 ;
        RECT -32.980 1395.370 -29.980 1395.380 ;
        RECT 2949.600 1395.370 2952.600 1395.380 ;
        RECT -32.980 1218.380 -29.980 1218.390 ;
        RECT 2949.600 1218.380 2952.600 1218.390 ;
        RECT -32.980 1215.380 2952.600 1218.380 ;
        RECT -32.980 1215.370 -29.980 1215.380 ;
        RECT 2949.600 1215.370 2952.600 1215.380 ;
        RECT -32.980 1038.380 -29.980 1038.390 ;
        RECT 2949.600 1038.380 2952.600 1038.390 ;
        RECT -32.980 1035.380 2952.600 1038.380 ;
        RECT -32.980 1035.370 -29.980 1035.380 ;
        RECT 2949.600 1035.370 2952.600 1035.380 ;
        RECT -32.980 858.380 -29.980 858.390 ;
        RECT 2949.600 858.380 2952.600 858.390 ;
        RECT -32.980 855.380 2952.600 858.380 ;
        RECT -32.980 855.370 -29.980 855.380 ;
        RECT 2949.600 855.370 2952.600 855.380 ;
        RECT -32.980 678.380 -29.980 678.390 ;
        RECT 2949.600 678.380 2952.600 678.390 ;
        RECT -32.980 675.380 2952.600 678.380 ;
        RECT -32.980 675.370 -29.980 675.380 ;
        RECT 2949.600 675.370 2952.600 675.380 ;
        RECT -32.980 498.380 -29.980 498.390 ;
        RECT 2949.600 498.380 2952.600 498.390 ;
        RECT -32.980 495.380 2952.600 498.380 ;
        RECT -32.980 495.370 -29.980 495.380 ;
        RECT 2949.600 495.370 2952.600 495.380 ;
        RECT -32.980 318.380 -29.980 318.390 ;
        RECT 2949.600 318.380 2952.600 318.390 ;
        RECT -32.980 315.380 2952.600 318.380 ;
        RECT -32.980 315.370 -29.980 315.380 ;
        RECT 2949.600 315.370 2952.600 315.380 ;
        RECT -32.980 138.380 -29.980 138.390 ;
        RECT 2949.600 138.380 2952.600 138.390 ;
        RECT -32.980 135.380 2952.600 138.380 ;
        RECT -32.980 135.370 -29.980 135.380 ;
        RECT 2949.600 135.370 2952.600 135.380 ;
        RECT -32.980 -24.620 -29.980 -24.610 ;
        RECT 2949.600 -24.620 2952.600 -24.610 ;
        RECT -32.980 -27.620 2952.600 -24.620 ;
        RECT -32.980 -27.630 -29.980 -27.620 ;
        RECT 2949.600 -27.630 2952.600 -27.620 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -42.180 -36.820 -39.180 3556.500 ;
        RECT 2958.800 -36.820 2961.800 3556.500 ;
      LAYER via4 ;
        RECT -41.270 3555.210 -40.090 3556.390 ;
        RECT -41.270 3553.610 -40.090 3554.790 ;
        RECT -41.270 3395.090 -40.090 3396.270 ;
        RECT -41.270 3393.490 -40.090 3394.670 ;
        RECT -41.270 3215.090 -40.090 3216.270 ;
        RECT -41.270 3213.490 -40.090 3214.670 ;
        RECT -41.270 3035.090 -40.090 3036.270 ;
        RECT -41.270 3033.490 -40.090 3034.670 ;
        RECT -41.270 2855.090 -40.090 2856.270 ;
        RECT -41.270 2853.490 -40.090 2854.670 ;
        RECT -41.270 2675.090 -40.090 2676.270 ;
        RECT -41.270 2673.490 -40.090 2674.670 ;
        RECT -41.270 2495.090 -40.090 2496.270 ;
        RECT -41.270 2493.490 -40.090 2494.670 ;
        RECT -41.270 2315.090 -40.090 2316.270 ;
        RECT -41.270 2313.490 -40.090 2314.670 ;
        RECT -41.270 2135.090 -40.090 2136.270 ;
        RECT -41.270 2133.490 -40.090 2134.670 ;
        RECT -41.270 1955.090 -40.090 1956.270 ;
        RECT -41.270 1953.490 -40.090 1954.670 ;
        RECT -41.270 1775.090 -40.090 1776.270 ;
        RECT -41.270 1773.490 -40.090 1774.670 ;
        RECT -41.270 1595.090 -40.090 1596.270 ;
        RECT -41.270 1593.490 -40.090 1594.670 ;
        RECT -41.270 1415.090 -40.090 1416.270 ;
        RECT -41.270 1413.490 -40.090 1414.670 ;
        RECT -41.270 1235.090 -40.090 1236.270 ;
        RECT -41.270 1233.490 -40.090 1234.670 ;
        RECT -41.270 1055.090 -40.090 1056.270 ;
        RECT -41.270 1053.490 -40.090 1054.670 ;
        RECT -41.270 875.090 -40.090 876.270 ;
        RECT -41.270 873.490 -40.090 874.670 ;
        RECT -41.270 695.090 -40.090 696.270 ;
        RECT -41.270 693.490 -40.090 694.670 ;
        RECT -41.270 515.090 -40.090 516.270 ;
        RECT -41.270 513.490 -40.090 514.670 ;
        RECT -41.270 335.090 -40.090 336.270 ;
        RECT -41.270 333.490 -40.090 334.670 ;
        RECT -41.270 155.090 -40.090 156.270 ;
        RECT -41.270 153.490 -40.090 154.670 ;
        RECT -41.270 -35.110 -40.090 -33.930 ;
        RECT -41.270 -36.710 -40.090 -35.530 ;
        RECT 2959.710 3555.210 2960.890 3556.390 ;
        RECT 2959.710 3553.610 2960.890 3554.790 ;
        RECT 2959.710 3395.090 2960.890 3396.270 ;
        RECT 2959.710 3393.490 2960.890 3394.670 ;
        RECT 2959.710 3215.090 2960.890 3216.270 ;
        RECT 2959.710 3213.490 2960.890 3214.670 ;
        RECT 2959.710 3035.090 2960.890 3036.270 ;
        RECT 2959.710 3033.490 2960.890 3034.670 ;
        RECT 2959.710 2855.090 2960.890 2856.270 ;
        RECT 2959.710 2853.490 2960.890 2854.670 ;
        RECT 2959.710 2675.090 2960.890 2676.270 ;
        RECT 2959.710 2673.490 2960.890 2674.670 ;
        RECT 2959.710 2495.090 2960.890 2496.270 ;
        RECT 2959.710 2493.490 2960.890 2494.670 ;
        RECT 2959.710 2315.090 2960.890 2316.270 ;
        RECT 2959.710 2313.490 2960.890 2314.670 ;
        RECT 2959.710 2135.090 2960.890 2136.270 ;
        RECT 2959.710 2133.490 2960.890 2134.670 ;
        RECT 2959.710 1955.090 2960.890 1956.270 ;
        RECT 2959.710 1953.490 2960.890 1954.670 ;
        RECT 2959.710 1775.090 2960.890 1776.270 ;
        RECT 2959.710 1773.490 2960.890 1774.670 ;
        RECT 2959.710 1595.090 2960.890 1596.270 ;
        RECT 2959.710 1593.490 2960.890 1594.670 ;
        RECT 2959.710 1415.090 2960.890 1416.270 ;
        RECT 2959.710 1413.490 2960.890 1414.670 ;
        RECT 2959.710 1235.090 2960.890 1236.270 ;
        RECT 2959.710 1233.490 2960.890 1234.670 ;
        RECT 2959.710 1055.090 2960.890 1056.270 ;
        RECT 2959.710 1053.490 2960.890 1054.670 ;
        RECT 2959.710 875.090 2960.890 876.270 ;
        RECT 2959.710 873.490 2960.890 874.670 ;
        RECT 2959.710 695.090 2960.890 696.270 ;
        RECT 2959.710 693.490 2960.890 694.670 ;
        RECT 2959.710 515.090 2960.890 516.270 ;
        RECT 2959.710 513.490 2960.890 514.670 ;
        RECT 2959.710 335.090 2960.890 336.270 ;
        RECT 2959.710 333.490 2960.890 334.670 ;
        RECT 2959.710 155.090 2960.890 156.270 ;
        RECT 2959.710 153.490 2960.890 154.670 ;
        RECT 2959.710 -35.110 2960.890 -33.930 ;
        RECT 2959.710 -36.710 2960.890 -35.530 ;
      LAYER met5 ;
        RECT -42.180 3556.500 -39.180 3556.510 ;
        RECT 2958.800 3556.500 2961.800 3556.510 ;
        RECT -42.180 3553.500 2961.800 3556.500 ;
        RECT -42.180 3553.490 -39.180 3553.500 ;
        RECT 2958.800 3553.490 2961.800 3553.500 ;
        RECT -42.180 3396.380 -39.180 3396.390 ;
        RECT 2958.800 3396.380 2961.800 3396.390 ;
        RECT -42.180 3393.380 2961.800 3396.380 ;
        RECT -42.180 3393.370 -39.180 3393.380 ;
        RECT 2958.800 3393.370 2961.800 3393.380 ;
        RECT -42.180 3216.380 -39.180 3216.390 ;
        RECT 2958.800 3216.380 2961.800 3216.390 ;
        RECT -42.180 3213.380 2961.800 3216.380 ;
        RECT -42.180 3213.370 -39.180 3213.380 ;
        RECT 2958.800 3213.370 2961.800 3213.380 ;
        RECT -42.180 3036.380 -39.180 3036.390 ;
        RECT 2958.800 3036.380 2961.800 3036.390 ;
        RECT -42.180 3033.380 2961.800 3036.380 ;
        RECT -42.180 3033.370 -39.180 3033.380 ;
        RECT 2958.800 3033.370 2961.800 3033.380 ;
        RECT -42.180 2856.380 -39.180 2856.390 ;
        RECT 2958.800 2856.380 2961.800 2856.390 ;
        RECT -42.180 2853.380 2961.800 2856.380 ;
        RECT -42.180 2853.370 -39.180 2853.380 ;
        RECT 2958.800 2853.370 2961.800 2853.380 ;
        RECT -42.180 2676.380 -39.180 2676.390 ;
        RECT 2958.800 2676.380 2961.800 2676.390 ;
        RECT -42.180 2673.380 2961.800 2676.380 ;
        RECT -42.180 2673.370 -39.180 2673.380 ;
        RECT 2958.800 2673.370 2961.800 2673.380 ;
        RECT -42.180 2496.380 -39.180 2496.390 ;
        RECT 2958.800 2496.380 2961.800 2496.390 ;
        RECT -42.180 2493.380 2961.800 2496.380 ;
        RECT -42.180 2493.370 -39.180 2493.380 ;
        RECT 2958.800 2493.370 2961.800 2493.380 ;
        RECT -42.180 2316.380 -39.180 2316.390 ;
        RECT 2958.800 2316.380 2961.800 2316.390 ;
        RECT -42.180 2313.380 2961.800 2316.380 ;
        RECT -42.180 2313.370 -39.180 2313.380 ;
        RECT 2958.800 2313.370 2961.800 2313.380 ;
        RECT -42.180 2136.380 -39.180 2136.390 ;
        RECT 2958.800 2136.380 2961.800 2136.390 ;
        RECT -42.180 2133.380 2961.800 2136.380 ;
        RECT -42.180 2133.370 -39.180 2133.380 ;
        RECT 2958.800 2133.370 2961.800 2133.380 ;
        RECT -42.180 1956.380 -39.180 1956.390 ;
        RECT 2958.800 1956.380 2961.800 1956.390 ;
        RECT -42.180 1953.380 2961.800 1956.380 ;
        RECT -42.180 1953.370 -39.180 1953.380 ;
        RECT 2958.800 1953.370 2961.800 1953.380 ;
        RECT -42.180 1776.380 -39.180 1776.390 ;
        RECT 2958.800 1776.380 2961.800 1776.390 ;
        RECT -42.180 1773.380 2961.800 1776.380 ;
        RECT -42.180 1773.370 -39.180 1773.380 ;
        RECT 2958.800 1773.370 2961.800 1773.380 ;
        RECT -42.180 1596.380 -39.180 1596.390 ;
        RECT 2958.800 1596.380 2961.800 1596.390 ;
        RECT -42.180 1593.380 2961.800 1596.380 ;
        RECT -42.180 1593.370 -39.180 1593.380 ;
        RECT 2958.800 1593.370 2961.800 1593.380 ;
        RECT -42.180 1416.380 -39.180 1416.390 ;
        RECT 2958.800 1416.380 2961.800 1416.390 ;
        RECT -42.180 1413.380 2961.800 1416.380 ;
        RECT -42.180 1413.370 -39.180 1413.380 ;
        RECT 2958.800 1413.370 2961.800 1413.380 ;
        RECT -42.180 1236.380 -39.180 1236.390 ;
        RECT 2958.800 1236.380 2961.800 1236.390 ;
        RECT -42.180 1233.380 2961.800 1236.380 ;
        RECT -42.180 1233.370 -39.180 1233.380 ;
        RECT 2958.800 1233.370 2961.800 1233.380 ;
        RECT -42.180 1056.380 -39.180 1056.390 ;
        RECT 2958.800 1056.380 2961.800 1056.390 ;
        RECT -42.180 1053.380 2961.800 1056.380 ;
        RECT -42.180 1053.370 -39.180 1053.380 ;
        RECT 2958.800 1053.370 2961.800 1053.380 ;
        RECT -42.180 876.380 -39.180 876.390 ;
        RECT 2958.800 876.380 2961.800 876.390 ;
        RECT -42.180 873.380 2961.800 876.380 ;
        RECT -42.180 873.370 -39.180 873.380 ;
        RECT 2958.800 873.370 2961.800 873.380 ;
        RECT -42.180 696.380 -39.180 696.390 ;
        RECT 2958.800 696.380 2961.800 696.390 ;
        RECT -42.180 693.380 2961.800 696.380 ;
        RECT -42.180 693.370 -39.180 693.380 ;
        RECT 2958.800 693.370 2961.800 693.380 ;
        RECT -42.180 516.380 -39.180 516.390 ;
        RECT 2958.800 516.380 2961.800 516.390 ;
        RECT -42.180 513.380 2961.800 516.380 ;
        RECT -42.180 513.370 -39.180 513.380 ;
        RECT 2958.800 513.370 2961.800 513.380 ;
        RECT -42.180 336.380 -39.180 336.390 ;
        RECT 2958.800 336.380 2961.800 336.390 ;
        RECT -42.180 333.380 2961.800 336.380 ;
        RECT -42.180 333.370 -39.180 333.380 ;
        RECT 2958.800 333.370 2961.800 333.380 ;
        RECT -42.180 156.380 -39.180 156.390 ;
        RECT 2958.800 156.380 2961.800 156.390 ;
        RECT -42.180 153.380 2961.800 156.380 ;
        RECT -42.180 153.370 -39.180 153.380 ;
        RECT 2958.800 153.370 2961.800 153.380 ;
        RECT -42.180 -33.820 -39.180 -33.810 ;
        RECT 2958.800 -33.820 2961.800 -33.810 ;
        RECT -42.180 -36.820 2961.800 -33.820 ;
        RECT -42.180 -36.830 -39.180 -36.820 ;
        RECT 2958.800 -36.830 2961.800 -36.820 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 10.520 15.795 2849.180 3394.205 ;
      LAYER li1 ;
        RECT 2850.765 2334.185 2850.935 2341.495 ;
        RECT 2850.765 2313.785 2850.935 2326.875 ;
        RECT 2849.845 1883.345 2850.015 1914.115 ;
        RECT 2850.765 1605.565 2850.935 1652.655 ;
        RECT 2851.685 1573.605 2851.855 1605.735 ;
        RECT 2852.605 1546.065 2852.775 1573.775 ;
        RECT 2850.305 1501.185 2850.475 1514.615 ;
        RECT 2851.225 1514.445 2851.395 1545.895 ;
        RECT 2851.225 1440.665 2851.395 1475.855 ;
        RECT 2852.145 1349.545 2852.315 1440.835 ;
        RECT 2850.305 1252.305 2850.475 1332.035 ;
        RECT 2849.845 1025.865 2850.015 1143.675 ;
        RECT 2851.685 1143.505 2851.855 1236.495 ;
        RECT 2849.845 1012.945 2850.015 1024.675 ;
        RECT 2849.845 887.145 2850.015 962.455 ;
        RECT 2850.305 670.905 2850.475 845.495 ;
        RECT 2852.605 845.325 2852.775 887.315 ;
        RECT 2850.765 283.305 2850.935 383.775 ;
        RECT 2849.385 211.565 2850.015 211.735 ;
        RECT 2849.385 90.695 2849.555 211.565 ;
        RECT 2849.385 90.525 2850.015 90.695 ;
        RECT 2849.845 40.545 2850.015 90.525 ;
        RECT 1689.725 4.845 1689.895 8.755 ;
        RECT 1744.925 5.865 1745.095 8.755 ;
      LAYER mcon ;
        RECT 2850.765 2341.325 2850.935 2341.495 ;
        RECT 2850.765 2326.705 2850.935 2326.875 ;
        RECT 2849.845 1913.945 2850.015 1914.115 ;
        RECT 2850.765 1652.485 2850.935 1652.655 ;
        RECT 2851.685 1605.565 2851.855 1605.735 ;
        RECT 2852.605 1573.605 2852.775 1573.775 ;
        RECT 2851.225 1545.725 2851.395 1545.895 ;
        RECT 2850.305 1514.445 2850.475 1514.615 ;
        RECT 2851.225 1475.685 2851.395 1475.855 ;
        RECT 2852.145 1440.665 2852.315 1440.835 ;
        RECT 2850.305 1331.865 2850.475 1332.035 ;
        RECT 2851.685 1236.325 2851.855 1236.495 ;
        RECT 2849.845 1143.505 2850.015 1143.675 ;
        RECT 2849.845 1024.505 2850.015 1024.675 ;
        RECT 2849.845 962.285 2850.015 962.455 ;
        RECT 2852.605 887.145 2852.775 887.315 ;
        RECT 2850.305 845.325 2850.475 845.495 ;
        RECT 2850.765 383.605 2850.935 383.775 ;
        RECT 2849.845 211.565 2850.015 211.735 ;
        RECT 1689.725 8.585 1689.895 8.755 ;
        RECT 1744.925 8.585 1745.095 8.755 ;
      LAYER met1 ;
        RECT 10.520 9.460 2849.180 3394.360 ;
      LAYER met1 ;
        RECT 2849.770 2341.480 2850.090 2341.540 ;
        RECT 2850.705 2341.480 2850.995 2341.525 ;
        RECT 2849.770 2341.340 2850.995 2341.480 ;
        RECT 2849.770 2341.280 2850.090 2341.340 ;
        RECT 2850.705 2341.295 2850.995 2341.340 ;
        RECT 2850.230 2334.340 2850.550 2334.400 ;
        RECT 2850.705 2334.340 2850.995 2334.385 ;
        RECT 2850.230 2334.200 2850.995 2334.340 ;
        RECT 2850.230 2334.140 2850.550 2334.200 ;
        RECT 2850.705 2334.155 2850.995 2334.200 ;
        RECT 2850.230 2326.860 2850.550 2326.920 ;
        RECT 2850.705 2326.860 2850.995 2326.905 ;
        RECT 2850.230 2326.720 2850.995 2326.860 ;
        RECT 2850.230 2326.660 2850.550 2326.720 ;
        RECT 2850.705 2326.675 2850.995 2326.720 ;
        RECT 2850.230 2313.940 2850.550 2314.000 ;
        RECT 2850.705 2313.940 2850.995 2313.985 ;
        RECT 2850.230 2313.800 2850.995 2313.940 ;
        RECT 2850.230 2313.740 2850.550 2313.800 ;
        RECT 2850.705 2313.755 2850.995 2313.800 ;
        RECT 2850.230 1973.260 2850.550 1973.320 ;
        RECT 2851.150 1973.260 2851.470 1973.320 ;
        RECT 2850.230 1973.120 2851.470 1973.260 ;
        RECT 2850.230 1973.060 2850.550 1973.120 ;
        RECT 2851.150 1973.060 2851.470 1973.120 ;
        RECT 2849.770 1941.980 2850.090 1942.040 ;
        RECT 2851.150 1941.980 2851.470 1942.040 ;
        RECT 2849.770 1941.840 2851.470 1941.980 ;
        RECT 2849.770 1941.780 2850.090 1941.840 ;
        RECT 2851.150 1941.780 2851.470 1941.840 ;
        RECT 2849.770 1914.100 2850.090 1914.160 ;
        RECT 2849.575 1913.960 2850.090 1914.100 ;
        RECT 2849.770 1913.900 2850.090 1913.960 ;
        RECT 2849.770 1883.500 2850.090 1883.560 ;
        RECT 2849.575 1883.360 2850.090 1883.500 ;
        RECT 2849.770 1883.300 2850.090 1883.360 ;
        RECT 2850.230 1811.760 2850.550 1811.820 ;
        RECT 2851.150 1811.760 2851.470 1811.820 ;
        RECT 2850.230 1811.620 2851.470 1811.760 ;
        RECT 2850.230 1811.560 2850.550 1811.620 ;
        RECT 2851.150 1811.560 2851.470 1811.620 ;
        RECT 2850.690 1790.480 2851.010 1790.740 ;
        RECT 2850.780 1789.720 2850.920 1790.480 ;
        RECT 2850.690 1789.460 2851.010 1789.720 ;
        RECT 2849.770 1652.640 2850.090 1652.700 ;
        RECT 2850.705 1652.640 2850.995 1652.685 ;
        RECT 2849.770 1652.500 2850.995 1652.640 ;
        RECT 2849.770 1652.440 2850.090 1652.500 ;
        RECT 2850.705 1652.455 2850.995 1652.500 ;
        RECT 2850.705 1605.720 2850.995 1605.765 ;
        RECT 2851.625 1605.720 2851.915 1605.765 ;
        RECT 2850.705 1605.580 2851.915 1605.720 ;
        RECT 2850.705 1605.535 2850.995 1605.580 ;
        RECT 2851.625 1605.535 2851.915 1605.580 ;
        RECT 2851.625 1573.760 2851.915 1573.805 ;
        RECT 2852.545 1573.760 2852.835 1573.805 ;
        RECT 2851.625 1573.620 2852.835 1573.760 ;
        RECT 2851.625 1573.575 2851.915 1573.620 ;
        RECT 2852.545 1573.575 2852.835 1573.620 ;
        RECT 2852.545 1546.220 2852.835 1546.265 ;
        RECT 2851.240 1546.080 2852.835 1546.220 ;
        RECT 2851.240 1545.925 2851.380 1546.080 ;
        RECT 2852.545 1546.035 2852.835 1546.080 ;
        RECT 2851.165 1545.695 2851.455 1545.925 ;
        RECT 2850.245 1514.600 2850.535 1514.645 ;
        RECT 2851.165 1514.600 2851.455 1514.645 ;
        RECT 2850.245 1514.460 2851.455 1514.600 ;
        RECT 2850.245 1514.415 2850.535 1514.460 ;
        RECT 2851.165 1514.415 2851.455 1514.460 ;
        RECT 2850.245 1501.340 2850.535 1501.385 ;
        RECT 2851.610 1501.340 2851.930 1501.400 ;
        RECT 2850.245 1501.200 2851.930 1501.340 ;
        RECT 2850.245 1501.155 2850.535 1501.200 ;
        RECT 2851.610 1501.140 2851.930 1501.200 ;
        RECT 2851.165 1475.840 2851.455 1475.885 ;
        RECT 2851.610 1475.840 2851.930 1475.900 ;
        RECT 2851.165 1475.700 2851.930 1475.840 ;
        RECT 2851.165 1475.655 2851.455 1475.700 ;
        RECT 2851.610 1475.640 2851.930 1475.700 ;
        RECT 2851.165 1440.820 2851.455 1440.865 ;
        RECT 2852.085 1440.820 2852.375 1440.865 ;
        RECT 2851.165 1440.680 2852.375 1440.820 ;
        RECT 2851.165 1440.635 2851.455 1440.680 ;
        RECT 2852.085 1440.635 2852.375 1440.680 ;
        RECT 2849.770 1349.700 2850.090 1349.760 ;
        RECT 2852.085 1349.700 2852.375 1349.745 ;
        RECT 2849.770 1349.560 2852.375 1349.700 ;
        RECT 2849.770 1349.500 2850.090 1349.560 ;
        RECT 2852.085 1349.515 2852.375 1349.560 ;
        RECT 2849.770 1332.020 2850.090 1332.080 ;
        RECT 2850.245 1332.020 2850.535 1332.065 ;
        RECT 2849.770 1331.880 2850.535 1332.020 ;
        RECT 2849.770 1331.820 2850.090 1331.880 ;
        RECT 2850.245 1331.835 2850.535 1331.880 ;
        RECT 2849.770 1252.460 2850.090 1252.520 ;
        RECT 2850.245 1252.460 2850.535 1252.505 ;
        RECT 2849.770 1252.320 2850.535 1252.460 ;
        RECT 2849.770 1252.260 2850.090 1252.320 ;
        RECT 2850.245 1252.275 2850.535 1252.320 ;
        RECT 2849.770 1236.480 2850.090 1236.540 ;
        RECT 2851.625 1236.480 2851.915 1236.525 ;
        RECT 2849.770 1236.340 2851.915 1236.480 ;
        RECT 2849.770 1236.280 2850.090 1236.340 ;
        RECT 2851.625 1236.295 2851.915 1236.340 ;
        RECT 2849.785 1143.660 2850.075 1143.705 ;
        RECT 2851.625 1143.660 2851.915 1143.705 ;
        RECT 2849.785 1143.520 2851.915 1143.660 ;
        RECT 2849.785 1143.475 2850.075 1143.520 ;
        RECT 2851.625 1143.475 2851.915 1143.520 ;
        RECT 2849.785 1026.020 2850.075 1026.065 ;
        RECT 2849.400 1025.880 2850.075 1026.020 ;
        RECT 2849.400 1024.660 2849.540 1025.880 ;
        RECT 2849.785 1025.835 2850.075 1025.880 ;
        RECT 2849.785 1024.660 2850.075 1024.705 ;
        RECT 2849.400 1024.520 2850.075 1024.660 ;
        RECT 2849.785 1024.475 2850.075 1024.520 ;
        RECT 2849.770 1013.100 2850.090 1013.160 ;
        RECT 2849.575 1012.960 2850.090 1013.100 ;
        RECT 2849.770 1012.900 2850.090 1012.960 ;
        RECT 2849.770 962.440 2850.090 962.500 ;
        RECT 2849.770 962.300 2850.285 962.440 ;
        RECT 2849.770 962.240 2850.090 962.300 ;
        RECT 2849.785 887.300 2850.075 887.345 ;
        RECT 2852.545 887.300 2852.835 887.345 ;
        RECT 2849.785 887.160 2852.835 887.300 ;
        RECT 2849.785 887.115 2850.075 887.160 ;
        RECT 2852.545 887.115 2852.835 887.160 ;
        RECT 2850.245 845.480 2850.535 845.525 ;
        RECT 2852.545 845.480 2852.835 845.525 ;
        RECT 2850.245 845.340 2852.835 845.480 ;
        RECT 2850.245 845.295 2850.535 845.340 ;
        RECT 2852.545 845.295 2852.835 845.340 ;
        RECT 2849.770 671.060 2850.090 671.120 ;
        RECT 2850.245 671.060 2850.535 671.105 ;
        RECT 2849.770 670.920 2850.535 671.060 ;
        RECT 2849.770 670.860 2850.090 670.920 ;
        RECT 2850.245 670.875 2850.535 670.920 ;
        RECT 2849.770 383.760 2850.090 383.820 ;
        RECT 2850.705 383.760 2850.995 383.805 ;
        RECT 2849.770 383.620 2850.995 383.760 ;
        RECT 2849.770 383.560 2850.090 383.620 ;
        RECT 2850.705 383.575 2850.995 383.620 ;
        RECT 2849.770 283.460 2850.090 283.520 ;
        RECT 2850.705 283.460 2850.995 283.505 ;
        RECT 2849.770 283.320 2850.995 283.460 ;
        RECT 2849.770 283.260 2850.090 283.320 ;
        RECT 2850.705 283.275 2850.995 283.320 ;
        RECT 2849.770 211.720 2850.090 211.780 ;
        RECT 2849.575 211.580 2850.090 211.720 ;
        RECT 2849.770 211.520 2850.090 211.580 ;
        RECT 2849.770 40.700 2850.090 40.760 ;
        RECT 2849.575 40.560 2850.090 40.700 ;
        RECT 2849.770 40.500 2850.090 40.560 ;
        RECT 1689.665 8.740 1689.955 8.785 ;
        RECT 1744.865 8.740 1745.155 8.785 ;
        RECT 1689.665 8.600 1745.155 8.740 ;
        RECT 1689.665 8.555 1689.955 8.600 ;
        RECT 1744.865 8.555 1745.155 8.600 ;
        RECT 1789.930 6.360 1790.250 6.420 ;
        RECT 1826.270 6.360 1826.590 6.420 ;
        RECT 1789.930 6.220 1826.590 6.360 ;
        RECT 1789.930 6.160 1790.250 6.220 ;
        RECT 1826.270 6.160 1826.590 6.220 ;
        RECT 1744.865 6.020 1745.155 6.065 ;
        RECT 1770.150 6.020 1770.470 6.080 ;
        RECT 1744.865 5.880 1770.470 6.020 ;
        RECT 1744.865 5.835 1745.155 5.880 ;
        RECT 1770.150 5.820 1770.470 5.880 ;
        RECT 1658.370 5.000 1658.690 5.060 ;
        RECT 1648.340 4.860 1658.690 5.000 ;
        RECT 1644.110 4.660 1644.430 4.720 ;
        RECT 1648.340 4.660 1648.480 4.860 ;
        RECT 1658.370 4.800 1658.690 4.860 ;
        RECT 1679.070 5.000 1679.390 5.060 ;
        RECT 1689.665 5.000 1689.955 5.045 ;
        RECT 1679.070 4.860 1689.955 5.000 ;
        RECT 1679.070 4.800 1679.390 4.860 ;
        RECT 1689.665 4.815 1689.955 4.860 ;
        RECT 1644.110 4.520 1648.480 4.660 ;
        RECT 1644.110 4.460 1644.430 4.520 ;
        RECT 2030.510 3.980 2030.830 4.040 ;
        RECT 2035.110 3.980 2035.430 4.040 ;
        RECT 2030.510 3.840 2035.430 3.980 ;
        RECT 2030.510 3.780 2030.830 3.840 ;
        RECT 2035.110 3.780 2035.430 3.840 ;
      LAYER via ;
        RECT 2849.800 2341.280 2850.060 2341.540 ;
        RECT 2850.260 2334.140 2850.520 2334.400 ;
        RECT 2850.260 2326.660 2850.520 2326.920 ;
        RECT 2850.260 2313.740 2850.520 2314.000 ;
        RECT 2850.260 1973.060 2850.520 1973.320 ;
        RECT 2851.180 1973.060 2851.440 1973.320 ;
        RECT 2849.800 1941.780 2850.060 1942.040 ;
        RECT 2851.180 1941.780 2851.440 1942.040 ;
        RECT 2849.800 1913.900 2850.060 1914.160 ;
        RECT 2849.800 1883.300 2850.060 1883.560 ;
        RECT 2850.260 1811.560 2850.520 1811.820 ;
        RECT 2851.180 1811.560 2851.440 1811.820 ;
        RECT 2850.720 1790.480 2850.980 1790.740 ;
        RECT 2850.720 1789.460 2850.980 1789.720 ;
        RECT 2849.800 1652.440 2850.060 1652.700 ;
        RECT 2851.640 1501.140 2851.900 1501.400 ;
        RECT 2851.640 1475.640 2851.900 1475.900 ;
        RECT 2849.800 1349.500 2850.060 1349.760 ;
        RECT 2849.800 1331.820 2850.060 1332.080 ;
        RECT 2849.800 1252.260 2850.060 1252.520 ;
        RECT 2849.800 1236.280 2850.060 1236.540 ;
        RECT 2849.800 1012.900 2850.060 1013.160 ;
        RECT 2849.800 962.240 2850.060 962.500 ;
        RECT 2849.800 670.860 2850.060 671.120 ;
        RECT 2849.800 383.560 2850.060 383.820 ;
        RECT 2849.800 283.260 2850.060 283.520 ;
        RECT 2849.800 211.520 2850.060 211.780 ;
        RECT 2849.800 40.500 2850.060 40.760 ;
        RECT 1789.960 6.160 1790.220 6.420 ;
        RECT 1826.300 6.160 1826.560 6.420 ;
        RECT 1770.180 5.820 1770.440 6.080 ;
        RECT 1644.140 4.460 1644.400 4.720 ;
        RECT 1658.400 4.800 1658.660 5.060 ;
        RECT 1679.100 4.800 1679.360 5.060 ;
        RECT 2030.540 3.780 2030.800 4.040 ;
        RECT 2035.140 3.780 2035.400 4.040 ;
      LAYER met2 ;
        RECT 19.350 3400.720 53.570 3401.000 ;
        RECT 54.410 3400.720 151.550 3401.000 ;
        RECT 152.390 3400.720 249.990 3401.000 ;
        RECT 250.830 3400.720 347.970 3401.000 ;
        RECT 348.810 3400.720 446.410 3401.000 ;
        RECT 447.250 3400.720 544.850 3401.000 ;
        RECT 545.690 3400.720 642.830 3401.000 ;
        RECT 643.670 3400.720 741.270 3401.000 ;
        RECT 742.110 3400.720 839.710 3401.000 ;
        RECT 840.550 3400.720 937.690 3401.000 ;
        RECT 938.530 3400.720 1036.130 3401.000 ;
        RECT 1036.970 3400.720 1134.570 3401.000 ;
        RECT 1135.410 3400.720 1232.550 3401.000 ;
        RECT 1233.390 3400.720 1330.990 3401.000 ;
        RECT 1331.830 3400.720 1429.430 3401.000 ;
        RECT 1430.270 3400.720 1527.410 3401.000 ;
        RECT 1528.250 3400.720 1625.850 3401.000 ;
        RECT 1626.690 3400.720 1724.290 3401.000 ;
        RECT 1725.130 3400.720 1822.270 3401.000 ;
        RECT 1823.110 3400.720 1920.710 3401.000 ;
        RECT 1921.550 3400.720 2019.150 3401.000 ;
        RECT 2019.990 3400.720 2117.130 3401.000 ;
        RECT 2117.970 3400.720 2215.570 3401.000 ;
        RECT 2216.410 3400.720 2314.010 3401.000 ;
        RECT 2314.850 3400.720 2411.990 3401.000 ;
        RECT 2412.830 3400.720 2510.430 3401.000 ;
        RECT 2511.270 3400.720 2608.870 3401.000 ;
        RECT 2609.710 3400.720 2706.850 3401.000 ;
        RECT 2707.690 3400.720 2805.290 3401.000 ;
        RECT 2806.130 3400.720 2840.810 3401.000 ;
        RECT 19.350 15.600 2840.810 3400.720 ;
      LAYER met2 ;
        RECT 2851.630 2518.450 2851.910 2518.565 ;
        RECT 2848.480 2518.310 2851.910 2518.450 ;
        RECT 2848.480 2341.650 2848.620 2518.310 ;
        RECT 2851.630 2518.195 2851.910 2518.310 ;
        RECT 2848.480 2341.570 2850.000 2341.650 ;
        RECT 2848.480 2341.510 2850.060 2341.570 ;
        RECT 2849.800 2341.250 2850.060 2341.510 ;
        RECT 2850.260 2334.110 2850.520 2334.430 ;
        RECT 2850.320 2326.950 2850.460 2334.110 ;
        RECT 2850.260 2326.630 2850.520 2326.950 ;
        RECT 2850.260 2313.710 2850.520 2314.030 ;
        RECT 2850.320 2307.650 2850.460 2313.710 ;
        RECT 2849.400 2307.510 2850.460 2307.650 ;
        RECT 2849.400 2287.250 2849.540 2307.510 ;
        RECT 2848.480 2287.110 2849.540 2287.250 ;
        RECT 2848.480 1997.570 2848.620 2287.110 ;
        RECT 2848.480 1997.430 2849.080 1997.570 ;
        RECT 2848.940 1981.930 2849.080 1997.430 ;
        RECT 2848.940 1981.790 2850.460 1981.930 ;
        RECT 2850.320 1973.350 2850.460 1981.790 ;
        RECT 2850.260 1973.030 2850.520 1973.350 ;
        RECT 2851.180 1973.030 2851.440 1973.350 ;
        RECT 2851.240 1942.070 2851.380 1973.030 ;
        RECT 2849.800 1941.810 2850.060 1942.070 ;
        RECT 2848.940 1941.750 2850.060 1941.810 ;
        RECT 2851.180 1941.750 2851.440 1942.070 ;
        RECT 2848.940 1941.670 2850.000 1941.750 ;
        RECT 2848.940 1914.610 2849.080 1941.670 ;
        RECT 2848.940 1914.470 2850.000 1914.610 ;
        RECT 2849.860 1914.190 2850.000 1914.470 ;
        RECT 2849.800 1913.870 2850.060 1914.190 ;
        RECT 2849.800 1883.500 2850.060 1883.590 ;
        RECT 2848.940 1883.360 2850.060 1883.500 ;
        RECT 2848.940 1881.970 2849.080 1883.360 ;
        RECT 2849.800 1883.270 2850.060 1883.360 ;
        RECT 2848.480 1881.830 2849.080 1881.970 ;
        RECT 2848.480 1847.970 2848.620 1881.830 ;
        RECT 2848.480 1847.830 2850.460 1847.970 ;
        RECT 2850.320 1811.850 2850.460 1847.830 ;
        RECT 2850.260 1811.530 2850.520 1811.850 ;
        RECT 2851.180 1811.530 2851.440 1811.850 ;
        RECT 2851.240 1810.570 2851.380 1811.530 ;
        RECT 2850.780 1810.430 2851.380 1810.570 ;
        RECT 2850.780 1790.770 2850.920 1810.430 ;
        RECT 2850.720 1790.450 2850.980 1790.770 ;
        RECT 2850.720 1789.430 2850.980 1789.750 ;
        RECT 2850.780 1739.340 2850.920 1789.430 ;
        RECT 2848.480 1739.200 2850.920 1739.340 ;
        RECT 2848.480 1701.600 2848.620 1739.200 ;
        RECT 2848.480 1701.460 2849.540 1701.600 ;
        RECT 2849.400 1679.330 2849.540 1701.460 ;
        RECT 2848.480 1679.190 2849.540 1679.330 ;
        RECT 2848.480 1653.490 2848.620 1679.190 ;
        RECT 2848.480 1653.350 2850.000 1653.490 ;
        RECT 2849.860 1652.730 2850.000 1653.350 ;
        RECT 2849.800 1652.410 2850.060 1652.730 ;
        RECT 2851.640 1501.110 2851.900 1501.430 ;
        RECT 2851.700 1475.930 2851.840 1501.110 ;
        RECT 2851.640 1475.610 2851.900 1475.930 ;
        RECT 2849.800 1349.530 2850.060 1349.790 ;
        RECT 2848.480 1349.470 2850.060 1349.530 ;
        RECT 2848.480 1349.390 2850.000 1349.470 ;
        RECT 2848.480 1335.250 2848.620 1349.390 ;
        RECT 2848.480 1335.110 2850.000 1335.250 ;
        RECT 2849.860 1332.110 2850.000 1335.110 ;
        RECT 2849.800 1331.790 2850.060 1332.110 ;
        RECT 2849.800 1252.290 2850.060 1252.550 ;
        RECT 2848.940 1252.230 2850.060 1252.290 ;
        RECT 2848.940 1252.150 2850.000 1252.230 ;
        RECT 2848.940 1241.410 2849.080 1252.150 ;
        RECT 2848.940 1241.270 2850.000 1241.410 ;
        RECT 2849.860 1236.570 2850.000 1241.270 ;
        RECT 2849.800 1236.250 2850.060 1236.570 ;
        RECT 2849.800 1012.930 2850.060 1013.190 ;
        RECT 2848.480 1012.870 2850.060 1012.930 ;
        RECT 2848.480 1012.790 2850.000 1012.870 ;
        RECT 2848.480 963.970 2848.620 1012.790 ;
        RECT 2848.480 963.830 2849.080 963.970 ;
        RECT 2848.940 963.290 2849.080 963.830 ;
        RECT 2848.940 963.150 2850.000 963.290 ;
        RECT 2849.860 962.530 2850.000 963.150 ;
        RECT 2849.800 962.210 2850.060 962.530 ;
        RECT 2849.800 671.060 2850.060 671.150 ;
        RECT 2848.480 670.920 2850.060 671.060 ;
        RECT 2848.480 385.290 2848.620 670.920 ;
        RECT 2849.800 670.830 2850.060 670.920 ;
        RECT 2848.480 385.150 2849.080 385.290 ;
        RECT 2848.940 383.930 2849.080 385.150 ;
        RECT 2848.940 383.850 2850.000 383.930 ;
        RECT 2848.940 383.790 2850.060 383.850 ;
        RECT 2849.800 383.530 2850.060 383.790 ;
        RECT 2848.480 283.830 2850.000 283.970 ;
        RECT 2848.480 215.970 2848.620 283.830 ;
        RECT 2849.860 283.550 2850.000 283.830 ;
        RECT 2849.800 283.230 2850.060 283.550 ;
        RECT 2848.480 215.830 2850.000 215.970 ;
        RECT 2849.860 211.810 2850.000 215.830 ;
        RECT 2849.800 211.490 2850.060 211.810 ;
        RECT 2849.800 40.530 2850.060 40.790 ;
      LAYER met2 ;
        RECT 19.350 15.340 621.560 15.600 ;
        RECT 621.820 15.340 889.740 15.600 ;
        RECT 890.000 15.340 1341.920 15.600 ;
        RECT 1342.180 15.340 2840.810 15.600 ;
        RECT 19.350 9.280 2840.810 15.340 ;
        RECT 19.350 9.000 28.270 9.280 ;
        RECT 29.110 9.000 75.650 9.280 ;
        RECT 76.490 9.000 123.030 9.280 ;
        RECT 123.870 9.000 170.410 9.280 ;
        RECT 171.250 9.000 218.250 9.280 ;
        RECT 219.090 9.000 265.630 9.280 ;
        RECT 266.470 9.000 313.010 9.280 ;
        RECT 313.850 9.000 360.390 9.280 ;
        RECT 361.230 9.000 408.230 9.280 ;
        RECT 409.070 9.000 455.610 9.280 ;
        RECT 456.450 9.000 502.990 9.280 ;
        RECT 503.830 9.000 550.370 9.280 ;
        RECT 551.210 9.000 598.210 9.280 ;
        RECT 599.050 9.000 645.590 9.280 ;
        RECT 646.430 9.000 692.970 9.280 ;
        RECT 693.810 9.000 740.810 9.280 ;
        RECT 741.650 9.000 788.190 9.280 ;
        RECT 789.030 9.000 835.570 9.280 ;
        RECT 836.410 9.000 882.950 9.280 ;
        RECT 883.790 9.000 930.790 9.280 ;
        RECT 931.630 9.000 978.170 9.280 ;
        RECT 979.010 9.000 1025.550 9.280 ;
        RECT 1026.390 9.000 1072.930 9.280 ;
        RECT 1073.770 9.000 1120.770 9.280 ;
        RECT 1121.610 9.000 1168.150 9.280 ;
        RECT 1168.990 9.000 1215.530 9.280 ;
        RECT 1216.370 9.000 1262.910 9.280 ;
        RECT 1263.750 9.000 1310.750 9.280 ;
        RECT 1311.590 9.000 1358.130 9.280 ;
        RECT 1358.970 9.000 1405.510 9.280 ;
        RECT 1406.350 9.000 1453.350 9.280 ;
        RECT 1454.190 9.000 1500.730 9.280 ;
        RECT 1501.570 9.000 1548.110 9.280 ;
        RECT 1548.950 9.000 1595.490 9.280 ;
        RECT 1596.330 9.000 1643.330 9.280 ;
        RECT 1644.170 9.000 1690.710 9.280 ;
        RECT 1691.550 9.000 1738.090 9.280 ;
        RECT 1738.930 9.000 1785.470 9.280 ;
        RECT 1786.310 9.000 1833.310 9.280 ;
        RECT 1834.150 9.000 1880.690 9.280 ;
        RECT 1881.530 9.000 1928.070 9.280 ;
        RECT 1928.910 9.000 1975.450 9.280 ;
        RECT 1976.290 9.000 2023.290 9.280 ;
        RECT 2024.130 9.000 2070.670 9.280 ;
        RECT 2071.510 9.000 2118.050 9.280 ;
        RECT 2118.890 9.000 2165.890 9.280 ;
        RECT 2166.730 9.000 2213.270 9.280 ;
        RECT 2214.110 9.000 2260.650 9.280 ;
        RECT 2261.490 9.000 2308.030 9.280 ;
        RECT 2308.870 9.000 2355.870 9.280 ;
        RECT 2356.710 9.000 2403.250 9.280 ;
        RECT 2404.090 9.000 2450.630 9.280 ;
        RECT 2451.470 9.000 2498.010 9.280 ;
        RECT 2498.850 9.000 2545.850 9.280 ;
        RECT 2546.690 9.000 2593.230 9.280 ;
        RECT 2594.070 9.000 2640.610 9.280 ;
        RECT 2641.450 9.000 2687.990 9.280 ;
        RECT 2688.830 9.000 2735.830 9.280 ;
        RECT 2736.670 9.000 2783.210 9.280 ;
        RECT 2784.050 9.000 2830.590 9.280 ;
        RECT 2831.430 9.000 2840.810 9.280 ;
      LAYER met2 ;
        RECT 2848.020 40.470 2850.060 40.530 ;
        RECT 2848.020 40.390 2850.000 40.470 ;
        RECT 2848.020 8.685 2848.160 40.390 ;
        RECT 1608.710 8.315 1608.990 8.685 ;
        RECT 1901.730 8.315 1902.010 8.685 ;
        RECT 2847.950 8.315 2848.230 8.685 ;
        RECT 1608.780 5.170 1608.920 8.315 ;
        RECT 1789.960 6.130 1790.220 6.450 ;
        RECT 1826.300 6.130 1826.560 6.450 ;
        RECT 1610.550 5.850 1610.830 5.965 ;
        RECT 1610.160 5.710 1610.830 5.850 ;
        RECT 1610.160 5.170 1610.300 5.710 ;
        RECT 1610.550 5.595 1610.830 5.710 ;
        RECT 1644.130 5.595 1644.410 5.965 ;
        RECT 1659.770 5.850 1660.050 5.965 ;
        RECT 1659.380 5.710 1660.050 5.850 ;
        RECT 1608.780 5.030 1610.300 5.170 ;
        RECT 1644.200 4.750 1644.340 5.595 ;
        RECT 1658.400 4.770 1658.660 5.090 ;
        RECT 1644.140 4.430 1644.400 4.750 ;
        RECT 1658.460 4.490 1658.600 4.770 ;
        RECT 1659.380 4.490 1659.520 5.710 ;
        RECT 1659.770 5.595 1660.050 5.710 ;
        RECT 1679.090 5.595 1679.370 5.965 ;
        RECT 1770.180 5.790 1770.440 6.110 ;
        RECT 1679.160 5.090 1679.300 5.595 ;
        RECT 1679.100 4.770 1679.360 5.090 ;
        RECT 1658.460 4.350 1659.520 4.490 ;
        RECT 1770.240 3.925 1770.380 5.790 ;
        RECT 1790.020 4.490 1790.160 6.130 ;
        RECT 1788.180 4.350 1790.160 4.490 ;
        RECT 1788.180 3.925 1788.320 4.350 ;
        RECT 1770.170 3.555 1770.450 3.925 ;
        RECT 1788.110 3.555 1788.390 3.925 ;
        RECT 1826.360 3.245 1826.500 6.130 ;
        RECT 1901.800 3.245 1901.940 8.315 ;
        RECT 2035.130 7.635 2035.410 8.005 ;
        RECT 2075.610 7.635 2075.890 8.005 ;
        RECT 2035.200 4.070 2035.340 7.635 ;
        RECT 2030.540 3.925 2030.800 4.070 ;
        RECT 2030.530 3.555 2030.810 3.925 ;
        RECT 2035.140 3.750 2035.400 4.070 ;
        RECT 2075.680 3.245 2075.820 7.635 ;
        RECT 1826.290 2.875 1826.570 3.245 ;
        RECT 1901.730 2.875 1902.010 3.245 ;
        RECT 2075.610 2.875 2075.890 3.245 ;
        RECT 2139.090 2.875 2139.370 3.245 ;
        RECT 2139.160 1.885 2139.300 2.875 ;
        RECT 2139.090 1.515 2139.370 1.885 ;
      LAYER via2 ;
        RECT 2851.630 2518.240 2851.910 2518.520 ;
        RECT 1608.710 8.360 1608.990 8.640 ;
        RECT 1901.730 8.360 1902.010 8.640 ;
        RECT 2847.950 8.360 2848.230 8.640 ;
        RECT 1610.550 5.640 1610.830 5.920 ;
        RECT 1644.130 5.640 1644.410 5.920 ;
        RECT 1659.770 5.640 1660.050 5.920 ;
        RECT 1679.090 5.640 1679.370 5.920 ;
        RECT 1770.170 3.600 1770.450 3.880 ;
        RECT 1788.110 3.600 1788.390 3.880 ;
        RECT 2035.130 7.680 2035.410 7.960 ;
        RECT 2075.610 7.680 2075.890 7.960 ;
        RECT 2030.530 3.600 2030.810 3.880 ;
        RECT 1826.290 2.920 1826.570 3.200 ;
        RECT 1901.730 2.920 1902.010 3.200 ;
        RECT 2075.610 2.920 2075.890 3.200 ;
        RECT 2139.090 2.920 2139.370 3.200 ;
        RECT 2139.090 1.560 2139.370 1.840 ;
      LAYER met3 ;
        RECT 9.000 3348.920 2851.000 3400.745 ;
        RECT 9.400 3347.520 2851.000 3348.920 ;
        RECT 9.000 3338.040 2851.000 3347.520 ;
        RECT 9.000 3336.640 2850.600 3338.040 ;
        RECT 9.000 3235.360 2851.000 3336.640 ;
        RECT 9.400 3233.960 2851.000 3235.360 ;
        RECT 9.000 3202.040 2851.000 3233.960 ;
        RECT 9.000 3200.640 2850.600 3202.040 ;
        RECT 9.000 3122.480 2851.000 3200.640 ;
        RECT 9.400 3121.080 2851.000 3122.480 ;
        RECT 9.000 3066.040 2851.000 3121.080 ;
        RECT 9.000 3064.640 2850.600 3066.040 ;
        RECT 9.000 3008.920 2851.000 3064.640 ;
        RECT 9.400 3007.520 2851.000 3008.920 ;
        RECT 9.000 2930.040 2851.000 3007.520 ;
        RECT 9.000 2928.640 2850.600 2930.040 ;
        RECT 9.000 2895.360 2851.000 2928.640 ;
        RECT 9.400 2893.960 2851.000 2895.360 ;
        RECT 9.000 2794.040 2851.000 2893.960 ;
        RECT 9.000 2792.640 2850.600 2794.040 ;
        RECT 9.000 2782.480 2851.000 2792.640 ;
        RECT 9.400 2781.080 2851.000 2782.480 ;
        RECT 9.000 2668.920 2851.000 2781.080 ;
        RECT 9.400 2667.520 2851.000 2668.920 ;
        RECT 9.000 2658.040 2851.000 2667.520 ;
        RECT 9.000 2656.640 2850.600 2658.040 ;
        RECT 9.000 2555.360 2851.000 2656.640 ;
        RECT 9.400 2553.960 2851.000 2555.360 ;
        RECT 9.000 2522.040 2851.000 2553.960 ;
        RECT 9.000 2520.640 2850.600 2522.040 ;
      LAYER met3 ;
        RECT 2851.000 2521.040 2855.000 2521.640 ;
      LAYER met3 ;
        RECT 9.000 2442.480 2851.000 2520.640 ;
      LAYER met3 ;
        RECT 2851.390 2518.545 2851.690 2521.040 ;
        RECT 2851.390 2518.230 2851.935 2518.545 ;
        RECT 2851.605 2518.215 2851.935 2518.230 ;
      LAYER met3 ;
        RECT 9.400 2441.080 2851.000 2442.480 ;
        RECT 9.000 2386.040 2851.000 2441.080 ;
        RECT 9.000 2384.640 2850.600 2386.040 ;
        RECT 9.000 2328.920 2851.000 2384.640 ;
        RECT 9.400 2327.520 2851.000 2328.920 ;
        RECT 9.000 2250.040 2851.000 2327.520 ;
        RECT 9.000 2248.640 2850.600 2250.040 ;
        RECT 9.000 2215.360 2851.000 2248.640 ;
        RECT 9.400 2213.960 2851.000 2215.360 ;
        RECT 9.000 2114.040 2851.000 2213.960 ;
        RECT 9.000 2112.640 2850.600 2114.040 ;
        RECT 9.000 2102.480 2851.000 2112.640 ;
        RECT 9.400 2101.080 2851.000 2102.480 ;
        RECT 9.000 1988.920 2851.000 2101.080 ;
        RECT 9.400 1987.520 2851.000 1988.920 ;
        RECT 9.000 1978.040 2851.000 1987.520 ;
        RECT 9.000 1976.640 2850.600 1978.040 ;
        RECT 9.000 1875.360 2851.000 1976.640 ;
        RECT 9.400 1873.960 2851.000 1875.360 ;
        RECT 9.000 1842.040 2851.000 1873.960 ;
        RECT 9.000 1840.640 2850.600 1842.040 ;
        RECT 9.000 1762.480 2851.000 1840.640 ;
        RECT 9.400 1761.080 2851.000 1762.480 ;
        RECT 9.000 1706.040 2851.000 1761.080 ;
        RECT 9.000 1704.640 2850.600 1706.040 ;
        RECT 9.000 1648.920 2851.000 1704.640 ;
        RECT 9.400 1647.520 2851.000 1648.920 ;
        RECT 9.000 1570.040 2851.000 1647.520 ;
        RECT 9.000 1568.640 2850.600 1570.040 ;
        RECT 9.000 1535.360 2851.000 1568.640 ;
        RECT 9.400 1533.960 2851.000 1535.360 ;
        RECT 9.000 1434.040 2851.000 1533.960 ;
        RECT 9.000 1432.640 2850.600 1434.040 ;
        RECT 9.000 1422.480 2851.000 1432.640 ;
        RECT 9.400 1421.080 2851.000 1422.480 ;
        RECT 9.000 1308.920 2851.000 1421.080 ;
        RECT 9.400 1307.520 2851.000 1308.920 ;
        RECT 9.000 1298.040 2851.000 1307.520 ;
        RECT 9.000 1296.640 2850.600 1298.040 ;
        RECT 9.000 1195.360 2851.000 1296.640 ;
        RECT 9.400 1193.960 2851.000 1195.360 ;
        RECT 9.000 1162.040 2851.000 1193.960 ;
        RECT 9.000 1160.640 2850.600 1162.040 ;
        RECT 9.000 1082.480 2851.000 1160.640 ;
        RECT 9.400 1081.080 2851.000 1082.480 ;
        RECT 9.000 1026.040 2851.000 1081.080 ;
        RECT 9.000 1024.640 2850.600 1026.040 ;
        RECT 9.000 968.920 2851.000 1024.640 ;
        RECT 9.400 967.520 2851.000 968.920 ;
        RECT 9.000 892.640 2851.000 967.520 ;
        RECT 9.000 892.360 2846.180 892.640 ;
        RECT 2846.390 892.360 2851.000 892.640 ;
        RECT 9.000 890.040 2851.000 892.360 ;
        RECT 9.000 888.640 2850.600 890.040 ;
        RECT 9.000 855.360 2851.000 888.640 ;
        RECT 9.400 853.960 2851.000 855.360 ;
        RECT 9.000 754.040 2851.000 853.960 ;
        RECT 9.000 752.640 2850.600 754.040 ;
        RECT 9.000 742.480 2851.000 752.640 ;
        RECT 9.400 741.080 2851.000 742.480 ;
        RECT 9.000 628.920 2851.000 741.080 ;
        RECT 9.400 627.520 2851.000 628.920 ;
        RECT 9.000 618.040 2851.000 627.520 ;
        RECT 9.000 616.640 2850.600 618.040 ;
        RECT 9.000 515.360 2851.000 616.640 ;
        RECT 9.400 513.960 2851.000 515.360 ;
        RECT 9.000 482.040 2851.000 513.960 ;
        RECT 9.000 480.640 2850.600 482.040 ;
        RECT 9.000 402.480 2851.000 480.640 ;
        RECT 9.400 401.080 2851.000 402.480 ;
        RECT 9.000 346.040 2851.000 401.080 ;
        RECT 9.000 344.640 2850.600 346.040 ;
        RECT 9.000 288.920 2851.000 344.640 ;
        RECT 9.400 287.520 2851.000 288.920 ;
        RECT 9.000 210.040 2851.000 287.520 ;
        RECT 9.000 208.640 2850.600 210.040 ;
        RECT 9.000 201.760 2851.000 208.640 ;
        RECT 9.000 201.480 19.020 201.760 ;
        RECT 19.230 201.480 2851.000 201.760 ;
        RECT 9.000 175.360 2851.000 201.480 ;
        RECT 9.400 173.960 2851.000 175.360 ;
        RECT 9.000 74.040 2851.000 173.960 ;
        RECT 9.000 72.640 2850.600 74.040 ;
        RECT 9.000 66.440 2851.000 72.640 ;
        RECT 9.000 66.160 100.370 66.440 ;
      LAYER met3 ;
        RECT 100.370 66.160 100.580 66.440 ;
      LAYER met3 ;
        RECT 100.580 66.160 2851.000 66.440 ;
        RECT 9.000 62.480 2851.000 66.160 ;
        RECT 9.400 61.080 2851.000 62.480 ;
        RECT 9.000 39.920 2851.000 61.080 ;
        RECT 9.000 39.640 99.980 39.920 ;
        RECT 100.190 39.640 2851.000 39.920 ;
        RECT 9.000 32.440 2851.000 39.640 ;
        RECT 9.000 32.160 1128.470 32.440 ;
      LAYER met3 ;
        RECT 1128.470 32.160 1128.750 32.440 ;
      LAYER met3 ;
        RECT 1128.750 32.160 2851.000 32.440 ;
        RECT 9.000 25.640 2851.000 32.160 ;
        RECT 9.000 25.360 1128.930 25.640 ;
      LAYER met3 ;
        RECT 1128.930 25.360 1129.140 25.640 ;
      LAYER met3 ;
        RECT 1129.140 25.360 2851.000 25.640 ;
        RECT 9.000 9.255 2851.000 25.360 ;
      LAYER met3 ;
        RECT 1553.230 8.650 1553.610 8.660 ;
        RECT 1608.685 8.650 1609.015 8.665 ;
        RECT 1553.230 8.350 1609.015 8.650 ;
        RECT 1553.230 8.340 1553.610 8.350 ;
        RECT 1608.685 8.335 1609.015 8.350 ;
        RECT 1901.705 8.650 1902.035 8.665 ;
        RECT 2847.925 8.660 2848.255 8.665 ;
        RECT 1928.590 8.650 1928.970 8.660 ;
        RECT 2847.670 8.650 2848.255 8.660 ;
        RECT 1901.705 8.350 1928.970 8.650 ;
        RECT 2847.470 8.350 2848.255 8.650 ;
        RECT 1901.705 8.335 1902.035 8.350 ;
        RECT 1928.590 8.340 1928.970 8.350 ;
        RECT 2847.670 8.340 2848.255 8.350 ;
        RECT 2847.925 8.335 2848.255 8.340 ;
        RECT 2035.105 7.970 2035.435 7.985 ;
        RECT 2075.585 7.970 2075.915 7.985 ;
        RECT 2035.105 7.670 2075.915 7.970 ;
        RECT 2035.105 7.655 2035.435 7.670 ;
        RECT 2075.585 7.655 2075.915 7.670 ;
        RECT 2797.070 7.290 2797.450 7.300 ;
        RECT 2800.750 7.290 2801.130 7.300 ;
        RECT 2797.070 6.990 2801.130 7.290 ;
        RECT 2797.070 6.980 2797.450 6.990 ;
        RECT 2800.750 6.980 2801.130 6.990 ;
        RECT 1610.525 5.930 1610.855 5.945 ;
        RECT 1641.550 5.930 1641.930 5.940 ;
        RECT 1610.525 5.630 1641.930 5.930 ;
        RECT 1610.525 5.615 1610.855 5.630 ;
        RECT 1641.550 5.620 1641.930 5.630 ;
        RECT 1642.470 5.930 1642.850 5.940 ;
        RECT 1644.105 5.930 1644.435 5.945 ;
        RECT 1642.470 5.630 1644.435 5.930 ;
        RECT 1642.470 5.620 1642.850 5.630 ;
        RECT 1644.105 5.615 1644.435 5.630 ;
        RECT 1659.745 5.930 1660.075 5.945 ;
        RECT 1679.065 5.930 1679.395 5.945 ;
        RECT 1659.745 5.630 1679.395 5.930 ;
        RECT 1659.745 5.615 1660.075 5.630 ;
        RECT 1679.065 5.615 1679.395 5.630 ;
        RECT 2418.950 5.930 2419.330 5.940 ;
        RECT 2570.750 5.930 2571.130 5.940 ;
        RECT 2418.950 5.630 2571.130 5.930 ;
        RECT 2418.950 5.620 2419.330 5.630 ;
        RECT 2570.750 5.620 2571.130 5.630 ;
        RECT 1770.145 3.890 1770.475 3.905 ;
        RECT 1788.085 3.890 1788.415 3.905 ;
        RECT 1770.145 3.590 1788.415 3.890 ;
        RECT 1770.145 3.575 1770.475 3.590 ;
        RECT 1788.085 3.575 1788.415 3.590 ;
        RECT 1929.510 3.890 1929.890 3.900 ;
        RECT 2030.505 3.890 2030.835 3.905 ;
        RECT 1929.510 3.590 2030.835 3.890 ;
        RECT 1929.510 3.580 1929.890 3.590 ;
        RECT 2030.505 3.575 2030.835 3.590 ;
        RECT 1826.265 3.210 1826.595 3.225 ;
        RECT 1901.705 3.210 1902.035 3.225 ;
        RECT 1826.265 2.910 1902.035 3.210 ;
        RECT 1826.265 2.895 1826.595 2.910 ;
        RECT 1901.705 2.895 1902.035 2.910 ;
        RECT 2075.585 3.210 2075.915 3.225 ;
        RECT 2139.065 3.210 2139.395 3.225 ;
        RECT 2075.585 2.910 2139.395 3.210 ;
        RECT 2075.585 2.895 2075.915 2.910 ;
        RECT 2139.065 2.895 2139.395 2.910 ;
        RECT 2139.065 1.850 2139.395 1.865 ;
        RECT 2214.710 1.850 2215.090 1.860 ;
        RECT 2139.065 1.550 2215.090 1.850 ;
        RECT 2139.065 1.535 2139.395 1.550 ;
        RECT 2214.710 1.540 2215.090 1.550 ;
      LAYER via3 ;
        RECT 1553.260 8.340 1553.580 8.660 ;
        RECT 1928.620 8.340 1928.940 8.660 ;
        RECT 2847.700 8.340 2848.020 8.660 ;
        RECT 2797.100 6.980 2797.420 7.300 ;
        RECT 2800.780 6.980 2801.100 7.300 ;
        RECT 1641.580 5.620 1641.900 5.940 ;
        RECT 1642.500 5.620 1642.820 5.940 ;
        RECT 2418.980 5.620 2419.300 5.940 ;
        RECT 2570.780 5.620 2571.100 5.940 ;
        RECT 1929.540 3.580 1929.860 3.900 ;
        RECT 2214.740 1.540 2215.060 1.860 ;
      LAYER met4 ;
        RECT 26.040 66.890 2792.440 3394.360 ;
        RECT 26.040 65.710 100.150 66.890 ;
        RECT 101.330 65.710 2792.440 66.890 ;
        RECT 26.040 39.945 2792.440 65.710 ;
        RECT 26.040 39.690 99.655 39.945 ;
        RECT 99.985 39.690 2792.440 39.945 ;
        RECT 26.040 38.510 99.230 39.690 ;
        RECT 100.410 38.510 2792.440 39.690 ;
        RECT 26.040 32.890 2792.440 38.510 ;
        RECT 26.040 31.710 1128.710 32.890 ;
        RECT 1129.890 31.710 2792.440 32.890 ;
        RECT 26.040 26.090 2792.440 31.710 ;
        RECT 26.040 24.910 1128.710 26.090 ;
        RECT 1129.890 24.910 2792.440 26.090 ;
        RECT 26.040 19.290 2792.440 24.910 ;
        RECT 26.040 18.110 621.100 19.290 ;
        RECT 622.280 18.110 889.280 19.290 ;
        RECT 890.460 18.110 1341.460 19.290 ;
      LAYER met4 ;
        RECT 1341.460 18.110 1342.640 19.290 ;
      LAYER met4 ;
        RECT 1342.640 18.110 2792.440 19.290 ;
      LAYER met4 ;
        RECT 2796.670 18.110 2797.850 19.290 ;
        RECT 2800.350 18.110 2801.530 19.290 ;
        RECT 2847.270 18.110 2848.450 19.290 ;
      LAYER met4 ;
        RECT 26.040 15.890 2792.440 18.110 ;
        RECT 26.040 15.640 74.390 15.890 ;
        RECT 75.570 15.640 144.310 15.890 ;
        RECT 145.490 15.640 261.150 15.890 ;
        RECT 262.330 15.640 374.310 15.890 ;
        RECT 375.490 15.640 381.670 15.890 ;
        RECT 382.850 15.640 392.710 15.890 ;
        RECT 393.890 15.640 411.110 15.890 ;
        RECT 412.290 15.640 457.110 15.890 ;
        RECT 458.290 15.640 473.670 15.890 ;
        RECT 474.850 15.640 478.270 15.890 ;
        RECT 479.450 15.640 483.790 15.890 ;
        RECT 484.970 15.640 513.230 15.890 ;
        RECT 514.410 15.640 626.390 15.890 ;
        RECT 627.570 15.640 630.070 15.890 ;
        RECT 631.250 15.640 635.590 15.890 ;
        RECT 636.770 15.640 678.830 15.890 ;
        RECT 680.010 15.640 682.510 15.890 ;
        RECT 683.690 15.640 729.430 15.890 ;
        RECT 730.610 15.640 768.070 15.890 ;
        RECT 769.250 15.640 771.750 15.890 ;
        RECT 772.930 15.640 776.350 15.890 ;
        RECT 777.530 15.640 780.030 15.890 ;
        RECT 781.210 15.640 790.150 15.890 ;
        RECT 791.330 15.640 970.470 15.890 ;
        RECT 971.650 15.640 977.830 15.890 ;
        RECT 979.010 15.640 1004.510 15.890 ;
        RECT 1005.690 15.640 1120.430 15.890 ;
        RECT 1121.610 15.640 1125.030 15.890 ;
        RECT 1126.210 15.640 1134.230 15.890 ;
        RECT 1135.410 15.640 1138.830 15.890 ;
        RECT 1140.010 15.640 1143.430 15.890 ;
        RECT 1144.610 15.640 1266.710 15.890 ;
        RECT 1267.890 15.640 1300.750 15.890 ;
        RECT 1301.930 15.640 1471.870 15.890 ;
        RECT 1473.050 15.640 1550.070 15.890 ;
      LAYER met4 ;
        RECT 1550.070 14.710 1551.250 15.890 ;
      LAYER met4 ;
        RECT 1551.250 15.640 1555.590 15.890 ;
        RECT 1556.770 15.640 1683.470 15.890 ;
        RECT 1684.650 15.640 1744.190 15.890 ;
        RECT 1745.370 15.640 1770.870 15.890 ;
        RECT 1772.050 15.640 1862.180 15.890 ;
        RECT 1863.360 15.640 2096.550 15.890 ;
        RECT 2097.730 15.640 2134.270 15.890 ;
        RECT 2135.450 15.640 2214.310 15.890 ;
      LAYER met4 ;
        RECT 2214.310 14.710 2215.490 15.890 ;
      LAYER met4 ;
        RECT 2215.490 15.640 2418.550 15.890 ;
      LAYER met4 ;
        RECT 2418.550 14.710 2419.730 15.890 ;
      LAYER met4 ;
        RECT 2419.730 15.640 2565.750 15.890 ;
        RECT 2566.930 15.640 2572.190 15.890 ;
      LAYER met4 ;
        RECT 2572.190 14.710 2573.370 15.890 ;
      LAYER met4 ;
        RECT 2573.370 15.640 2792.440 15.890 ;
      LAYER met4 ;
        RECT 1550.510 7.970 1550.810 14.710 ;
        RECT 1553.255 8.335 1553.585 8.665 ;
        RECT 1928.615 8.650 1928.945 8.665 ;
        RECT 1928.615 8.350 1929.850 8.650 ;
        RECT 1928.615 8.335 1928.945 8.350 ;
        RECT 1553.270 7.970 1553.570 8.335 ;
        RECT 1550.510 7.670 1553.570 7.970 ;
        RECT 1641.575 5.930 1641.905 5.945 ;
        RECT 1642.495 5.930 1642.825 5.945 ;
        RECT 1641.575 5.630 1642.825 5.930 ;
        RECT 1641.575 5.615 1641.905 5.630 ;
        RECT 1642.495 5.615 1642.825 5.630 ;
        RECT 1929.550 3.905 1929.850 8.350 ;
        RECT 1929.535 3.575 1929.865 3.905 ;
        RECT 2214.750 1.865 2215.050 14.710 ;
        RECT 2418.990 5.945 2419.290 14.710 ;
        RECT 2572.630 12.050 2572.930 14.710 ;
        RECT 2570.790 11.750 2572.930 12.050 ;
        RECT 2570.790 5.945 2571.090 11.750 ;
        RECT 2797.110 7.305 2797.410 18.110 ;
        RECT 2800.790 7.305 2801.090 18.110 ;
        RECT 2847.710 8.665 2848.010 18.110 ;
        RECT 2847.695 8.335 2848.025 8.665 ;
        RECT 2797.095 6.975 2797.425 7.305 ;
        RECT 2800.775 6.975 2801.105 7.305 ;
        RECT 2418.975 5.615 2419.305 5.945 ;
        RECT 2570.775 5.615 2571.105 5.945 ;
        RECT 2214.735 1.535 2215.065 1.865 ;
      LAYER met5 ;
        RECT 10.520 3306.380 2849.180 3326.460 ;
        RECT 10.520 3288.380 2849.180 3303.380 ;
        RECT 10.520 3270.380 2849.180 3285.380 ;
        RECT 10.520 3252.380 2849.180 3267.380 ;
        RECT 10.520 3216.380 2849.180 3249.380 ;
        RECT 10.520 3198.380 2849.180 3213.380 ;
        RECT 10.520 3180.380 2849.180 3195.380 ;
        RECT 10.520 3162.380 2849.180 3177.380 ;
        RECT 10.520 3126.380 2849.180 3159.380 ;
        RECT 10.520 3108.380 2849.180 3123.380 ;
        RECT 10.520 3090.380 2849.180 3105.380 ;
        RECT 10.520 3072.380 2849.180 3087.380 ;
        RECT 10.520 3036.380 2849.180 3069.380 ;
        RECT 10.520 3018.380 2849.180 3033.380 ;
        RECT 10.520 3000.380 2849.180 3015.380 ;
        RECT 10.520 2982.380 2849.180 2997.380 ;
        RECT 10.520 2946.380 2849.180 2979.380 ;
        RECT 10.520 2928.380 2849.180 2943.380 ;
        RECT 10.520 2910.380 2849.180 2925.380 ;
        RECT 10.520 2892.380 2849.180 2907.380 ;
        RECT 10.520 2856.380 2849.180 2889.380 ;
        RECT 10.520 2838.380 2849.180 2853.380 ;
        RECT 10.520 2820.380 2849.180 2835.380 ;
        RECT 10.520 2802.380 2849.180 2817.380 ;
        RECT 10.520 2766.380 2849.180 2799.380 ;
        RECT 10.520 2748.380 2849.180 2763.380 ;
        RECT 10.520 2730.380 2849.180 2745.380 ;
        RECT 10.520 2712.380 2849.180 2727.380 ;
        RECT 10.520 2676.380 2849.180 2709.380 ;
        RECT 10.520 2658.380 2849.180 2673.380 ;
        RECT 10.520 2640.380 2849.180 2655.380 ;
        RECT 10.520 2622.380 2849.180 2637.380 ;
        RECT 10.520 2586.380 2849.180 2619.380 ;
        RECT 10.520 2568.380 2849.180 2583.380 ;
        RECT 10.520 2550.380 2849.180 2565.380 ;
        RECT 10.520 2532.380 2849.180 2547.380 ;
        RECT 10.520 2496.380 2849.180 2529.380 ;
        RECT 10.520 2478.380 2849.180 2493.380 ;
        RECT 10.520 2460.380 2849.180 2475.380 ;
        RECT 10.520 2442.380 2849.180 2457.380 ;
        RECT 10.520 2406.380 2849.180 2439.380 ;
        RECT 10.520 2388.380 2849.180 2403.380 ;
        RECT 10.520 2370.380 2849.180 2385.380 ;
        RECT 10.520 2352.380 2849.180 2367.380 ;
        RECT 10.520 2316.380 2849.180 2349.380 ;
        RECT 10.520 2298.380 2849.180 2313.380 ;
        RECT 10.520 2280.380 2849.180 2295.380 ;
        RECT 10.520 2262.380 2849.180 2277.380 ;
        RECT 10.520 2226.380 2849.180 2259.380 ;
        RECT 10.520 2208.380 2849.180 2223.380 ;
        RECT 10.520 2190.380 2849.180 2205.380 ;
        RECT 10.520 2172.380 2849.180 2187.380 ;
        RECT 10.520 2136.380 2849.180 2169.380 ;
        RECT 10.520 2118.380 2849.180 2133.380 ;
        RECT 10.520 2100.380 2849.180 2115.380 ;
        RECT 10.520 2082.380 2849.180 2097.380 ;
        RECT 10.520 2046.380 2849.180 2079.380 ;
        RECT 10.520 2028.380 2849.180 2043.380 ;
        RECT 10.520 2010.380 2849.180 2025.380 ;
        RECT 10.520 1992.380 2849.180 2007.380 ;
        RECT 10.520 1956.380 2849.180 1989.380 ;
        RECT 10.520 1938.380 2849.180 1953.380 ;
        RECT 10.520 1920.380 2849.180 1935.380 ;
        RECT 10.520 1902.380 2849.180 1917.380 ;
        RECT 10.520 1866.380 2849.180 1899.380 ;
        RECT 10.520 1848.380 2849.180 1863.380 ;
        RECT 10.520 1830.380 2849.180 1845.380 ;
        RECT 10.520 1812.380 2849.180 1827.380 ;
        RECT 10.520 1776.380 2849.180 1809.380 ;
        RECT 10.520 1758.380 2849.180 1773.380 ;
        RECT 10.520 1740.380 2849.180 1755.380 ;
        RECT 10.520 1722.380 2849.180 1737.380 ;
        RECT 10.520 1686.380 2849.180 1719.380 ;
        RECT 10.520 1668.380 2849.180 1683.380 ;
        RECT 10.520 1650.380 2849.180 1665.380 ;
        RECT 10.520 1632.380 2849.180 1647.380 ;
        RECT 10.520 1596.380 2849.180 1629.380 ;
        RECT 10.520 1578.380 2849.180 1593.380 ;
        RECT 10.520 1560.380 2849.180 1575.380 ;
        RECT 10.520 1542.380 2849.180 1557.380 ;
        RECT 10.520 1506.380 2849.180 1539.380 ;
        RECT 10.520 1488.380 2849.180 1503.380 ;
        RECT 10.520 1470.380 2849.180 1485.380 ;
        RECT 10.520 1452.380 2849.180 1467.380 ;
        RECT 10.520 1416.380 2849.180 1449.380 ;
        RECT 10.520 1398.380 2849.180 1413.380 ;
        RECT 10.520 1380.380 2849.180 1395.380 ;
        RECT 10.520 1362.380 2849.180 1377.380 ;
        RECT 10.520 1326.380 2849.180 1359.380 ;
        RECT 10.520 1308.380 2849.180 1323.380 ;
        RECT 10.520 1290.380 2849.180 1305.380 ;
        RECT 10.520 1272.380 2849.180 1287.380 ;
        RECT 10.520 1236.380 2849.180 1269.380 ;
        RECT 10.520 1218.380 2849.180 1233.380 ;
        RECT 10.520 1200.380 2849.180 1215.380 ;
        RECT 10.520 1182.380 2849.180 1197.380 ;
        RECT 10.520 1146.380 2849.180 1179.380 ;
        RECT 10.520 1128.380 2849.180 1143.380 ;
        RECT 10.520 1110.380 2849.180 1125.380 ;
        RECT 10.520 1092.380 2849.180 1107.380 ;
        RECT 10.520 1056.380 2849.180 1089.380 ;
        RECT 10.520 1038.380 2849.180 1053.380 ;
        RECT 10.520 1020.380 2849.180 1035.380 ;
        RECT 10.520 1002.380 2849.180 1017.380 ;
        RECT 10.520 966.380 2849.180 999.380 ;
        RECT 10.520 948.380 2849.180 963.380 ;
        RECT 10.520 930.380 2849.180 945.380 ;
        RECT 10.520 912.380 2849.180 927.380 ;
        RECT 10.520 876.380 2849.180 909.380 ;
        RECT 10.520 858.380 2849.180 873.380 ;
        RECT 10.520 840.380 2849.180 855.380 ;
        RECT 10.520 822.380 2849.180 837.380 ;
        RECT 10.520 786.380 2849.180 819.380 ;
        RECT 10.520 768.380 2849.180 783.380 ;
        RECT 10.520 750.380 2849.180 765.380 ;
        RECT 10.520 732.380 2849.180 747.380 ;
        RECT 10.520 696.380 2849.180 729.380 ;
        RECT 10.520 678.380 2849.180 693.380 ;
        RECT 10.520 660.380 2849.180 675.380 ;
        RECT 10.520 642.380 2849.180 657.380 ;
        RECT 10.520 606.380 2849.180 639.380 ;
        RECT 10.520 588.380 2849.180 603.380 ;
        RECT 10.520 570.380 2849.180 585.380 ;
        RECT 10.520 552.380 2849.180 567.380 ;
        RECT 10.520 516.380 2849.180 549.380 ;
        RECT 10.520 498.380 2849.180 513.380 ;
        RECT 10.520 480.380 2849.180 495.380 ;
        RECT 10.520 462.380 2849.180 477.380 ;
        RECT 10.520 426.380 2849.180 459.380 ;
        RECT 10.520 408.380 2849.180 423.380 ;
        RECT 10.520 390.380 2849.180 405.380 ;
        RECT 10.520 372.380 2849.180 387.380 ;
        RECT 10.520 336.380 2849.180 369.380 ;
        RECT 10.520 318.380 2849.180 333.380 ;
        RECT 10.520 300.380 2849.180 315.380 ;
        RECT 10.520 282.380 2849.180 297.380 ;
        RECT 10.520 246.380 2849.180 279.380 ;
        RECT 10.520 228.380 2849.180 243.380 ;
        RECT 10.520 210.380 2849.180 225.380 ;
        RECT 10.520 192.380 2849.180 207.380 ;
        RECT 10.520 184.670 2849.180 189.380 ;
      LAYER met5 ;
        RECT 10.520 108.080 2849.180 109.680 ;
        RECT 1380.580 21.300 1398.740 22.900 ;
        RECT 1380.580 19.500 1382.180 21.300 ;
        RECT 1341.250 17.900 1382.180 19.500 ;
        RECT 1397.140 19.500 1398.740 21.300 ;
        RECT 2654.780 21.300 2664.660 22.900 ;
        RECT 1397.140 17.900 1551.460 19.500 ;
        RECT 1549.860 14.500 1551.460 17.900 ;
        RECT 2364.060 17.900 2419.940 19.500 ;
        RECT 2364.060 16.100 2365.660 17.900 ;
        RECT 2214.100 14.500 2365.660 16.100 ;
        RECT 2418.340 14.500 2419.940 17.900 ;
        RECT 2654.780 16.100 2656.380 21.300 ;
        RECT 2571.980 14.500 2656.380 16.100 ;
        RECT 2663.060 16.100 2664.660 21.300 ;
        RECT 2682.380 21.300 2706.060 22.900 ;
        RECT 2682.380 16.100 2683.980 21.300 ;
        RECT 2663.060 14.500 2683.980 16.100 ;
        RECT 2704.460 16.100 2706.060 21.300 ;
        RECT 2723.780 21.300 2747.460 22.900 ;
        RECT 2723.780 16.100 2725.380 21.300 ;
        RECT 2704.460 14.500 2725.380 16.100 ;
        RECT 2745.860 16.100 2747.460 21.300 ;
        RECT 2765.180 21.300 2791.620 22.900 ;
        RECT 2765.180 16.100 2766.780 21.300 ;
        RECT 2790.020 19.500 2791.620 21.300 ;
        RECT 2790.020 17.900 2798.060 19.500 ;
        RECT 2800.140 17.900 2848.660 19.500 ;
        RECT 2745.860 14.500 2766.780 16.100 ;
  END
END user_project_wrapper
END LIBRARY


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga
  CLASS BLOCK ;
  FOREIGN fpga ;
  ORIGIN 0.000 0.000 ;
  SIZE 2745.000 BY 3320.000 ;
  PIN gpio_east[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 59.200 2745.000 59.800 ;
    END
  END gpio_east[0]
  PIN gpio_east[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 177.520 2745.000 178.120 ;
    END
  END gpio_east[1]
  PIN gpio_east[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 295.840 2745.000 296.440 ;
    END
  END gpio_east[2]
  PIN gpio_east[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 414.840 2745.000 415.440 ;
    END
  END gpio_east[3]
  PIN gpio_east[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 533.160 2745.000 533.760 ;
    END
  END gpio_east[4]
  PIN gpio_east[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 651.480 2745.000 652.080 ;
    END
  END gpio_east[5]
  PIN gpio_east[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 770.480 2745.000 771.080 ;
    END
  END gpio_east[6]
  PIN gpio_east[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 888.800 2745.000 889.400 ;
    END
  END gpio_east[7]
  PIN gpio_east[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 1007.120 2745.000 1007.720 ;
    END
  END gpio_east[8]
  PIN gpio_east[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 1126.120 2745.000 1126.720 ;
    END
  END gpio_east[9]
  PIN gpio_north[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 44.250 3316.000 44.530 3320.000 ;
    END
  END gpio_north[0]
  PIN gpio_north[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 132.570 3316.000 132.850 3320.000 ;
    END
  END gpio_north[1]
  PIN gpio_north[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 220.890 3316.000 221.170 3320.000 ;
    END
  END gpio_north[2]
  PIN gpio_north[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 309.670 3316.000 309.950 3320.000 ;
    END
  END gpio_north[3]
  PIN gpio_north[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 397.990 3316.000 398.270 3320.000 ;
    END
  END gpio_north[4]
  PIN gpio_north[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 486.770 3316.000 487.050 3320.000 ;
    END
  END gpio_north[5]
  PIN gpio_north[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 575.090 3316.000 575.370 3320.000 ;
    END
  END gpio_north[6]
  PIN gpio_north[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 663.870 3316.000 664.150 3320.000 ;
    END
  END gpio_north[7]
  PIN gpio_north[8]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 752.190 3316.000 752.470 3320.000 ;
    END
  END gpio_north[8]
  PIN gpio_north[9]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 840.970 3316.000 841.250 3320.000 ;
    END
  END gpio_north[9]
  PIN gpio_south[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END gpio_south[0]
  PIN gpio_south[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END gpio_south[1]
  PIN gpio_south[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 4.000 ;
    END
  END gpio_south[2]
  PIN gpio_south[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 159.710 0.000 159.990 4.000 ;
    END
  END gpio_south[3]
  PIN gpio_south[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.530 4.000 ;
    END
  END gpio_south[4]
  PIN gpio_south[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END gpio_south[5]
  PIN gpio_south[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 4.000 ;
    END
  END gpio_south[6]
  PIN gpio_south[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 342.790 0.000 343.070 4.000 ;
    END
  END gpio_south[7]
  PIN gpio_west[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END gpio_west[0]
  PIN gpio_west[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END gpio_west[1]
  PIN gpio_west[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.200 4.000 331.800 ;
    END
  END gpio_west[2]
  PIN gpio_west[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END gpio_west[3]
  PIN gpio_west[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 597.080 4.000 597.680 ;
    END
  END gpio_west[4]
  PIN gpio_west[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 729.680 4.000 730.280 ;
    END
  END gpio_west[5]
  PIN gpio_west[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 862.280 4.000 862.880 ;
    END
  END gpio_west[6]
  PIN gpio_west[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 994.880 4.000 995.480 ;
    END
  END gpio_west[7]
  PIN gpio_west[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1128.160 4.000 1128.760 ;
    END
  END gpio_west[8]
  PIN gpio_west[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1260.760 4.000 1261.360 ;
    END
  END gpio_west[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1852.510 0.000 1852.790 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1898.050 0.000 1898.330 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1393.360 4.000 1393.960 ;
    END
  END wbs_ack_o
  PIN wbs_addr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1526.640 4.000 1527.240 ;
    END
  END wbs_addr_i[0]
  PIN wbs_addr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 1600.080 2745.000 1600.680 ;
    END
  END wbs_addr_i[10]
  PIN wbs_addr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2035.130 0.000 2035.410 4.000 ;
    END
  END wbs_addr_i[11]
  PIN wbs_addr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1791.840 4.000 1792.440 ;
    END
  END wbs_addr_i[12]
  PIN wbs_addr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2081.130 0.000 2081.410 4.000 ;
    END
  END wbs_addr_i[13]
  PIN wbs_addr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2126.670 0.000 2126.950 4.000 ;
    END
  END wbs_addr_i[14]
  PIN wbs_addr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2172.670 0.000 2172.950 4.000 ;
    END
  END wbs_addr_i[15]
  PIN wbs_addr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 1719.080 2745.000 1719.680 ;
    END
  END wbs_addr_i[16]
  PIN wbs_addr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1195.170 3316.000 1195.450 3320.000 ;
    END
  END wbs_addr_i[17]
  PIN wbs_addr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1283.490 3316.000 1283.770 3320.000 ;
    END
  END wbs_addr_i[18]
  PIN wbs_addr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 1837.400 2745.000 1838.000 ;
    END
  END wbs_addr_i[19]
  PIN wbs_addr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1659.240 4.000 1659.840 ;
    END
  END wbs_addr_i[1]
  PIN wbs_addr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2218.210 0.000 2218.490 4.000 ;
    END
  END wbs_addr_i[20]
  PIN wbs_addr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 1955.720 2745.000 1956.320 ;
    END
  END wbs_addr_i[21]
  PIN wbs_addr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1924.440 4.000 1925.040 ;
    END
  END wbs_addr_i[22]
  PIN wbs_addr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1372.270 3316.000 1372.550 3320.000 ;
    END
  END wbs_addr_i[23]
  PIN wbs_addr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1460.590 3316.000 1460.870 3320.000 ;
    END
  END wbs_addr_i[24]
  PIN wbs_addr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 2074.720 2745.000 2075.320 ;
    END
  END wbs_addr_i[25]
  PIN wbs_addr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1549.370 3316.000 1549.650 3320.000 ;
    END
  END wbs_addr_i[26]
  PIN wbs_addr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 2193.040 2745.000 2193.640 ;
    END
  END wbs_addr_i[27]
  PIN wbs_addr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2264.210 0.000 2264.490 4.000 ;
    END
  END wbs_addr_i[28]
  PIN wbs_addr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 2311.360 2745.000 2311.960 ;
    END
  END wbs_addr_i[29]
  PIN wbs_addr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 1244.440 2745.000 1245.040 ;
    END
  END wbs_addr_i[2]
  PIN wbs_addr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1637.690 3316.000 1637.970 3320.000 ;
    END
  END wbs_addr_i[30]
  PIN wbs_addr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 2430.360 2745.000 2430.960 ;
    END
  END wbs_addr_i[31]
  PIN wbs_addr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 1362.760 2745.000 1363.360 ;
    END
  END wbs_addr_i[3]
  PIN wbs_addr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 1481.760 2745.000 1482.360 ;
    END
  END wbs_addr_i[4]
  PIN wbs_addr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 929.290 3316.000 929.570 3320.000 ;
    END
  END wbs_addr_i[5]
  PIN wbs_addr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1943.590 0.000 1943.870 4.000 ;
    END
  END wbs_addr_i[6]
  PIN wbs_addr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1018.070 3316.000 1018.350 3320.000 ;
    END
  END wbs_addr_i[7]
  PIN wbs_addr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1989.590 0.000 1989.870 4.000 ;
    END
  END wbs_addr_i[8]
  PIN wbs_addr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1106.390 3316.000 1106.670 3320.000 ;
    END
  END wbs_addr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 2548.680 2745.000 2549.280 ;
    END
  END wbs_cyc_i
  PIN wbs_data_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1726.470 3316.000 1726.750 3320.000 ;
    END
  END wbs_data_i[0]
  PIN wbs_data_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1991.890 3316.000 1992.170 3320.000 ;
    END
  END wbs_data_i[10]
  PIN wbs_data_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2080.670 3316.000 2080.950 3320.000 ;
    END
  END wbs_data_i[11]
  PIN wbs_data_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2190.320 4.000 2190.920 ;
    END
  END wbs_data_i[12]
  PIN wbs_data_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2168.990 3316.000 2169.270 3320.000 ;
    END
  END wbs_data_i[13]
  PIN wbs_data_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2538.370 0.000 2538.650 4.000 ;
    END
  END wbs_data_i[14]
  PIN wbs_data_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 2786.000 2745.000 2786.600 ;
    END
  END wbs_data_i[15]
  PIN wbs_data_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2257.770 3316.000 2258.050 3320.000 ;
    END
  END wbs_data_i[16]
  PIN wbs_data_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2346.090 3316.000 2346.370 3320.000 ;
    END
  END wbs_data_i[17]
  PIN wbs_data_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 2904.320 2745.000 2904.920 ;
    END
  END wbs_data_i[18]
  PIN wbs_data_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 3022.640 2745.000 3023.240 ;
    END
  END wbs_data_i[19]
  PIN wbs_data_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1814.790 3316.000 1815.070 3320.000 ;
    END
  END wbs_data_i[1]
  PIN wbs_data_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2322.920 4.000 2323.520 ;
    END
  END wbs_data_i[20]
  PIN wbs_data_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2456.200 4.000 2456.800 ;
    END
  END wbs_data_i[21]
  PIN wbs_data_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2588.800 4.000 2589.400 ;
    END
  END wbs_data_i[22]
  PIN wbs_data_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 3141.640 2745.000 3142.240 ;
    END
  END wbs_data_i[23]
  PIN wbs_data_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2434.870 3316.000 2435.150 3320.000 ;
    END
  END wbs_data_i[24]
  PIN wbs_data_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2721.400 4.000 2722.000 ;
    END
  END wbs_data_i[25]
  PIN wbs_data_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2523.190 3316.000 2523.470 3320.000 ;
    END
  END wbs_data_i[26]
  PIN wbs_data_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 3259.960 2745.000 3260.560 ;
    END
  END wbs_data_i[27]
  PIN wbs_data_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2611.970 3316.000 2612.250 3320.000 ;
    END
  END wbs_data_i[28]
  PIN wbs_data_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2584.370 0.000 2584.650 4.000 ;
    END
  END wbs_data_i[29]
  PIN wbs_data_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2309.750 0.000 2310.030 4.000 ;
    END
  END wbs_data_i[2]
  PIN wbs_data_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2854.000 4.000 2854.600 ;
    END
  END wbs_data_i[30]
  PIN wbs_data_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2629.910 0.000 2630.190 4.000 ;
    END
  END wbs_data_i[31]
  PIN wbs_data_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2057.720 4.000 2058.320 ;
    END
  END wbs_data_i[3]
  PIN wbs_data_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1903.570 3316.000 1903.850 3320.000 ;
    END
  END wbs_data_i[4]
  PIN wbs_data_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2355.290 0.000 2355.570 4.000 ;
    END
  END wbs_data_i[5]
  PIN wbs_data_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2401.290 0.000 2401.570 4.000 ;
    END
  END wbs_data_i[6]
  PIN wbs_data_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2741.000 2667.000 2745.000 2667.600 ;
    END
  END wbs_data_i[7]
  PIN wbs_data_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2446.830 0.000 2447.110 4.000 ;
    END
  END wbs_data_i[8]
  PIN wbs_data_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2492.830 0.000 2493.110 4.000 ;
    END
  END wbs_data_i[9]
  PIN wbs_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 388.330 0.000 388.610 4.000 ;
    END
  END wbs_data_o[0]
  PIN wbs_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 846.030 0.000 846.310 4.000 ;
    END
  END wbs_data_o[10]
  PIN wbs_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 891.570 0.000 891.850 4.000 ;
    END
  END wbs_data_o[11]
  PIN wbs_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 937.570 0.000 937.850 4.000 ;
    END
  END wbs_data_o[12]
  PIN wbs_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 983.110 0.000 983.390 4.000 ;
    END
  END wbs_data_o[13]
  PIN wbs_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1028.650 0.000 1028.930 4.000 ;
    END
  END wbs_data_o[14]
  PIN wbs_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1074.650 0.000 1074.930 4.000 ;
    END
  END wbs_data_o[15]
  PIN wbs_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1120.190 0.000 1120.470 4.000 ;
    END
  END wbs_data_o[16]
  PIN wbs_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1166.190 0.000 1166.470 4.000 ;
    END
  END wbs_data_o[17]
  PIN wbs_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1211.730 0.000 1212.010 4.000 ;
    END
  END wbs_data_o[18]
  PIN wbs_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1257.730 0.000 1258.010 4.000 ;
    END
  END wbs_data_o[19]
  PIN wbs_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 434.330 0.000 434.610 4.000 ;
    END
  END wbs_data_o[1]
  PIN wbs_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1303.270 0.000 1303.550 4.000 ;
    END
  END wbs_data_o[20]
  PIN wbs_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1349.270 0.000 1349.550 4.000 ;
    END
  END wbs_data_o[21]
  PIN wbs_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1394.810 0.000 1395.090 4.000 ;
    END
  END wbs_data_o[22]
  PIN wbs_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1440.350 0.000 1440.630 4.000 ;
    END
  END wbs_data_o[23]
  PIN wbs_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1486.350 0.000 1486.630 4.000 ;
    END
  END wbs_data_o[24]
  PIN wbs_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1531.890 0.000 1532.170 4.000 ;
    END
  END wbs_data_o[25]
  PIN wbs_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1577.890 0.000 1578.170 4.000 ;
    END
  END wbs_data_o[26]
  PIN wbs_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1623.430 0.000 1623.710 4.000 ;
    END
  END wbs_data_o[27]
  PIN wbs_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1669.430 0.000 1669.710 4.000 ;
    END
  END wbs_data_o[28]
  PIN wbs_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1714.970 0.000 1715.250 4.000 ;
    END
  END wbs_data_o[29]
  PIN wbs_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 479.870 0.000 480.150 4.000 ;
    END
  END wbs_data_o[2]
  PIN wbs_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1760.970 0.000 1761.250 4.000 ;
    END
  END wbs_data_o[30]
  PIN wbs_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1806.510 0.000 1806.790 4.000 ;
    END
  END wbs_data_o[31]
  PIN wbs_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 525.410 0.000 525.690 4.000 ;
    END
  END wbs_data_o[3]
  PIN wbs_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 571.410 0.000 571.690 4.000 ;
    END
  END wbs_data_o[4]
  PIN wbs_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 616.950 0.000 617.230 4.000 ;
    END
  END wbs_data_o[5]
  PIN wbs_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 662.950 0.000 663.230 4.000 ;
    END
  END wbs_data_o[6]
  PIN wbs_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 708.490 0.000 708.770 4.000 ;
    END
  END wbs_data_o[7]
  PIN wbs_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 754.490 0.000 754.770 4.000 ;
    END
  END wbs_data_o[8]
  PIN wbs_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 800.030 0.000 800.310 4.000 ;
    END
  END wbs_data_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2675.910 0.000 2676.190 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2721.450 0.000 2721.730 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2700.290 3316.000 2700.570 3320.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2987.280 4.000 2987.880 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3119.880 4.000 3120.480 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3252.480 4.000 3253.080 ;
    END
  END wbs_we_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 2739.300 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 64.785 2739.300 66.385 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2739.300 3307.605 ;
      LAYER met1 ;
        RECT 5.520 10.640 2739.300 3315.640 ;
      LAYER met2 ;
        RECT 13.440 3315.720 43.970 3316.000 ;
        RECT 44.810 3315.720 132.290 3316.000 ;
        RECT 133.130 3315.720 220.610 3316.000 ;
        RECT 221.450 3315.720 309.390 3316.000 ;
        RECT 310.230 3315.720 397.710 3316.000 ;
        RECT 398.550 3315.720 486.490 3316.000 ;
        RECT 487.330 3315.720 574.810 3316.000 ;
        RECT 575.650 3315.720 663.590 3316.000 ;
        RECT 664.430 3315.720 751.910 3316.000 ;
        RECT 752.750 3315.720 840.690 3316.000 ;
        RECT 841.530 3315.720 929.010 3316.000 ;
        RECT 929.850 3315.720 1017.790 3316.000 ;
        RECT 1018.630 3315.720 1106.110 3316.000 ;
        RECT 1106.950 3315.720 1194.890 3316.000 ;
        RECT 1195.730 3315.720 1283.210 3316.000 ;
        RECT 1284.050 3315.720 1371.990 3316.000 ;
        RECT 1372.830 3315.720 1460.310 3316.000 ;
        RECT 1461.150 3315.720 1549.090 3316.000 ;
        RECT 1549.930 3315.720 1637.410 3316.000 ;
        RECT 1638.250 3315.720 1726.190 3316.000 ;
        RECT 1727.030 3315.720 1814.510 3316.000 ;
        RECT 1815.350 3315.720 1903.290 3316.000 ;
        RECT 1904.130 3315.720 1991.610 3316.000 ;
        RECT 1992.450 3315.720 2080.390 3316.000 ;
        RECT 2081.230 3315.720 2168.710 3316.000 ;
        RECT 2169.550 3315.720 2257.490 3316.000 ;
        RECT 2258.330 3315.720 2345.810 3316.000 ;
        RECT 2346.650 3315.720 2434.590 3316.000 ;
        RECT 2435.430 3315.720 2522.910 3316.000 ;
        RECT 2523.750 3315.720 2611.690 3316.000 ;
        RECT 2612.530 3315.720 2700.010 3316.000 ;
        RECT 2700.850 3315.720 2725.410 3316.000 ;
        RECT 13.440 4.280 2725.410 3315.720 ;
        RECT 13.440 4.000 22.350 4.280 ;
        RECT 23.190 4.000 67.890 4.280 ;
        RECT 68.730 4.000 113.430 4.280 ;
        RECT 114.270 4.000 159.430 4.280 ;
        RECT 160.270 4.000 204.970 4.280 ;
        RECT 205.810 4.000 250.970 4.280 ;
        RECT 251.810 4.000 296.510 4.280 ;
        RECT 297.350 4.000 342.510 4.280 ;
        RECT 343.350 4.000 388.050 4.280 ;
        RECT 388.890 4.000 434.050 4.280 ;
        RECT 434.890 4.000 479.590 4.280 ;
        RECT 480.430 4.000 525.130 4.280 ;
        RECT 525.970 4.000 571.130 4.280 ;
        RECT 571.970 4.000 616.670 4.280 ;
        RECT 617.510 4.000 662.670 4.280 ;
        RECT 663.510 4.000 708.210 4.280 ;
        RECT 709.050 4.000 754.210 4.280 ;
        RECT 755.050 4.000 799.750 4.280 ;
        RECT 800.590 4.000 845.750 4.280 ;
        RECT 846.590 4.000 891.290 4.280 ;
        RECT 892.130 4.000 937.290 4.280 ;
        RECT 938.130 4.000 982.830 4.280 ;
        RECT 983.670 4.000 1028.370 4.280 ;
        RECT 1029.210 4.000 1074.370 4.280 ;
        RECT 1075.210 4.000 1119.910 4.280 ;
        RECT 1120.750 4.000 1165.910 4.280 ;
        RECT 1166.750 4.000 1211.450 4.280 ;
        RECT 1212.290 4.000 1257.450 4.280 ;
        RECT 1258.290 4.000 1302.990 4.280 ;
        RECT 1303.830 4.000 1348.990 4.280 ;
        RECT 1349.830 4.000 1394.530 4.280 ;
        RECT 1395.370 4.000 1440.070 4.280 ;
        RECT 1440.910 4.000 1486.070 4.280 ;
        RECT 1486.910 4.000 1531.610 4.280 ;
        RECT 1532.450 4.000 1577.610 4.280 ;
        RECT 1578.450 4.000 1623.150 4.280 ;
        RECT 1623.990 4.000 1669.150 4.280 ;
        RECT 1669.990 4.000 1714.690 4.280 ;
        RECT 1715.530 4.000 1760.690 4.280 ;
        RECT 1761.530 4.000 1806.230 4.280 ;
        RECT 1807.070 4.000 1852.230 4.280 ;
        RECT 1853.070 4.000 1897.770 4.280 ;
        RECT 1898.610 4.000 1943.310 4.280 ;
        RECT 1944.150 4.000 1989.310 4.280 ;
        RECT 1990.150 4.000 2034.850 4.280 ;
        RECT 2035.690 4.000 2080.850 4.280 ;
        RECT 2081.690 4.000 2126.390 4.280 ;
        RECT 2127.230 4.000 2172.390 4.280 ;
        RECT 2173.230 4.000 2217.930 4.280 ;
        RECT 2218.770 4.000 2263.930 4.280 ;
        RECT 2264.770 4.000 2309.470 4.280 ;
        RECT 2310.310 4.000 2355.010 4.280 ;
        RECT 2355.850 4.000 2401.010 4.280 ;
        RECT 2401.850 4.000 2446.550 4.280 ;
        RECT 2447.390 4.000 2492.550 4.280 ;
        RECT 2493.390 4.000 2538.090 4.280 ;
        RECT 2538.930 4.000 2584.090 4.280 ;
        RECT 2584.930 4.000 2629.630 4.280 ;
        RECT 2630.470 4.000 2675.630 4.280 ;
        RECT 2676.470 4.000 2721.170 4.280 ;
        RECT 2722.010 4.000 2725.410 4.280 ;
      LAYER met3 ;
        RECT 4.000 3260.960 2741.000 3307.685 ;
        RECT 4.000 3259.560 2740.600 3260.960 ;
        RECT 4.000 3253.480 2741.000 3259.560 ;
        RECT 4.400 3252.080 2741.000 3253.480 ;
        RECT 4.000 3142.640 2741.000 3252.080 ;
        RECT 4.000 3141.240 2740.600 3142.640 ;
        RECT 4.000 3120.880 2741.000 3141.240 ;
        RECT 4.400 3119.480 2741.000 3120.880 ;
        RECT 4.000 3023.640 2741.000 3119.480 ;
        RECT 4.000 3022.240 2740.600 3023.640 ;
        RECT 4.000 2988.280 2741.000 3022.240 ;
        RECT 4.400 2986.880 2741.000 2988.280 ;
        RECT 4.000 2905.320 2741.000 2986.880 ;
        RECT 4.000 2903.920 2740.600 2905.320 ;
        RECT 4.000 2855.000 2741.000 2903.920 ;
        RECT 4.400 2853.600 2741.000 2855.000 ;
        RECT 4.000 2787.000 2741.000 2853.600 ;
        RECT 4.000 2785.600 2740.600 2787.000 ;
        RECT 4.000 2722.400 2741.000 2785.600 ;
        RECT 4.400 2721.000 2741.000 2722.400 ;
        RECT 4.000 2668.000 2741.000 2721.000 ;
        RECT 4.000 2666.600 2740.600 2668.000 ;
        RECT 4.000 2589.800 2741.000 2666.600 ;
        RECT 4.400 2588.400 2741.000 2589.800 ;
        RECT 4.000 2549.680 2741.000 2588.400 ;
        RECT 4.000 2548.280 2740.600 2549.680 ;
        RECT 4.000 2457.200 2741.000 2548.280 ;
        RECT 4.400 2455.800 2741.000 2457.200 ;
        RECT 4.000 2431.360 2741.000 2455.800 ;
        RECT 4.000 2429.960 2740.600 2431.360 ;
        RECT 4.000 2323.920 2741.000 2429.960 ;
        RECT 4.400 2322.520 2741.000 2323.920 ;
        RECT 4.000 2312.360 2741.000 2322.520 ;
        RECT 4.000 2310.960 2740.600 2312.360 ;
        RECT 4.000 2194.040 2741.000 2310.960 ;
        RECT 4.000 2192.640 2740.600 2194.040 ;
        RECT 4.000 2191.320 2741.000 2192.640 ;
        RECT 4.400 2189.920 2741.000 2191.320 ;
        RECT 4.000 2075.720 2741.000 2189.920 ;
        RECT 4.000 2074.320 2740.600 2075.720 ;
        RECT 4.000 2058.720 2741.000 2074.320 ;
        RECT 4.400 2057.320 2741.000 2058.720 ;
        RECT 4.000 1956.720 2741.000 2057.320 ;
        RECT 4.000 1955.320 2740.600 1956.720 ;
        RECT 4.000 1925.440 2741.000 1955.320 ;
        RECT 4.400 1924.040 2741.000 1925.440 ;
        RECT 4.000 1838.400 2741.000 1924.040 ;
        RECT 4.000 1837.000 2740.600 1838.400 ;
        RECT 4.000 1792.840 2741.000 1837.000 ;
        RECT 4.400 1791.440 2741.000 1792.840 ;
        RECT 4.000 1720.080 2741.000 1791.440 ;
        RECT 4.000 1718.680 2740.600 1720.080 ;
        RECT 4.000 1660.240 2741.000 1718.680 ;
        RECT 4.400 1658.840 2741.000 1660.240 ;
        RECT 4.000 1601.080 2741.000 1658.840 ;
        RECT 4.000 1599.680 2740.600 1601.080 ;
        RECT 4.000 1527.640 2741.000 1599.680 ;
        RECT 4.400 1526.240 2741.000 1527.640 ;
        RECT 4.000 1482.760 2741.000 1526.240 ;
        RECT 4.000 1481.360 2740.600 1482.760 ;
        RECT 4.000 1394.360 2741.000 1481.360 ;
        RECT 4.400 1392.960 2741.000 1394.360 ;
        RECT 4.000 1363.760 2741.000 1392.960 ;
        RECT 4.000 1362.360 2740.600 1363.760 ;
        RECT 4.000 1261.760 2741.000 1362.360 ;
        RECT 4.400 1260.360 2741.000 1261.760 ;
        RECT 4.000 1245.440 2741.000 1260.360 ;
        RECT 4.000 1244.040 2740.600 1245.440 ;
        RECT 4.000 1129.160 2741.000 1244.040 ;
        RECT 4.400 1127.760 2741.000 1129.160 ;
        RECT 4.000 1127.120 2741.000 1127.760 ;
        RECT 4.000 1125.720 2740.600 1127.120 ;
        RECT 4.000 1008.120 2741.000 1125.720 ;
        RECT 4.000 1006.720 2740.600 1008.120 ;
        RECT 4.000 995.880 2741.000 1006.720 ;
        RECT 4.400 994.480 2741.000 995.880 ;
        RECT 4.000 889.800 2741.000 994.480 ;
        RECT 4.000 888.400 2740.600 889.800 ;
        RECT 4.000 863.280 2741.000 888.400 ;
        RECT 4.400 861.880 2741.000 863.280 ;
        RECT 4.000 771.480 2741.000 861.880 ;
        RECT 4.000 770.080 2740.600 771.480 ;
        RECT 4.000 730.680 2741.000 770.080 ;
        RECT 4.400 729.280 2741.000 730.680 ;
        RECT 4.000 652.480 2741.000 729.280 ;
        RECT 4.000 651.080 2740.600 652.480 ;
        RECT 4.000 598.080 2741.000 651.080 ;
        RECT 4.400 596.680 2741.000 598.080 ;
        RECT 4.000 534.160 2741.000 596.680 ;
        RECT 4.000 532.760 2740.600 534.160 ;
        RECT 4.000 464.800 2741.000 532.760 ;
        RECT 4.400 463.400 2741.000 464.800 ;
        RECT 4.000 415.840 2741.000 463.400 ;
        RECT 4.000 414.440 2740.600 415.840 ;
        RECT 4.000 332.200 2741.000 414.440 ;
        RECT 4.400 330.800 2741.000 332.200 ;
        RECT 4.000 296.840 2741.000 330.800 ;
        RECT 4.000 295.440 2740.600 296.840 ;
        RECT 4.000 199.600 2741.000 295.440 ;
        RECT 4.400 198.200 2741.000 199.600 ;
        RECT 4.000 178.520 2741.000 198.200 ;
        RECT 4.000 177.120 2740.600 178.520 ;
        RECT 4.000 67.000 2741.000 177.120 ;
        RECT 4.400 65.600 2741.000 67.000 ;
        RECT 4.000 60.200 2741.000 65.600 ;
        RECT 4.000 58.800 2740.600 60.200 ;
        RECT 4.000 4.255 2741.000 58.800 ;
      LAYER met4 ;
        RECT 18.905 10.640 2706.705 3307.760 ;
      LAYER met5 ;
        RECT 5.520 92.700 2739.300 3283.165 ;
  END
END fpga
END LIBRARY


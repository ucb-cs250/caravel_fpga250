magic
tech sky130A
magscale 1 2
timestamp 1608149048
<< locali >>
rect 16589 3519 16623 3825
rect 26157 3519 26191 3825
rect 35909 2907 35943 3825
rect 45477 2975 45511 3825
rect 55229 3179 55263 3825
rect 64797 3247 64831 3825
rect 69673 3315 69707 4029
rect 69765 3247 69799 4029
rect 74549 3859 74583 4097
rect 84117 3859 84151 4097
rect 102517 3927 102551 4165
rect 102609 3383 102643 3893
rect 102701 3383 102735 3689
<< viali >>
rect 102517 4165 102551 4199
rect 74549 4097 74583 4131
rect 69673 4029 69707 4063
rect 16589 3825 16623 3859
rect 16589 3485 16623 3519
rect 26157 3825 26191 3859
rect 26157 3485 26191 3519
rect 35909 3825 35943 3859
rect 45477 3825 45511 3859
rect 55229 3825 55263 3859
rect 64797 3825 64831 3859
rect 69673 3281 69707 3315
rect 69765 4029 69799 4063
rect 64797 3213 64831 3247
rect 74549 3825 74583 3859
rect 84117 4097 84151 4131
rect 102517 3893 102551 3927
rect 102609 3893 102643 3927
rect 84117 3825 84151 3859
rect 102609 3349 102643 3383
rect 102701 3689 102735 3723
rect 102701 3349 102735 3383
rect 69765 3213 69799 3247
rect 55229 3145 55263 3179
rect 45477 2941 45511 2975
rect 35909 2873 35943 2907
<< metal1 >>
rect 144822 700680 144828 700732
rect 144880 700720 144886 700732
rect 170306 700720 170312 700732
rect 144880 700692 170312 700720
rect 144880 700680 144886 700692
rect 170306 700680 170312 700692
rect 170364 700680 170370 700732
rect 105446 700612 105452 700664
rect 105504 700652 105510 700664
rect 106182 700652 106188 700664
rect 105504 700624 106188 700652
rect 105504 700612 105510 700624
rect 106182 700612 106188 700624
rect 106240 700612 106246 700664
rect 124122 700612 124128 700664
rect 124180 700652 124186 700664
rect 235166 700652 235172 700664
rect 124180 700624 235172 700652
rect 124180 700612 124186 700624
rect 235166 700612 235172 700624
rect 235224 700612 235230 700664
rect 102042 700544 102048 700596
rect 102100 700584 102106 700596
rect 300118 700584 300124 700596
rect 102100 700556 300124 700584
rect 102100 700544 102106 700556
rect 300118 700544 300124 700556
rect 300176 700544 300182 700596
rect 81342 700476 81348 700528
rect 81400 700516 81406 700528
rect 364978 700516 364984 700528
rect 81400 700488 364984 700516
rect 81400 700476 81406 700488
rect 364978 700476 364984 700488
rect 365036 700476 365042 700528
rect 40494 700408 40500 700460
rect 40552 700448 40558 700460
rect 41322 700448 41328 700460
rect 40552 700420 41328 700448
rect 40552 700408 40558 700420
rect 41322 700408 41328 700420
rect 41380 700408 41386 700460
rect 60642 700408 60648 700460
rect 60700 700448 60706 700460
rect 429838 700448 429844 700460
rect 60700 700420 429844 700448
rect 60700 700408 60706 700420
rect 429838 700408 429844 700420
rect 429896 700408 429902 700460
rect 38562 700340 38568 700392
rect 38620 700380 38626 700392
rect 494790 700380 494796 700392
rect 38620 700352 494796 700380
rect 38620 700340 38626 700352
rect 494790 700340 494796 700352
rect 494848 700340 494854 700392
rect 17862 700272 17868 700324
rect 17920 700312 17926 700324
rect 559650 700312 559656 700324
rect 17920 700284 559656 700312
rect 17920 700272 17926 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 123018 689732 123024 689784
rect 123076 689772 123082 689784
rect 124122 689772 124128 689784
rect 123076 689744 124128 689772
rect 123076 689732 123082 689744
rect 124122 689732 124128 689744
rect 124180 689732 124186 689784
rect 144086 689732 144092 689784
rect 144144 689772 144150 689784
rect 144822 689772 144828 689784
rect 144144 689744 144828 689772
rect 144144 689732 144150 689744
rect 144822 689732 144828 689744
rect 144880 689732 144886 689784
rect 59630 689664 59636 689716
rect 59688 689704 59694 689716
rect 60642 689704 60648 689716
rect 59688 689676 60648 689704
rect 59688 689664 59694 689676
rect 60642 689664 60648 689676
rect 60700 689664 60706 689716
rect 106182 689664 106188 689716
rect 106240 689704 106246 689716
rect 165246 689704 165252 689716
rect 106240 689676 165252 689704
rect 106240 689664 106246 689676
rect 165246 689664 165252 689676
rect 165304 689664 165310 689716
rect 41322 689596 41328 689648
rect 41380 689636 41386 689648
rect 186314 689636 186320 689648
rect 41380 689608 186320 689636
rect 41380 689596 41386 689608
rect 186314 689596 186320 689608
rect 186372 689596 186378 689648
rect 2682 689528 2688 689580
rect 2740 689568 2746 689580
rect 228542 689568 228548 689580
rect 2740 689540 228548 689568
rect 2740 689528 2746 689540
rect 228542 689528 228548 689540
rect 228600 689528 228606 689580
rect 8110 689460 8116 689512
rect 8168 689500 8174 689512
rect 249702 689500 249708 689512
rect 8168 689472 249708 689500
rect 8168 689460 8174 689472
rect 249702 689460 249708 689472
rect 249760 689460 249766 689512
rect 9214 689392 9220 689444
rect 9272 689432 9278 689444
rect 270770 689432 270776 689444
rect 9272 689404 270776 689432
rect 9272 689392 9278 689404
rect 270770 689392 270776 689404
rect 270828 689392 270834 689444
rect 9674 689324 9680 689376
rect 9732 689364 9738 689376
rect 291930 689364 291936 689376
rect 9732 689336 291936 689364
rect 9732 689324 9738 689336
rect 291930 689324 291936 689336
rect 291988 689324 291994 689376
rect 9582 689256 9588 689308
rect 9640 689296 9646 689308
rect 312998 689296 313004 689308
rect 9640 689268 313004 689296
rect 9640 689256 9646 689268
rect 312998 689256 313004 689268
rect 313056 689256 313062 689308
rect 9030 689188 9036 689240
rect 9088 689228 9094 689240
rect 334158 689228 334164 689240
rect 9088 689200 334164 689228
rect 9088 689188 9094 689200
rect 334158 689188 334164 689200
rect 334216 689188 334222 689240
rect 8202 689120 8208 689172
rect 8260 689160 8266 689172
rect 355226 689160 355232 689172
rect 8260 689132 355232 689160
rect 8260 689120 8266 689132
rect 355226 689120 355232 689132
rect 355284 689120 355290 689172
rect 207474 689052 207480 689104
rect 207532 689092 207538 689104
rect 576118 689092 576124 689104
rect 207532 689064 576124 689092
rect 207532 689052 207538 689064
rect 576118 689052 576124 689064
rect 576176 689052 576182 689104
rect 4062 688984 4068 689036
rect 4120 689024 4126 689036
rect 376386 689024 376392 689036
rect 4120 688996 376392 689024
rect 4120 688984 4126 688996
rect 376386 688984 376392 688996
rect 376444 688984 376450 689036
rect 8938 688916 8944 688968
rect 8996 688956 9002 688968
rect 397454 688956 397460 688968
rect 8996 688928 397460 688956
rect 8996 688916 9002 688928
rect 397454 688916 397460 688928
rect 397512 688916 397518 688968
rect 9306 688848 9312 688900
rect 9364 688888 9370 688900
rect 418614 688888 418620 688900
rect 9364 688860 418620 688888
rect 9364 688848 9370 688860
rect 418614 688848 418620 688860
rect 418672 688848 418678 688900
rect 9122 688780 9128 688832
rect 9180 688820 9186 688832
rect 439682 688820 439688 688832
rect 9180 688792 439688 688820
rect 9180 688780 9186 688792
rect 439682 688780 439688 688792
rect 439740 688780 439746 688832
rect 9398 688712 9404 688764
rect 9456 688752 9462 688764
rect 460842 688752 460848 688764
rect 9456 688724 460848 688752
rect 9456 688712 9462 688724
rect 460842 688712 460848 688724
rect 460900 688712 460906 688764
rect 9490 688644 9496 688696
rect 9548 688684 9554 688696
rect 481910 688684 481916 688696
rect 9548 688656 481916 688684
rect 9548 688644 9554 688656
rect 481910 688644 481916 688656
rect 481968 688644 481974 688696
rect 3142 681708 3148 681760
rect 3200 681748 3206 681760
rect 6178 681748 6184 681760
rect 3200 681720 6184 681748
rect 3200 681708 3206 681720
rect 6178 681708 6184 681720
rect 6236 681708 6242 681760
rect 3970 567196 3976 567248
rect 4028 567236 4034 567248
rect 6270 567236 6276 567248
rect 4028 567208 6276 567236
rect 4028 567196 4034 567208
rect 6270 567196 6276 567208
rect 6328 567196 6334 567248
rect 3510 509260 3516 509312
rect 3568 509300 3574 509312
rect 7558 509300 7564 509312
rect 3568 509272 7564 509300
rect 3568 509260 3574 509272
rect 7558 509260 7564 509272
rect 7616 509260 7622 509312
rect 576118 487092 576124 487144
rect 576176 487132 576182 487144
rect 579706 487132 579712 487144
rect 576176 487104 579712 487132
rect 576176 487092 576182 487104
rect 579706 487092 579712 487104
rect 579764 487092 579770 487144
rect 578142 238212 578148 238264
rect 578200 238252 578206 238264
rect 580626 238252 580632 238264
rect 578200 238224 580632 238252
rect 578200 238212 578206 238224
rect 580626 238212 580632 238224
rect 580684 238212 580690 238264
rect 578142 213868 578148 213920
rect 578200 213908 578206 213920
rect 580718 213908 580724 213920
rect 578200 213880 580724 213908
rect 578200 213868 578206 213880
rect 580718 213868 580724 213880
rect 580776 213868 580782 213920
rect 578142 189796 578148 189848
rect 578200 189836 578206 189848
rect 580810 189836 580816 189848
rect 578200 189808 580816 189836
rect 578200 189796 578206 189808
rect 580810 189796 580816 189808
rect 580868 189796 580874 189848
rect 3326 181092 3332 181144
rect 3384 181132 3390 181144
rect 4154 181132 4160 181144
rect 3384 181104 4160 181132
rect 3384 181092 3390 181104
rect 4154 181092 4160 181104
rect 4212 181092 4218 181144
rect 578142 165452 578148 165504
rect 578200 165492 578206 165504
rect 580902 165492 580908 165504
rect 578200 165464 580908 165492
rect 578200 165452 578206 165464
rect 580902 165452 580908 165464
rect 580960 165452 580966 165504
rect 3234 121388 3240 121440
rect 3292 121428 3298 121440
rect 4154 121428 4160 121440
rect 3292 121400 4160 121428
rect 3292 121388 3298 121400
rect 4154 121388 4160 121400
rect 4212 121388 4218 121440
rect 578142 116900 578148 116952
rect 578200 116940 578206 116952
rect 580626 116940 580632 116952
rect 578200 116912 580632 116940
rect 578200 116900 578206 116912
rect 580626 116900 580632 116912
rect 580684 116900 580690 116952
rect 578142 92420 578148 92472
rect 578200 92460 578206 92472
rect 580718 92460 580724 92472
rect 578200 92432 580724 92460
rect 578200 92420 578206 92432
rect 580718 92420 580724 92432
rect 580776 92420 580782 92472
rect 578142 68348 578148 68400
rect 578200 68388 578206 68400
rect 580626 68388 580632 68400
rect 578200 68360 580632 68388
rect 578200 68348 578206 68360
rect 580626 68348 580632 68360
rect 580684 68348 580690 68400
rect 578142 44004 578148 44056
rect 578200 44044 578206 44056
rect 580626 44044 580632 44056
rect 578200 44016 580632 44044
rect 578200 44004 578206 44016
rect 580626 44004 580632 44016
rect 580684 44004 580690 44056
rect 52730 6808 52736 6860
rect 52788 6848 52794 6860
rect 580534 6848 580540 6860
rect 52788 6820 580540 6848
rect 52788 6808 52794 6820
rect 580534 6808 580540 6820
rect 580592 6808 580598 6860
rect 62942 6740 62948 6792
rect 63000 6780 63006 6792
rect 580442 6780 580448 6792
rect 63000 6752 580448 6780
rect 63000 6740 63006 6752
rect 580442 6740 580448 6752
rect 580500 6740 580506 6792
rect 73062 6672 73068 6724
rect 73120 6712 73126 6724
rect 580350 6712 580356 6724
rect 73120 6684 580356 6712
rect 73120 6672 73126 6684
rect 580350 6672 580356 6684
rect 580408 6672 580414 6724
rect 83274 6604 83280 6656
rect 83332 6644 83338 6656
rect 580258 6644 580264 6656
rect 83332 6616 580264 6644
rect 83332 6604 83338 6616
rect 580258 6604 580264 6616
rect 580316 6604 580322 6656
rect 4522 6536 4528 6588
rect 4580 6576 4586 6588
rect 90910 6576 90916 6588
rect 4580 6548 90916 6576
rect 4580 6536 4586 6548
rect 90910 6536 90916 6548
rect 90968 6536 90974 6588
rect 92106 6536 92112 6588
rect 92164 6576 92170 6588
rect 578326 6576 578332 6588
rect 92164 6548 578332 6576
rect 92164 6536 92170 6548
rect 578326 6536 578332 6548
rect 578384 6536 578390 6588
rect 84930 6468 84936 6520
rect 84988 6508 84994 6520
rect 578418 6508 578424 6520
rect 84988 6480 578424 6508
rect 84988 6468 84994 6480
rect 578418 6468 578424 6480
rect 578476 6468 578482 6520
rect 81434 6400 81440 6452
rect 81492 6440 81498 6452
rect 578510 6440 578516 6452
rect 81492 6412 578516 6440
rect 81492 6400 81498 6412
rect 578510 6400 578516 6412
rect 578568 6400 578574 6452
rect 56410 6332 56416 6384
rect 56468 6372 56474 6384
rect 578602 6372 578608 6384
rect 56468 6344 578608 6372
rect 56468 6332 56474 6344
rect 578602 6332 578608 6344
rect 578660 6332 578666 6384
rect 52822 6264 52828 6316
rect 52880 6304 52886 6316
rect 578694 6304 578700 6316
rect 52880 6276 578700 6304
rect 52880 6264 52886 6276
rect 578694 6264 578700 6276
rect 578752 6264 578758 6316
rect 33870 6196 33876 6248
rect 33928 6236 33934 6248
rect 579430 6236 579436 6248
rect 33928 6208 579436 6236
rect 33928 6196 33934 6208
rect 579430 6196 579436 6208
rect 579488 6196 579494 6248
rect 30282 6128 30288 6180
rect 30340 6168 30346 6180
rect 579522 6168 579528 6180
rect 30340 6140 579528 6168
rect 30340 6128 30346 6140
rect 579522 6128 579528 6140
rect 579580 6128 579586 6180
rect 4430 6060 4436 6112
rect 4488 6100 4494 6112
rect 87322 6100 87328 6112
rect 4488 6072 87328 6100
rect 4488 6060 4494 6072
rect 87322 6060 87328 6072
rect 87380 6060 87386 6112
rect 94498 6060 94504 6112
rect 94556 6100 94562 6112
rect 579338 6100 579344 6112
rect 94556 6072 579344 6100
rect 94556 6060 94562 6072
rect 579338 6060 579344 6072
rect 579396 6060 579402 6112
rect 4706 5992 4712 6044
rect 4764 6032 4770 6044
rect 105170 6032 105176 6044
rect 4764 6004 105176 6032
rect 4764 5992 4770 6004
rect 105170 5992 105176 6004
rect 105228 5992 105234 6044
rect 108758 5992 108764 6044
rect 108816 6032 108822 6044
rect 579246 6032 579252 6044
rect 108816 6004 579252 6032
rect 108816 5992 108822 6004
rect 579246 5992 579252 6004
rect 579304 5992 579310 6044
rect 4614 5924 4620 5976
rect 4672 5964 4678 5976
rect 101582 5964 101588 5976
rect 4672 5936 101588 5964
rect 4672 5924 4678 5936
rect 101582 5924 101588 5936
rect 101640 5924 101646 5976
rect 112346 5924 112352 5976
rect 112404 5964 112410 5976
rect 579154 5964 579160 5976
rect 112404 5936 579160 5964
rect 112404 5924 112410 5936
rect 579154 5924 579160 5936
rect 579212 5924 579218 5976
rect 4798 5856 4804 5908
rect 4856 5896 4862 5908
rect 115934 5896 115940 5908
rect 4856 5868 115940 5896
rect 4856 5856 4862 5868
rect 115934 5856 115940 5868
rect 115992 5856 115998 5908
rect 119430 5856 119436 5908
rect 119488 5896 119494 5908
rect 579062 5896 579068 5908
rect 119488 5868 579068 5896
rect 119488 5856 119494 5868
rect 579062 5856 579068 5868
rect 579120 5856 579126 5908
rect 4890 5788 4896 5840
rect 4948 5828 4954 5840
rect 123018 5828 123024 5840
rect 4948 5800 123024 5828
rect 4948 5788 4954 5800
rect 123018 5788 123024 5800
rect 123076 5788 123082 5840
rect 5166 5720 5172 5772
rect 5224 5760 5230 5772
rect 117130 5760 117136 5772
rect 5224 5732 117136 5760
rect 5224 5720 5230 5732
rect 117130 5720 117136 5732
rect 117188 5720 117194 5772
rect 7558 5448 7564 5500
rect 7616 5488 7622 5500
rect 42518 5488 42524 5500
rect 7616 5460 42524 5488
rect 7616 5448 7622 5460
rect 42518 5448 42524 5460
rect 42576 5448 42582 5500
rect 89714 5448 89720 5500
rect 89772 5488 89778 5500
rect 307202 5488 307208 5500
rect 89772 5460 307208 5488
rect 89772 5448 89778 5460
rect 307202 5448 307208 5460
rect 307260 5448 307266 5500
rect 6270 5380 6276 5432
rect 6328 5420 6334 5432
rect 32398 5420 32404 5432
rect 6328 5392 32404 5420
rect 6328 5380 6334 5392
rect 32398 5380 32404 5392
rect 32456 5380 32462 5432
rect 96890 5380 96896 5432
rect 96948 5420 96954 5432
rect 327534 5420 327540 5432
rect 96948 5392 327540 5420
rect 96948 5380 96954 5392
rect 327534 5380 327540 5392
rect 327592 5380 327598 5432
rect 3418 5312 3424 5364
rect 3476 5352 3482 5364
rect 22186 5352 22192 5364
rect 3476 5324 22192 5352
rect 3476 5312 3482 5324
rect 22186 5312 22192 5324
rect 22244 5312 22250 5364
rect 103974 5312 103980 5364
rect 104032 5352 104038 5364
rect 347958 5352 347964 5364
rect 104032 5324 347964 5352
rect 104032 5312 104038 5324
rect 347958 5312 347964 5324
rect 348016 5312 348022 5364
rect 6178 5244 6184 5296
rect 6236 5284 6242 5296
rect 12066 5284 12072 5296
rect 6236 5256 12072 5284
rect 6236 5244 6242 5256
rect 12066 5244 12072 5256
rect 12124 5244 12130 5296
rect 24302 5244 24308 5296
rect 24360 5284 24366 5296
rect 124030 5284 124036 5296
rect 24360 5256 124036 5284
rect 24360 5244 24366 5256
rect 124030 5244 124036 5256
rect 124088 5244 124094 5296
rect 124122 5244 124128 5296
rect 124180 5284 124186 5296
rect 398834 5284 398840 5296
rect 124180 5256 398840 5284
rect 124180 5244 124186 5256
rect 398834 5244 398840 5256
rect 398892 5244 398898 5296
rect 65978 5176 65984 5228
rect 66036 5216 66042 5228
rect 459922 5216 459928 5228
rect 66036 5188 459928 5216
rect 66036 5176 66042 5188
rect 459922 5176 459928 5188
rect 459980 5176 459986 5228
rect 69474 5108 69480 5160
rect 69532 5148 69538 5160
rect 470042 5148 470048 5160
rect 69532 5120 470048 5148
rect 69532 5108 69538 5120
rect 470042 5108 470048 5120
rect 470100 5108 470106 5160
rect 98086 5040 98092 5092
rect 98144 5080 98150 5092
rect 500586 5080 500592 5092
rect 98144 5052 500592 5080
rect 98144 5040 98150 5052
rect 500586 5040 500592 5052
rect 500644 5040 500650 5092
rect 48130 4972 48136 5024
rect 48188 5012 48194 5024
rect 449710 5012 449716 5024
rect 48188 4984 449716 5012
rect 48188 4972 48194 4984
rect 449710 4972 449716 4984
rect 449768 4972 449774 5024
rect 4246 4904 4252 4956
rect 4304 4944 4310 4956
rect 51626 4944 51632 4956
rect 4304 4916 51632 4944
rect 4304 4904 4310 4916
rect 51626 4904 51632 4916
rect 51684 4904 51690 4956
rect 83826 4904 83832 4956
rect 83884 4944 83890 4956
rect 490466 4944 490472 4956
rect 83884 4916 490472 4944
rect 83884 4904 83890 4916
rect 490466 4904 490472 4916
rect 490524 4904 490530 4956
rect 4338 4836 4344 4888
rect 4396 4876 4402 4888
rect 55214 4876 55220 4888
rect 4396 4848 55220 4876
rect 4396 4836 4402 4848
rect 55214 4836 55220 4848
rect 55272 4836 55278 4888
rect 73062 4836 73068 4888
rect 73120 4876 73126 4888
rect 480254 4876 480260 4888
rect 73120 4848 480260 4876
rect 73120 4836 73126 4848
rect 480254 4836 480260 4848
rect 480312 4836 480318 4888
rect 566 4768 572 4820
rect 624 4808 630 4820
rect 419166 4808 419172 4820
rect 624 4780 419172 4808
rect 624 4768 630 4780
rect 419166 4768 419172 4780
rect 419224 4768 419230 4820
rect 82630 4700 82636 4752
rect 82688 4740 82694 4752
rect 286870 4740 286876 4752
rect 82688 4712 286876 4740
rect 82688 4700 82694 4712
rect 286870 4700 286876 4712
rect 286928 4700 286934 4752
rect 75454 4632 75460 4684
rect 75512 4672 75518 4684
rect 266538 4672 266544 4684
rect 75512 4644 266544 4672
rect 75512 4632 75518 4644
rect 266538 4632 266544 4644
rect 266596 4632 266602 4684
rect 68278 4564 68284 4616
rect 68336 4604 68342 4616
rect 246114 4604 246120 4616
rect 68336 4576 246120 4604
rect 68336 4564 68342 4576
rect 246114 4564 246120 4576
rect 246172 4564 246178 4616
rect 46934 4496 46940 4548
rect 46992 4536 46998 4548
rect 185026 4536 185032 4548
rect 46992 4508 185032 4536
rect 46992 4496 46998 4508
rect 185026 4496 185032 4508
rect 185084 4496 185090 4548
rect 39758 4428 39764 4480
rect 39816 4468 39822 4480
rect 164694 4468 164700 4480
rect 39816 4440 164700 4468
rect 39816 4428 39822 4440
rect 164694 4428 164700 4440
rect 164752 4428 164758 4480
rect 19518 4360 19524 4412
rect 19576 4400 19582 4412
rect 113082 4400 113088 4412
rect 19576 4372 113088 4400
rect 19576 4360 19582 4372
rect 113082 4360 113088 4372
rect 113140 4360 113146 4412
rect 113910 4360 113916 4412
rect 113968 4400 113974 4412
rect 225782 4400 225788 4412
rect 113968 4372 225788 4400
rect 113968 4360 113974 4372
rect 225782 4360 225788 4372
rect 225840 4360 225846 4412
rect 32674 4292 32680 4344
rect 32732 4332 32738 4344
rect 144362 4332 144368 4344
rect 32732 4304 144368 4332
rect 32732 4292 32738 4304
rect 144362 4292 144368 4304
rect 144420 4292 144426 4344
rect 29086 4224 29092 4276
rect 29144 4264 29150 4276
rect 134150 4264 134156 4276
rect 29144 4236 134156 4264
rect 29144 4224 29150 4236
rect 134150 4224 134156 4236
rect 134208 4224 134214 4276
rect 102505 4199 102563 4205
rect 102505 4165 102517 4199
rect 102551 4196 102563 4199
rect 103606 4196 103612 4208
rect 102551 4168 103612 4196
rect 102551 4165 102563 4168
rect 102505 4159 102563 4165
rect 103606 4156 103612 4168
rect 103664 4156 103670 4208
rect 110414 4156 110420 4208
rect 110472 4196 110478 4208
rect 205450 4196 205456 4208
rect 110472 4168 205456 4196
rect 110472 4156 110478 4168
rect 205450 4156 205456 4168
rect 205508 4156 205514 4208
rect 6914 4088 6920 4140
rect 6972 4128 6978 4140
rect 70670 4128 70676 4140
rect 6972 4100 70676 4128
rect 6972 4088 6978 4100
rect 70670 4088 70676 4100
rect 70728 4088 70734 4140
rect 74537 4131 74595 4137
rect 74537 4097 74549 4131
rect 74583 4128 74595 4131
rect 84105 4131 84163 4137
rect 84105 4128 84117 4131
rect 74583 4100 84117 4128
rect 74583 4097 74595 4100
rect 74537 4091 74595 4097
rect 84105 4097 84117 4100
rect 84151 4097 84163 4131
rect 84105 4091 84163 4097
rect 100478 4088 100484 4140
rect 100536 4128 100542 4140
rect 337746 4128 337752 4140
rect 100536 4100 337752 4128
rect 100536 4088 100542 4100
rect 337746 4088 337752 4100
rect 337804 4088 337810 4140
rect 4982 4020 4988 4072
rect 5040 4060 5046 4072
rect 8846 4060 8852 4072
rect 5040 4032 8852 4060
rect 5040 4020 5046 4032
rect 8846 4020 8852 4032
rect 8904 4020 8910 4072
rect 9030 4020 9036 4072
rect 9088 4060 9094 4072
rect 69661 4063 69719 4069
rect 69661 4060 69673 4063
rect 9088 4032 69673 4060
rect 9088 4020 9094 4032
rect 69661 4029 69673 4032
rect 69707 4029 69719 4063
rect 69661 4023 69719 4029
rect 69753 4063 69811 4069
rect 69753 4029 69765 4063
rect 69799 4060 69811 4063
rect 113910 4060 113916 4072
rect 69799 4032 113916 4060
rect 69799 4029 69811 4032
rect 69753 4023 69811 4029
rect 113910 4020 113916 4032
rect 113968 4020 113974 4072
rect 358078 4060 358084 4072
rect 117884 4032 358084 4060
rect 8202 3952 8208 4004
rect 8260 3992 8266 4004
rect 80238 3992 80244 4004
rect 8260 3964 80244 3992
rect 8260 3952 8266 3964
rect 80238 3952 80244 3964
rect 80296 3952 80302 4004
rect 107562 3952 107568 4004
rect 107620 3992 107626 4004
rect 117884 3992 117912 4032
rect 358078 4020 358084 4032
rect 358136 4020 358142 4072
rect 368290 3992 368296 4004
rect 107620 3964 117912 3992
rect 117976 3964 368296 3992
rect 107620 3952 107626 3964
rect 6822 3884 6828 3936
rect 6880 3924 6886 3936
rect 88518 3924 88524 3936
rect 6880 3896 88524 3924
rect 6880 3884 6886 3896
rect 88518 3884 88524 3896
rect 88576 3884 88582 3936
rect 102505 3927 102563 3933
rect 102505 3924 102517 3927
rect 98656 3896 102517 3924
rect 14826 3816 14832 3868
rect 14884 3856 14890 3868
rect 16577 3859 16635 3865
rect 16577 3856 16589 3859
rect 14884 3828 16589 3856
rect 14884 3816 14890 3828
rect 16577 3825 16589 3828
rect 16623 3825 16635 3859
rect 16577 3819 16635 3825
rect 26145 3859 26203 3865
rect 26145 3825 26157 3859
rect 26191 3856 26203 3859
rect 35897 3859 35955 3865
rect 35897 3856 35909 3859
rect 26191 3828 35909 3856
rect 26191 3825 26203 3828
rect 26145 3819 26203 3825
rect 35897 3825 35909 3828
rect 35943 3825 35955 3859
rect 35897 3819 35955 3825
rect 45465 3859 45523 3865
rect 45465 3825 45477 3859
rect 45511 3856 45523 3859
rect 55217 3859 55275 3865
rect 55217 3856 55229 3859
rect 45511 3828 55229 3856
rect 45511 3825 45523 3828
rect 45465 3819 45523 3825
rect 55217 3825 55229 3828
rect 55263 3825 55275 3859
rect 55217 3819 55275 3825
rect 64785 3859 64843 3865
rect 64785 3825 64797 3859
rect 64831 3856 64843 3859
rect 74537 3859 74595 3865
rect 74537 3856 74549 3859
rect 64831 3828 74549 3856
rect 64831 3825 64843 3828
rect 64785 3819 64843 3825
rect 74537 3825 74549 3828
rect 74583 3825 74595 3859
rect 74537 3819 74595 3825
rect 84105 3859 84163 3865
rect 84105 3825 84117 3859
rect 84151 3856 84163 3859
rect 98656 3856 98684 3896
rect 102505 3893 102517 3896
rect 102551 3893 102563 3927
rect 102505 3887 102563 3893
rect 102597 3927 102655 3933
rect 102597 3893 102609 3927
rect 102643 3924 102655 3927
rect 110414 3924 110420 3936
rect 102643 3896 110420 3924
rect 102643 3893 102655 3896
rect 102597 3887 102655 3893
rect 110414 3884 110420 3896
rect 110472 3884 110478 3936
rect 111150 3884 111156 3936
rect 111208 3924 111214 3936
rect 117976 3924 118004 3964
rect 368290 3952 368296 3964
rect 368348 3952 368354 4004
rect 378502 3924 378508 3936
rect 111208 3896 118004 3924
rect 118068 3896 378508 3924
rect 111208 3884 111214 3896
rect 84151 3828 98684 3856
rect 84151 3825 84163 3828
rect 84105 3819 84163 3825
rect 113542 3816 113548 3868
rect 113600 3856 113606 3868
rect 114554 3856 114560 3868
rect 113600 3828 114560 3856
rect 113600 3816 113606 3828
rect 114554 3816 114560 3828
rect 114612 3816 114618 3868
rect 114738 3816 114744 3868
rect 114796 3856 114802 3868
rect 118068 3856 118096 3896
rect 378502 3884 378508 3896
rect 378560 3884 378566 3936
rect 114796 3828 118096 3856
rect 114796 3816 114802 3828
rect 118234 3816 118240 3868
rect 118292 3856 118298 3868
rect 388622 3856 388628 3868
rect 118292 3828 388628 3856
rect 118292 3816 118298 3828
rect 388622 3816 388628 3828
rect 388680 3816 388686 3868
rect 5258 3748 5264 3800
rect 5316 3788 5322 3800
rect 120626 3788 120632 3800
rect 5316 3760 120632 3788
rect 5316 3748 5322 3760
rect 120626 3748 120632 3760
rect 120684 3748 120690 3800
rect 121822 3748 121828 3800
rect 121880 3788 121886 3800
rect 124122 3788 124128 3800
rect 121880 3760 124128 3788
rect 121880 3748 121886 3760
rect 124122 3748 124128 3760
rect 124180 3748 124186 3800
rect 125410 3748 125416 3800
rect 125468 3788 125474 3800
rect 409046 3788 409052 3800
rect 125468 3760 409052 3788
rect 125468 3748 125474 3760
rect 409046 3748 409052 3760
rect 409104 3748 409110 3800
rect 10042 3680 10048 3732
rect 10100 3720 10106 3732
rect 93118 3720 93124 3732
rect 10100 3692 93124 3720
rect 10100 3680 10106 3692
rect 93118 3680 93124 3692
rect 93176 3680 93182 3732
rect 93302 3680 93308 3732
rect 93360 3720 93366 3732
rect 102689 3723 102747 3729
rect 102689 3720 102701 3723
rect 93360 3692 102701 3720
rect 93360 3680 93366 3692
rect 102689 3689 102701 3692
rect 102735 3689 102747 3723
rect 102689 3683 102747 3689
rect 102778 3680 102784 3732
rect 102836 3720 102842 3732
rect 551554 3720 551560 3732
rect 102836 3692 551560 3720
rect 102836 3680 102842 3692
rect 551554 3680 551560 3692
rect 551612 3680 551618 3732
rect 9582 3612 9588 3664
rect 9640 3652 9646 3664
rect 62390 3652 62396 3664
rect 9640 3624 62396 3652
rect 9640 3612 9646 3624
rect 62390 3612 62396 3624
rect 62448 3612 62454 3664
rect 63586 3612 63592 3664
rect 63644 3652 63650 3664
rect 541342 3652 541348 3664
rect 63644 3624 541348 3652
rect 63644 3612 63650 3624
rect 541342 3612 541348 3624
rect 541400 3612 541406 3664
rect 5350 3544 5356 3596
rect 5408 3584 5414 3596
rect 11238 3584 11244 3596
rect 5408 3556 11244 3584
rect 5408 3544 5414 3556
rect 11238 3544 11244 3556
rect 11296 3544 11302 3596
rect 13630 3544 13636 3596
rect 13688 3584 13694 3596
rect 510798 3584 510804 3596
rect 13688 3556 510804 3584
rect 13688 3544 13694 3556
rect 510798 3544 510804 3556
rect 510856 3544 510862 3596
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 2682 3516 2688 3528
rect 1728 3488 2688 3516
rect 1728 3476 1734 3488
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 5442 3476 5448 3528
rect 5500 3516 5506 3528
rect 16022 3516 16028 3528
rect 5500 3488 16028 3516
rect 5500 3476 5506 3488
rect 16022 3476 16028 3488
rect 16080 3476 16086 3528
rect 16577 3519 16635 3525
rect 16577 3485 16589 3519
rect 16623 3516 16635 3519
rect 26145 3519 26203 3525
rect 26145 3516 26157 3519
rect 16623 3488 26157 3516
rect 16623 3485 16635 3488
rect 16577 3479 16635 3485
rect 26145 3485 26157 3488
rect 26191 3485 26203 3519
rect 26145 3479 26203 3485
rect 31478 3476 31484 3528
rect 31536 3516 31542 3528
rect 578878 3516 578884 3528
rect 31536 3488 578884 3516
rect 31536 3476 31542 3488
rect 578878 3476 578884 3488
rect 578936 3476 578942 3528
rect 6546 3408 6552 3460
rect 6604 3448 6610 3460
rect 26694 3448 26700 3460
rect 6604 3420 26700 3448
rect 6604 3408 6610 3420
rect 26694 3408 26700 3420
rect 26752 3408 26758 3460
rect 27890 3408 27896 3460
rect 27948 3448 27954 3460
rect 578970 3448 578976 3460
rect 27948 3420 578976 3448
rect 27948 3408 27954 3420
rect 578970 3408 578976 3420
rect 579028 3408 579034 3460
rect 6730 3340 6736 3392
rect 6788 3380 6794 3392
rect 49326 3380 49332 3392
rect 6788 3352 49332 3380
rect 6788 3340 6794 3352
rect 49326 3340 49332 3352
rect 49384 3340 49390 3392
rect 54018 3340 54024 3392
rect 54076 3380 54082 3392
rect 102597 3383 102655 3389
rect 102597 3380 102609 3383
rect 54076 3352 102609 3380
rect 54076 3340 54082 3352
rect 102597 3349 102609 3352
rect 102643 3349 102655 3383
rect 102597 3343 102655 3349
rect 102689 3383 102747 3389
rect 102689 3349 102701 3383
rect 102735 3380 102747 3383
rect 317414 3380 317420 3392
rect 102735 3352 317420 3380
rect 102735 3349 102747 3352
rect 102689 3343 102747 3349
rect 317414 3340 317420 3352
rect 317472 3340 317478 3392
rect 9122 3272 9128 3324
rect 9180 3312 9186 3324
rect 59998 3312 60004 3324
rect 9180 3284 60004 3312
rect 9180 3272 9186 3284
rect 59998 3272 60004 3284
rect 60056 3272 60062 3324
rect 61194 3272 61200 3324
rect 61252 3312 61258 3324
rect 69661 3315 69719 3321
rect 61252 3284 69612 3312
rect 61252 3272 61258 3284
rect 9674 3204 9680 3256
rect 9732 3244 9738 3256
rect 58802 3244 58808 3256
rect 9732 3216 58808 3244
rect 9732 3204 9738 3216
rect 58802 3204 58808 3216
rect 58860 3204 58866 3256
rect 64785 3247 64843 3253
rect 64785 3213 64797 3247
rect 64831 3213 64843 3247
rect 69584 3244 69612 3284
rect 69661 3281 69673 3315
rect 69707 3312 69719 3315
rect 76650 3312 76656 3324
rect 69707 3284 76656 3312
rect 69707 3281 69719 3284
rect 69661 3275 69719 3281
rect 76650 3272 76656 3284
rect 76708 3272 76714 3324
rect 86126 3272 86132 3324
rect 86184 3312 86190 3324
rect 297082 3312 297088 3324
rect 86184 3284 297088 3312
rect 86184 3272 86190 3284
rect 297082 3272 297088 3284
rect 297140 3272 297146 3324
rect 69753 3247 69811 3253
rect 69753 3244 69765 3247
rect 69584 3216 69765 3244
rect 64785 3207 64843 3213
rect 69753 3213 69765 3216
rect 69799 3213 69811 3247
rect 69753 3207 69811 3213
rect 5074 3136 5080 3188
rect 5132 3176 5138 3188
rect 45738 3176 45744 3188
rect 5132 3148 45744 3176
rect 5132 3136 5138 3148
rect 45738 3136 45744 3148
rect 45796 3136 45802 3188
rect 55217 3179 55275 3185
rect 55217 3145 55229 3179
rect 55263 3176 55275 3179
rect 64800 3176 64828 3207
rect 79042 3204 79048 3256
rect 79100 3244 79106 3256
rect 276658 3244 276664 3256
rect 79100 3216 276664 3244
rect 79100 3204 79106 3216
rect 276658 3204 276664 3216
rect 276716 3204 276722 3256
rect 55263 3148 64828 3176
rect 55263 3145 55275 3148
rect 55217 3139 55275 3145
rect 71866 3136 71872 3188
rect 71924 3176 71930 3188
rect 256326 3176 256332 3188
rect 71924 3148 256332 3176
rect 71924 3136 71930 3148
rect 256326 3136 256332 3148
rect 256384 3136 256390 3188
rect 7006 3068 7012 3120
rect 7064 3108 7070 3120
rect 44542 3108 44548 3120
rect 7064 3080 44548 3108
rect 7064 3068 7070 3080
rect 44542 3068 44548 3080
rect 44600 3068 44606 3120
rect 64782 3068 64788 3120
rect 64840 3108 64846 3120
rect 235994 3108 236000 3120
rect 64840 3080 236000 3108
rect 64840 3068 64846 3080
rect 235994 3068 236000 3080
rect 236052 3068 236058 3120
rect 6638 3000 6644 3052
rect 6696 3040 6702 3052
rect 40954 3040 40960 3052
rect 6696 3012 40960 3040
rect 6696 3000 6702 3012
rect 40954 3000 40960 3012
rect 41012 3000 41018 3052
rect 57606 3000 57612 3052
rect 57664 3040 57670 3052
rect 215570 3040 215576 3052
rect 57664 3012 215576 3040
rect 57664 3000 57670 3012
rect 215570 3000 215576 3012
rect 215628 3000 215634 3052
rect 7098 2932 7104 2984
rect 7156 2972 7162 2984
rect 37366 2972 37372 2984
rect 7156 2944 37372 2972
rect 7156 2932 7162 2944
rect 37366 2932 37372 2944
rect 37424 2932 37430 2984
rect 45465 2975 45523 2981
rect 45465 2972 45477 2975
rect 37476 2944 45477 2972
rect 9214 2864 9220 2916
rect 9272 2904 9278 2916
rect 21910 2904 21916 2916
rect 9272 2876 21916 2904
rect 9272 2864 9278 2876
rect 21910 2864 21916 2876
rect 21968 2864 21974 2916
rect 35897 2907 35955 2913
rect 35897 2873 35909 2907
rect 35943 2904 35955 2907
rect 37476 2904 37504 2944
rect 45465 2941 45477 2944
rect 45511 2941 45523 2975
rect 45465 2935 45523 2941
rect 50522 2932 50528 2984
rect 50580 2972 50586 2984
rect 195238 2972 195244 2984
rect 50580 2944 195244 2972
rect 50580 2932 50586 2944
rect 195238 2932 195244 2944
rect 195296 2932 195302 2984
rect 35943 2876 37504 2904
rect 35943 2873 35955 2876
rect 35897 2867 35955 2873
rect 43346 2864 43352 2916
rect 43404 2904 43410 2916
rect 174906 2904 174912 2916
rect 43404 2876 174912 2904
rect 43404 2864 43410 2876
rect 174906 2864 174912 2876
rect 174964 2864 174970 2916
rect 8110 2796 8116 2848
rect 8168 2836 8174 2848
rect 17218 2836 17224 2848
rect 8168 2808 17224 2836
rect 8168 2796 8174 2808
rect 17218 2796 17224 2808
rect 17276 2796 17282 2848
rect 36170 2796 36176 2848
rect 36228 2836 36234 2848
rect 154574 2836 154580 2848
rect 36228 2808 154580 2836
rect 36228 2796 36234 2808
rect 154574 2796 154580 2808
rect 154632 2796 154638 2848
<< via1 >>
rect 144828 700680 144880 700732
rect 170312 700680 170364 700732
rect 105452 700612 105504 700664
rect 106188 700612 106240 700664
rect 124128 700612 124180 700664
rect 235172 700612 235224 700664
rect 102048 700544 102100 700596
rect 300124 700544 300176 700596
rect 81348 700476 81400 700528
rect 364984 700476 365036 700528
rect 40500 700408 40552 700460
rect 41328 700408 41380 700460
rect 60648 700408 60700 700460
rect 429844 700408 429896 700460
rect 38568 700340 38620 700392
rect 494796 700340 494848 700392
rect 17868 700272 17920 700324
rect 559656 700272 559708 700324
rect 123024 689732 123076 689784
rect 124128 689732 124180 689784
rect 144092 689732 144144 689784
rect 144828 689732 144880 689784
rect 59636 689664 59688 689716
rect 60648 689664 60700 689716
rect 106188 689664 106240 689716
rect 165252 689664 165304 689716
rect 41328 689596 41380 689648
rect 186320 689596 186372 689648
rect 2688 689528 2740 689580
rect 228548 689528 228600 689580
rect 8116 689460 8168 689512
rect 249708 689460 249760 689512
rect 9220 689392 9272 689444
rect 270776 689392 270828 689444
rect 9680 689324 9732 689376
rect 291936 689324 291988 689376
rect 9588 689256 9640 689308
rect 313004 689256 313056 689308
rect 9036 689188 9088 689240
rect 334164 689188 334216 689240
rect 8208 689120 8260 689172
rect 355232 689120 355284 689172
rect 207480 689052 207532 689104
rect 576124 689052 576176 689104
rect 4068 688984 4120 689036
rect 376392 688984 376444 689036
rect 8944 688916 8996 688968
rect 397460 688916 397512 688968
rect 9312 688848 9364 688900
rect 418620 688848 418672 688900
rect 9128 688780 9180 688832
rect 439688 688780 439740 688832
rect 9404 688712 9456 688764
rect 460848 688712 460900 688764
rect 9496 688644 9548 688696
rect 481916 688644 481968 688696
rect 3148 681708 3200 681760
rect 6184 681708 6236 681760
rect 3976 567196 4028 567248
rect 6276 567196 6328 567248
rect 3516 509260 3568 509312
rect 7564 509260 7616 509312
rect 576124 487092 576176 487144
rect 579712 487092 579764 487144
rect 578148 238212 578200 238264
rect 580632 238212 580684 238264
rect 578148 213868 578200 213920
rect 580724 213868 580776 213920
rect 578148 189796 578200 189848
rect 580816 189796 580868 189848
rect 3332 181092 3384 181144
rect 4160 181092 4212 181144
rect 578148 165452 578200 165504
rect 580908 165452 580960 165504
rect 3240 121388 3292 121440
rect 4160 121388 4212 121440
rect 578148 116900 578200 116952
rect 580632 116900 580684 116952
rect 578148 92420 578200 92472
rect 580724 92420 580776 92472
rect 578148 68348 578200 68400
rect 580632 68348 580684 68400
rect 578148 44004 578200 44056
rect 580632 44004 580684 44056
rect 52736 6808 52788 6860
rect 580540 6808 580592 6860
rect 62948 6740 63000 6792
rect 580448 6740 580500 6792
rect 73068 6672 73120 6724
rect 580356 6672 580408 6724
rect 83280 6604 83332 6656
rect 580264 6604 580316 6656
rect 4528 6536 4580 6588
rect 90916 6536 90968 6588
rect 92112 6536 92164 6588
rect 578332 6536 578384 6588
rect 84936 6468 84988 6520
rect 578424 6468 578476 6520
rect 81440 6400 81492 6452
rect 578516 6400 578568 6452
rect 56416 6332 56468 6384
rect 578608 6332 578660 6384
rect 52828 6264 52880 6316
rect 578700 6264 578752 6316
rect 33876 6196 33928 6248
rect 579436 6196 579488 6248
rect 30288 6128 30340 6180
rect 579528 6128 579580 6180
rect 4436 6060 4488 6112
rect 87328 6060 87380 6112
rect 94504 6060 94556 6112
rect 579344 6060 579396 6112
rect 4712 5992 4764 6044
rect 105176 5992 105228 6044
rect 108764 5992 108816 6044
rect 579252 5992 579304 6044
rect 4620 5924 4672 5976
rect 101588 5924 101640 5976
rect 112352 5924 112404 5976
rect 579160 5924 579212 5976
rect 4804 5856 4856 5908
rect 115940 5856 115992 5908
rect 119436 5856 119488 5908
rect 579068 5856 579120 5908
rect 4896 5788 4948 5840
rect 123024 5788 123076 5840
rect 5172 5720 5224 5772
rect 117136 5720 117188 5772
rect 7564 5448 7616 5500
rect 42524 5448 42576 5500
rect 89720 5448 89772 5500
rect 307208 5448 307260 5500
rect 6276 5380 6328 5432
rect 32404 5380 32456 5432
rect 96896 5380 96948 5432
rect 327540 5380 327592 5432
rect 3424 5312 3476 5364
rect 22192 5312 22244 5364
rect 103980 5312 104032 5364
rect 347964 5312 348016 5364
rect 6184 5244 6236 5296
rect 12072 5244 12124 5296
rect 24308 5244 24360 5296
rect 124036 5244 124088 5296
rect 124128 5244 124180 5296
rect 398840 5244 398892 5296
rect 65984 5176 66036 5228
rect 459928 5176 459980 5228
rect 69480 5108 69532 5160
rect 470048 5108 470100 5160
rect 98092 5040 98144 5092
rect 500592 5040 500644 5092
rect 48136 4972 48188 5024
rect 449716 4972 449768 5024
rect 4252 4904 4304 4956
rect 51632 4904 51684 4956
rect 83832 4904 83884 4956
rect 490472 4904 490524 4956
rect 4344 4836 4396 4888
rect 55220 4836 55272 4888
rect 73068 4836 73120 4888
rect 480260 4836 480312 4888
rect 572 4768 624 4820
rect 419172 4768 419224 4820
rect 82636 4700 82688 4752
rect 286876 4700 286928 4752
rect 75460 4632 75512 4684
rect 266544 4632 266596 4684
rect 68284 4564 68336 4616
rect 246120 4564 246172 4616
rect 46940 4496 46992 4548
rect 185032 4496 185084 4548
rect 39764 4428 39816 4480
rect 164700 4428 164752 4480
rect 19524 4360 19576 4412
rect 113088 4360 113140 4412
rect 113916 4360 113968 4412
rect 225788 4360 225840 4412
rect 32680 4292 32732 4344
rect 144368 4292 144420 4344
rect 29092 4224 29144 4276
rect 134156 4224 134208 4276
rect 103612 4156 103664 4208
rect 110420 4156 110472 4208
rect 205456 4156 205508 4208
rect 6920 4088 6972 4140
rect 70676 4088 70728 4140
rect 100484 4088 100536 4140
rect 337752 4088 337804 4140
rect 4988 4020 5040 4072
rect 8852 4020 8904 4072
rect 9036 4020 9088 4072
rect 113916 4020 113968 4072
rect 8208 3952 8260 4004
rect 80244 3952 80296 4004
rect 107568 3952 107620 4004
rect 358084 4020 358136 4072
rect 6828 3884 6880 3936
rect 88524 3884 88576 3936
rect 14832 3816 14884 3868
rect 110420 3884 110472 3936
rect 111156 3884 111208 3936
rect 368296 3952 368348 4004
rect 113548 3816 113600 3868
rect 114560 3816 114612 3868
rect 114744 3816 114796 3868
rect 378508 3884 378560 3936
rect 118240 3816 118292 3868
rect 388628 3816 388680 3868
rect 5264 3748 5316 3800
rect 120632 3748 120684 3800
rect 121828 3748 121880 3800
rect 124128 3748 124180 3800
rect 125416 3748 125468 3800
rect 409052 3748 409104 3800
rect 10048 3680 10100 3732
rect 93124 3680 93176 3732
rect 93308 3680 93360 3732
rect 102784 3680 102836 3732
rect 551560 3680 551612 3732
rect 9588 3612 9640 3664
rect 62396 3612 62448 3664
rect 63592 3612 63644 3664
rect 541348 3612 541400 3664
rect 5356 3544 5408 3596
rect 11244 3544 11296 3596
rect 13636 3544 13688 3596
rect 510804 3544 510856 3596
rect 1676 3476 1728 3528
rect 2688 3476 2740 3528
rect 5448 3476 5500 3528
rect 16028 3476 16080 3528
rect 31484 3476 31536 3528
rect 578884 3476 578936 3528
rect 6552 3408 6604 3460
rect 26700 3408 26752 3460
rect 27896 3408 27948 3460
rect 578976 3408 579028 3460
rect 6736 3340 6788 3392
rect 49332 3340 49384 3392
rect 54024 3340 54076 3392
rect 317420 3340 317472 3392
rect 9128 3272 9180 3324
rect 60004 3272 60056 3324
rect 61200 3272 61252 3324
rect 9680 3204 9732 3256
rect 58808 3204 58860 3256
rect 76656 3272 76708 3324
rect 86132 3272 86184 3324
rect 297088 3272 297140 3324
rect 5080 3136 5132 3188
rect 45744 3136 45796 3188
rect 79048 3204 79100 3256
rect 276664 3204 276716 3256
rect 71872 3136 71924 3188
rect 256332 3136 256384 3188
rect 7012 3068 7064 3120
rect 44548 3068 44600 3120
rect 64788 3068 64840 3120
rect 236000 3068 236052 3120
rect 6644 3000 6696 3052
rect 40960 3000 41012 3052
rect 57612 3000 57664 3052
rect 215576 3000 215628 3052
rect 7104 2932 7156 2984
rect 37372 2932 37424 2984
rect 9220 2864 9272 2916
rect 21916 2864 21968 2916
rect 50528 2932 50580 2984
rect 195244 2932 195296 2984
rect 43352 2864 43404 2916
rect 174912 2864 174964 2916
rect 8116 2796 8168 2848
rect 17224 2796 17276 2848
rect 36176 2796 36228 2848
rect 154580 2796 154632 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 40512 700466 40540 703520
rect 105464 700670 105492 703520
rect 170324 700738 170352 703520
rect 144828 700732 144880 700738
rect 144828 700674 144880 700680
rect 170312 700732 170364 700738
rect 170312 700674 170364 700680
rect 105452 700664 105504 700670
rect 105452 700606 105504 700612
rect 106188 700664 106240 700670
rect 106188 700606 106240 700612
rect 124128 700664 124180 700670
rect 124128 700606 124180 700612
rect 102048 700596 102100 700602
rect 102048 700538 102100 700544
rect 81348 700528 81400 700534
rect 81348 700470 81400 700476
rect 40500 700460 40552 700466
rect 40500 700402 40552 700408
rect 41328 700460 41380 700466
rect 41328 700402 41380 700408
rect 60648 700460 60700 700466
rect 60648 700402 60700 700408
rect 38568 700392 38620 700398
rect 38568 700334 38620 700340
rect 17868 700324 17920 700330
rect 17868 700266 17920 700272
rect 2688 689580 2740 689586
rect 2688 689522 2740 689528
rect 572 4820 624 4826
rect 572 4762 624 4768
rect 584 480 612 4762
rect 2700 3534 2728 689522
rect 8116 689512 8168 689518
rect 8116 689454 8168 689460
rect 4068 689036 4120 689042
rect 4068 688978 4120 688984
rect 3146 682272 3202 682281
rect 3146 682207 3202 682216
rect 3160 681766 3188 682207
rect 3148 681760 3200 681766
rect 3148 681702 3200 681708
rect 3422 624880 3478 624889
rect 3422 624815 3478 624824
rect 3238 208176 3294 208185
rect 3238 208111 3294 208120
rect 3146 165064 3202 165073
rect 3146 164999 3202 165008
rect 3160 141545 3188 164999
rect 3146 141536 3202 141545
rect 3146 141471 3202 141480
rect 3252 121446 3280 208111
rect 3332 181144 3384 181150
rect 3332 181086 3384 181092
rect 3240 121440 3292 121446
rect 3240 121382 3292 121388
rect 3344 78985 3372 181086
rect 3330 78976 3386 78985
rect 3330 78911 3386 78920
rect 2870 5400 2926 5409
rect 3436 5370 3464 624815
rect 3974 567352 4030 567361
rect 3974 567287 4030 567296
rect 3988 567254 4016 567287
rect 3976 567248 4028 567254
rect 3976 567190 4028 567196
rect 3514 509960 3570 509969
rect 3514 509895 3570 509904
rect 3528 509318 3556 509895
rect 3516 509312 3568 509318
rect 3516 509254 3568 509260
rect 3514 452432 3570 452441
rect 3514 452367 3570 452376
rect 3528 17921 3556 452367
rect 3606 395040 3662 395049
rect 3606 394975 3662 394984
rect 3620 38321 3648 394975
rect 3698 337512 3754 337521
rect 3698 337447 3754 337456
rect 3712 59129 3740 337447
rect 3790 294400 3846 294409
rect 3790 294335 3846 294344
rect 3804 79665 3832 294335
rect 3974 251288 4030 251297
rect 3974 251223 4030 251232
rect 3882 202056 3938 202065
rect 3882 201991 3938 202000
rect 3790 79656 3846 79665
rect 3790 79591 3846 79600
rect 3698 59120 3754 59129
rect 3698 59055 3754 59064
rect 3606 38312 3662 38321
rect 3606 38247 3662 38256
rect 3896 35873 3924 201991
rect 3988 100337 4016 251223
rect 3974 100328 4030 100337
rect 3974 100263 4030 100272
rect 3882 35864 3938 35873
rect 3882 35799 3938 35808
rect 3514 17912 3570 17921
rect 3514 17847 3570 17856
rect 2870 5335 2926 5344
rect 3424 5364 3476 5370
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 1688 480 1716 3470
rect 2884 480 2912 5335
rect 3424 5306 3476 5312
rect 4080 480 4108 688978
rect 6184 681760 6236 681766
rect 6184 681702 6236 681708
rect 5446 676424 5502 676433
rect 5446 676359 5502 676368
rect 5354 655616 5410 655625
rect 5354 655551 5410 655560
rect 5262 614136 5318 614145
rect 5262 614071 5318 614080
rect 5170 593600 5226 593609
rect 5170 593535 5226 593544
rect 5078 511184 5134 511193
rect 5078 511119 5134 511128
rect 4986 490512 5042 490521
rect 4986 490447 5042 490456
rect 4894 469976 4950 469985
rect 4894 469911 4950 469920
rect 4802 449984 4858 449993
rect 4802 449919 4858 449928
rect 4710 429312 4766 429321
rect 4710 429247 4766 429256
rect 4618 408640 4674 408649
rect 4618 408575 4674 408584
rect 4526 387832 4582 387841
rect 4526 387767 4582 387776
rect 4434 367296 4490 367305
rect 4434 367231 4490 367240
rect 4342 346488 4398 346497
rect 4342 346423 4398 346432
rect 4250 325816 4306 325825
rect 4250 325751 4306 325760
rect 4158 181520 4214 181529
rect 4158 181455 4214 181464
rect 4172 181150 4200 181455
rect 4160 181144 4212 181150
rect 4160 181086 4212 181092
rect 4158 160848 4214 160857
rect 4158 160783 4214 160792
rect 4172 122097 4200 160783
rect 4158 122088 4214 122097
rect 4158 122023 4214 122032
rect 4160 121440 4212 121446
rect 4160 121382 4212 121388
rect 4172 120873 4200 121382
rect 4158 120864 4214 120873
rect 4158 120799 4214 120808
rect 4264 4962 4292 325751
rect 4252 4956 4304 4962
rect 4252 4898 4304 4904
rect 4356 4894 4384 346423
rect 4448 6118 4476 367231
rect 4540 6594 4568 387767
rect 4528 6588 4580 6594
rect 4528 6530 4580 6536
rect 4436 6112 4488 6118
rect 4436 6054 4488 6060
rect 4632 5982 4660 408575
rect 4724 6050 4752 429247
rect 4712 6044 4764 6050
rect 4712 5986 4764 5992
rect 4620 5976 4672 5982
rect 4620 5918 4672 5924
rect 4816 5914 4844 449919
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 4908 5846 4936 469911
rect 4896 5840 4948 5846
rect 4896 5782 4948 5788
rect 4344 4888 4396 4894
rect 4344 4830 4396 4836
rect 5000 4078 5028 490447
rect 4988 4072 5040 4078
rect 4988 4014 5040 4020
rect 5092 3194 5120 511119
rect 5184 5778 5212 593535
rect 5172 5772 5224 5778
rect 5172 5714 5224 5720
rect 5276 3806 5304 614071
rect 5264 3800 5316 3806
rect 5264 3742 5316 3748
rect 5368 3602 5396 655551
rect 5356 3596 5408 3602
rect 5356 3538 5408 3544
rect 5460 3534 5488 676359
rect 6196 5302 6224 681702
rect 6826 573336 6882 573345
rect 6826 573271 6882 573280
rect 6276 567248 6328 567254
rect 6276 567190 6328 567196
rect 6288 5438 6316 567190
rect 6734 532128 6790 532137
rect 6734 532063 6790 532072
rect 6642 284880 6698 284889
rect 6642 284815 6698 284824
rect 6550 243672 6606 243681
rect 6550 243607 6606 243616
rect 6276 5432 6328 5438
rect 6276 5374 6328 5380
rect 6184 5296 6236 5302
rect 6184 5238 6236 5244
rect 6458 4856 6514 4865
rect 6458 4791 6514 4800
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5262 3360 5318 3369
rect 5262 3295 5318 3304
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 5276 480 5304 3295
rect 6472 480 6500 4791
rect 6564 3466 6592 243607
rect 6552 3460 6604 3466
rect 6552 3402 6604 3408
rect 6656 3058 6684 284815
rect 6748 3398 6776 532063
rect 6840 3942 6868 573271
rect 6918 552392 6974 552401
rect 6918 552327 6974 552336
rect 6932 4146 6960 552327
rect 7564 509312 7616 509318
rect 7564 509254 7616 509260
rect 7010 305144 7066 305153
rect 7010 305079 7066 305088
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 7024 3126 7052 305079
rect 7102 263936 7158 263945
rect 7102 263871 7158 263880
rect 7012 3120 7064 3126
rect 7012 3062 7064 3068
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 7116 2990 7144 263871
rect 7194 222728 7250 222737
rect 7194 222663 7250 222672
rect 7208 3210 7236 222663
rect 7576 5506 7604 509254
rect 7564 5500 7616 5506
rect 7564 5442 7616 5448
rect 7208 3182 7696 3210
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 7668 480 7696 3182
rect 8128 2854 8156 689454
rect 9220 689444 9272 689450
rect 9220 689386 9272 689392
rect 9036 689240 9088 689246
rect 9036 689182 9088 689188
rect 8208 689172 8260 689178
rect 8208 689114 8260 689120
rect 8220 4010 8248 689114
rect 8944 688968 8996 688974
rect 8944 688910 8996 688916
rect 8852 4072 8904 4078
rect 8852 4014 8904 4020
rect 8208 4004 8260 4010
rect 8208 3946 8260 3952
rect 8116 2848 8168 2854
rect 8116 2790 8168 2796
rect 8864 480 8892 4014
rect 8956 3505 8984 688910
rect 9048 4078 9076 689182
rect 9128 688832 9180 688838
rect 9128 688774 9180 688780
rect 9036 4072 9088 4078
rect 9036 4014 9088 4020
rect 8942 3496 8998 3505
rect 8942 3431 8998 3440
rect 9140 3330 9168 688774
rect 9128 3324 9180 3330
rect 9128 3266 9180 3272
rect 9232 2922 9260 689386
rect 9680 689376 9732 689382
rect 9680 689318 9732 689324
rect 9588 689308 9640 689314
rect 9588 689250 9640 689256
rect 9312 688900 9364 688906
rect 9312 688842 9364 688848
rect 9324 3641 9352 688842
rect 9404 688764 9456 688770
rect 9404 688706 9456 688712
rect 9416 4049 9444 688706
rect 9496 688696 9548 688702
rect 9496 688638 9548 688644
rect 9402 4040 9458 4049
rect 9402 3975 9458 3984
rect 9508 3913 9536 688638
rect 9494 3904 9550 3913
rect 9494 3839 9550 3848
rect 9600 3670 9628 689250
rect 9588 3664 9640 3670
rect 9310 3632 9366 3641
rect 9588 3606 9640 3612
rect 9310 3567 9366 3576
rect 9692 3262 9720 689318
rect 17880 686882 17908 700266
rect 17526 686854 17908 686882
rect 38580 686868 38608 700334
rect 41340 689654 41368 700402
rect 60660 689722 60688 700402
rect 59636 689716 59688 689722
rect 59636 689658 59688 689664
rect 60648 689716 60700 689722
rect 60648 689658 60700 689664
rect 41328 689648 41380 689654
rect 41328 689590 41380 689596
rect 59648 686868 59676 689658
rect 81360 686746 81388 700470
rect 102060 686882 102088 700538
rect 106200 689722 106228 700606
rect 124140 689790 124168 700606
rect 144840 689790 144868 700674
rect 235184 700670 235212 703520
rect 235172 700664 235224 700670
rect 235172 700606 235224 700612
rect 300136 700602 300164 703520
rect 300124 700596 300176 700602
rect 300124 700538 300176 700544
rect 364996 700534 365024 703520
rect 364984 700528 365036 700534
rect 364984 700470 365036 700476
rect 429856 700466 429884 703520
rect 429844 700460 429896 700466
rect 429844 700402 429896 700408
rect 494808 700398 494836 703520
rect 494796 700392 494848 700398
rect 494796 700334 494848 700340
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 123024 689784 123076 689790
rect 123024 689726 123076 689732
rect 124128 689784 124180 689790
rect 124128 689726 124180 689732
rect 144092 689784 144144 689790
rect 144092 689726 144144 689732
rect 144828 689784 144880 689790
rect 144828 689726 144880 689732
rect 106188 689716 106240 689722
rect 106188 689658 106240 689664
rect 101890 686854 102088 686882
rect 123036 686868 123064 689726
rect 144104 686868 144132 689726
rect 165252 689716 165304 689722
rect 165252 689658 165304 689664
rect 165264 686868 165292 689658
rect 186320 689648 186372 689654
rect 186320 689590 186372 689596
rect 186332 686868 186360 689590
rect 228548 689580 228600 689586
rect 228548 689522 228600 689528
rect 207480 689104 207532 689110
rect 207480 689046 207532 689052
rect 207492 686868 207520 689046
rect 228560 686868 228588 689522
rect 249708 689512 249760 689518
rect 249708 689454 249760 689460
rect 249720 686868 249748 689454
rect 270776 689444 270828 689450
rect 270776 689386 270828 689392
rect 270788 686868 270816 689386
rect 291936 689376 291988 689382
rect 291936 689318 291988 689324
rect 291948 686868 291976 689318
rect 313004 689308 313056 689314
rect 313004 689250 313056 689256
rect 313016 686868 313044 689250
rect 334164 689240 334216 689246
rect 334164 689182 334216 689188
rect 334176 686868 334204 689182
rect 355232 689172 355284 689178
rect 355232 689114 355284 689120
rect 355244 686868 355272 689114
rect 576124 689104 576176 689110
rect 503074 689072 503130 689081
rect 376392 689036 376444 689042
rect 576124 689046 576176 689052
rect 503074 689007 503130 689016
rect 376392 688978 376444 688984
rect 376404 686868 376432 688978
rect 397460 688968 397512 688974
rect 397460 688910 397512 688916
rect 397472 686868 397500 688910
rect 418620 688900 418672 688906
rect 418620 688842 418672 688848
rect 418632 686868 418660 688842
rect 439688 688832 439740 688838
rect 439688 688774 439740 688780
rect 439700 686868 439728 688774
rect 460848 688764 460900 688770
rect 460848 688706 460900 688712
rect 460860 686868 460888 688706
rect 481916 688696 481968 688702
rect 481916 688638 481968 688644
rect 481928 686868 481956 688638
rect 503088 686868 503116 689007
rect 545302 688936 545358 688945
rect 545302 688871 545358 688880
rect 524142 688800 524198 688809
rect 524142 688735 524198 688744
rect 524156 686868 524184 688735
rect 545316 686868 545344 688871
rect 566370 688664 566426 688673
rect 566370 688599 566426 688608
rect 566384 686868 566412 688599
rect 80822 686718 81388 686746
rect 576136 487150 576164 689046
rect 580262 674656 580318 674665
rect 580262 674591 580318 674600
rect 578238 601760 578294 601769
rect 578238 601695 578294 601704
rect 576124 487144 576176 487150
rect 576124 487086 576176 487092
rect 578148 238264 578200 238270
rect 578146 238232 578148 238241
rect 578200 238232 578202 238241
rect 578146 238167 578202 238176
rect 578148 213920 578200 213926
rect 578146 213888 578148 213897
rect 578200 213888 578202 213897
rect 578146 213823 578202 213832
rect 578148 189848 578200 189854
rect 578146 189816 578148 189825
rect 578200 189816 578202 189825
rect 578146 189751 578202 189760
rect 578148 165504 578200 165510
rect 578146 165472 578148 165481
rect 578200 165472 578202 165481
rect 578146 165407 578202 165416
rect 578148 116952 578200 116958
rect 578146 116920 578148 116929
rect 578200 116920 578202 116929
rect 578146 116855 578202 116864
rect 578148 92472 578200 92478
rect 578146 92440 578148 92449
rect 578200 92440 578202 92449
rect 578146 92375 578202 92384
rect 578148 68400 578200 68406
rect 578146 68368 578148 68377
rect 578200 68368 578202 68377
rect 578146 68303 578202 68312
rect 578148 44056 578200 44062
rect 578146 44024 578148 44033
rect 578200 44024 578202 44033
rect 578146 43959 578202 43968
rect 109958 7712 110014 7721
rect 109958 7647 110014 7656
rect 106370 7576 106426 7585
rect 106370 7511 106426 7520
rect 93136 7126 93518 7154
rect 12084 5302 12112 7004
rect 12438 5536 12494 5545
rect 12438 5471 12494 5480
rect 12072 5296 12124 5302
rect 12072 5238 12124 5244
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 9680 3256 9732 3262
rect 9680 3198 9732 3204
rect 9220 2916 9272 2922
rect 9220 2858 9272 2864
rect 10060 480 10088 3674
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 11256 480 11284 3538
rect 12452 480 12480 5471
rect 22204 5370 22232 7004
rect 30288 6180 30340 6186
rect 30288 6122 30340 6128
rect 22192 5364 22244 5370
rect 22192 5306 22244 5312
rect 24308 5296 24360 5302
rect 24308 5238 24360 5244
rect 19524 4412 19576 4418
rect 19524 4354 19576 4360
rect 14832 3868 14884 3874
rect 14832 3810 14884 3816
rect 13636 3596 13688 3602
rect 13636 3538 13688 3544
rect 13648 480 13676 3538
rect 14844 480 14872 3810
rect 16028 3528 16080 3534
rect 16028 3470 16080 3476
rect 18326 3496 18382 3505
rect 16040 480 16068 3470
rect 18326 3431 18382 3440
rect 17224 2848 17276 2854
rect 17224 2790 17276 2796
rect 17236 480 17264 2790
rect 18340 480 18368 3431
rect 19536 480 19564 4354
rect 23110 3632 23166 3641
rect 23110 3567 23166 3576
rect 20718 3496 20774 3505
rect 20718 3431 20774 3440
rect 20732 480 20760 3431
rect 21916 2916 21968 2922
rect 21916 2858 21968 2864
rect 21928 480 21956 2858
rect 23124 480 23152 3567
rect 24320 480 24348 5238
rect 29092 4276 29144 4282
rect 29092 4218 29144 4224
rect 25502 3632 25558 3641
rect 25502 3567 25558 3576
rect 25516 480 25544 3567
rect 26700 3460 26752 3466
rect 26700 3402 26752 3408
rect 27896 3460 27948 3466
rect 27896 3402 27948 3408
rect 26712 480 26740 3402
rect 27908 480 27936 3402
rect 29104 480 29132 4218
rect 30300 480 30328 6122
rect 32416 5438 32444 7004
rect 33876 6248 33928 6254
rect 33876 6190 33928 6196
rect 32404 5432 32456 5438
rect 32404 5374 32456 5380
rect 32680 4344 32732 4350
rect 32680 4286 32732 4292
rect 31484 3528 31536 3534
rect 31484 3470 31536 3476
rect 31496 480 31524 3470
rect 32692 480 32720 4286
rect 33888 480 33916 6190
rect 42536 5506 42564 7004
rect 52748 6866 52776 7004
rect 52736 6860 52788 6866
rect 52736 6802 52788 6808
rect 62960 6798 62988 7004
rect 62948 6792 63000 6798
rect 62948 6734 63000 6740
rect 73080 6730 73108 7004
rect 73068 6724 73120 6730
rect 73068 6666 73120 6672
rect 83292 6662 83320 7004
rect 83280 6656 83332 6662
rect 83280 6598 83332 6604
rect 90916 6588 90968 6594
rect 90916 6530 90968 6536
rect 92112 6588 92164 6594
rect 92112 6530 92164 6536
rect 84936 6520 84988 6526
rect 84936 6462 84988 6468
rect 81440 6452 81492 6458
rect 81440 6394 81492 6400
rect 56416 6384 56468 6390
rect 56416 6326 56468 6332
rect 52828 6316 52880 6322
rect 52828 6258 52880 6264
rect 42524 5500 42576 5506
rect 42524 5442 42576 5448
rect 34978 5128 35034 5137
rect 34978 5063 35034 5072
rect 34992 480 35020 5063
rect 48136 5024 48188 5030
rect 38566 4992 38622 5001
rect 48136 4966 48188 4972
rect 38566 4927 38622 4936
rect 37372 2984 37424 2990
rect 37372 2926 37424 2932
rect 36176 2848 36228 2854
rect 36176 2790 36228 2796
rect 36188 480 36216 2790
rect 37384 480 37412 2926
rect 38580 480 38608 4927
rect 46940 4548 46992 4554
rect 46940 4490 46992 4496
rect 39764 4480 39816 4486
rect 39764 4422 39816 4428
rect 39776 480 39804 4422
rect 42154 3768 42210 3777
rect 42154 3703 42210 3712
rect 40960 3052 41012 3058
rect 40960 2994 41012 3000
rect 40972 480 41000 2994
rect 42168 480 42196 3703
rect 45744 3188 45796 3194
rect 45744 3130 45796 3136
rect 44548 3120 44600 3126
rect 44548 3062 44600 3068
rect 43352 2916 43404 2922
rect 43352 2858 43404 2864
rect 43364 480 43392 2858
rect 44560 480 44588 3062
rect 45756 480 45784 3130
rect 46952 480 46980 4490
rect 48148 480 48176 4966
rect 51632 4956 51684 4962
rect 51632 4898 51684 4904
rect 49332 3392 49384 3398
rect 49332 3334 49384 3340
rect 49344 480 49372 3334
rect 50528 2984 50580 2990
rect 50528 2926 50580 2932
rect 50540 480 50568 2926
rect 51644 480 51672 4898
rect 52840 480 52868 6258
rect 55220 4888 55272 4894
rect 55220 4830 55272 4836
rect 54024 3392 54076 3398
rect 54024 3334 54076 3340
rect 54036 480 54064 3334
rect 55232 480 55260 4830
rect 56428 480 56456 6326
rect 65984 5228 66036 5234
rect 65984 5170 66036 5176
rect 62396 3664 62448 3670
rect 62396 3606 62448 3612
rect 63592 3664 63644 3670
rect 63592 3606 63644 3612
rect 60004 3324 60056 3330
rect 60004 3266 60056 3272
rect 61200 3324 61252 3330
rect 61200 3266 61252 3272
rect 58808 3256 58860 3262
rect 58808 3198 58860 3204
rect 57612 3052 57664 3058
rect 57612 2994 57664 3000
rect 57624 480 57652 2994
rect 58820 480 58848 3198
rect 60016 480 60044 3266
rect 61212 480 61240 3266
rect 62408 480 62436 3606
rect 63604 480 63632 3606
rect 64788 3120 64840 3126
rect 64788 3062 64840 3068
rect 64800 480 64828 3062
rect 65996 480 66024 5170
rect 69480 5160 69532 5166
rect 69480 5102 69532 5108
rect 68284 4616 68336 4622
rect 68284 4558 68336 4564
rect 67178 4040 67234 4049
rect 67178 3975 67234 3984
rect 67192 480 67220 3975
rect 68296 480 68324 4558
rect 69492 480 69520 5102
rect 73068 4888 73120 4894
rect 73068 4830 73120 4836
rect 70676 4140 70728 4146
rect 70676 4082 70728 4088
rect 70688 480 70716 4082
rect 71872 3188 71924 3194
rect 71872 3130 71924 3136
rect 71884 480 71912 3130
rect 73080 480 73108 4830
rect 75460 4684 75512 4690
rect 75460 4626 75512 4632
rect 74262 3904 74318 3913
rect 74262 3839 74318 3848
rect 74276 480 74304 3839
rect 75472 480 75500 4626
rect 80244 4004 80296 4010
rect 80244 3946 80296 3952
rect 77850 3904 77906 3913
rect 77850 3839 77906 3848
rect 76656 3324 76708 3330
rect 76656 3266 76708 3272
rect 76668 480 76696 3266
rect 77864 480 77892 3839
rect 79048 3256 79100 3262
rect 79048 3198 79100 3204
rect 79060 480 79088 3198
rect 80256 480 80284 3946
rect 81452 480 81480 6394
rect 83832 4956 83884 4962
rect 83832 4898 83884 4904
rect 82636 4752 82688 4758
rect 82636 4694 82688 4700
rect 82648 480 82676 4694
rect 83844 480 83872 4898
rect 84948 480 84976 6462
rect 87328 6112 87380 6118
rect 87328 6054 87380 6060
rect 86132 3324 86184 3330
rect 86132 3266 86184 3272
rect 86144 480 86172 3266
rect 87340 480 87368 6054
rect 89720 5500 89772 5506
rect 89720 5442 89772 5448
rect 88524 3936 88576 3942
rect 88524 3878 88576 3884
rect 88536 480 88564 3878
rect 89732 480 89760 5442
rect 90928 480 90956 6530
rect 92124 480 92152 6530
rect 93136 3738 93164 7126
rect 94504 6112 94556 6118
rect 94504 6054 94556 6060
rect 93124 3732 93176 3738
rect 93124 3674 93176 3680
rect 93308 3732 93360 3738
rect 93308 3674 93360 3680
rect 93320 480 93348 3674
rect 94516 480 94544 6054
rect 101588 5976 101640 5982
rect 101588 5918 101640 5924
rect 96896 5432 96948 5438
rect 96896 5374 96948 5380
rect 95698 4040 95754 4049
rect 95698 3975 95754 3984
rect 95712 480 95740 3975
rect 96908 480 96936 5374
rect 98092 5092 98144 5098
rect 98092 5034 98144 5040
rect 98104 480 98132 5034
rect 100484 4140 100536 4146
rect 100484 4082 100536 4088
rect 99286 3224 99342 3233
rect 99286 3159 99342 3168
rect 99300 480 99328 3159
rect 100496 480 100524 4082
rect 101600 480 101628 5918
rect 103624 4214 103652 7004
rect 105176 6044 105228 6050
rect 105176 5986 105228 5992
rect 103980 5364 104032 5370
rect 103980 5306 104032 5312
rect 103612 4208 103664 4214
rect 103612 4150 103664 4156
rect 102784 3732 102836 3738
rect 102784 3674 102836 3680
rect 102796 480 102824 3674
rect 103992 480 104020 5306
rect 105188 480 105216 5986
rect 106384 480 106412 7511
rect 108764 6044 108816 6050
rect 108764 5986 108816 5992
rect 107568 4004 107620 4010
rect 107568 3946 107620 3952
rect 107580 480 107608 3946
rect 108776 480 108804 5986
rect 109972 480 110000 7647
rect 113192 7126 113850 7154
rect 112352 5976 112404 5982
rect 112352 5918 112404 5924
rect 110420 4208 110472 4214
rect 110420 4150 110472 4156
rect 110432 3942 110460 4150
rect 110420 3936 110472 3942
rect 110420 3878 110472 3884
rect 111156 3936 111208 3942
rect 111156 3878 111208 3884
rect 111168 480 111196 3878
rect 112364 480 112392 5918
rect 113192 4570 113220 7126
rect 115940 5908 115992 5914
rect 115940 5850 115992 5856
rect 119436 5908 119488 5914
rect 119436 5850 119488 5856
rect 114558 5264 114614 5273
rect 114558 5199 114614 5208
rect 113100 4542 113220 4570
rect 113100 4418 113128 4542
rect 113088 4412 113140 4418
rect 113088 4354 113140 4360
rect 113916 4412 113968 4418
rect 113916 4354 113968 4360
rect 113928 4078 113956 4354
rect 113916 4072 113968 4078
rect 113916 4014 113968 4020
rect 114572 3874 114600 5199
rect 113548 3868 113600 3874
rect 113548 3810 113600 3816
rect 114560 3868 114612 3874
rect 114560 3810 114612 3816
rect 114744 3868 114796 3874
rect 114744 3810 114796 3816
rect 113560 480 113588 3810
rect 114756 480 114784 3810
rect 115952 480 115980 5850
rect 117136 5772 117188 5778
rect 117136 5714 117188 5720
rect 117148 480 117176 5714
rect 118240 3868 118292 3874
rect 118240 3810 118292 3816
rect 118252 480 118280 3810
rect 119448 480 119476 5850
rect 123024 5840 123076 5846
rect 123024 5782 123076 5788
rect 120632 3800 120684 3806
rect 120632 3742 120684 3748
rect 121828 3800 121880 3806
rect 121828 3742 121880 3748
rect 120644 480 120672 3742
rect 121840 480 121868 3742
rect 123036 480 123064 5782
rect 124048 5302 124076 7004
rect 124036 5296 124088 5302
rect 124036 5238 124088 5244
rect 124128 5296 124180 5302
rect 124128 5238 124180 5244
rect 124140 3806 124168 5238
rect 134168 4282 134196 7004
rect 144380 4350 144408 7004
rect 144368 4344 144420 4350
rect 144368 4286 144420 4292
rect 134156 4276 134208 4282
rect 134156 4218 134208 4224
rect 124128 3800 124180 3806
rect 124128 3742 124180 3748
rect 125416 3800 125468 3806
rect 125416 3742 125468 3748
rect 124218 3088 124274 3097
rect 124218 3023 124274 3032
rect 124232 480 124260 3023
rect 125428 480 125456 3742
rect 154592 2854 154620 7004
rect 164712 4486 164740 7004
rect 164700 4480 164752 4486
rect 164700 4422 164752 4428
rect 174924 2922 174952 7004
rect 185044 4554 185072 7004
rect 185032 4548 185084 4554
rect 185032 4490 185084 4496
rect 195256 2990 195284 7004
rect 205468 4214 205496 7004
rect 205456 4208 205508 4214
rect 205456 4150 205508 4156
rect 215588 3058 215616 7004
rect 225800 4418 225828 7004
rect 225788 4412 225840 4418
rect 225788 4354 225840 4360
rect 236012 3126 236040 7004
rect 246132 4622 246160 7004
rect 246120 4616 246172 4622
rect 246120 4558 246172 4564
rect 256344 3194 256372 7004
rect 266556 4690 266584 7004
rect 266544 4684 266596 4690
rect 266544 4626 266596 4632
rect 276676 3262 276704 7004
rect 286888 4758 286916 7004
rect 286876 4752 286928 4758
rect 286876 4694 286928 4700
rect 297100 3330 297128 7004
rect 307220 5506 307248 7004
rect 307208 5500 307260 5506
rect 307208 5442 307260 5448
rect 317432 3398 317460 7004
rect 327552 5438 327580 7004
rect 327540 5432 327592 5438
rect 327540 5374 327592 5380
rect 337764 4146 337792 7004
rect 347976 5370 348004 7004
rect 347964 5364 348016 5370
rect 347964 5306 348016 5312
rect 337752 4140 337804 4146
rect 337752 4082 337804 4088
rect 358096 4078 358124 7004
rect 358084 4072 358136 4078
rect 358084 4014 358136 4020
rect 368308 4010 368336 7004
rect 368296 4004 368348 4010
rect 368296 3946 368348 3952
rect 378520 3942 378548 7004
rect 378508 3936 378560 3942
rect 378508 3878 378560 3884
rect 388640 3874 388668 7004
rect 398852 5302 398880 7004
rect 398840 5296 398892 5302
rect 398840 5238 398892 5244
rect 388628 3868 388680 3874
rect 388628 3810 388680 3816
rect 409064 3806 409092 7004
rect 419184 4826 419212 7004
rect 429396 5409 429424 7004
rect 439608 5545 439636 7004
rect 439594 5536 439650 5545
rect 439594 5471 439650 5480
rect 429382 5400 429438 5409
rect 429382 5335 429438 5344
rect 449728 5030 449756 7004
rect 459940 5234 459968 7004
rect 459928 5228 459980 5234
rect 459928 5170 459980 5176
rect 470060 5166 470088 7004
rect 470048 5160 470100 5166
rect 470048 5102 470100 5108
rect 449716 5024 449768 5030
rect 449716 4966 449768 4972
rect 480272 4894 480300 7004
rect 490484 4962 490512 7004
rect 500604 5098 500632 7004
rect 500592 5092 500644 5098
rect 500592 5034 500644 5040
rect 490472 4956 490524 4962
rect 490472 4898 490524 4904
rect 480260 4888 480312 4894
rect 480260 4830 480312 4836
rect 419172 4820 419224 4826
rect 419172 4762 419224 4768
rect 409052 3800 409104 3806
rect 409052 3742 409104 3748
rect 510816 3602 510844 7004
rect 521028 5137 521056 7004
rect 521014 5128 521070 5137
rect 521014 5063 521070 5072
rect 531148 5001 531176 7004
rect 531134 4992 531190 5001
rect 531134 4927 531190 4936
rect 541360 3670 541388 7004
rect 551572 3738 551600 7004
rect 561692 5273 561720 7004
rect 561678 5264 561734 5273
rect 561678 5199 561734 5208
rect 571904 4865 571932 7004
rect 571890 4856 571946 4865
rect 571890 4791 571946 4800
rect 578252 4049 578280 601695
rect 578330 577280 578386 577289
rect 578330 577215 578386 577224
rect 578344 6594 578372 577215
rect 578422 553480 578478 553489
rect 578422 553415 578478 553424
rect 578332 6588 578384 6594
rect 578332 6530 578384 6536
rect 578436 6526 578464 553415
rect 578514 528864 578570 528873
rect 578514 528799 578570 528808
rect 578424 6520 578476 6526
rect 578424 6462 578476 6468
rect 578528 6458 578556 528799
rect 578606 504248 578662 504257
rect 578606 504183 578662 504192
rect 578516 6452 578568 6458
rect 578516 6394 578568 6400
rect 578620 6390 578648 504183
rect 579712 487144 579764 487150
rect 579712 487086 579764 487092
rect 579724 486849 579752 487086
rect 579710 486840 579766 486849
rect 579710 486775 579766 486784
rect 578698 480448 578754 480457
rect 578698 480383 578754 480392
rect 578608 6384 578660 6390
rect 578608 6326 578660 6332
rect 578712 6322 578740 480383
rect 578790 455696 578846 455705
rect 578790 455631 578846 455640
rect 578700 6316 578752 6322
rect 578700 6258 578752 6264
rect 578238 4040 578294 4049
rect 578238 3975 578294 3984
rect 578804 3777 578832 455631
rect 578882 431352 578938 431361
rect 578882 431287 578938 431296
rect 578790 3768 578846 3777
rect 551560 3732 551612 3738
rect 578790 3703 578846 3712
rect 551560 3674 551612 3680
rect 541348 3664 541400 3670
rect 541348 3606 541400 3612
rect 510804 3596 510856 3602
rect 510804 3538 510856 3544
rect 578896 3534 578924 431287
rect 578974 407144 579030 407153
rect 578974 407079 579030 407088
rect 578884 3528 578936 3534
rect 578884 3470 578936 3476
rect 578988 3466 579016 407079
rect 579066 382800 579122 382809
rect 579066 382735 579122 382744
rect 579080 5914 579108 382735
rect 579158 358864 579214 358873
rect 579158 358799 579214 358808
rect 579172 5982 579200 358799
rect 579250 334248 579306 334257
rect 579250 334183 579306 334192
rect 579264 6050 579292 334183
rect 579342 309904 579398 309913
rect 579342 309839 579398 309848
rect 579356 6118 579384 309839
rect 579434 285696 579490 285705
rect 579434 285631 579490 285640
rect 579448 6254 579476 285631
rect 579526 261352 579582 261361
rect 579526 261287 579582 261296
rect 579436 6248 579488 6254
rect 579436 6190 579488 6196
rect 579540 6186 579568 261287
rect 580170 252240 580226 252249
rect 580170 252175 580226 252184
rect 580184 140729 580212 252175
rect 580170 140720 580226 140729
rect 580170 140655 580226 140664
rect 579618 18592 579674 18601
rect 579618 18527 579674 18536
rect 579632 17649 579660 18527
rect 579618 17640 579674 17649
rect 579618 17575 579674 17584
rect 580276 6662 580304 674591
rect 580354 627736 580410 627745
rect 580354 627671 580410 627680
rect 580368 6730 580396 627671
rect 580446 580816 580502 580825
rect 580446 580751 580502 580760
rect 580460 6798 580488 580751
rect 580538 533896 580594 533905
rect 580538 533831 580594 533840
rect 580552 6866 580580 533831
rect 580630 439920 580686 439929
rect 580630 439855 580686 439864
rect 580644 238270 580672 439855
rect 580722 393000 580778 393009
rect 580722 392935 580778 392944
rect 580632 238264 580684 238270
rect 580632 238206 580684 238212
rect 580736 213926 580764 392935
rect 580814 346080 580870 346089
rect 580814 346015 580870 346024
rect 580724 213920 580776 213926
rect 580724 213862 580776 213868
rect 580630 205320 580686 205329
rect 580630 205255 580686 205264
rect 580644 116958 580672 205255
rect 580828 189854 580856 346015
rect 580906 299160 580962 299169
rect 580906 299095 580962 299104
rect 580816 189848 580868 189854
rect 580816 189790 580868 189796
rect 580920 165510 580948 299095
rect 580908 165504 580960 165510
rect 580908 165446 580960 165452
rect 580722 158400 580778 158409
rect 580722 158335 580778 158344
rect 580632 116952 580684 116958
rect 580632 116894 580684 116900
rect 580630 111480 580686 111489
rect 580630 111415 580686 111424
rect 580644 68406 580672 111415
rect 580736 92478 580764 158335
rect 580724 92472 580776 92478
rect 580724 92414 580776 92420
rect 580632 68400 580684 68406
rect 580632 68342 580684 68348
rect 580630 64560 580686 64569
rect 580630 64495 580686 64504
rect 580644 44062 580672 64495
rect 580632 44056 580684 44062
rect 580632 43998 580684 44004
rect 580540 6860 580592 6866
rect 580540 6802 580592 6808
rect 580448 6792 580500 6798
rect 580448 6734 580500 6740
rect 580356 6724 580408 6730
rect 580356 6666 580408 6672
rect 580264 6656 580316 6662
rect 580264 6598 580316 6604
rect 579528 6180 579580 6186
rect 579528 6122 579580 6128
rect 579344 6112 579396 6118
rect 579344 6054 579396 6060
rect 579252 6044 579304 6050
rect 579252 5986 579304 5992
rect 579160 5976 579212 5982
rect 579160 5918 579212 5924
rect 579068 5908 579120 5914
rect 579068 5850 579120 5856
rect 578976 3460 579028 3466
rect 578976 3402 579028 3408
rect 317420 3392 317472 3398
rect 317420 3334 317472 3340
rect 297088 3324 297140 3330
rect 297088 3266 297140 3272
rect 276664 3256 276716 3262
rect 276664 3198 276716 3204
rect 256332 3188 256384 3194
rect 256332 3130 256384 3136
rect 236000 3120 236052 3126
rect 236000 3062 236052 3068
rect 215576 3052 215628 3058
rect 215576 2994 215628 3000
rect 195244 2984 195296 2990
rect 195244 2926 195296 2932
rect 174912 2916 174964 2922
rect 174912 2858 174964 2864
rect 154580 2848 154632 2854
rect 154580 2790 154632 2796
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3146 682216 3202 682272
rect 3422 624824 3478 624880
rect 3238 208120 3294 208176
rect 3146 165008 3202 165064
rect 3146 141480 3202 141536
rect 3330 78920 3386 78976
rect 2870 5344 2926 5400
rect 3974 567296 4030 567352
rect 3514 509904 3570 509960
rect 3514 452376 3570 452432
rect 3606 394984 3662 395040
rect 3698 337456 3754 337512
rect 3790 294344 3846 294400
rect 3974 251232 4030 251288
rect 3882 202000 3938 202056
rect 3790 79600 3846 79656
rect 3698 59064 3754 59120
rect 3606 38256 3662 38312
rect 3974 100272 4030 100328
rect 3882 35808 3938 35864
rect 3514 17856 3570 17912
rect 5446 676368 5502 676424
rect 5354 655560 5410 655616
rect 5262 614080 5318 614136
rect 5170 593544 5226 593600
rect 5078 511128 5134 511184
rect 4986 490456 5042 490512
rect 4894 469920 4950 469976
rect 4802 449928 4858 449984
rect 4710 429256 4766 429312
rect 4618 408584 4674 408640
rect 4526 387776 4582 387832
rect 4434 367240 4490 367296
rect 4342 346432 4398 346488
rect 4250 325760 4306 325816
rect 4158 181464 4214 181520
rect 4158 160792 4214 160848
rect 4158 122032 4214 122088
rect 4158 120808 4214 120864
rect 6826 573280 6882 573336
rect 6734 532072 6790 532128
rect 6642 284824 6698 284880
rect 6550 243616 6606 243672
rect 6458 4800 6514 4856
rect 5262 3304 5318 3360
rect 6918 552336 6974 552392
rect 7010 305088 7066 305144
rect 7102 263880 7158 263936
rect 7194 222672 7250 222728
rect 8942 3440 8998 3496
rect 9402 3984 9458 4040
rect 9494 3848 9550 3904
rect 9310 3576 9366 3632
rect 503074 689016 503130 689072
rect 545302 688880 545358 688936
rect 524142 688744 524198 688800
rect 566370 688608 566426 688664
rect 580262 674600 580318 674656
rect 578238 601704 578294 601760
rect 578146 238212 578148 238232
rect 578148 238212 578200 238232
rect 578200 238212 578202 238232
rect 578146 238176 578202 238212
rect 578146 213868 578148 213888
rect 578148 213868 578200 213888
rect 578200 213868 578202 213888
rect 578146 213832 578202 213868
rect 578146 189796 578148 189816
rect 578148 189796 578200 189816
rect 578200 189796 578202 189816
rect 578146 189760 578202 189796
rect 578146 165452 578148 165472
rect 578148 165452 578200 165472
rect 578200 165452 578202 165472
rect 578146 165416 578202 165452
rect 578146 116900 578148 116920
rect 578148 116900 578200 116920
rect 578200 116900 578202 116920
rect 578146 116864 578202 116900
rect 578146 92420 578148 92440
rect 578148 92420 578200 92440
rect 578200 92420 578202 92440
rect 578146 92384 578202 92420
rect 578146 68348 578148 68368
rect 578148 68348 578200 68368
rect 578200 68348 578202 68368
rect 578146 68312 578202 68348
rect 578146 44004 578148 44024
rect 578148 44004 578200 44024
rect 578200 44004 578202 44024
rect 578146 43968 578202 44004
rect 109958 7656 110014 7712
rect 106370 7520 106426 7576
rect 12438 5480 12494 5536
rect 18326 3440 18382 3496
rect 23110 3576 23166 3632
rect 20718 3440 20774 3496
rect 25502 3576 25558 3632
rect 34978 5072 35034 5128
rect 38566 4936 38622 4992
rect 42154 3712 42210 3768
rect 67178 3984 67234 4040
rect 74262 3848 74318 3904
rect 77850 3848 77906 3904
rect 95698 3984 95754 4040
rect 99286 3168 99342 3224
rect 114558 5208 114614 5264
rect 124218 3032 124274 3088
rect 439594 5480 439650 5536
rect 429382 5344 429438 5400
rect 521014 5072 521070 5128
rect 531134 4936 531190 4992
rect 561678 5208 561734 5264
rect 571890 4800 571946 4856
rect 578330 577224 578386 577280
rect 578422 553424 578478 553480
rect 578514 528808 578570 528864
rect 578606 504192 578662 504248
rect 579710 486784 579766 486840
rect 578698 480392 578754 480448
rect 578790 455640 578846 455696
rect 578238 3984 578294 4040
rect 578882 431296 578938 431352
rect 578790 3712 578846 3768
rect 578974 407088 579030 407144
rect 579066 382744 579122 382800
rect 579158 358808 579214 358864
rect 579250 334192 579306 334248
rect 579342 309848 579398 309904
rect 579434 285640 579490 285696
rect 579526 261296 579582 261352
rect 580170 252184 580226 252240
rect 580170 140664 580226 140720
rect 579618 18536 579674 18592
rect 579618 17584 579674 17640
rect 580354 627680 580410 627736
rect 580446 580760 580502 580816
rect 580538 533840 580594 533896
rect 580630 439864 580686 439920
rect 580722 392944 580778 393000
rect 580814 346024 580870 346080
rect 580630 205264 580686 205320
rect 580906 299104 580962 299160
rect 580722 158344 580778 158400
rect 580630 111424 580686 111480
rect 580630 64504 580686 64560
<< metal3 >>
rect 583520 697900 584960 698140
rect -960 696540 480 696780
rect 503069 689074 503135 689077
rect 569902 689074 569908 689076
rect 503069 689072 569908 689074
rect 503069 689016 503074 689072
rect 503130 689016 569908 689072
rect 503069 689014 569908 689016
rect 503069 689011 503135 689014
rect 569902 689012 569908 689014
rect 569972 689012 569978 689076
rect 545297 688938 545363 688941
rect 570270 688938 570276 688940
rect 545297 688936 570276 688938
rect 545297 688880 545302 688936
rect 545358 688880 570276 688936
rect 545297 688878 570276 688880
rect 545297 688875 545363 688878
rect 570270 688876 570276 688878
rect 570340 688876 570346 688940
rect 524137 688802 524203 688805
rect 570086 688802 570092 688804
rect 524137 688800 570092 688802
rect 524137 688744 524142 688800
rect 524198 688744 570092 688800
rect 524137 688742 570092 688744
rect 524137 688739 524203 688742
rect 570086 688740 570092 688742
rect 570156 688740 570162 688804
rect 566365 688666 566431 688669
rect 571374 688666 571380 688668
rect 566365 688664 571380 688666
rect 566365 688608 566370 688664
rect 566426 688608 571380 688664
rect 566365 688606 571380 688608
rect 566365 688603 566431 688606
rect 571374 688604 571380 688606
rect 571444 688604 571450 688668
rect 583520 686204 584960 686444
rect -960 682274 480 682364
rect 3141 682274 3207 682277
rect -960 682272 3207 682274
rect -960 682216 3146 682272
rect 3202 682216 3207 682272
rect -960 682214 3207 682216
rect -960 682124 480 682214
rect 3141 682211 3207 682214
rect 5441 676426 5507 676429
rect 7054 676426 7114 676600
rect 5441 676424 7114 676426
rect 5441 676368 5446 676424
rect 5502 676368 7114 676424
rect 5441 676366 7114 676368
rect 5441 676363 5507 676366
rect 578182 674930 578188 674932
rect 576902 674870 578188 674930
rect 576902 674832 576962 674870
rect 578182 674868 578188 674870
rect 578252 674868 578258 674932
rect 580257 674658 580323 674661
rect 583520 674658 584960 674748
rect 580257 674656 584960 674658
rect 580257 674600 580262 674656
rect 580318 674600 584960 674656
rect 580257 674598 584960 674600
rect 580257 674595 580323 674598
rect 583520 674508 584960 674598
rect -960 667844 480 668084
rect 583520 662676 584960 662916
rect 5349 655618 5415 655621
rect 7054 655618 7114 655928
rect 5349 655616 7114 655618
rect 5349 655560 5354 655616
rect 5410 655560 7114 655616
rect 5349 655558 7114 655560
rect 5349 655555 5415 655558
rect -960 653428 480 653668
rect 583520 650980 584960 651220
rect 576902 650042 576962 650488
rect 578366 650042 578372 650044
rect 576902 649982 578372 650042
rect 578366 649980 578372 649982
rect 578436 649980 578442 650044
rect 583520 639284 584960 639524
rect -960 639012 480 639252
rect 5390 634884 5396 634948
rect 5460 634946 5466 634948
rect 7054 634946 7114 635392
rect 5460 634886 7114 634946
rect 5460 634884 5466 634886
rect 580349 627738 580415 627741
rect 583520 627738 584960 627828
rect 580349 627736 584960 627738
rect 580349 627680 580354 627736
rect 580410 627680 584960 627736
rect 580349 627678 584960 627680
rect 580349 627675 580415 627678
rect 583520 627588 584960 627678
rect 576902 625698 576962 626280
rect 578550 625698 578556 625700
rect 576902 625638 578556 625698
rect 578550 625636 578556 625638
rect 578620 625636 578626 625700
rect -960 624882 480 624972
rect 3417 624882 3483 624885
rect -960 624880 3483 624882
rect -960 624824 3422 624880
rect 3478 624824 3483 624880
rect -960 624822 3483 624824
rect -960 624732 480 624822
rect 3417 624819 3483 624822
rect 583520 615756 584960 615996
rect 5257 614138 5323 614141
rect 7054 614138 7114 614720
rect 5257 614136 7114 614138
rect 5257 614080 5262 614136
rect 5318 614080 7114 614136
rect 5257 614078 7114 614080
rect 5257 614075 5323 614078
rect -960 610316 480 610556
rect 583520 604060 584960 604300
rect 576902 601762 576962 601936
rect 578233 601762 578299 601765
rect 576902 601760 578299 601762
rect 576902 601704 578238 601760
rect 578294 601704 578299 601760
rect 576902 601702 578299 601704
rect 578233 601699 578299 601702
rect -960 595900 480 596140
rect 5165 593602 5231 593605
rect 7054 593602 7114 594184
rect 5165 593600 7114 593602
rect 5165 593544 5170 593600
rect 5226 593544 7114 593600
rect 5165 593542 7114 593544
rect 5165 593539 5231 593542
rect 583520 592364 584960 592604
rect -960 581620 480 581860
rect 580441 580818 580507 580821
rect 583520 580818 584960 580908
rect 580441 580816 584960 580818
rect 580441 580760 580446 580816
rect 580502 580760 584960 580816
rect 580441 580758 584960 580760
rect 580441 580755 580507 580758
rect 583520 580668 584960 580758
rect 576902 577282 576962 577728
rect 578325 577282 578391 577285
rect 576902 577280 578391 577282
rect 576902 577224 578330 577280
rect 578386 577224 578391 577280
rect 576902 577222 578391 577224
rect 578325 577219 578391 577222
rect 6821 573338 6887 573341
rect 7054 573338 7114 573512
rect 6821 573336 7114 573338
rect 6821 573280 6826 573336
rect 6882 573280 7114 573336
rect 6821 573278 7114 573280
rect 6821 573275 6887 573278
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 3969 567354 4035 567357
rect -960 567352 4035 567354
rect -960 567296 3974 567352
rect 4030 567296 4035 567352
rect -960 567294 4035 567296
rect -960 567204 480 567294
rect 3969 567291 4035 567294
rect 583520 557140 584960 557380
rect 578417 553482 578483 553485
rect 576902 553480 578483 553482
rect 576902 553424 578422 553480
rect 578478 553424 578483 553480
rect 576902 553422 578483 553424
rect 576902 553384 576962 553422
rect 578417 553419 578483 553422
rect -960 552924 480 553164
rect 6913 552394 6979 552397
rect 7054 552394 7114 552976
rect 6913 552392 7114 552394
rect 6913 552336 6918 552392
rect 6974 552336 7114 552392
rect 6913 552334 7114 552336
rect 6913 552331 6979 552334
rect 583520 545444 584960 545684
rect -960 538508 480 538748
rect 580533 533898 580599 533901
rect 583520 533898 584960 533988
rect 580533 533896 584960 533898
rect 580533 533840 580538 533896
rect 580594 533840 584960 533896
rect 580533 533838 584960 533840
rect 580533 533835 580599 533838
rect 583520 533748 584960 533838
rect 6686 532274 7084 532334
rect 6686 532133 6746 532274
rect 6686 532128 6795 532133
rect 6686 532072 6734 532128
rect 6790 532072 6795 532128
rect 6686 532070 6795 532072
rect 6729 532067 6795 532070
rect 576902 528866 576962 529176
rect 578509 528866 578575 528869
rect 576902 528864 578575 528866
rect 576902 528808 578514 528864
rect 578570 528808 578575 528864
rect 576902 528806 578575 528808
rect 578509 528803 578575 528806
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 5073 511186 5139 511189
rect 7054 511186 7114 511768
rect 5073 511184 7114 511186
rect 5073 511128 5078 511184
rect 5134 511128 7114 511184
rect 5073 511126 7114 511128
rect 5073 511123 5139 511126
rect 583520 510220 584960 510460
rect -960 509962 480 510052
rect 3509 509962 3575 509965
rect -960 509960 3575 509962
rect -960 509904 3514 509960
rect 3570 509904 3575 509960
rect -960 509902 3575 509904
rect -960 509812 480 509902
rect 3509 509899 3575 509902
rect 576902 504250 576962 504832
rect 578601 504250 578667 504253
rect 576902 504248 578667 504250
rect 576902 504192 578606 504248
rect 578662 504192 578667 504248
rect 576902 504190 578667 504192
rect 578601 504187 578667 504190
rect 583520 498524 584960 498764
rect -960 495396 480 495636
rect 4981 490514 5047 490517
rect 7054 490514 7114 491096
rect 4981 490512 7114 490514
rect 4981 490456 4986 490512
rect 5042 490456 7114 490512
rect 4981 490454 7114 490456
rect 4981 490451 5047 490454
rect 579705 486842 579771 486845
rect 583520 486842 584960 486932
rect 579705 486840 584960 486842
rect 579705 486784 579710 486840
rect 579766 486784 584960 486840
rect 579705 486782 584960 486784
rect 579705 486779 579771 486782
rect 583520 486692 584960 486782
rect -960 480980 480 481220
rect 576902 480450 576962 480488
rect 578693 480450 578759 480453
rect 576902 480448 578759 480450
rect 576902 480392 578698 480448
rect 578754 480392 578759 480448
rect 576902 480390 578759 480392
rect 578693 480387 578759 480390
rect 583520 474996 584960 475236
rect 4889 469978 4955 469981
rect 7054 469978 7114 470560
rect 4889 469976 7114 469978
rect 4889 469920 4894 469976
rect 4950 469920 7114 469976
rect 4889 469918 7114 469920
rect 4889 469915 4955 469918
rect -960 466700 480 466940
rect 583520 463300 584960 463540
rect 576902 455698 576962 456280
rect 578785 455698 578851 455701
rect 576902 455696 578851 455698
rect 576902 455640 578790 455696
rect 578846 455640 578851 455696
rect 576902 455638 578851 455640
rect 578785 455635 578851 455638
rect -960 452434 480 452524
rect 3509 452434 3575 452437
rect -960 452432 3575 452434
rect -960 452376 3514 452432
rect 3570 452376 3575 452432
rect -960 452374 3575 452376
rect -960 452284 480 452374
rect 3509 452371 3575 452374
rect 583520 451604 584960 451844
rect 4797 449986 4863 449989
rect 4797 449984 7114 449986
rect 4797 449928 4802 449984
rect 4858 449928 7114 449984
rect 4797 449926 7114 449928
rect 4797 449923 4863 449926
rect 7054 449888 7114 449926
rect 580625 439922 580691 439925
rect 583520 439922 584960 440012
rect 580625 439920 584960 439922
rect 580625 439864 580630 439920
rect 580686 439864 584960 439920
rect 580625 439862 584960 439864
rect 580625 439859 580691 439862
rect 583520 439772 584960 439862
rect -960 437868 480 438108
rect 576902 431354 576962 431936
rect 578877 431354 578943 431357
rect 576902 431352 578943 431354
rect 576902 431296 578882 431352
rect 578938 431296 578943 431352
rect 576902 431294 578943 431296
rect 578877 431291 578943 431294
rect 4705 429314 4771 429317
rect 7054 429314 7114 429352
rect 4705 429312 7114 429314
rect 4705 429256 4710 429312
rect 4766 429256 7114 429312
rect 4705 429254 7114 429256
rect 4705 429251 4771 429254
rect 583520 428076 584960 428316
rect -960 423588 480 423828
rect 583520 416380 584960 416620
rect -960 409172 480 409412
rect 4613 408642 4679 408645
rect 7054 408642 7114 408680
rect 4613 408640 7114 408642
rect 4613 408584 4618 408640
rect 4674 408584 7114 408640
rect 4613 408582 7114 408584
rect 4613 408579 4679 408582
rect 576902 407146 576962 407728
rect 578969 407146 579035 407149
rect 576902 407144 579035 407146
rect 576902 407088 578974 407144
rect 579030 407088 579035 407144
rect 576902 407086 579035 407088
rect 578969 407083 579035 407086
rect 583520 404684 584960 404924
rect -960 395042 480 395132
rect 3601 395042 3667 395045
rect -960 395040 3667 395042
rect -960 394984 3606 395040
rect 3662 394984 3667 395040
rect -960 394982 3667 394984
rect -960 394892 480 394982
rect 3601 394979 3667 394982
rect 580717 393002 580783 393005
rect 583520 393002 584960 393092
rect 580717 393000 584960 393002
rect 580717 392944 580722 393000
rect 580778 392944 584960 393000
rect 580717 392942 584960 392944
rect 580717 392939 580783 392942
rect 583520 392852 584960 392942
rect 4521 387834 4587 387837
rect 7054 387834 7114 388144
rect 4521 387832 7114 387834
rect 4521 387776 4526 387832
rect 4582 387776 7114 387832
rect 4521 387774 7114 387776
rect 4521 387771 4587 387774
rect 576902 382802 576962 383384
rect 579061 382802 579127 382805
rect 576902 382800 579127 382802
rect 576902 382744 579066 382800
rect 579122 382744 579127 382800
rect 576902 382742 579127 382744
rect 579061 382739 579127 382742
rect 583520 381156 584960 381396
rect -960 380476 480 380716
rect 583520 369460 584960 369700
rect 4429 367298 4495 367301
rect 7054 367298 7114 367472
rect 4429 367296 7114 367298
rect 4429 367240 4434 367296
rect 4490 367240 7114 367296
rect 4429 367238 7114 367240
rect 4429 367235 4495 367238
rect -960 366060 480 366300
rect 576902 358866 576962 359176
rect 579153 358866 579219 358869
rect 576902 358864 579219 358866
rect 576902 358808 579158 358864
rect 579214 358808 579219 358864
rect 576902 358806 579219 358808
rect 579153 358803 579219 358806
rect 583520 357764 584960 358004
rect -960 351780 480 352020
rect 4337 346490 4403 346493
rect 7054 346490 7114 346936
rect 4337 346488 7114 346490
rect 4337 346432 4342 346488
rect 4398 346432 7114 346488
rect 4337 346430 7114 346432
rect 4337 346427 4403 346430
rect 580809 346082 580875 346085
rect 583520 346082 584960 346172
rect 580809 346080 584960 346082
rect 580809 346024 580814 346080
rect 580870 346024 584960 346080
rect 580809 346022 584960 346024
rect 580809 346019 580875 346022
rect 583520 345932 584960 346022
rect -960 337514 480 337604
rect 3693 337514 3759 337517
rect -960 337512 3759 337514
rect -960 337456 3698 337512
rect 3754 337456 3759 337512
rect -960 337454 3759 337456
rect -960 337364 480 337454
rect 3693 337451 3759 337454
rect 576902 334250 576962 334832
rect 579245 334250 579311 334253
rect 576902 334248 579311 334250
rect 576902 334192 579250 334248
rect 579306 334192 579311 334248
rect 583520 334236 584960 334476
rect 576902 334190 579311 334192
rect 579245 334187 579311 334190
rect 4245 325818 4311 325821
rect 7054 325818 7114 326264
rect 4245 325816 7114 325818
rect 4245 325760 4250 325816
rect 4306 325760 7114 325816
rect 4245 325758 7114 325760
rect 4245 325755 4311 325758
rect -960 322948 480 323188
rect 583520 322540 584960 322780
rect 583520 310708 584960 310948
rect 576902 309906 576962 310488
rect 579337 309906 579403 309909
rect 576902 309904 579403 309906
rect 576902 309848 579342 309904
rect 579398 309848 579403 309904
rect 576902 309846 579403 309848
rect 579337 309843 579403 309846
rect -960 308668 480 308908
rect 7054 305149 7114 305728
rect 7005 305144 7114 305149
rect 7005 305088 7010 305144
rect 7066 305088 7114 305144
rect 7005 305086 7114 305088
rect 7005 305083 7071 305086
rect 580901 299162 580967 299165
rect 583520 299162 584960 299252
rect 580901 299160 584960 299162
rect 580901 299104 580906 299160
rect 580962 299104 584960 299160
rect 580901 299102 584960 299104
rect 580901 299099 580967 299102
rect 583520 299012 584960 299102
rect -960 294402 480 294492
rect 3785 294402 3851 294405
rect -960 294400 3851 294402
rect -960 294344 3790 294400
rect 3846 294344 3851 294400
rect -960 294342 3851 294344
rect -960 294252 480 294342
rect 3785 294339 3851 294342
rect 583520 287316 584960 287556
rect 576902 285698 576962 286280
rect 579429 285698 579495 285701
rect 576902 285696 579495 285698
rect 576902 285640 579434 285696
rect 579490 285640 579495 285696
rect 576902 285638 579495 285640
rect 579429 285635 579495 285638
rect 6637 284882 6703 284885
rect 7054 284882 7114 285056
rect 6637 284880 7114 284882
rect 6637 284824 6642 284880
rect 6698 284824 7114 284880
rect 6637 284822 7114 284824
rect 6637 284819 6703 284822
rect -960 279972 480 280212
rect 583520 275620 584960 275860
rect -960 265556 480 265796
rect 7054 263941 7114 264520
rect 7054 263936 7163 263941
rect 7054 263880 7102 263936
rect 7158 263880 7163 263936
rect 7054 263878 7163 263880
rect 7097 263875 7163 263878
rect 583520 263788 584960 264028
rect 576902 261354 576962 261936
rect 579521 261354 579587 261357
rect 576902 261352 579587 261354
rect 576902 261296 579526 261352
rect 579582 261296 579587 261352
rect 576902 261294 579587 261296
rect 579521 261291 579587 261294
rect 580165 252242 580231 252245
rect 583520 252242 584960 252332
rect 580165 252240 584960 252242
rect 580165 252184 580170 252240
rect 580226 252184 584960 252240
rect 580165 252182 584960 252184
rect 580165 252179 580231 252182
rect 583520 252092 584960 252182
rect -960 251290 480 251380
rect 3969 251290 4035 251293
rect -960 251288 4035 251290
rect -960 251232 3974 251288
rect 4030 251232 4035 251288
rect -960 251230 4035 251232
rect -960 251140 480 251230
rect 3969 251227 4035 251230
rect 6545 243674 6611 243677
rect 7054 243674 7114 243848
rect 6545 243672 7114 243674
rect 6545 243616 6550 243672
rect 6606 243616 7114 243672
rect 6545 243614 7114 243616
rect 6545 243611 6611 243614
rect 583520 240396 584960 240636
rect 578141 238234 578207 238237
rect 576902 238232 578207 238234
rect 576902 238176 578146 238232
rect 578202 238176 578207 238232
rect 576902 238174 578207 238176
rect 576902 237728 576962 238174
rect 578141 238171 578207 238174
rect -960 236860 480 237100
rect 583520 228700 584960 228940
rect 7238 222733 7298 223312
rect 7189 222728 7298 222733
rect -960 222444 480 222684
rect 7189 222672 7194 222728
rect 7250 222672 7298 222728
rect 7189 222670 7298 222672
rect 7189 222667 7255 222670
rect 583520 216868 584960 217108
rect 578141 213890 578207 213893
rect 576902 213888 578207 213890
rect 576902 213832 578146 213888
rect 578202 213832 578207 213888
rect 576902 213830 578207 213832
rect 576902 213384 576962 213830
rect 578141 213827 578207 213830
rect -960 208178 480 208268
rect 3233 208178 3299 208181
rect -960 208176 3299 208178
rect -960 208120 3238 208176
rect 3294 208120 3299 208176
rect -960 208118 3299 208120
rect -960 208028 480 208118
rect 3233 208115 3299 208118
rect 580625 205322 580691 205325
rect 583520 205322 584960 205412
rect 580625 205320 584960 205322
rect 580625 205264 580630 205320
rect 580686 205264 584960 205320
rect 580625 205262 584960 205264
rect 580625 205259 580691 205262
rect 583520 205172 584960 205262
rect 3877 202058 3943 202061
rect 7054 202058 7114 202640
rect 3877 202056 7114 202058
rect 3877 202000 3882 202056
rect 3938 202000 7114 202056
rect 3877 201998 7114 202000
rect 3877 201995 3943 201998
rect -960 193748 480 193988
rect 583520 193476 584960 193716
rect 578141 189818 578207 189821
rect 576902 189816 578207 189818
rect 576902 189760 578146 189816
rect 578202 189760 578207 189816
rect 576902 189758 578207 189760
rect 576902 189176 576962 189758
rect 578141 189755 578207 189758
rect 4153 181522 4219 181525
rect 7054 181522 7114 182104
rect 583520 181780 584960 182020
rect 4153 181520 7114 181522
rect 4153 181464 4158 181520
rect 4214 181464 7114 181520
rect 4153 181462 7114 181464
rect 4153 181459 4219 181462
rect -960 179332 480 179572
rect 583520 169948 584960 170188
rect 578141 165474 578207 165477
rect 576902 165472 578207 165474
rect 576902 165416 578146 165472
rect 578202 165416 578207 165472
rect 576902 165414 578207 165416
rect -960 165066 480 165156
rect 3141 165066 3207 165069
rect -960 165064 3207 165066
rect -960 165008 3146 165064
rect 3202 165008 3207 165064
rect -960 165006 3207 165008
rect -960 164916 480 165006
rect 3141 165003 3207 165006
rect 576902 164832 576962 165414
rect 578141 165411 578207 165414
rect 4153 160850 4219 160853
rect 7054 160850 7114 161432
rect 4153 160848 7114 160850
rect 4153 160792 4158 160848
rect 4214 160792 7114 160848
rect 4153 160790 7114 160792
rect 4153 160787 4219 160790
rect 580717 158402 580783 158405
rect 583520 158402 584960 158492
rect 580717 158400 584960 158402
rect 580717 158344 580722 158400
rect 580778 158344 584960 158400
rect 580717 158342 584960 158344
rect 580717 158339 580783 158342
rect 583520 158252 584960 158342
rect -960 150636 480 150876
rect 583520 146556 584960 146796
rect 3141 141538 3207 141541
rect 3141 141536 7114 141538
rect 3141 141480 3146 141536
rect 3202 141480 7114 141536
rect 3141 141478 7114 141480
rect 3141 141475 3207 141478
rect 7054 140896 7114 141478
rect 580165 140722 580231 140725
rect 576902 140720 580231 140722
rect 576902 140664 580170 140720
rect 580226 140664 580231 140720
rect 576902 140662 580231 140664
rect 576902 140488 576962 140662
rect 580165 140659 580231 140662
rect -960 136220 480 136460
rect 583520 134724 584960 134964
rect 583520 123028 584960 123268
rect -960 122090 480 122180
rect 4153 122090 4219 122093
rect -960 122088 4219 122090
rect -960 122032 4158 122088
rect 4214 122032 4219 122088
rect -960 122030 4219 122032
rect -960 121940 480 122030
rect 4153 122027 4219 122030
rect 4153 120866 4219 120869
rect 4153 120864 7114 120866
rect 4153 120808 4158 120864
rect 4214 120808 7114 120864
rect 4153 120806 7114 120808
rect 4153 120803 4219 120806
rect 7054 120224 7114 120806
rect 578141 116922 578207 116925
rect 576902 116920 578207 116922
rect 576902 116864 578146 116920
rect 578202 116864 578207 116920
rect 576902 116862 578207 116864
rect 576902 116280 576962 116862
rect 578141 116859 578207 116862
rect 580625 111482 580691 111485
rect 583520 111482 584960 111572
rect 580625 111480 584960 111482
rect 580625 111424 580630 111480
rect 580686 111424 584960 111480
rect 580625 111422 584960 111424
rect 580625 111419 580691 111422
rect 583520 111332 584960 111422
rect -960 107524 480 107764
rect 3969 100330 4035 100333
rect 3969 100328 7114 100330
rect 3969 100272 3974 100328
rect 4030 100272 7114 100328
rect 3969 100270 7114 100272
rect 3969 100267 4035 100270
rect 7054 99688 7114 100270
rect 583520 99636 584960 99876
rect -960 93108 480 93348
rect 578141 92442 578207 92445
rect 576902 92440 578207 92442
rect 576902 92384 578146 92440
rect 578202 92384 578207 92440
rect 576902 92382 578207 92384
rect 576902 91936 576962 92382
rect 578141 92379 578207 92382
rect 583520 87804 584960 88044
rect 3785 79658 3851 79661
rect 3785 79656 7114 79658
rect 3785 79600 3790 79656
rect 3846 79600 7114 79656
rect 3785 79598 7114 79600
rect 3785 79595 3851 79598
rect -960 78978 480 79068
rect 7054 79016 7114 79598
rect 3325 78978 3391 78981
rect -960 78976 3391 78978
rect -960 78920 3330 78976
rect 3386 78920 3391 78976
rect -960 78918 3391 78920
rect -960 78828 480 78918
rect 3325 78915 3391 78918
rect 583520 76108 584960 76348
rect 578141 68370 578207 68373
rect 576902 68368 578207 68370
rect 576902 68312 578146 68368
rect 578202 68312 578207 68368
rect 576902 68310 578207 68312
rect 576902 67728 576962 68310
rect 578141 68307 578207 68310
rect -960 64412 480 64652
rect 580625 64562 580691 64565
rect 583520 64562 584960 64652
rect 580625 64560 584960 64562
rect 580625 64504 580630 64560
rect 580686 64504 584960 64560
rect 580625 64502 584960 64504
rect 580625 64499 580691 64502
rect 583520 64412 584960 64502
rect 3693 59122 3759 59125
rect 3693 59120 7114 59122
rect 3693 59064 3698 59120
rect 3754 59064 7114 59120
rect 3693 59062 7114 59064
rect 3693 59059 3759 59062
rect 7054 58480 7114 59062
rect 583520 52716 584960 52956
rect -960 49996 480 50236
rect 578141 44026 578207 44029
rect 576902 44024 578207 44026
rect 576902 43968 578146 44024
rect 578202 43968 578207 44024
rect 576902 43966 578207 43968
rect 576902 43384 576962 43966
rect 578141 43963 578207 43966
rect 583520 40884 584960 41124
rect 3601 38314 3667 38317
rect 3601 38312 7114 38314
rect 3601 38256 3606 38312
rect 3662 38256 7114 38312
rect 3601 38254 7114 38256
rect 3601 38251 3667 38254
rect 7054 37808 7114 38254
rect -960 35866 480 35956
rect 3877 35866 3943 35869
rect -960 35864 3943 35866
rect -960 35808 3882 35864
rect 3938 35808 3943 35864
rect -960 35806 3943 35808
rect -960 35716 480 35806
rect 3877 35803 3943 35806
rect 583520 29188 584960 29428
rect -960 21300 480 21540
rect 576902 18594 576962 19176
rect 579613 18594 579679 18597
rect 576902 18592 579679 18594
rect 576902 18536 579618 18592
rect 579674 18536 579679 18592
rect 576902 18534 579679 18536
rect 579613 18531 579679 18534
rect 3509 17914 3575 17917
rect 3509 17912 7114 17914
rect 3509 17856 3514 17912
rect 3570 17856 7114 17912
rect 3509 17854 7114 17856
rect 3509 17851 3575 17854
rect 7054 17272 7114 17854
rect 579613 17642 579679 17645
rect 583520 17642 584960 17732
rect 579613 17640 584960 17642
rect 579613 17584 579618 17640
rect 579674 17584 584960 17640
rect 579613 17582 584960 17584
rect 579613 17579 579679 17582
rect 583520 17492 584960 17582
rect 109953 7714 110019 7717
rect 570270 7714 570276 7716
rect 109953 7712 570276 7714
rect 109953 7656 109958 7712
rect 110014 7656 570276 7712
rect 109953 7654 570276 7656
rect 109953 7651 110019 7654
rect 570270 7652 570276 7654
rect 570340 7652 570346 7716
rect 106365 7578 106431 7581
rect 570086 7578 570092 7580
rect 106365 7576 570092 7578
rect 106365 7520 106370 7576
rect 106426 7520 570092 7576
rect 106365 7518 570092 7520
rect 106365 7515 106431 7518
rect 570086 7516 570092 7518
rect 570156 7516 570162 7580
rect -960 7020 480 7260
rect 583520 5796 584960 6036
rect 12433 5538 12499 5541
rect 439589 5538 439655 5541
rect 12433 5536 439655 5538
rect 12433 5480 12438 5536
rect 12494 5480 439594 5536
rect 439650 5480 439655 5536
rect 12433 5478 439655 5480
rect 12433 5475 12499 5478
rect 439589 5475 439655 5478
rect 2865 5402 2931 5405
rect 429377 5402 429443 5405
rect 2865 5400 429443 5402
rect 2865 5344 2870 5400
rect 2926 5344 429382 5400
rect 429438 5344 429443 5400
rect 2865 5342 429443 5344
rect 2865 5339 2931 5342
rect 429377 5339 429443 5342
rect 114553 5266 114619 5269
rect 561673 5266 561739 5269
rect 114553 5264 561739 5266
rect 114553 5208 114558 5264
rect 114614 5208 561678 5264
rect 561734 5208 561739 5264
rect 114553 5206 561739 5208
rect 114553 5203 114619 5206
rect 561673 5203 561739 5206
rect 34973 5130 35039 5133
rect 521009 5130 521075 5133
rect 34973 5128 521075 5130
rect 34973 5072 34978 5128
rect 35034 5072 521014 5128
rect 521070 5072 521075 5128
rect 34973 5070 521075 5072
rect 34973 5067 35039 5070
rect 521009 5067 521075 5070
rect 38561 4994 38627 4997
rect 531129 4994 531195 4997
rect 38561 4992 531195 4994
rect 38561 4936 38566 4992
rect 38622 4936 531134 4992
rect 531190 4936 531195 4992
rect 38561 4934 531195 4936
rect 38561 4931 38627 4934
rect 531129 4931 531195 4934
rect 6453 4858 6519 4861
rect 571885 4858 571951 4861
rect 6453 4856 571951 4858
rect 6453 4800 6458 4856
rect 6514 4800 571890 4856
rect 571946 4800 571951 4856
rect 6453 4798 571951 4800
rect 6453 4795 6519 4798
rect 571885 4795 571951 4798
rect 9397 4042 9463 4045
rect 67173 4042 67239 4045
rect 9397 4040 67239 4042
rect 9397 3984 9402 4040
rect 9458 3984 67178 4040
rect 67234 3984 67239 4040
rect 9397 3982 67239 3984
rect 9397 3979 9463 3982
rect 67173 3979 67239 3982
rect 95693 4042 95759 4045
rect 578233 4042 578299 4045
rect 95693 4040 578299 4042
rect 95693 3984 95698 4040
rect 95754 3984 578238 4040
rect 578294 3984 578299 4040
rect 95693 3982 578299 3984
rect 95693 3979 95759 3982
rect 578233 3979 578299 3982
rect 9489 3906 9555 3909
rect 74257 3906 74323 3909
rect 9489 3904 74323 3906
rect 9489 3848 9494 3904
rect 9550 3848 74262 3904
rect 74318 3848 74323 3904
rect 9489 3846 74323 3848
rect 9489 3843 9555 3846
rect 74257 3843 74323 3846
rect 77845 3906 77911 3909
rect 569902 3906 569908 3908
rect 77845 3904 569908 3906
rect 77845 3848 77850 3904
rect 77906 3848 569908 3904
rect 77845 3846 569908 3848
rect 77845 3843 77911 3846
rect 569902 3844 569908 3846
rect 569972 3844 569978 3908
rect 42149 3770 42215 3773
rect 578785 3770 578851 3773
rect 42149 3768 578851 3770
rect 42149 3712 42154 3768
rect 42210 3712 578790 3768
rect 578846 3712 578851 3768
rect 42149 3710 578851 3712
rect 42149 3707 42215 3710
rect 578785 3707 578851 3710
rect 9305 3634 9371 3637
rect 23105 3634 23171 3637
rect 9305 3632 23171 3634
rect 9305 3576 9310 3632
rect 9366 3576 23110 3632
rect 23166 3576 23171 3632
rect 9305 3574 23171 3576
rect 9305 3571 9371 3574
rect 23105 3571 23171 3574
rect 25497 3634 25563 3637
rect 571374 3634 571380 3636
rect 25497 3632 571380 3634
rect 25497 3576 25502 3632
rect 25558 3576 571380 3632
rect 25497 3574 571380 3576
rect 25497 3571 25563 3574
rect 571374 3572 571380 3574
rect 571444 3572 571450 3636
rect 8937 3498 9003 3501
rect 18321 3498 18387 3501
rect 8937 3496 18387 3498
rect 8937 3440 8942 3496
rect 8998 3440 18326 3496
rect 18382 3440 18387 3496
rect 8937 3438 18387 3440
rect 8937 3435 9003 3438
rect 18321 3435 18387 3438
rect 20713 3498 20779 3501
rect 578366 3498 578372 3500
rect 20713 3496 578372 3498
rect 20713 3440 20718 3496
rect 20774 3440 578372 3496
rect 20713 3438 578372 3440
rect 20713 3435 20779 3438
rect 578366 3436 578372 3438
rect 578436 3436 578442 3500
rect 5257 3362 5323 3365
rect 578182 3362 578188 3364
rect 5257 3360 578188 3362
rect 5257 3304 5262 3360
rect 5318 3304 578188 3360
rect 5257 3302 578188 3304
rect 5257 3299 5323 3302
rect 578182 3300 578188 3302
rect 578252 3300 578258 3364
rect 99281 3226 99347 3229
rect 578550 3226 578556 3228
rect 99281 3224 578556 3226
rect 99281 3168 99286 3224
rect 99342 3168 578556 3224
rect 99281 3166 578556 3168
rect 99281 3163 99347 3166
rect 578550 3164 578556 3166
rect 578620 3164 578626 3228
rect 5390 3028 5396 3092
rect 5460 3090 5466 3092
rect 124213 3090 124279 3093
rect 5460 3088 124279 3090
rect 5460 3032 124218 3088
rect 124274 3032 124279 3088
rect 5460 3030 124279 3032
rect 5460 3028 5466 3030
rect 124213 3027 124279 3030
<< via3 >>
rect 569908 689012 569972 689076
rect 570276 688876 570340 688940
rect 570092 688740 570156 688804
rect 571380 688604 571444 688668
rect 578188 674868 578252 674932
rect 578372 649980 578436 650044
rect 5396 634884 5460 634948
rect 578556 625636 578620 625700
rect 570276 7652 570340 7716
rect 570092 7516 570156 7580
rect 569908 3844 569972 3908
rect 571380 3572 571444 3636
rect 578372 3436 578436 3500
rect 578188 3300 578252 3364
rect 578556 3164 578620 3228
rect 5396 3028 5460 3092
<< metal4 >>
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 -1286 -2336 705222
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 -346 -1396 704282
rect 23424 704838 24024 705800
rect 23424 704602 23606 704838
rect 23842 704602 24024 704838
rect 23424 704518 24024 704602
rect 23424 704282 23606 704518
rect 23842 704282 24024 704518
rect 5395 634948 5461 634949
rect 5395 634884 5396 634948
rect 5460 634884 5461 634948
rect 5395 634883 5461 634884
rect 5398 3093 5458 634883
rect 5395 3092 5461 3093
rect 5395 3028 5396 3092
rect 5460 3028 5461 3092
rect 5395 3027 5461 3028
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 23424 -346 24024 704282
rect 23424 -582 23606 -346
rect 23842 -582 24024 -346
rect 23424 -666 24024 -582
rect 23424 -902 23606 -666
rect 23842 -902 24024 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 23424 -1864 24024 -902
rect 99424 705778 100024 705800
rect 99424 705542 99606 705778
rect 99842 705542 100024 705778
rect 99424 705458 100024 705542
rect 99424 705222 99606 705458
rect 99842 705222 100024 705458
rect 99424 -1286 100024 705222
rect 99424 -1522 99606 -1286
rect 99842 -1522 100024 -1286
rect 99424 -1606 100024 -1522
rect 99424 -1842 99606 -1606
rect 99842 -1842 100024 -1606
rect 99424 -1864 100024 -1842
rect 175424 704838 176024 705800
rect 175424 704602 175606 704838
rect 175842 704602 176024 704838
rect 175424 704518 176024 704602
rect 175424 704282 175606 704518
rect 175842 704282 176024 704518
rect 175424 -346 176024 704282
rect 175424 -582 175606 -346
rect 175842 -582 176024 -346
rect 175424 -666 176024 -582
rect 175424 -902 175606 -666
rect 175842 -902 176024 -666
rect 175424 -1864 176024 -902
rect 251424 705778 252024 705800
rect 251424 705542 251606 705778
rect 251842 705542 252024 705778
rect 251424 705458 252024 705542
rect 251424 705222 251606 705458
rect 251842 705222 252024 705458
rect 251424 -1286 252024 705222
rect 251424 -1522 251606 -1286
rect 251842 -1522 252024 -1286
rect 251424 -1606 252024 -1522
rect 251424 -1842 251606 -1606
rect 251842 -1842 252024 -1606
rect 251424 -1864 252024 -1842
rect 327424 704838 328024 705800
rect 327424 704602 327606 704838
rect 327842 704602 328024 704838
rect 327424 704518 328024 704602
rect 327424 704282 327606 704518
rect 327842 704282 328024 704518
rect 327424 -346 328024 704282
rect 327424 -582 327606 -346
rect 327842 -582 328024 -346
rect 327424 -666 328024 -582
rect 327424 -902 327606 -666
rect 327842 -902 328024 -666
rect 327424 -1864 328024 -902
rect 403424 705778 404024 705800
rect 403424 705542 403606 705778
rect 403842 705542 404024 705778
rect 403424 705458 404024 705542
rect 403424 705222 403606 705458
rect 403842 705222 404024 705458
rect 403424 -1286 404024 705222
rect 403424 -1522 403606 -1286
rect 403842 -1522 404024 -1286
rect 403424 -1606 404024 -1522
rect 403424 -1842 403606 -1606
rect 403842 -1842 404024 -1606
rect 403424 -1864 404024 -1842
rect 479424 704838 480024 705800
rect 479424 704602 479606 704838
rect 479842 704602 480024 704838
rect 479424 704518 480024 704602
rect 479424 704282 479606 704518
rect 479842 704282 480024 704518
rect 479424 -346 480024 704282
rect 479424 -582 479606 -346
rect 479842 -582 480024 -346
rect 479424 -666 480024 -582
rect 479424 -902 479606 -666
rect 479842 -902 480024 -666
rect 479424 -1864 480024 -902
rect 555424 705778 556024 705800
rect 555424 705542 555606 705778
rect 555842 705542 556024 705778
rect 555424 705458 556024 705542
rect 555424 705222 555606 705458
rect 555842 705222 556024 705458
rect 555424 -1286 556024 705222
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 569907 689076 569973 689077
rect 569907 689012 569908 689076
rect 569972 689012 569973 689076
rect 569907 689011 569973 689012
rect 569910 3909 569970 689011
rect 570275 688940 570341 688941
rect 570275 688876 570276 688940
rect 570340 688876 570341 688940
rect 570275 688875 570341 688876
rect 570091 688804 570157 688805
rect 570091 688740 570092 688804
rect 570156 688740 570157 688804
rect 570091 688739 570157 688740
rect 570094 7581 570154 688739
rect 570278 7717 570338 688875
rect 571379 688668 571445 688669
rect 571379 688604 571380 688668
rect 571444 688604 571445 688668
rect 571379 688603 571445 688604
rect 570275 7716 570341 7717
rect 570275 7652 570276 7716
rect 570340 7652 570341 7716
rect 570275 7651 570341 7652
rect 570091 7580 570157 7581
rect 570091 7516 570092 7580
rect 570156 7516 570157 7580
rect 570091 7515 570157 7516
rect 569907 3908 569973 3909
rect 569907 3844 569908 3908
rect 569972 3844 569973 3908
rect 569907 3843 569973 3844
rect 571382 3637 571442 688603
rect 578187 674932 578253 674933
rect 578187 674868 578188 674932
rect 578252 674868 578253 674932
rect 578187 674867 578253 674868
rect 571379 3636 571445 3637
rect 571379 3572 571380 3636
rect 571444 3572 571445 3636
rect 571379 3571 571445 3572
rect 578190 3365 578250 674867
rect 578371 650044 578437 650045
rect 578371 649980 578372 650044
rect 578436 649980 578437 650044
rect 578371 649979 578437 649980
rect 578374 3501 578434 649979
rect 578555 625700 578621 625701
rect 578555 625636 578556 625700
rect 578620 625636 578621 625700
rect 578555 625635 578621 625636
rect 578371 3500 578437 3501
rect 578371 3436 578372 3500
rect 578436 3436 578437 3500
rect 578371 3435 578437 3436
rect 578187 3364 578253 3365
rect 578187 3300 578188 3364
rect 578252 3300 578253 3364
rect 578187 3299 578253 3300
rect 578558 3229 578618 625635
rect 578555 3228 578621 3229
rect 578555 3164 578556 3228
rect 578620 3164 578621 3228
rect 578555 3163 578621 3164
rect 585320 -346 585920 704282
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 555424 -1522 555606 -1286
rect 555842 -1522 556024 -1286
rect 555424 -1606 556024 -1522
rect 555424 -1842 555606 -1606
rect 555842 -1842 556024 -1606
rect 555424 -1864 556024 -1842
rect 586260 -1286 586860 705222
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
<< via4 >>
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect 23606 704602 23842 704838
rect 23606 704282 23842 704518
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 23606 -582 23842 -346
rect 23606 -902 23842 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 99606 705542 99842 705778
rect 99606 705222 99842 705458
rect 99606 -1522 99842 -1286
rect 99606 -1842 99842 -1606
rect 175606 704602 175842 704838
rect 175606 704282 175842 704518
rect 175606 -582 175842 -346
rect 175606 -902 175842 -666
rect 251606 705542 251842 705778
rect 251606 705222 251842 705458
rect 251606 -1522 251842 -1286
rect 251606 -1842 251842 -1606
rect 327606 704602 327842 704838
rect 327606 704282 327842 704518
rect 327606 -582 327842 -346
rect 327606 -902 327842 -666
rect 403606 705542 403842 705778
rect 403606 705222 403842 705458
rect 403606 -1522 403842 -1286
rect 403606 -1842 403842 -1606
rect 479606 704602 479842 704838
rect 479606 704282 479842 704518
rect 479606 -582 479842 -346
rect 479606 -902 479842 -666
rect 555606 705542 555842 705778
rect 555606 705222 555842 705458
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 555606 -1522 555842 -1286
rect 555606 -1842 555842 -1606
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
<< metal5 >>
rect -2936 705800 -2336 705802
rect 99424 705800 100024 705802
rect 251424 705800 252024 705802
rect 403424 705800 404024 705802
rect 555424 705800 556024 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 99606 705778
rect 99842 705542 251606 705778
rect 251842 705542 403606 705778
rect 403842 705542 555606 705778
rect 555842 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 99606 705458
rect 99842 705222 251606 705458
rect 251842 705222 403606 705458
rect 403842 705222 555606 705458
rect 555842 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 99424 705198 100024 705200
rect 251424 705198 252024 705200
rect 403424 705198 404024 705200
rect 555424 705198 556024 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 23424 704860 24024 704862
rect 175424 704860 176024 704862
rect 327424 704860 328024 704862
rect 479424 704860 480024 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 23606 704838
rect 23842 704602 175606 704838
rect 175842 704602 327606 704838
rect 327842 704602 479606 704838
rect 479842 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 23606 704518
rect 23842 704282 175606 704518
rect 175842 704282 327606 704518
rect 327842 704282 479606 704518
rect 479842 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 23424 704258 24024 704260
rect 175424 704258 176024 704260
rect 327424 704258 328024 704260
rect 479424 704258 480024 704260
rect 585320 704258 585920 704260
rect -1996 -324 -1396 -322
rect 23424 -324 24024 -322
rect 175424 -324 176024 -322
rect 327424 -324 328024 -322
rect 479424 -324 480024 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 23606 -346
rect 23842 -582 175606 -346
rect 175842 -582 327606 -346
rect 327842 -582 479606 -346
rect 479842 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 23606 -666
rect 23842 -902 175606 -666
rect 175842 -902 327606 -666
rect 327842 -902 479606 -666
rect 479842 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 23424 -926 24024 -924
rect 175424 -926 176024 -924
rect 327424 -926 328024 -924
rect 479424 -926 480024 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 99424 -1264 100024 -1262
rect 251424 -1264 252024 -1262
rect 403424 -1264 404024 -1262
rect 555424 -1264 556024 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 99606 -1286
rect 99842 -1522 251606 -1286
rect 251842 -1522 403606 -1286
rect 403842 -1522 555606 -1286
rect 555842 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 99606 -1606
rect 99842 -1842 251606 -1606
rect 251842 -1842 403606 -1606
rect 403842 -1842 555606 -1606
rect 555842 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 99424 -1866 100024 -1864
rect 251424 -1866 252024 -1864
rect 403424 -1866 404024 -1864
rect 555424 -1866 556024 -1864
rect 586260 -1866 586860 -1864
use fpga  fpga250
timestamp 1608149048
transform 1 0 7000 0 1 7000
box 0 0 570000 680000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 637 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1608157735
<< locali >>
rect 27077 16439 27111 16541
rect 50813 16439 50847 16745
rect 19993 16031 20027 16201
rect 39773 16031 39807 16133
rect 34897 15895 34931 15997
rect 21649 15487 21683 15589
rect 23489 15555 23523 15657
rect 29745 15555 29779 15657
rect 25881 15419 25915 15521
rect 38301 15351 38335 15453
rect 25605 14943 25639 15045
rect 19349 14807 19383 14909
rect 30573 14807 30607 14909
rect 31125 14875 31159 15045
rect 34069 14943 34103 15113
rect 46489 14807 46523 14909
rect 51549 14875 51583 15113
rect 6653 14263 6687 14433
rect 10701 14263 10735 14569
rect 6837 13855 6871 14025
rect 12081 13923 12115 14025
rect 25973 13787 26007 13889
rect 31033 13787 31067 13957
rect 43269 13787 43303 14025
rect 49801 13719 49835 13957
rect 50905 13855 50939 14025
rect 7573 13379 7607 13481
rect 7665 13175 7699 13277
rect 15669 13175 15703 13481
rect 21281 13175 21315 13277
rect 39037 13175 39071 13413
rect 42257 13311 42291 13413
rect 43085 13175 43119 13345
rect 44005 13243 44039 13345
rect 47869 13175 47903 13481
rect 48513 13379 48547 13481
rect 3157 12631 3191 12937
rect 27813 12767 27847 12869
rect 4445 12631 4479 12733
rect 29745 12631 29779 12869
rect 50905 12631 50939 12801
rect 54401 12631 54435 12733
rect 17693 12291 17727 12393
rect 22017 12087 22051 12325
rect 27997 12087 28031 12393
rect 31711 12325 31803 12359
rect 31769 12291 31803 12325
rect 41613 12087 41647 12393
rect 46305 12087 46339 12325
rect 11989 11543 12023 11713
rect 15393 11679 15427 11781
rect 42441 11679 42475 11849
rect 21833 11067 21867 11305
rect 22109 11135 22143 11305
rect 53021 11203 53055 11305
rect 34529 10455 34563 10557
rect 40601 10455 40635 10625
rect 8033 10115 8067 10217
rect 24777 9911 24811 10013
rect 22051 9605 22143 9639
rect 15393 9503 15427 9605
rect 22109 9571 22143 9605
rect 16221 9367 16255 9469
rect 34989 9367 35023 9469
rect 42349 9367 42383 9605
rect 7849 8959 7883 9129
rect 49341 8823 49375 8993
rect 7941 8347 7975 8449
rect 8033 8415 8067 8517
rect 18061 8415 18095 8517
rect 21373 8279 21407 8381
rect 24133 8347 24167 8517
rect 29929 8279 29963 8517
rect 34529 8279 34563 8381
rect 37841 8279 37875 8381
rect 40141 8347 40175 8517
rect 42717 8483 42751 8585
rect 51365 8415 51399 8517
rect 52929 8415 52963 8517
rect 10517 7735 10551 7905
rect 24777 7735 24811 8041
rect 36369 7803 36403 7905
rect 48053 7735 48087 8041
rect 12909 7259 12943 7497
rect 25053 7191 25087 7497
rect 28457 7259 28491 7497
rect 50629 7327 50663 7497
rect 17601 6647 17635 6953
rect 46397 6647 46431 6953
rect 51549 6783 51583 6953
rect 11713 6103 11747 6409
rect 19165 6239 19199 6341
rect 34437 6307 34471 6409
rect 27445 6103 27479 6205
rect 39589 6171 39623 6341
rect 45017 6307 45051 6409
rect 47041 6171 47075 6341
rect 47501 6239 47535 6341
rect 50997 6307 51031 6409
rect 55229 6103 55263 6341
rect 18521 5559 18555 5661
rect 18981 5559 19015 5797
rect 31309 5627 31343 5865
rect 42809 5627 42843 5797
rect 18889 5219 18923 5321
rect 24041 5015 24075 5321
rect 24501 5015 24535 5185
rect 31217 5015 31251 5253
rect 34437 5151 34471 5321
rect 32965 5015 32999 5117
rect 35449 5015 35483 5253
rect 39405 5015 39439 5321
rect 41429 5219 41463 5321
rect 7665 4675 7699 4777
rect 19625 4471 19659 4777
rect 22385 4471 22419 4641
rect 31585 4607 31619 4709
rect 38853 4471 38887 4777
rect 38945 4607 38979 4777
rect 28825 3995 28859 4165
rect 32413 3927 32447 4233
rect 47317 4131 47351 4233
rect 49157 4063 49191 4165
rect 50905 3927 50939 4029
rect 57897 3587 57931 3689
rect 35357 3383 35391 3485
rect 47501 3383 47535 3553
rect 10241 2975 10275 3145
rect 11621 2907 11655 3145
rect 21465 2975 21499 3145
rect 25605 2839 25639 3077
rect 35633 3043 35667 3145
rect 42717 3043 42751 3145
rect 30297 2839 30331 2941
rect 34069 2839 34103 3009
rect 10701 2499 10735 2601
rect 12173 2295 12207 2601
rect 14749 2431 14783 2601
rect 14657 2295 14691 2397
rect 50905 2295 50939 2465
rect 9597 1955 9631 2057
<< viali >>
rect 14381 17289 14415 17323
rect 23489 17289 23523 17323
rect 28549 17289 28583 17323
rect 42533 17289 42567 17323
rect 48421 17289 48455 17323
rect 53941 17289 53975 17323
rect 20453 17221 20487 17255
rect 33793 17221 33827 17255
rect 49985 17221 50019 17255
rect 12449 17153 12483 17187
rect 12817 17153 12851 17187
rect 19257 17153 19291 17187
rect 26709 17153 26743 17187
rect 29745 17153 29779 17187
rect 31033 17153 31067 17187
rect 34805 17153 34839 17187
rect 40325 17153 40359 17187
rect 40969 17153 41003 17187
rect 46673 17153 46707 17187
rect 50997 17153 51031 17187
rect 13093 17085 13127 17119
rect 18797 17085 18831 17119
rect 19165 17085 19199 17119
rect 22569 17085 22603 17119
rect 22753 17085 22787 17119
rect 22937 17085 22971 17119
rect 23765 17085 23799 17119
rect 27169 17085 27203 17119
rect 27445 17085 27479 17119
rect 30205 17085 30239 17119
rect 30573 17085 30607 17119
rect 30665 17085 30699 17119
rect 33977 17085 34011 17119
rect 34161 17085 34195 17119
rect 34345 17085 34379 17119
rect 35173 17085 35207 17119
rect 39497 17085 39531 17119
rect 39681 17085 39715 17119
rect 39865 17085 39899 17119
rect 41153 17085 41187 17119
rect 41429 17085 41463 17119
rect 46857 17085 46891 17119
rect 47133 17085 47167 17119
rect 50169 17085 50203 17119
rect 50353 17085 50387 17119
rect 50537 17085 50571 17119
rect 53113 17085 53147 17119
rect 53481 17085 53515 17119
rect 53573 17085 53607 17119
rect 18337 17017 18371 17051
rect 19625 17017 19659 17051
rect 22109 17017 22143 17051
rect 31401 17017 31435 17051
rect 39037 17017 39071 17051
rect 52653 17017 52687 17051
rect 20085 16949 20119 16983
rect 20729 16949 20763 16983
rect 21373 16949 21407 16983
rect 21741 16949 21775 16983
rect 29377 16949 29411 16983
rect 38945 16949 38979 16983
rect 43085 16949 43119 16983
rect 51457 16949 51491 16983
rect 54309 16949 54343 16983
rect 12633 16745 12667 16779
rect 17141 16745 17175 16779
rect 19625 16745 19659 16779
rect 22477 16745 22511 16779
rect 24961 16745 24995 16779
rect 36001 16745 36035 16779
rect 41613 16745 41647 16779
rect 48789 16745 48823 16779
rect 50353 16745 50387 16779
rect 50813 16745 50847 16779
rect 54125 16745 54159 16779
rect 8217 16609 8251 16643
rect 8401 16609 8435 16643
rect 8585 16609 8619 16643
rect 11069 16609 11103 16643
rect 13185 16609 13219 16643
rect 18061 16609 18095 16643
rect 18245 16609 18279 16643
rect 21373 16609 21407 16643
rect 23581 16609 23615 16643
rect 30297 16609 30331 16643
rect 30665 16609 30699 16643
rect 34069 16609 34103 16643
rect 34437 16609 34471 16643
rect 47501 16609 47535 16643
rect 47685 16609 47719 16643
rect 47869 16609 47903 16643
rect 48973 16609 49007 16643
rect 11345 16541 11379 16575
rect 15761 16541 15795 16575
rect 16037 16541 16071 16575
rect 18521 16541 18555 16575
rect 21097 16541 21131 16575
rect 23857 16541 23891 16575
rect 27077 16541 27111 16575
rect 27353 16541 27387 16575
rect 27629 16541 27663 16575
rect 30757 16541 30791 16575
rect 32137 16541 32171 16575
rect 32413 16541 32447 16575
rect 34621 16541 34655 16575
rect 34897 16541 34931 16575
rect 37749 16541 37783 16575
rect 38025 16541 38059 16575
rect 39129 16541 39163 16575
rect 40233 16541 40267 16575
rect 40509 16541 40543 16575
rect 49249 16541 49283 16575
rect 8033 16473 8067 16507
rect 30113 16473 30147 16507
rect 42533 16473 42567 16507
rect 42901 16473 42935 16507
rect 47317 16473 47351 16507
rect 54769 16609 54803 16643
rect 51825 16541 51859 16575
rect 52101 16541 52135 16575
rect 9045 16405 9079 16439
rect 9505 16405 9539 16439
rect 10885 16405 10919 16439
rect 14289 16405 14323 16439
rect 20361 16405 20395 16439
rect 23121 16405 23155 16439
rect 27077 16405 27111 16439
rect 27169 16405 27203 16439
rect 28733 16405 28767 16439
rect 29561 16405 29595 16439
rect 31125 16405 31159 16439
rect 33517 16405 33551 16439
rect 37381 16405 37415 16439
rect 39957 16405 39991 16439
rect 42165 16405 42199 16439
rect 46581 16405 46615 16439
rect 46949 16405 46983 16439
rect 48329 16405 48363 16439
rect 50813 16405 50847 16439
rect 50905 16405 50939 16439
rect 53205 16405 53239 16439
rect 53757 16405 53791 16439
rect 8217 16201 8251 16235
rect 9873 16201 9907 16235
rect 11253 16201 11287 16235
rect 11805 16201 11839 16235
rect 12265 16201 12299 16235
rect 14657 16201 14691 16235
rect 16129 16201 16163 16235
rect 16773 16201 16807 16235
rect 19993 16201 20027 16235
rect 21465 16201 21499 16235
rect 49709 16201 49743 16235
rect 52193 16201 52227 16235
rect 52745 16201 52779 16235
rect 54677 16201 54711 16235
rect 8585 16065 8619 16099
rect 10333 16065 10367 16099
rect 16313 16065 16347 16099
rect 17785 16065 17819 16099
rect 19349 16065 19383 16099
rect 22477 16133 22511 16167
rect 25421 16133 25455 16167
rect 27537 16133 27571 16167
rect 30665 16133 30699 16167
rect 33701 16133 33735 16167
rect 39773 16133 39807 16167
rect 39957 16133 39991 16167
rect 43453 16133 43487 16167
rect 46397 16133 46431 16167
rect 47225 16133 47259 16167
rect 49985 16133 50019 16167
rect 23121 16065 23155 16099
rect 24409 16065 24443 16099
rect 24685 16065 24719 16099
rect 25053 16065 25087 16099
rect 26709 16065 26743 16099
rect 28365 16065 28399 16099
rect 33333 16065 33367 16099
rect 41889 16065 41923 16099
rect 47593 16065 47627 16099
rect 53573 16065 53607 16099
rect 8309 15997 8343 16031
rect 10885 15997 10919 16031
rect 11069 15997 11103 16031
rect 13829 15997 13863 16031
rect 14197 15997 14231 16031
rect 14289 15997 14323 16031
rect 16589 15997 16623 16031
rect 18521 15997 18555 16031
rect 18889 15997 18923 16031
rect 18981 15997 19015 16031
rect 19993 15997 20027 16031
rect 20085 15997 20119 16031
rect 20361 15997 20395 16031
rect 23673 15997 23707 16031
rect 23949 15997 23983 16031
rect 25237 15997 25271 16031
rect 25789 15997 25823 16031
rect 27169 15997 27203 16031
rect 27721 15997 27755 16031
rect 27905 15997 27939 16031
rect 29009 15997 29043 16031
rect 29285 15997 29319 16031
rect 29561 15997 29595 16031
rect 32873 15997 32907 16031
rect 33241 15997 33275 16031
rect 34069 15997 34103 16031
rect 34897 15997 34931 16031
rect 36461 15997 36495 16031
rect 37197 15997 37231 16031
rect 37381 15997 37415 16031
rect 39037 15997 39071 16031
rect 39221 15997 39255 16031
rect 39405 15997 39439 16031
rect 39773 15997 39807 16031
rect 40325 15997 40359 16031
rect 40509 15997 40543 16031
rect 42165 15997 42199 16031
rect 46213 15997 46247 16031
rect 46765 15997 46799 16031
rect 47317 15997 47351 16031
rect 49801 15997 49835 16031
rect 50353 15997 50387 16031
rect 51549 15997 51583 16031
rect 51733 15997 51767 16031
rect 52009 15997 52043 16031
rect 53297 15997 53331 16031
rect 10701 15929 10735 15963
rect 10977 15929 11011 15963
rect 13369 15929 13403 15963
rect 16497 15929 16531 15963
rect 17417 15929 17451 15963
rect 18061 15929 18095 15963
rect 22109 15929 22143 15963
rect 23857 15929 23891 15963
rect 27813 15929 27847 15963
rect 32413 15929 32447 15963
rect 38577 15929 38611 15963
rect 51917 15929 51951 15963
rect 7389 15861 7423 15895
rect 7849 15861 7883 15895
rect 15025 15861 15059 15895
rect 15761 15861 15795 15895
rect 19809 15861 19843 15895
rect 23489 15861 23523 15895
rect 28641 15861 28675 15895
rect 31217 15861 31251 15895
rect 31953 15861 31987 15895
rect 32229 15861 32263 15895
rect 34621 15861 34655 15895
rect 34897 15861 34931 15895
rect 35081 15861 35115 15895
rect 35541 15861 35575 15895
rect 36001 15861 36035 15895
rect 37565 15861 37599 15895
rect 38117 15861 38151 15895
rect 38485 15861 38519 15895
rect 40693 15861 40727 15895
rect 41061 15861 41095 15895
rect 41613 15861 41647 15895
rect 48697 15861 48731 15895
rect 49341 15861 49375 15895
rect 50721 15861 50755 15895
rect 51181 15861 51215 15895
rect 53205 15861 53239 15895
rect 57529 15861 57563 15895
rect 6929 15657 6963 15691
rect 9137 15657 9171 15691
rect 15485 15657 15519 15691
rect 19165 15657 19199 15691
rect 23489 15657 23523 15691
rect 24041 15657 24075 15691
rect 24409 15657 24443 15691
rect 29745 15657 29779 15691
rect 30389 15657 30423 15691
rect 31125 15657 31159 15691
rect 31585 15657 31619 15691
rect 31953 15657 31987 15691
rect 33701 15657 33735 15691
rect 34805 15657 34839 15691
rect 40141 15657 40175 15691
rect 40877 15657 40911 15691
rect 47225 15657 47259 15691
rect 48605 15657 48639 15691
rect 49985 15657 50019 15691
rect 52469 15657 52503 15691
rect 54033 15657 54067 15691
rect 8217 15589 8251 15623
rect 8769 15589 8803 15623
rect 13645 15589 13679 15623
rect 14473 15589 14507 15623
rect 17601 15589 17635 15623
rect 17877 15589 17911 15623
rect 18429 15589 18463 15623
rect 18705 15589 18739 15623
rect 20361 15589 20395 15623
rect 21465 15589 21499 15623
rect 21649 15589 21683 15623
rect 8309 15521 8343 15555
rect 10333 15521 10367 15555
rect 10977 15521 11011 15555
rect 13461 15521 13495 15555
rect 13737 15521 13771 15555
rect 15301 15521 15335 15555
rect 17233 15521 17267 15555
rect 17969 15521 18003 15555
rect 19533 15521 19567 15555
rect 19809 15521 19843 15555
rect 20729 15521 20763 15555
rect 26065 15589 26099 15623
rect 27169 15589 27203 15623
rect 27721 15589 27755 15623
rect 27997 15589 28031 15623
rect 28549 15589 28583 15623
rect 30665 15589 30699 15623
rect 32321 15589 32355 15623
rect 33977 15589 34011 15623
rect 34529 15589 34563 15623
rect 47501 15589 47535 15623
rect 48053 15589 48087 15623
rect 49157 15589 49191 15623
rect 52653 15589 52687 15623
rect 23489 15521 23523 15555
rect 24225 15521 24259 15555
rect 25881 15521 25915 15555
rect 27077 15521 27111 15555
rect 27261 15521 27295 15555
rect 29009 15521 29043 15555
rect 29193 15521 29227 15555
rect 29377 15521 29411 15555
rect 29745 15521 29779 15555
rect 30941 15521 30975 15555
rect 32413 15521 32447 15555
rect 34069 15521 34103 15555
rect 35357 15521 35391 15555
rect 36553 15521 36587 15555
rect 41889 15521 41923 15555
rect 42073 15521 42107 15555
rect 42257 15521 42291 15555
rect 46213 15521 46247 15555
rect 46857 15521 46891 15555
rect 47593 15521 47627 15555
rect 49249 15521 49283 15555
rect 51273 15521 51307 15555
rect 51641 15521 51675 15555
rect 53113 15521 53147 15555
rect 53481 15521 53515 15555
rect 53573 15521 53607 15555
rect 56885 15521 56919 15555
rect 57069 15521 57103 15555
rect 57253 15521 57287 15555
rect 5365 15453 5399 15487
rect 5641 15453 5675 15487
rect 11253 15453 11287 15487
rect 19993 15453 20027 15487
rect 21649 15453 21683 15487
rect 21741 15453 21775 15487
rect 22017 15453 22051 15487
rect 26893 15453 26927 15487
rect 28365 15453 28399 15487
rect 29929 15453 29963 15487
rect 32137 15453 32171 15487
rect 38301 15453 38335 15487
rect 38577 15453 38611 15487
rect 38853 15453 38887 15487
rect 50813 15453 50847 15487
rect 51733 15453 51767 15487
rect 56149 15453 56183 15487
rect 56425 15453 56459 15487
rect 58081 15453 58115 15487
rect 8033 15385 8067 15419
rect 13001 15385 13035 15419
rect 16681 15385 16715 15419
rect 25881 15385 25915 15419
rect 35541 15385 35575 15419
rect 36737 15385 36771 15419
rect 41245 15385 41279 15419
rect 41705 15385 41739 15419
rect 46397 15385 46431 15419
rect 7665 15317 7699 15351
rect 10609 15317 10643 15351
rect 12541 15317 12575 15351
rect 13277 15317 13311 15351
rect 13921 15317 13955 15351
rect 16313 15317 16347 15351
rect 17693 15317 17727 15351
rect 21097 15317 21131 15351
rect 23305 15317 23339 15351
rect 23673 15317 23707 15351
rect 25605 15317 25639 15351
rect 32597 15317 32631 15351
rect 33333 15317 33367 15351
rect 33793 15317 33827 15351
rect 35173 15317 35207 15351
rect 36185 15317 36219 15351
rect 37197 15317 37231 15351
rect 37473 15317 37507 15351
rect 38301 15317 38335 15351
rect 38393 15317 38427 15351
rect 40509 15317 40543 15351
rect 42901 15317 42935 15351
rect 43545 15317 43579 15351
rect 43913 15317 43947 15351
rect 47317 15317 47351 15351
rect 48973 15317 49007 15351
rect 49433 15317 49467 15351
rect 50353 15317 50387 15351
rect 52193 15317 52227 15351
rect 55689 15317 55723 15351
rect 57805 15317 57839 15351
rect 4537 15113 4571 15147
rect 6193 15113 6227 15147
rect 7205 15113 7239 15147
rect 22753 15113 22787 15147
rect 28273 15113 28307 15147
rect 29009 15113 29043 15147
rect 29285 15113 29319 15147
rect 29745 15113 29779 15147
rect 30297 15113 30331 15147
rect 31309 15113 31343 15147
rect 31769 15113 31803 15147
rect 32045 15113 32079 15147
rect 32873 15113 32907 15147
rect 34069 15113 34103 15147
rect 36829 15113 36863 15147
rect 38393 15113 38427 15147
rect 39865 15113 39899 15147
rect 42349 15113 42383 15147
rect 43913 15113 43947 15147
rect 49985 15113 50019 15147
rect 51365 15113 51399 15147
rect 51549 15113 51583 15147
rect 51917 15113 51951 15147
rect 53849 15113 53883 15147
rect 56885 15113 56919 15147
rect 58909 15113 58943 15147
rect 8861 15045 8895 15079
rect 11069 15045 11103 15079
rect 14105 15045 14139 15079
rect 14473 15045 14507 15079
rect 15577 15045 15611 15079
rect 16405 15045 16439 15079
rect 17509 15045 17543 15079
rect 21005 15045 21039 15079
rect 21373 15045 21407 15079
rect 23121 15045 23155 15079
rect 25605 15045 25639 15079
rect 25697 15045 25731 15079
rect 27077 15045 27111 15079
rect 27905 15045 27939 15079
rect 31125 15045 31159 15079
rect 32505 15045 32539 15079
rect 33241 15045 33275 15079
rect 9781 14977 9815 15011
rect 13737 14977 13771 15011
rect 15209 14977 15243 15011
rect 18797 14977 18831 15011
rect 20545 14977 20579 15011
rect 22385 14977 22419 15011
rect 24409 14977 24443 15011
rect 25053 14977 25087 15011
rect 27997 14977 28031 15011
rect 28733 14977 28767 15011
rect 5273 14909 5307 14943
rect 5365 14909 5399 14943
rect 5457 14909 5491 14943
rect 7297 14909 7331 14943
rect 7573 14909 7607 14943
rect 10241 14909 10275 14943
rect 10425 14909 10459 14943
rect 10563 14909 10597 14943
rect 12449 14909 12483 14943
rect 12909 14909 12943 14943
rect 13277 14909 13311 14943
rect 13369 14909 13403 14943
rect 14289 14909 14323 14943
rect 14933 14909 14967 14943
rect 15393 14909 15427 14943
rect 16865 14909 16899 14943
rect 18061 14909 18095 14943
rect 18337 14909 18371 14943
rect 19349 14909 19383 14943
rect 20085 14909 20119 14943
rect 20453 14909 20487 14943
rect 21925 14909 21959 14943
rect 22293 14909 22327 14943
rect 23673 14909 23707 14943
rect 23949 14909 23983 14943
rect 25605 14909 25639 14943
rect 25881 14909 25915 14943
rect 25973 14909 26007 14943
rect 27629 14909 27663 14943
rect 27776 14909 27810 14943
rect 29561 14909 29595 14943
rect 30573 14909 30607 14943
rect 30849 14909 30883 14943
rect 4905 14841 4939 14875
rect 5917 14841 5951 14875
rect 9229 14841 9263 14875
rect 11897 14841 11931 14875
rect 18245 14841 18279 14875
rect 19625 14841 19659 14875
rect 21465 14841 21499 14875
rect 23857 14841 23891 14875
rect 24685 14841 24719 14875
rect 26433 14841 26467 14875
rect 27537 14841 27571 14875
rect 29469 14841 29503 14875
rect 35725 15045 35759 15079
rect 41337 15045 41371 15079
rect 46765 15045 46799 15079
rect 47593 15045 47627 15079
rect 49433 15045 49467 15079
rect 49525 15045 49559 15079
rect 34713 14977 34747 15011
rect 37381 14977 37415 15011
rect 39589 14977 39623 15011
rect 42809 14977 42843 15011
rect 43637 14977 43671 15011
rect 48973 14977 49007 15011
rect 31861 14909 31895 14943
rect 33425 14909 33459 14943
rect 33609 14909 33643 14943
rect 33793 14909 33827 14943
rect 34069 14909 34103 14943
rect 35081 14909 35115 14943
rect 35449 14909 35483 14943
rect 36737 14909 36771 14943
rect 38853 14909 38887 14943
rect 39037 14909 39071 14943
rect 39129 14909 39163 14943
rect 41521 14909 41555 14943
rect 41889 14909 41923 14943
rect 41981 14909 42015 14943
rect 42901 14909 42935 14943
rect 43085 14909 43119 14943
rect 43177 14909 43211 14943
rect 46489 14909 46523 14943
rect 46581 14909 46615 14943
rect 47133 14909 47167 14943
rect 48145 14909 48179 14943
rect 48329 14909 48363 14943
rect 48513 14909 48547 14943
rect 49801 14909 49835 14943
rect 30941 14841 30975 14875
rect 31125 14841 31159 14875
rect 34253 14841 34287 14875
rect 34897 14841 34931 14875
rect 36553 14841 36587 14875
rect 38761 14841 38795 14875
rect 40325 14841 40359 14875
rect 46305 14841 46339 14875
rect 52653 15045 52687 15079
rect 52837 15045 52871 15079
rect 54217 15045 54251 15079
rect 52377 14977 52411 15011
rect 53573 14977 53607 15011
rect 51733 14909 51767 14943
rect 53021 14909 53055 14943
rect 53113 14909 53147 14943
rect 55689 14909 55723 14943
rect 55873 14909 55907 14943
rect 55965 14909 55999 14943
rect 57345 14909 57379 14943
rect 57621 14909 57655 14943
rect 47685 14841 47719 14875
rect 49709 14841 49743 14875
rect 50997 14841 51031 14875
rect 51549 14841 51583 14875
rect 55597 14841 55631 14875
rect 56425 14841 56459 14875
rect 6561 14773 6595 14807
rect 11437 14773 11471 14807
rect 12265 14773 12299 14807
rect 16037 14773 16071 14807
rect 16773 14773 16807 14807
rect 17049 14773 17083 14807
rect 17877 14773 17911 14807
rect 19165 14773 19199 14807
rect 19349 14773 19383 14807
rect 19533 14773 19567 14807
rect 30573 14773 30607 14807
rect 30665 14773 30699 14807
rect 36369 14773 36403 14807
rect 37749 14773 37783 14807
rect 40693 14773 40727 14807
rect 46489 14773 46523 14807
rect 50537 14773 50571 14807
rect 10701 14569 10735 14603
rect 10885 14569 10919 14603
rect 14197 14569 14231 14603
rect 18889 14569 18923 14603
rect 20545 14569 20579 14603
rect 32413 14569 32447 14603
rect 34161 14569 34195 14603
rect 42717 14569 42751 14603
rect 42993 14569 43027 14603
rect 47133 14569 47167 14603
rect 53205 14569 53239 14603
rect 55965 14569 55999 14603
rect 58449 14569 58483 14603
rect 8769 14501 8803 14535
rect 5825 14433 5859 14467
rect 6009 14433 6043 14467
rect 6101 14433 6135 14467
rect 6653 14433 6687 14467
rect 7849 14433 7883 14467
rect 8217 14433 8251 14467
rect 8309 14433 8343 14467
rect 9689 14433 9723 14467
rect 9873 14433 9907 14467
rect 7389 14365 7423 14399
rect 10241 14365 10275 14399
rect 13185 14501 13219 14535
rect 23857 14501 23891 14535
rect 27721 14501 27755 14535
rect 29377 14501 29411 14535
rect 30941 14501 30975 14535
rect 35449 14501 35483 14535
rect 37565 14501 37599 14535
rect 38117 14501 38151 14535
rect 40877 14501 40911 14535
rect 41797 14501 41831 14535
rect 42349 14501 42383 14535
rect 49525 14501 49559 14535
rect 11253 14433 11287 14467
rect 13461 14433 13495 14467
rect 14013 14433 14047 14467
rect 15301 14433 15335 14467
rect 18521 14433 18555 14467
rect 19625 14433 19659 14467
rect 19993 14433 20027 14467
rect 24869 14433 24903 14467
rect 25145 14433 25179 14467
rect 26617 14433 26651 14467
rect 27169 14433 27203 14467
rect 28457 14433 28491 14467
rect 29745 14433 29779 14467
rect 30205 14433 30239 14467
rect 35541 14433 35575 14467
rect 37933 14433 37967 14467
rect 38209 14433 38243 14467
rect 39957 14433 39991 14467
rect 40141 14433 40175 14467
rect 40325 14433 40359 14467
rect 41889 14433 41923 14467
rect 43361 14433 43395 14467
rect 45477 14433 45511 14467
rect 45569 14433 45603 14467
rect 48513 14433 48547 14467
rect 48973 14433 49007 14467
rect 52653 14433 52687 14467
rect 57345 14433 57379 14467
rect 11529 14365 11563 14399
rect 11805 14365 11839 14399
rect 16865 14365 16899 14399
rect 17141 14365 17175 14399
rect 21833 14365 21867 14399
rect 22109 14365 22143 14399
rect 25053 14365 25087 14399
rect 25605 14365 25639 14399
rect 27868 14365 27902 14399
rect 28089 14365 28123 14399
rect 30573 14365 30607 14399
rect 32781 14365 32815 14399
rect 33057 14365 33091 14399
rect 35265 14365 35299 14399
rect 38945 14365 38979 14399
rect 39313 14365 39347 14399
rect 39497 14365 39531 14399
rect 41613 14365 41647 14399
rect 44649 14365 44683 14399
rect 45017 14365 45051 14399
rect 45845 14365 45879 14399
rect 47501 14365 47535 14399
rect 50169 14365 50203 14399
rect 50445 14365 50479 14399
rect 51549 14365 51583 14399
rect 54585 14365 54619 14399
rect 54861 14365 54895 14399
rect 56517 14365 56551 14399
rect 57069 14365 57103 14399
rect 31585 14297 31619 14331
rect 34805 14297 34839 14331
rect 44281 14297 44315 14331
rect 52101 14297 52135 14331
rect 5641 14229 5675 14263
rect 6285 14229 6319 14263
rect 6653 14229 6687 14263
rect 6929 14229 6963 14263
rect 9321 14229 9355 14263
rect 10701 14229 10735 14263
rect 13921 14229 13955 14263
rect 14749 14229 14783 14263
rect 15485 14229 15519 14263
rect 15945 14229 15979 14263
rect 16313 14229 16347 14263
rect 16773 14229 16807 14263
rect 19257 14229 19291 14263
rect 21097 14229 21131 14263
rect 21465 14229 21499 14263
rect 23397 14229 23431 14263
rect 24225 14229 24259 14263
rect 25881 14229 25915 14263
rect 26249 14229 26283 14263
rect 26801 14229 26835 14263
rect 27537 14229 27571 14263
rect 27997 14229 28031 14263
rect 28825 14229 28859 14263
rect 30370 14229 30404 14263
rect 30481 14229 30515 14263
rect 31953 14229 31987 14263
rect 35081 14229 35115 14263
rect 35725 14229 35759 14263
rect 36277 14229 36311 14263
rect 36737 14229 36771 14263
rect 37013 14229 37047 14263
rect 38393 14229 38427 14263
rect 41429 14229 41463 14263
rect 43545 14229 43579 14263
rect 43913 14229 43947 14263
rect 48237 14229 48271 14263
rect 49157 14229 49191 14263
rect 49893 14229 49927 14263
rect 52837 14229 52871 14263
rect 53665 14229 53699 14263
rect 56885 14229 56919 14263
rect 59001 14229 59035 14263
rect 4905 14025 4939 14059
rect 6561 14025 6595 14059
rect 6837 14025 6871 14059
rect 7481 14025 7515 14059
rect 7573 14025 7607 14059
rect 8033 14025 8067 14059
rect 8585 14025 8619 14059
rect 8953 14025 8987 14059
rect 10793 14025 10827 14059
rect 11253 14025 11287 14059
rect 12081 14025 12115 14059
rect 12633 14025 12667 14059
rect 16405 14025 16439 14059
rect 20177 14025 20211 14059
rect 22569 14025 22603 14059
rect 27169 14025 27203 14059
rect 28089 14025 28123 14059
rect 29009 14025 29043 14059
rect 29837 14025 29871 14059
rect 33609 14025 33643 14059
rect 36001 14025 36035 14059
rect 36369 14025 36403 14059
rect 39313 14025 39347 14059
rect 41705 14025 41739 14059
rect 42625 14025 42659 14059
rect 43269 14025 43303 14059
rect 44005 14025 44039 14059
rect 45845 14025 45879 14059
rect 47501 14025 47535 14059
rect 48329 14025 48363 14059
rect 49065 14025 49099 14059
rect 49893 14025 49927 14059
rect 50077 14025 50111 14059
rect 50905 14025 50939 14059
rect 51089 14025 51123 14059
rect 51917 14025 51951 14059
rect 53021 14025 53055 14059
rect 56149 14025 56183 14059
rect 57069 14025 57103 14059
rect 58725 14025 58759 14059
rect 5917 13889 5951 13923
rect 14105 13957 14139 13991
rect 16129 13957 16163 13991
rect 19349 13957 19383 13991
rect 23857 13957 23891 13991
rect 27537 13957 27571 13991
rect 27905 13957 27939 13991
rect 31033 13957 31067 13991
rect 36645 13957 36679 13991
rect 38301 13957 38335 13991
rect 38761 13957 38795 13991
rect 39129 13957 39163 13991
rect 42257 13957 42291 13991
rect 9137 13889 9171 13923
rect 10701 13889 10735 13923
rect 12081 13889 12115 13923
rect 12173 13889 12207 13923
rect 13369 13889 13403 13923
rect 13737 13889 13771 13923
rect 14749 13889 14783 13923
rect 16865 13889 16899 13923
rect 17233 13889 17267 13923
rect 18061 13889 18095 13923
rect 23305 13889 23339 13923
rect 24869 13889 24903 13923
rect 25973 13889 26007 13923
rect 26065 13889 26099 13923
rect 26249 13889 26283 13923
rect 26801 13889 26835 13923
rect 27997 13889 28031 13923
rect 28733 13889 28767 13923
rect 30481 13889 30515 13923
rect 3893 13821 3927 13855
rect 3985 13821 4019 13855
rect 4169 13821 4203 13855
rect 4537 13821 4571 13855
rect 5273 13821 5307 13855
rect 5365 13821 5399 13855
rect 5549 13821 5583 13855
rect 6285 13821 6319 13855
rect 6837 13821 6871 13855
rect 7021 13821 7055 13855
rect 7757 13821 7791 13855
rect 7849 13821 7883 13855
rect 9229 13821 9263 13855
rect 10977 13821 11011 13855
rect 11069 13821 11103 13855
rect 11897 13821 11931 13855
rect 12817 13821 12851 13855
rect 12909 13821 12943 13855
rect 14841 13821 14875 13855
rect 15209 13821 15243 13855
rect 15301 13821 15335 13855
rect 15761 13821 15795 13855
rect 16221 13821 16255 13855
rect 18521 13821 18555 13855
rect 18705 13821 18739 13855
rect 18889 13821 18923 13855
rect 19901 13821 19935 13855
rect 20085 13821 20119 13855
rect 20729 13821 20763 13855
rect 21281 13821 21315 13855
rect 21741 13821 21775 13855
rect 21925 13821 21959 13855
rect 22109 13821 22143 13855
rect 23673 13821 23707 13855
rect 24225 13821 24259 13855
rect 24961 13821 24995 13855
rect 25421 13821 25455 13855
rect 26341 13821 26375 13855
rect 27629 13821 27663 13855
rect 27776 13821 27810 13855
rect 29929 13821 29963 13855
rect 30021 13821 30055 13855
rect 31493 13889 31527 13923
rect 33241 13889 33275 13923
rect 35633 13889 35667 13923
rect 37473 13889 37507 13923
rect 38025 13889 38059 13923
rect 39221 13889 39255 13923
rect 40049 13889 40083 13923
rect 40509 13889 40543 13923
rect 43085 13889 43119 13923
rect 32229 13821 32263 13855
rect 32781 13821 32815 13855
rect 33057 13821 33091 13855
rect 33885 13821 33919 13855
rect 34345 13821 34379 13855
rect 37289 13821 37323 13855
rect 37565 13821 37599 13855
rect 39000 13821 39034 13855
rect 40601 13821 40635 13855
rect 41061 13821 41095 13855
rect 41981 13821 42015 13855
rect 42128 13821 42162 13855
rect 42320 13821 42354 13855
rect 43821 13957 43855 13991
rect 44925 13957 44959 13991
rect 47777 13957 47811 13991
rect 49801 13957 49835 13991
rect 43913 13889 43947 13923
rect 48200 13889 48234 13923
rect 48421 13889 48455 13923
rect 48513 13889 48547 13923
rect 49617 13889 49651 13923
rect 43545 13821 43579 13855
rect 43692 13821 43726 13855
rect 46581 13821 46615 13855
rect 46765 13821 46799 13855
rect 46949 13821 46983 13855
rect 9689 13753 9723 13787
rect 14197 13753 14231 13787
rect 21189 13753 21223 13787
rect 22937 13753 22971 13787
rect 24685 13753 24719 13787
rect 25697 13753 25731 13787
rect 25973 13753 26007 13787
rect 30757 13753 30791 13787
rect 31033 13753 31067 13787
rect 31217 13753 31251 13787
rect 32137 13753 32171 13787
rect 34621 13753 34655 13787
rect 34897 13753 34931 13787
rect 35265 13753 35299 13787
rect 38853 13753 38887 13787
rect 43269 13753 43303 13787
rect 44557 13753 44591 13787
rect 46121 13753 46155 13787
rect 48053 13753 48087 13787
rect 54309 13957 54343 13991
rect 55137 13957 55171 13991
rect 57621 13957 57655 13991
rect 50261 13821 50295 13855
rect 50353 13821 50387 13855
rect 50813 13821 50847 13855
rect 50905 13821 50939 13855
rect 51733 13821 51767 13855
rect 52653 13821 52687 13855
rect 52837 13821 52871 13855
rect 53389 13821 53423 13855
rect 54769 13821 54803 13855
rect 55321 13821 55355 13855
rect 55505 13821 55539 13855
rect 55689 13821 55723 13855
rect 56517 13821 56551 13855
rect 57805 13821 57839 13855
rect 57989 13821 58023 13855
rect 58173 13821 58207 13855
rect 59001 13821 59035 13855
rect 10057 13685 10091 13719
rect 17877 13685 17911 13719
rect 19717 13685 19751 13719
rect 35081 13685 35115 13719
rect 35173 13685 35207 13719
rect 43361 13685 43395 13719
rect 45569 13685 45603 13719
rect 49801 13685 49835 13719
rect 51457 13685 51491 13719
rect 52285 13685 52319 13719
rect 6101 13481 6135 13515
rect 7573 13481 7607 13515
rect 7757 13481 7791 13515
rect 8953 13481 8987 13515
rect 15669 13481 15703 13515
rect 16405 13481 16439 13515
rect 25145 13481 25179 13515
rect 25513 13481 25547 13515
rect 26249 13481 26283 13515
rect 27813 13481 27847 13515
rect 28181 13481 28215 13515
rect 28549 13481 28583 13515
rect 28917 13481 28951 13515
rect 29285 13481 29319 13515
rect 29745 13481 29779 13515
rect 30481 13481 30515 13515
rect 31125 13481 31159 13515
rect 36645 13481 36679 13515
rect 41613 13481 41647 13515
rect 42349 13481 42383 13515
rect 42809 13481 42843 13515
rect 44189 13481 44223 13515
rect 46673 13481 46707 13515
rect 47869 13481 47903 13515
rect 6285 13413 6319 13447
rect 10609 13413 10643 13447
rect 11713 13413 11747 13447
rect 4997 13345 5031 13379
rect 6929 13345 6963 13379
rect 7297 13345 7331 13379
rect 7573 13345 7607 13379
rect 9781 13345 9815 13379
rect 12173 13345 12207 13379
rect 12541 13345 12575 13379
rect 12633 13345 12667 13379
rect 13093 13345 13127 13379
rect 13829 13345 13863 13379
rect 14013 13345 14047 13379
rect 14749 13345 14783 13379
rect 15301 13345 15335 13379
rect 4905 13277 4939 13311
rect 5457 13277 5491 13311
rect 6837 13277 6871 13311
rect 7389 13277 7423 13311
rect 7665 13277 7699 13311
rect 9699 13277 9733 13311
rect 10241 13277 10275 13311
rect 14381 13277 14415 13311
rect 15025 13277 15059 13311
rect 11437 13209 11471 13243
rect 13461 13209 13495 13243
rect 15485 13209 15519 13243
rect 16773 13413 16807 13447
rect 27169 13413 27203 13447
rect 31585 13413 31619 13447
rect 33701 13413 33735 13447
rect 37565 13413 37599 13447
rect 39037 13413 39071 13447
rect 39589 13413 39623 13447
rect 40141 13413 40175 13447
rect 42257 13413 42291 13447
rect 45017 13413 45051 13447
rect 45385 13413 45419 13447
rect 45937 13413 45971 13447
rect 46305 13413 46339 13447
rect 47317 13413 47351 13447
rect 16589 13345 16623 13379
rect 17417 13345 17451 13379
rect 17785 13345 17819 13379
rect 17969 13345 18003 13379
rect 18981 13345 19015 13379
rect 19809 13345 19843 13379
rect 21097 13345 21131 13379
rect 21833 13345 21867 13379
rect 22017 13345 22051 13379
rect 22201 13345 22235 13379
rect 23121 13345 23155 13379
rect 24041 13345 24075 13379
rect 25329 13345 25363 13379
rect 28733 13345 28767 13379
rect 29837 13345 29871 13379
rect 30941 13345 30975 13379
rect 31953 13345 31987 13379
rect 32321 13345 32355 13379
rect 32413 13345 32447 13379
rect 33517 13345 33551 13379
rect 34253 13345 34287 13379
rect 34437 13345 34471 13379
rect 34621 13345 34655 13379
rect 36001 13345 36035 13379
rect 38117 13345 38151 13379
rect 15945 13277 15979 13311
rect 17325 13277 17359 13311
rect 19533 13277 19567 13311
rect 19993 13277 20027 13311
rect 20637 13277 20671 13311
rect 21281 13277 21315 13311
rect 23213 13277 23247 13311
rect 23765 13277 23799 13311
rect 24225 13277 24259 13311
rect 27537 13277 27571 13311
rect 34805 13277 34839 13311
rect 35081 13277 35115 13311
rect 36369 13277 36403 13311
rect 37013 13277 37047 13311
rect 38025 13277 38059 13311
rect 38577 13277 38611 13311
rect 20361 13209 20395 13243
rect 21649 13209 21683 13243
rect 22753 13209 22787 13243
rect 25881 13209 25915 13243
rect 27334 13209 27368 13243
rect 35449 13209 35483 13243
rect 39405 13345 39439 13379
rect 39681 13345 39715 13379
rect 40417 13345 40451 13379
rect 40969 13345 41003 13379
rect 42993 13345 43027 13379
rect 43085 13345 43119 13379
rect 43361 13345 43395 13379
rect 43453 13345 43487 13379
rect 43913 13345 43947 13379
rect 44005 13345 44039 13379
rect 44557 13345 44591 13379
rect 45477 13345 45511 13379
rect 46857 13345 46891 13379
rect 40877 13277 40911 13311
rect 41337 13277 41371 13311
rect 42257 13277 42291 13311
rect 41134 13209 41168 13243
rect 46765 13277 46799 13311
rect 44005 13209 44039 13243
rect 48513 13481 48547 13515
rect 49617 13481 49651 13515
rect 50261 13481 50295 13515
rect 54769 13481 54803 13515
rect 55505 13481 55539 13515
rect 57161 13481 57195 13515
rect 53757 13413 53791 13447
rect 57713 13413 57747 13447
rect 58081 13413 58115 13447
rect 58449 13413 58483 13447
rect 48329 13345 48363 13379
rect 48513 13345 48547 13379
rect 48973 13345 49007 13379
rect 51089 13345 51123 13379
rect 51365 13345 51399 13379
rect 52377 13345 52411 13379
rect 54585 13345 54619 13379
rect 58265 13345 58299 13379
rect 58541 13345 58575 13379
rect 49341 13277 49375 13311
rect 50537 13277 50571 13311
rect 51549 13277 51583 13311
rect 55137 13277 55171 13311
rect 55781 13277 55815 13311
rect 56057 13277 56091 13311
rect 53481 13209 53515 13243
rect 2421 13141 2455 13175
rect 3893 13141 3927 13175
rect 4721 13141 4755 13175
rect 5825 13141 5859 13175
rect 7665 13141 7699 13175
rect 8125 13141 8159 13175
rect 8493 13141 8527 13175
rect 9413 13141 9447 13175
rect 11161 13141 11195 13175
rect 15669 13141 15703 13175
rect 16313 13141 16347 13175
rect 18613 13141 18647 13175
rect 21281 13141 21315 13175
rect 24869 13141 24903 13175
rect 26709 13141 26743 13175
rect 27445 13141 27479 13175
rect 30021 13141 30055 13175
rect 32137 13141 32171 13175
rect 32597 13141 32631 13175
rect 33241 13141 33275 13175
rect 35817 13141 35851 13175
rect 36166 13141 36200 13175
rect 36277 13141 36311 13175
rect 39037 13141 39071 13175
rect 39221 13141 39255 13175
rect 41245 13141 41279 13175
rect 41981 13141 42015 13175
rect 43085 13141 43119 13175
rect 45201 13141 45235 13175
rect 47593 13141 47627 13175
rect 47869 13141 47903 13175
rect 48053 13141 48087 13175
rect 48145 13141 48179 13175
rect 48697 13141 48731 13175
rect 49111 13141 49145 13175
rect 49249 13141 49283 13175
rect 51825 13141 51859 13175
rect 52193 13141 52227 13175
rect 52561 13141 52595 13175
rect 53021 13141 53055 13175
rect 58725 13141 58759 13175
rect 59277 13141 59311 13175
rect 3157 12937 3191 12971
rect 4077 12937 4111 12971
rect 9781 12937 9815 12971
rect 11069 12937 11103 12971
rect 14565 12937 14599 12971
rect 17417 12937 17451 12971
rect 18521 12937 18555 12971
rect 22385 12937 22419 12971
rect 22937 12937 22971 12971
rect 23397 12937 23431 12971
rect 24225 12937 24259 12971
rect 25605 12937 25639 12971
rect 28089 12937 28123 12971
rect 28457 12937 28491 12971
rect 30941 12937 30975 12971
rect 32689 12937 32723 12971
rect 35173 12937 35207 12971
rect 38117 12937 38151 12971
rect 38577 12937 38611 12971
rect 39313 12937 39347 12971
rect 39865 12937 39899 12971
rect 40693 12937 40727 12971
rect 41061 12937 41095 12971
rect 41521 12937 41555 12971
rect 44557 12937 44591 12971
rect 45201 12937 45235 12971
rect 45661 12937 45695 12971
rect 47225 12937 47259 12971
rect 47593 12937 47627 12971
rect 48651 12937 48685 12971
rect 49157 12937 49191 12971
rect 50721 12937 50755 12971
rect 58265 12937 58299 12971
rect 2973 12801 3007 12835
rect 2421 12733 2455 12767
rect 2605 12733 2639 12767
rect 12725 12869 12759 12903
rect 14105 12869 14139 12903
rect 16405 12869 16439 12903
rect 24501 12869 24535 12903
rect 25973 12869 26007 12903
rect 27445 12869 27479 12903
rect 27813 12869 27847 12903
rect 29469 12869 29503 12903
rect 29745 12869 29779 12903
rect 29929 12869 29963 12903
rect 43545 12869 43579 12903
rect 46489 12869 46523 12903
rect 47087 12869 47121 12903
rect 48789 12869 48823 12903
rect 49893 12869 49927 12903
rect 50353 12869 50387 12903
rect 51089 12869 51123 12903
rect 52653 12869 52687 12903
rect 56057 12869 56091 12903
rect 56793 12869 56827 12903
rect 6653 12801 6687 12835
rect 7665 12801 7699 12835
rect 8769 12801 8803 12835
rect 9965 12801 9999 12835
rect 10701 12801 10735 12835
rect 12173 12801 12207 12835
rect 12817 12801 12851 12835
rect 13461 12801 13495 12835
rect 24685 12801 24719 12835
rect 25237 12801 25271 12835
rect 26341 12801 26375 12835
rect 3801 12733 3835 12767
rect 3985 12733 4019 12767
rect 4445 12733 4479 12767
rect 4997 12733 5031 12767
rect 5181 12733 5215 12767
rect 5457 12733 5491 12767
rect 5917 12733 5951 12767
rect 7205 12733 7239 12767
rect 8125 12733 8159 12767
rect 8309 12733 8343 12767
rect 8585 12733 8619 12767
rect 9137 12733 9171 12767
rect 10149 12733 10183 12767
rect 12596 12733 12630 12767
rect 14749 12733 14783 12767
rect 14841 12733 14875 12767
rect 15301 12733 15335 12767
rect 16037 12733 16071 12767
rect 16589 12733 16623 12767
rect 16957 12733 16991 12767
rect 17049 12733 17083 12767
rect 18245 12733 18279 12767
rect 18429 12733 18463 12767
rect 19625 12733 19659 12767
rect 19901 12733 19935 12767
rect 22293 12733 22327 12767
rect 23673 12733 23707 12767
rect 24777 12733 24811 12767
rect 26065 12733 26099 12767
rect 27813 12733 27847 12767
rect 29285 12733 29319 12767
rect 5365 12665 5399 12699
rect 6193 12665 6227 12699
rect 10333 12665 10367 12699
rect 11805 12665 11839 12699
rect 12449 12665 12483 12699
rect 14473 12665 14507 12699
rect 19533 12665 19567 12699
rect 21833 12665 21867 12699
rect 22109 12665 22143 12699
rect 23765 12665 23799 12699
rect 31769 12801 31803 12835
rect 33149 12801 33183 12835
rect 33701 12801 33735 12835
rect 36277 12801 36311 12835
rect 37565 12801 37599 12835
rect 43269 12801 43303 12835
rect 46765 12801 46799 12835
rect 47317 12801 47351 12835
rect 47961 12801 47995 12835
rect 48329 12801 48363 12835
rect 48881 12801 48915 12835
rect 49525 12801 49559 12835
rect 50445 12801 50479 12835
rect 50905 12801 50939 12835
rect 53849 12801 53883 12835
rect 55413 12801 55447 12835
rect 58633 12801 58667 12835
rect 58909 12801 58943 12835
rect 30205 12733 30239 12767
rect 31401 12733 31435 12767
rect 33241 12733 33275 12767
rect 33610 12733 33644 12767
rect 35081 12733 35115 12767
rect 36737 12733 36771 12767
rect 37013 12733 37047 12767
rect 37197 12733 37231 12767
rect 37749 12733 37783 12767
rect 39037 12733 39071 12767
rect 39170 12733 39204 12767
rect 40509 12733 40543 12767
rect 41613 12733 41647 12767
rect 41889 12733 41923 12767
rect 44465 12733 44499 12767
rect 45845 12733 45879 12767
rect 50224 12733 50258 12767
rect 30665 12665 30699 12699
rect 31217 12665 31251 12699
rect 32137 12665 32171 12699
rect 34069 12665 34103 12699
rect 34897 12665 34931 12699
rect 40325 12665 40359 12699
rect 43913 12665 43947 12699
rect 44281 12665 44315 12699
rect 46949 12665 46983 12699
rect 48513 12665 48547 12699
rect 50077 12665 50111 12699
rect 51917 12733 51951 12767
rect 53297 12733 53331 12767
rect 53389 12733 53423 12767
rect 54401 12733 54435 12767
rect 54677 12733 54711 12767
rect 54953 12733 54987 12767
rect 57345 12733 57379 12767
rect 57897 12733 57931 12767
rect 51457 12665 51491 12699
rect 51733 12665 51767 12699
rect 52929 12665 52963 12699
rect 54861 12665 54895 12699
rect 56425 12665 56459 12699
rect 3157 12597 3191 12631
rect 3341 12597 3375 12631
rect 4445 12597 4479 12631
rect 4721 12597 4755 12631
rect 7573 12597 7607 12631
rect 9505 12597 9539 12631
rect 10241 12597 10275 12631
rect 11345 12597 11379 12631
rect 13093 12597 13127 12631
rect 15669 12597 15703 12631
rect 17877 12597 17911 12631
rect 19073 12597 19107 12631
rect 21189 12597 21223 12631
rect 28733 12597 28767 12631
rect 29745 12597 29779 12631
rect 32413 12597 32447 12631
rect 34621 12597 34655 12631
rect 35817 12597 35851 12631
rect 36185 12597 36219 12631
rect 38945 12597 38979 12631
rect 50905 12597 50939 12631
rect 52009 12597 52043 12631
rect 54125 12597 54159 12631
rect 54401 12597 54435 12631
rect 54493 12597 54527 12631
rect 55689 12597 55723 12631
rect 57529 12597 57563 12631
rect 60013 12597 60047 12631
rect 6561 12393 6595 12427
rect 7297 12393 7331 12427
rect 8861 12393 8895 12427
rect 10241 12393 10275 12427
rect 11345 12393 11379 12427
rect 12081 12393 12115 12427
rect 12449 12393 12483 12427
rect 15577 12393 15611 12427
rect 17693 12393 17727 12427
rect 18061 12393 18095 12427
rect 19533 12393 19567 12427
rect 24501 12393 24535 12427
rect 24961 12393 24995 12427
rect 26249 12393 26283 12427
rect 27721 12393 27755 12427
rect 27997 12393 28031 12427
rect 33241 12393 33275 12427
rect 33517 12393 33551 12427
rect 35265 12393 35299 12427
rect 36369 12393 36403 12427
rect 37197 12393 37231 12427
rect 40233 12393 40267 12427
rect 40693 12393 40727 12427
rect 41613 12393 41647 12427
rect 41797 12393 41831 12427
rect 43085 12393 43119 12427
rect 58817 12393 58851 12427
rect 3157 12325 3191 12359
rect 8125 12325 8159 12359
rect 9321 12325 9355 12359
rect 13369 12325 13403 12359
rect 17233 12325 17267 12359
rect 20913 12325 20947 12359
rect 22017 12325 22051 12359
rect 22201 12325 22235 12359
rect 23489 12325 23523 12359
rect 2605 12257 2639 12291
rect 2789 12257 2823 12291
rect 5089 12257 5123 12291
rect 5457 12257 5491 12291
rect 7389 12257 7423 12291
rect 10701 12257 10735 12291
rect 11805 12257 11839 12291
rect 12265 12257 12299 12291
rect 14197 12257 14231 12291
rect 15025 12257 15059 12291
rect 15301 12257 15335 12291
rect 15485 12257 15519 12291
rect 16681 12257 16715 12291
rect 16865 12257 16899 12291
rect 17693 12257 17727 12291
rect 18245 12257 18279 12291
rect 18889 12257 18923 12291
rect 20637 12257 20671 12291
rect 21373 12257 21407 12291
rect 21741 12257 21775 12291
rect 21833 12257 21867 12291
rect 3525 12189 3559 12223
rect 4629 12189 4663 12223
rect 5549 12189 5583 12223
rect 7536 12189 7570 12223
rect 7757 12189 7791 12223
rect 8493 12189 8527 12223
rect 11069 12189 11103 12223
rect 13185 12189 13219 12223
rect 13921 12189 13955 12223
rect 14381 12189 14415 12223
rect 16129 12189 16163 12223
rect 16589 12189 16623 12223
rect 19257 12189 19291 12223
rect 10866 12121 10900 12155
rect 14749 12121 14783 12155
rect 17969 12121 18003 12155
rect 19027 12121 19061 12155
rect 20453 12121 20487 12155
rect 22937 12257 22971 12291
rect 23029 12257 23063 12291
rect 24961 12257 24995 12291
rect 25329 12257 25363 12291
rect 26694 12257 26728 12291
rect 26801 12257 26835 12291
rect 27261 12257 27295 12291
rect 27445 12257 27479 12291
rect 22753 12189 22787 12223
rect 31493 12325 31527 12359
rect 31677 12325 31711 12359
rect 33701 12325 33735 12359
rect 37749 12325 37783 12359
rect 28733 12257 28767 12291
rect 28825 12257 28859 12291
rect 29561 12257 29595 12291
rect 30113 12257 30147 12291
rect 30665 12257 30699 12291
rect 31769 12257 31803 12291
rect 32321 12257 32355 12291
rect 32413 12257 32447 12291
rect 34345 12257 34379 12291
rect 34713 12257 34747 12291
rect 34897 12257 34931 12291
rect 35725 12257 35759 12291
rect 38577 12257 38611 12291
rect 38761 12257 38795 12291
rect 39037 12257 39071 12291
rect 39681 12257 39715 12291
rect 40785 12257 40819 12291
rect 40932 12257 40966 12291
rect 31217 12189 31251 12223
rect 31953 12189 31987 12223
rect 32873 12189 32907 12223
rect 34253 12189 34287 12223
rect 36093 12189 36127 12223
rect 38301 12189 38335 12223
rect 41153 12189 41187 12223
rect 28273 12121 28307 12155
rect 29929 12121 29963 12155
rect 30297 12121 30331 12155
rect 35863 12121 35897 12155
rect 39589 12121 39623 12155
rect 41245 12121 41279 12155
rect 46121 12325 46155 12359
rect 46305 12325 46339 12359
rect 48789 12325 48823 12359
rect 50353 12325 50387 12359
rect 54861 12325 54895 12359
rect 55873 12325 55907 12359
rect 61025 12325 61059 12359
rect 43545 12257 43579 12291
rect 44097 12257 44131 12291
rect 42257 12189 42291 12223
rect 44189 12189 44223 12223
rect 44465 12189 44499 12223
rect 45569 12189 45603 12223
rect 46765 12257 46799 12291
rect 48053 12257 48087 12291
rect 49065 12257 49099 12291
rect 50721 12257 50755 12291
rect 51549 12257 51583 12291
rect 53205 12257 53239 12291
rect 54401 12257 54435 12291
rect 55137 12257 55171 12291
rect 57069 12257 57103 12291
rect 57805 12257 57839 12291
rect 60197 12257 60231 12291
rect 60289 12257 60323 12291
rect 46489 12189 46523 12223
rect 46673 12189 46707 12223
rect 47225 12189 47259 12223
rect 47501 12189 47535 12223
rect 48973 12189 49007 12223
rect 51273 12189 51307 12223
rect 51733 12189 51767 12223
rect 53113 12189 53147 12223
rect 53665 12189 53699 12223
rect 55505 12189 55539 12223
rect 58081 12189 58115 12223
rect 58449 12189 58483 12223
rect 52745 12121 52779 12155
rect 57345 12121 57379 12155
rect 6929 12053 6963 12087
rect 7665 12053 7699 12087
rect 10609 12053 10643 12087
rect 10977 12053 11011 12087
rect 12909 12053 12943 12087
rect 17509 12053 17543 12087
rect 18797 12053 18831 12087
rect 19165 12053 19199 12087
rect 19993 12053 20027 12087
rect 22017 12053 22051 12087
rect 22569 12053 22603 12087
rect 23765 12053 23799 12087
rect 24133 12053 24167 12087
rect 25881 12053 25915 12087
rect 27997 12053 28031 12087
rect 28549 12053 28583 12087
rect 29009 12053 29043 12087
rect 35633 12053 35667 12087
rect 36001 12053 36035 12087
rect 36829 12053 36863 12087
rect 39865 12053 39899 12087
rect 41061 12053 41095 12087
rect 41613 12053 41647 12087
rect 42533 12053 42567 12087
rect 46305 12053 46339 12087
rect 48421 12053 48455 12087
rect 49249 12053 49283 12087
rect 50077 12053 50111 12087
rect 52009 12053 52043 12087
rect 52377 12053 52411 12087
rect 53941 12053 53975 12087
rect 55275 12053 55309 12087
rect 55413 12053 55447 12087
rect 56241 12053 56275 12087
rect 56609 12053 56643 12087
rect 56885 12053 56919 12087
rect 59185 12053 59219 12087
rect 59737 12053 59771 12087
rect 60473 12053 60507 12087
rect 2881 11849 2915 11883
rect 4629 11849 4663 11883
rect 5825 11849 5859 11883
rect 6561 11849 6595 11883
rect 7941 11849 7975 11883
rect 8769 11849 8803 11883
rect 10333 11849 10367 11883
rect 12173 11849 12207 11883
rect 14289 11849 14323 11883
rect 15669 11849 15703 11883
rect 16773 11849 16807 11883
rect 17049 11849 17083 11883
rect 21833 11849 21867 11883
rect 23857 11849 23891 11883
rect 27445 11849 27479 11883
rect 29009 11849 29043 11883
rect 30481 11849 30515 11883
rect 33149 11849 33183 11883
rect 34345 11849 34379 11883
rect 35081 11849 35115 11883
rect 35541 11849 35575 11883
rect 36185 11849 36219 11883
rect 38945 11849 38979 11883
rect 39773 11849 39807 11883
rect 40233 11849 40267 11883
rect 40877 11849 40911 11883
rect 41245 11849 41279 11883
rect 42441 11849 42475 11883
rect 43085 11849 43119 11883
rect 48421 11849 48455 11883
rect 48789 11849 48823 11883
rect 49709 11849 49743 11883
rect 50537 11849 50571 11883
rect 51549 11849 51583 11883
rect 52239 11849 52273 11883
rect 52377 11849 52411 11883
rect 52561 11849 52595 11883
rect 53481 11849 53515 11883
rect 54585 11849 54619 11883
rect 56333 11849 56367 11883
rect 58449 11849 58483 11883
rect 7205 11781 7239 11815
rect 7573 11781 7607 11815
rect 11897 11781 11931 11815
rect 12725 11781 12759 11815
rect 15393 11781 15427 11815
rect 15945 11781 15979 11815
rect 21097 11781 21131 11815
rect 30849 11781 30883 11815
rect 36737 11781 36771 11815
rect 41613 11781 41647 11815
rect 3341 11713 3375 11747
rect 7665 11713 7699 11747
rect 8309 11713 8343 11747
rect 10701 11713 10735 11747
rect 10793 11713 10827 11747
rect 11989 11713 12023 11747
rect 3065 11645 3099 11679
rect 7444 11645 7478 11679
rect 8861 11645 8895 11679
rect 8953 11645 8987 11679
rect 10977 11645 11011 11679
rect 11069 11645 11103 11679
rect 7297 11577 7331 11611
rect 9413 11577 9447 11611
rect 11161 11577 11195 11611
rect 11529 11577 11563 11611
rect 25789 11713 25823 11747
rect 27169 11713 27203 11747
rect 31585 11713 31619 11747
rect 33885 11713 33919 11747
rect 37749 11713 37783 11747
rect 42257 11713 42291 11747
rect 44097 11781 44131 11815
rect 44465 11781 44499 11815
rect 52009 11781 52043 11815
rect 54401 11781 54435 11815
rect 55965 11781 55999 11815
rect 59553 11781 59587 11815
rect 42625 11713 42659 11747
rect 45477 11713 45511 11747
rect 47409 11713 47443 11747
rect 49433 11713 49467 11747
rect 52469 11713 52503 11747
rect 53113 11713 53147 11747
rect 54493 11713 54527 11747
rect 55137 11713 55171 11747
rect 55505 11713 55539 11747
rect 56057 11713 56091 11747
rect 56701 11713 56735 11747
rect 58725 11713 58759 11747
rect 13093 11645 13127 11679
rect 13369 11645 13403 11679
rect 14381 11645 14415 11679
rect 14473 11645 14507 11679
rect 15393 11645 15427 11679
rect 15761 11645 15795 11679
rect 16865 11645 16899 11679
rect 17417 11645 17451 11679
rect 18337 11645 18371 11679
rect 18429 11645 18463 11679
rect 19717 11645 19751 11679
rect 19993 11645 20027 11679
rect 22201 11645 22235 11679
rect 22293 11645 22327 11679
rect 23489 11645 23523 11679
rect 24317 11645 24351 11679
rect 25513 11645 25547 11679
rect 27997 11645 28031 11679
rect 28549 11645 28583 11679
rect 29285 11645 29319 11679
rect 29469 11645 29503 11679
rect 30665 11645 30699 11679
rect 31953 11645 31987 11679
rect 33057 11645 33091 11679
rect 33425 11645 33459 11679
rect 35725 11645 35759 11679
rect 35909 11645 35943 11679
rect 36001 11645 36035 11679
rect 37473 11645 37507 11679
rect 38853 11645 38887 11679
rect 41797 11645 41831 11679
rect 42165 11645 42199 11679
rect 42441 11645 42475 11679
rect 44649 11645 44683 11679
rect 44833 11645 44867 11679
rect 45017 11645 45051 11679
rect 46305 11645 46339 11679
rect 46857 11645 46891 11679
rect 46949 11645 46983 11679
rect 47685 11645 47719 11679
rect 49065 11645 49099 11679
rect 50261 11645 50295 11679
rect 50353 11645 50387 11679
rect 52101 11645 52135 11679
rect 54125 11645 54159 11679
rect 54272 11645 54306 11679
rect 55836 11645 55870 11679
rect 57069 11645 57103 11679
rect 57437 11645 57471 11679
rect 57805 11645 57839 11679
rect 58173 11645 58207 11679
rect 59093 11645 59127 11679
rect 59737 11645 59771 11679
rect 59921 11645 59955 11679
rect 60105 11645 60139 11679
rect 13921 11577 13955 11611
rect 14933 11577 14967 11611
rect 18889 11577 18923 11611
rect 22753 11577 22787 11611
rect 24133 11577 24167 11611
rect 24685 11577 24719 11611
rect 31309 11577 31343 11611
rect 31769 11577 31803 11611
rect 32321 11577 32355 11611
rect 33333 11577 33367 11611
rect 37105 11577 37139 11611
rect 37289 11577 37323 11611
rect 38669 11577 38703 11611
rect 45845 11577 45879 11611
rect 46765 11577 46799 11611
rect 48881 11577 48915 11611
rect 50077 11577 50111 11611
rect 51181 11577 51215 11611
rect 55689 11577 55723 11611
rect 61301 11577 61335 11611
rect 2513 11509 2547 11543
rect 5089 11509 5123 11543
rect 5549 11509 5583 11543
rect 9781 11509 9815 11543
rect 11989 11509 12023 11543
rect 12909 11509 12943 11543
rect 15209 11509 15243 11543
rect 16405 11509 16439 11543
rect 17785 11509 17819 11543
rect 19257 11509 19291 11543
rect 23029 11509 23063 11543
rect 25053 11509 25087 11543
rect 27813 11509 27847 11543
rect 28181 11509 28215 11543
rect 29561 11509 29595 11543
rect 30205 11509 30239 11543
rect 32689 11509 32723 11543
rect 38301 11509 38335 11543
rect 43729 11509 43763 11543
rect 54033 11509 54067 11543
rect 60565 11509 60599 11543
rect 61025 11509 61059 11543
rect 6009 11305 6043 11339
rect 7941 11305 7975 11339
rect 8401 11305 8435 11339
rect 10701 11305 10735 11339
rect 11161 11305 11195 11339
rect 14289 11305 14323 11339
rect 15117 11305 15151 11339
rect 17049 11305 17083 11339
rect 18797 11305 18831 11339
rect 21833 11305 21867 11339
rect 22017 11305 22051 11339
rect 22109 11305 22143 11339
rect 22569 11305 22603 11339
rect 22937 11305 22971 11339
rect 23305 11305 23339 11339
rect 26709 11305 26743 11339
rect 29561 11305 29595 11339
rect 31125 11305 31159 11339
rect 33241 11305 33275 11339
rect 33701 11305 33735 11339
rect 36093 11305 36127 11339
rect 37473 11305 37507 11339
rect 38301 11305 38335 11339
rect 51273 11305 51307 11339
rect 53021 11305 53055 11339
rect 53481 11305 53515 11339
rect 54217 11305 54251 11339
rect 54953 11305 54987 11339
rect 57805 11305 57839 11339
rect 59553 11305 59587 11339
rect 61577 11305 61611 11339
rect 8861 11237 8895 11271
rect 13185 11237 13219 11271
rect 15301 11237 15335 11271
rect 16037 11237 16071 11271
rect 19993 11237 20027 11271
rect 20729 11237 20763 11271
rect 20913 11237 20947 11271
rect 21649 11237 21683 11271
rect 7297 11169 7331 11203
rect 9689 11169 9723 11203
rect 9781 11169 9815 11203
rect 11989 11169 12023 11203
rect 12173 11169 12207 11203
rect 12357 11169 12391 11203
rect 13645 11169 13679 11203
rect 14657 11169 14691 11203
rect 17969 11169 18003 11203
rect 18429 11169 18463 11203
rect 19257 11169 19291 11203
rect 4629 11101 4663 11135
rect 4905 11101 4939 11135
rect 7444 11101 7478 11135
rect 7665 11101 7699 11135
rect 14013 11101 14047 11135
rect 15669 11101 15703 11135
rect 16773 11101 16807 11135
rect 17877 11101 17911 11135
rect 19625 11101 19659 11135
rect 21281 11101 21315 11135
rect 24317 11237 24351 11271
rect 25605 11237 25639 11271
rect 32965 11237 32999 11271
rect 35449 11237 35483 11271
rect 36277 11237 36311 11271
rect 36829 11237 36863 11271
rect 40141 11237 40175 11271
rect 47225 11237 47259 11271
rect 48053 11237 48087 11271
rect 49525 11237 49559 11271
rect 50905 11237 50939 11271
rect 52469 11237 52503 11271
rect 52837 11237 52871 11271
rect 57161 11237 57195 11271
rect 22477 11169 22511 11203
rect 23489 11169 23523 11203
rect 23673 11169 23707 11203
rect 24041 11169 24075 11203
rect 25053 11169 25087 11203
rect 25145 11169 25179 11203
rect 26249 11169 26283 11203
rect 26525 11169 26559 11203
rect 29929 11169 29963 11203
rect 30941 11169 30975 11203
rect 32505 11169 32539 11203
rect 34069 11169 34103 11203
rect 36461 11169 36495 11203
rect 38025 11169 38059 11203
rect 40417 11169 40451 11203
rect 41613 11169 41647 11203
rect 41797 11169 41831 11203
rect 41981 11169 42015 11203
rect 43361 11169 43395 11203
rect 44649 11169 44683 11203
rect 47593 11169 47627 11203
rect 49065 11169 49099 11203
rect 49985 11169 50019 11203
rect 50445 11169 50479 11203
rect 52009 11169 52043 11203
rect 53021 11169 53055 11203
rect 53297 11169 53331 11203
rect 53849 11169 53883 11203
rect 55137 11169 55171 11203
rect 55597 11169 55631 11203
rect 56425 11169 56459 11203
rect 58081 11169 58115 11203
rect 58725 11169 58759 11203
rect 59093 11169 59127 11203
rect 59921 11169 59955 11203
rect 60473 11169 60507 11203
rect 22109 11101 22143 11135
rect 27629 11101 27663 11135
rect 27905 11101 27939 11135
rect 32413 11101 32447 11135
rect 33793 11101 33827 11135
rect 38485 11101 38519 11135
rect 38761 11101 38795 11135
rect 41061 11101 41095 11135
rect 42901 11101 42935 11135
rect 44925 11101 44959 11135
rect 46029 11101 46063 11135
rect 46857 11101 46891 11135
rect 47501 11101 47535 11135
rect 48973 11101 49007 11135
rect 50353 11101 50387 11135
rect 51917 11101 51951 11135
rect 53205 11101 53239 11135
rect 55045 11101 55079 11135
rect 56793 11101 56827 11135
rect 59185 11101 59219 11135
rect 60197 11101 60231 11135
rect 3157 11033 3191 11067
rect 6837 11033 6871 11067
rect 11805 11033 11839 11067
rect 17785 11033 17819 11067
rect 19073 11033 19107 11067
rect 19395 11033 19429 11067
rect 21078 11033 21112 11067
rect 21833 11033 21867 11067
rect 24777 11033 24811 11067
rect 29009 11033 29043 11067
rect 31585 11033 31619 11067
rect 31953 11033 31987 11067
rect 35725 11033 35759 11067
rect 41429 11033 41463 11067
rect 43545 11033 43579 11067
rect 48421 11033 48455 11067
rect 58541 11033 58575 11067
rect 4261 10965 4295 10999
rect 7113 10965 7147 10999
rect 7573 10965 7607 10999
rect 9229 10965 9263 10999
rect 9965 10965 9999 10999
rect 12817 10965 12851 10999
rect 13810 10965 13844 10999
rect 13921 10965 13955 10999
rect 15466 10965 15500 10999
rect 15577 10965 15611 10999
rect 16313 10965 16347 10999
rect 19533 10965 19567 10999
rect 20361 10965 20395 10999
rect 21189 10965 21223 10999
rect 22293 10965 22327 10999
rect 24869 10965 24903 10999
rect 25973 10965 26007 10999
rect 27169 10965 27203 10999
rect 30389 10965 30423 10999
rect 30757 10965 30791 10999
rect 37105 10965 37139 10999
rect 42441 10965 42475 10999
rect 43913 10965 43947 10999
rect 44373 10965 44407 10999
rect 48789 10965 48823 10999
rect 51733 10965 51767 10999
rect 55965 10965 55999 10999
rect 56590 10965 56624 10999
rect 56701 10965 56735 10999
rect 5641 10761 5675 10795
rect 8125 10761 8159 10795
rect 8493 10761 8527 10795
rect 8953 10761 8987 10795
rect 9965 10761 9999 10795
rect 11253 10761 11287 10795
rect 15209 10761 15243 10795
rect 16589 10761 16623 10795
rect 19533 10761 19567 10795
rect 21557 10761 21591 10795
rect 21925 10761 21959 10795
rect 30205 10761 30239 10795
rect 30481 10761 30515 10795
rect 33885 10761 33919 10795
rect 36369 10761 36403 10795
rect 38393 10761 38427 10795
rect 44557 10761 44591 10795
rect 46397 10761 46431 10795
rect 47317 10761 47351 10795
rect 47869 10761 47903 10795
rect 50169 10761 50203 10795
rect 51457 10761 51491 10795
rect 55137 10761 55171 10795
rect 56149 10761 56183 10795
rect 56793 10761 56827 10795
rect 57621 10761 57655 10795
rect 61209 10761 61243 10795
rect 10241 10693 10275 10727
rect 12173 10693 12207 10727
rect 14473 10693 14507 10727
rect 15853 10693 15887 10727
rect 16221 10693 16255 10727
rect 17141 10693 17175 10727
rect 22937 10693 22971 10727
rect 23489 10693 23523 10727
rect 40233 10693 40267 10727
rect 43177 10693 43211 10727
rect 43729 10693 43763 10727
rect 48329 10693 48363 10727
rect 51917 10693 51951 10727
rect 60841 10693 60875 10727
rect 3801 10625 3835 10659
rect 10793 10625 10827 10659
rect 10977 10625 11011 10659
rect 12725 10625 12759 10659
rect 14105 10625 14139 10659
rect 14933 10625 14967 10659
rect 18061 10625 18095 10659
rect 18613 10625 18647 10659
rect 21005 10625 21039 10659
rect 22661 10625 22695 10659
rect 24317 10625 24351 10659
rect 25421 10625 25455 10659
rect 27997 10625 28031 10659
rect 28457 10625 28491 10659
rect 29285 10625 29319 10659
rect 29837 10625 29871 10659
rect 32229 10625 32263 10659
rect 35633 10625 35667 10659
rect 36461 10625 36495 10659
rect 36737 10625 36771 10659
rect 39405 10625 39439 10659
rect 40601 10625 40635 10659
rect 41613 10625 41647 10659
rect 42073 10625 42107 10659
rect 44281 10625 44315 10659
rect 45109 10625 45143 10659
rect 49341 10625 49375 10659
rect 51089 10625 51123 10659
rect 53021 10625 53055 10659
rect 57345 10625 57379 10659
rect 59553 10625 59587 10659
rect 4261 10557 4295 10591
rect 4537 10557 4571 10591
rect 6837 10557 6871 10591
rect 7297 10557 7331 10591
rect 7665 10557 7699 10591
rect 7757 10557 7791 10591
rect 8677 10557 8711 10591
rect 8769 10557 8803 10591
rect 11069 10557 11103 10591
rect 11805 10557 11839 10591
rect 12449 10557 12483 10591
rect 15025 10557 15059 10591
rect 18153 10557 18187 10591
rect 19625 10557 19659 10591
rect 19901 10557 19935 10591
rect 22293 10557 22327 10591
rect 23673 10557 23707 10591
rect 24869 10557 24903 10591
rect 24961 10557 24995 10591
rect 26249 10557 26283 10591
rect 26709 10557 26743 10591
rect 26985 10557 27019 10591
rect 27169 10557 27203 10591
rect 27353 10557 27387 10591
rect 27721 10557 27755 10591
rect 29377 10557 29411 10591
rect 30665 10557 30699 10591
rect 32328 10557 32362 10591
rect 32597 10557 32631 10591
rect 34529 10557 34563 10591
rect 35265 10557 35299 10591
rect 35909 10557 35943 10591
rect 38945 10557 38979 10591
rect 39129 10557 39163 10591
rect 39773 10557 39807 10591
rect 14841 10489 14875 10523
rect 18981 10489 19015 10523
rect 22109 10489 22143 10523
rect 26157 10489 26191 10523
rect 35081 10489 35115 10523
rect 40693 10557 40727 10591
rect 41245 10557 41279 10591
rect 41797 10557 41831 10591
rect 44373 10557 44407 10591
rect 46213 10557 46247 10591
rect 46765 10557 46799 10591
rect 47593 10557 47627 10591
rect 48513 10557 48547 10591
rect 48697 10557 48731 10591
rect 48881 10557 48915 10591
rect 49893 10557 49927 10591
rect 49985 10557 50019 10591
rect 50721 10557 50755 10591
rect 51733 10557 51767 10591
rect 53297 10557 53331 10591
rect 55873 10557 55907 10591
rect 55965 10557 55999 10591
rect 57437 10557 57471 10591
rect 58173 10557 58207 10591
rect 59277 10557 59311 10591
rect 4169 10421 4203 10455
rect 6285 10421 6319 10455
rect 6653 10421 6687 10455
rect 9597 10421 9631 10455
rect 17417 10421 17451 10455
rect 17877 10421 17911 10455
rect 23857 10421 23891 10455
rect 24777 10421 24811 10455
rect 25789 10421 25823 10455
rect 28825 10421 28859 10455
rect 30849 10421 30883 10455
rect 31309 10421 31343 10455
rect 31861 10421 31895 10455
rect 34345 10421 34379 10455
rect 34529 10421 34563 10455
rect 34713 10421 34747 10455
rect 38025 10421 38059 10455
rect 38761 10421 38795 10455
rect 40601 10421 40635 10455
rect 40877 10421 40911 10455
rect 44097 10421 44131 10455
rect 45477 10421 45511 10455
rect 45845 10421 45879 10455
rect 47409 10421 47443 10455
rect 49801 10421 49835 10455
rect 52285 10421 52319 10455
rect 52837 10421 52871 10455
rect 54401 10421 54435 10455
rect 55781 10421 55815 10455
rect 58817 10421 58851 10455
rect 59093 10421 59127 10455
rect 61577 10421 61611 10455
rect 61945 10421 61979 10455
rect 6745 10217 6779 10251
rect 8033 10217 8067 10251
rect 8677 10217 8711 10251
rect 13829 10217 13863 10251
rect 14197 10217 14231 10251
rect 14933 10217 14967 10251
rect 15853 10217 15887 10251
rect 20269 10217 20303 10251
rect 22937 10217 22971 10251
rect 24133 10217 24167 10251
rect 24869 10217 24903 10251
rect 26341 10217 26375 10251
rect 27077 10217 27111 10251
rect 32597 10217 32631 10251
rect 44097 10217 44131 10251
rect 46857 10217 46891 10251
rect 47961 10217 47995 10251
rect 48329 10217 48363 10251
rect 50905 10217 50939 10251
rect 53941 10217 53975 10251
rect 54401 10217 54435 10251
rect 54861 10217 54895 10251
rect 55781 10217 55815 10251
rect 56333 10217 56367 10251
rect 57253 10217 57287 10251
rect 57621 10217 57655 10251
rect 10241 10149 10275 10183
rect 13093 10149 13127 10183
rect 20913 10149 20947 10183
rect 24593 10149 24627 10183
rect 27813 10149 27847 10183
rect 29193 10149 29227 10183
rect 35633 10149 35667 10183
rect 39865 10149 39899 10183
rect 46029 10149 46063 10183
rect 51733 10149 51767 10183
rect 4445 10081 4479 10115
rect 6929 10081 6963 10115
rect 7389 10081 7423 10115
rect 7757 10081 7791 10115
rect 8033 10081 8067 10115
rect 9505 10081 9539 10115
rect 9781 10081 9815 10115
rect 11713 10081 11747 10115
rect 15301 10081 15335 10115
rect 17049 10081 17083 10115
rect 18337 10081 18371 10115
rect 18613 10081 18647 10115
rect 21373 10081 21407 10115
rect 21557 10081 21591 10115
rect 21741 10081 21775 10115
rect 22569 10081 22603 10115
rect 22753 10081 22787 10115
rect 23949 10081 23983 10115
rect 25145 10081 25179 10115
rect 25881 10081 25915 10115
rect 27353 10081 27387 10115
rect 28733 10081 28767 10115
rect 30021 10081 30055 10115
rect 31401 10081 31435 10115
rect 32137 10081 32171 10115
rect 32229 10081 32263 10115
rect 36093 10081 36127 10115
rect 36461 10081 36495 10115
rect 37289 10081 37323 10115
rect 38669 10081 38703 10115
rect 38853 10081 38887 10115
rect 39037 10081 39071 10115
rect 40417 10081 40451 10115
rect 40877 10081 40911 10115
rect 41797 10081 41831 10115
rect 44281 10081 44315 10115
rect 44833 10081 44867 10115
rect 45201 10081 45235 10115
rect 46673 10081 46707 10115
rect 47777 10081 47811 10115
rect 49065 10081 49099 10115
rect 49801 10081 49835 10115
rect 50537 10081 50571 10115
rect 51273 10081 51307 10115
rect 53021 10081 53055 10115
rect 53389 10081 53423 10115
rect 53481 10081 53515 10115
rect 55045 10081 55079 10115
rect 56517 10081 56551 10115
rect 58449 10081 58483 10115
rect 58817 10081 58851 10115
rect 60197 10081 60231 10115
rect 4721 10013 4755 10047
rect 5825 10013 5859 10047
rect 7849 10013 7883 10047
rect 8309 10013 8343 10047
rect 9689 10013 9723 10047
rect 11437 10013 11471 10047
rect 14565 10013 14599 10047
rect 16957 10013 16991 10047
rect 17509 10013 17543 10047
rect 22201 10013 22235 10047
rect 24777 10013 24811 10047
rect 25053 10013 25087 10047
rect 27261 10013 27295 10047
rect 28641 10013 28675 10047
rect 33149 10013 33183 10047
rect 33425 10013 33459 10047
rect 36553 10013 36587 10047
rect 40325 10013 40359 10047
rect 41153 10013 41187 10047
rect 41705 10013 41739 10047
rect 42533 10013 42567 10047
rect 45293 10013 45327 10047
rect 48973 10013 49007 10047
rect 51181 10013 51215 10047
rect 54953 10013 54987 10047
rect 56425 10013 56459 10047
rect 58357 10013 58391 10047
rect 58909 10013 58943 10047
rect 60473 10013 60507 10047
rect 15485 9945 15519 9979
rect 23397 9945 23431 9979
rect 30205 9945 30239 9979
rect 38485 9945 38519 9979
rect 44649 9945 44683 9979
rect 52377 9945 52411 9979
rect 52837 9945 52871 9979
rect 4261 9877 4295 9911
rect 6377 9877 6411 9911
rect 9137 9877 9171 9911
rect 10517 9877 10551 9911
rect 11069 9877 11103 9911
rect 13369 9877 13403 9911
rect 16313 9877 16347 9911
rect 16681 9877 16715 9911
rect 17785 9877 17819 9911
rect 18153 9877 18187 9911
rect 19717 9877 19751 9911
rect 20729 9877 20763 9911
rect 23857 9877 23891 9911
rect 24777 9877 24811 9911
rect 25329 9877 25363 9911
rect 28089 9877 28123 9911
rect 28457 9877 28491 9911
rect 29469 9877 29503 9911
rect 29929 9877 29963 9911
rect 30573 9877 30607 9911
rect 31033 9877 31067 9911
rect 31769 9877 31803 9911
rect 33057 9877 33091 9911
rect 34529 9877 34563 9911
rect 35265 9877 35299 9911
rect 36921 9877 36955 9911
rect 37933 9877 37967 9911
rect 39497 9877 39531 9911
rect 41521 9877 41555 9911
rect 41981 9877 42015 9911
rect 42901 9877 42935 9911
rect 43545 9877 43579 9911
rect 43913 9877 43947 9911
rect 46489 9877 46523 9911
rect 47225 9877 47259 9911
rect 47685 9877 47719 9911
rect 48697 9877 48731 9911
rect 49249 9877 49283 9911
rect 50169 9877 50203 9911
rect 50353 9877 50387 9911
rect 52009 9877 52043 9911
rect 55229 9877 55263 9911
rect 56701 9877 56735 9911
rect 57897 9877 57931 9911
rect 59369 9877 59403 9911
rect 59737 9877 59771 9911
rect 61761 9877 61795 9911
rect 5917 9673 5951 9707
rect 6285 9673 6319 9707
rect 11805 9673 11839 9707
rect 12265 9673 12299 9707
rect 14197 9673 14231 9707
rect 15025 9673 15059 9707
rect 16037 9673 16071 9707
rect 18981 9673 19015 9707
rect 22569 9673 22603 9707
rect 23213 9673 23247 9707
rect 27445 9673 27479 9707
rect 36369 9673 36403 9707
rect 39589 9673 39623 9707
rect 49617 9673 49651 9707
rect 54033 9673 54067 9707
rect 54401 9673 54435 9707
rect 55413 9673 55447 9707
rect 56425 9673 56459 9707
rect 58173 9673 58207 9707
rect 2973 9605 3007 9639
rect 5273 9605 5307 9639
rect 9229 9605 9263 9639
rect 12725 9605 12759 9639
rect 15117 9605 15151 9639
rect 15393 9605 15427 9639
rect 16497 9605 16531 9639
rect 19349 9605 19383 9639
rect 19809 9605 19843 9639
rect 22017 9605 22051 9639
rect 22753 9605 22787 9639
rect 23857 9605 23891 9639
rect 24593 9605 24627 9639
rect 26985 9605 27019 9639
rect 30113 9605 30147 9639
rect 31585 9605 31619 9639
rect 36737 9605 36771 9639
rect 37749 9605 37783 9639
rect 38485 9605 38519 9639
rect 39221 9605 39255 9639
rect 41061 9605 41095 9639
rect 42349 9605 42383 9639
rect 42441 9605 42475 9639
rect 44189 9605 44223 9639
rect 45293 9605 45327 9639
rect 45569 9605 45603 9639
rect 46673 9605 46707 9639
rect 47041 9605 47075 9639
rect 47501 9605 47535 9639
rect 50445 9605 50479 9639
rect 50721 9605 50755 9639
rect 51457 9605 51491 9639
rect 53665 9605 53699 9639
rect 56793 9605 56827 9639
rect 3801 9537 3835 9571
rect 3893 9537 3927 9571
rect 6837 9537 6871 9571
rect 8493 9537 8527 9571
rect 11529 9537 11563 9571
rect 13737 9537 13771 9571
rect 16589 9537 16623 9571
rect 17141 9537 17175 9571
rect 18705 9537 18739 9571
rect 21373 9537 21407 9571
rect 21925 9537 21959 9571
rect 22109 9537 22143 9571
rect 27537 9537 27571 9571
rect 28089 9537 28123 9571
rect 33517 9537 33551 9571
rect 2789 9469 2823 9503
rect 4169 9469 4203 9503
rect 7113 9469 7147 9503
rect 9321 9469 9355 9503
rect 9413 9469 9447 9503
rect 10977 9469 11011 9503
rect 11069 9469 11103 9503
rect 12909 9469 12943 9503
rect 13093 9469 13127 9503
rect 13277 9469 13311 9503
rect 14657 9469 14691 9503
rect 15301 9469 15335 9503
rect 15393 9469 15427 9503
rect 15485 9469 15519 9503
rect 16221 9469 16255 9503
rect 16681 9469 16715 9503
rect 17417 9469 17451 9503
rect 18153 9469 18187 9503
rect 18245 9469 18279 9503
rect 19993 9469 20027 9503
rect 20177 9469 20211 9503
rect 20361 9469 20395 9503
rect 21465 9469 21499 9503
rect 22937 9469 22971 9503
rect 24041 9469 24075 9503
rect 25053 9469 25087 9503
rect 25329 9469 25363 9503
rect 27629 9469 27663 9503
rect 28365 9469 28399 9503
rect 28733 9469 28767 9503
rect 29929 9469 29963 9503
rect 30573 9469 30607 9503
rect 31217 9469 31251 9503
rect 33425 9469 33459 9503
rect 33977 9469 34011 9503
rect 34161 9469 34195 9503
rect 34345 9469 34379 9503
rect 34989 9469 35023 9503
rect 35081 9469 35115 9503
rect 35173 9469 35207 9503
rect 35633 9469 35667 9503
rect 36921 9469 36955 9503
rect 37105 9469 37139 9503
rect 37289 9469 37323 9503
rect 38301 9469 38335 9503
rect 40325 9469 40359 9503
rect 41245 9469 41279 9503
rect 41429 9469 41463 9503
rect 41613 9469 41647 9503
rect 6653 9401 6687 9435
rect 9873 9401 9907 9435
rect 10241 9401 10275 9435
rect 20821 9401 20855 9435
rect 24133 9401 24167 9435
rect 29837 9401 29871 9435
rect 31677 9401 31711 9435
rect 38209 9401 38243 9435
rect 42901 9537 42935 9571
rect 48329 9537 48363 9571
rect 53113 9537 53147 9571
rect 54585 9537 54619 9571
rect 55137 9537 55171 9571
rect 58633 9537 58667 9571
rect 42625 9469 42659 9503
rect 45937 9469 45971 9503
rect 46857 9469 46891 9503
rect 48053 9469 48087 9503
rect 50537 9469 50571 9503
rect 51733 9469 51767 9503
rect 52009 9469 52043 9503
rect 54677 9469 54711 9503
rect 55965 9469 55999 9503
rect 58357 9469 58391 9503
rect 46397 9401 46431 9435
rect 50077 9401 50111 9435
rect 56057 9401 56091 9435
rect 3341 9333 3375 9367
rect 8861 9333 8895 9367
rect 10793 9333 10827 9367
rect 15669 9333 15703 9367
rect 16221 9333 16255 9367
rect 17785 9333 17819 9367
rect 21281 9333 21315 9367
rect 22293 9333 22327 9367
rect 24869 9333 24903 9367
rect 26433 9333 26467 9367
rect 30757 9333 30791 9367
rect 34989 9333 35023 9367
rect 35909 9333 35943 9367
rect 38853 9333 38887 9367
rect 42073 9333 42107 9367
rect 42349 9333 42383 9367
rect 44833 9333 44867 9367
rect 45753 9333 45787 9367
rect 47869 9333 47903 9367
rect 51181 9333 51215 9367
rect 55781 9333 55815 9367
rect 57805 9333 57839 9367
rect 59737 9333 59771 9367
rect 60473 9333 60507 9367
rect 60933 9333 60967 9367
rect 61301 9333 61335 9367
rect 7849 9129 7883 9163
rect 23581 9129 23615 9163
rect 33517 9129 33551 9163
rect 49157 9129 49191 9163
rect 61853 9129 61887 9163
rect 4813 9061 4847 9095
rect 6745 9061 6779 9095
rect 2605 8993 2639 9027
rect 2973 8993 3007 9027
rect 3065 8993 3099 9027
rect 5733 8993 5767 9027
rect 6653 8993 6687 9027
rect 7205 8993 7239 9027
rect 7573 8993 7607 9027
rect 9689 9061 9723 9095
rect 17785 9061 17819 9095
rect 18613 9061 18647 9095
rect 22845 9061 22879 9095
rect 24593 9061 24627 9095
rect 30481 9061 30515 9095
rect 33701 9061 33735 9095
rect 37933 9061 37967 9095
rect 38301 9061 38335 9095
rect 42349 9061 42383 9095
rect 43913 9061 43947 9095
rect 47777 9061 47811 9095
rect 49617 9061 49651 9095
rect 52653 9061 52687 9095
rect 54309 9061 54343 9095
rect 8769 8993 8803 9027
rect 9505 8993 9539 9027
rect 10149 8993 10183 9027
rect 10517 8993 10551 9027
rect 12357 8993 12391 9027
rect 13553 8993 13587 9027
rect 13737 8993 13771 9027
rect 15393 8993 15427 9027
rect 17025 8993 17059 9027
rect 17325 8993 17359 9027
rect 19073 8993 19107 9027
rect 19257 8993 19291 9027
rect 19441 8993 19475 9027
rect 21005 8993 21039 9027
rect 21465 8993 21499 9027
rect 22385 8993 22419 9027
rect 25053 8993 25087 9027
rect 25237 8993 25271 9027
rect 25421 8993 25455 9027
rect 27353 8993 27387 9027
rect 27813 8993 27847 9027
rect 28457 8993 28491 9027
rect 30021 8993 30055 9027
rect 31125 8993 31159 9027
rect 32413 8993 32447 9027
rect 34161 8993 34195 9027
rect 34529 8993 34563 9027
rect 35633 8993 35667 9027
rect 36369 8993 36403 9027
rect 41889 8993 41923 9027
rect 43453 8993 43487 9027
rect 47358 8993 47392 9027
rect 48053 8993 48087 9027
rect 48973 8993 49007 9027
rect 49341 8993 49375 9027
rect 50721 8993 50755 9027
rect 50905 8993 50939 9027
rect 51089 8993 51123 9027
rect 52193 8993 52227 9027
rect 53481 8993 53515 9027
rect 54677 8993 54711 9027
rect 58725 8993 58759 9027
rect 60657 8993 60691 9027
rect 61025 8993 61059 9027
rect 4905 8925 4939 8959
rect 5457 8925 5491 8959
rect 5917 8925 5951 8959
rect 7665 8925 7699 8959
rect 7849 8925 7883 8959
rect 8125 8925 8159 8959
rect 10609 8925 10643 8959
rect 11529 8925 11563 8959
rect 12081 8925 12115 8959
rect 12541 8925 12575 8959
rect 12909 8925 12943 8959
rect 13645 8925 13679 8959
rect 15301 8925 15335 8959
rect 17233 8925 17267 8959
rect 20637 8925 20671 8959
rect 20913 8925 20947 8959
rect 22293 8925 22327 8959
rect 23213 8925 23247 8959
rect 26525 8925 26559 8959
rect 27077 8925 27111 8959
rect 27537 8925 27571 8959
rect 28365 8925 28399 8959
rect 29929 8925 29963 8959
rect 30757 8925 30791 8959
rect 32321 8925 32355 8959
rect 32873 8925 32907 8959
rect 34621 8925 34655 8959
rect 35541 8925 35575 8959
rect 36093 8925 36127 8959
rect 38485 8925 38519 8959
rect 38761 8925 38795 8959
rect 41613 8925 41647 8959
rect 41797 8925 41831 8959
rect 43361 8925 43395 8959
rect 44741 8925 44775 8959
rect 45017 8925 45051 8959
rect 47225 8925 47259 8959
rect 2421 8857 2455 8891
rect 9045 8857 9079 8891
rect 11161 8857 11195 8891
rect 13369 8857 13403 8891
rect 14565 8857 14599 8891
rect 28181 8857 28215 8891
rect 40049 8857 40083 8891
rect 42993 8857 43027 8891
rect 46673 8857 46707 8891
rect 48789 8857 48823 8891
rect 52101 8925 52135 8959
rect 54585 8925 54619 8959
rect 56149 8925 56183 8959
rect 56425 8925 56459 8959
rect 58633 8925 58667 8959
rect 61117 8925 61151 8959
rect 61485 8925 61519 8959
rect 50537 8857 50571 8891
rect 53573 8857 53607 8891
rect 55413 8857 55447 8891
rect 58173 8857 58207 8891
rect 60473 8857 60507 8891
rect 4261 8789 4295 8823
rect 6285 8789 6319 8823
rect 13185 8789 13219 8823
rect 13921 8789 13955 8823
rect 15117 8789 15151 8823
rect 15577 8789 15611 8823
rect 16129 8789 16163 8823
rect 16773 8789 16807 8823
rect 16865 8789 16899 8823
rect 18245 8789 18279 8823
rect 19993 8789 20027 8823
rect 20361 8789 20395 8823
rect 21741 8789 21775 8823
rect 22109 8789 22143 8823
rect 24041 8789 24075 8823
rect 24409 8789 24443 8823
rect 25881 8789 25915 8823
rect 26249 8789 26283 8823
rect 28641 8789 28675 8823
rect 29285 8789 29319 8823
rect 29653 8789 29687 8823
rect 31585 8789 31619 8823
rect 31953 8789 31987 8823
rect 35081 8789 35115 8823
rect 36737 8789 36771 8823
rect 37197 8789 37231 8823
rect 40601 8789 40635 8823
rect 41245 8789 41279 8823
rect 42625 8789 42659 8823
rect 44281 8789 44315 8823
rect 44649 8789 44683 8823
rect 46305 8789 46339 8823
rect 47041 8789 47075 8823
rect 49341 8789 49375 8823
rect 50077 8789 50111 8823
rect 51549 8789 51583 8823
rect 52009 8789 52043 8823
rect 53021 8789 53055 8823
rect 54861 8789 54895 8823
rect 56057 8789 56091 8823
rect 57529 8789 57563 8823
rect 58449 8789 58483 8823
rect 58909 8789 58943 8823
rect 59461 8789 59495 8823
rect 59829 8789 59863 8823
rect 3065 8585 3099 8619
rect 8677 8585 8711 8619
rect 11897 8585 11931 8619
rect 12265 8585 12299 8619
rect 12633 8585 12667 8619
rect 15117 8585 15151 8619
rect 16037 8585 16071 8619
rect 16865 8585 16899 8619
rect 20177 8585 20211 8619
rect 21189 8585 21223 8619
rect 22845 8585 22879 8619
rect 24041 8585 24075 8619
rect 28457 8585 28491 8619
rect 30849 8585 30883 8619
rect 33057 8585 33091 8619
rect 33333 8585 33367 8619
rect 34621 8585 34655 8619
rect 36645 8585 36679 8619
rect 38761 8585 38795 8619
rect 42257 8585 42291 8619
rect 42717 8585 42751 8619
rect 48973 8585 49007 8619
rect 52745 8585 52779 8619
rect 53573 8585 53607 8619
rect 55321 8585 55355 8619
rect 57161 8585 57195 8619
rect 58633 8585 58667 8619
rect 61485 8585 61519 8619
rect 61853 8585 61887 8619
rect 3341 8517 3375 8551
rect 8033 8517 8067 8551
rect 8585 8517 8619 8551
rect 15669 8517 15703 8551
rect 18061 8517 18095 8551
rect 18383 8517 18417 8551
rect 24133 8517 24167 8551
rect 2697 8449 2731 8483
rect 4169 8449 4203 8483
rect 7849 8449 7883 8483
rect 7941 8449 7975 8483
rect 4261 8381 4295 8415
rect 4537 8381 4571 8415
rect 6837 8381 6871 8415
rect 7389 8381 7423 8415
rect 7665 8381 7699 8415
rect 8217 8449 8251 8483
rect 9413 8449 9447 8483
rect 14749 8449 14783 8483
rect 16589 8449 16623 8483
rect 18613 8449 18647 8483
rect 8033 8381 8067 8415
rect 8953 8381 8987 8415
rect 10609 8381 10643 8415
rect 11161 8381 11195 8415
rect 11253 8381 11287 8415
rect 14013 8381 14047 8415
rect 14289 8381 14323 8415
rect 14473 8381 14507 8415
rect 15485 8381 15519 8415
rect 16681 8381 16715 8415
rect 18061 8381 18095 8415
rect 18475 8381 18509 8415
rect 19257 8381 19291 8415
rect 20361 8381 20395 8415
rect 20729 8381 20763 8415
rect 21373 8381 21407 8415
rect 21465 8381 21499 8415
rect 21649 8381 21683 8415
rect 21741 8381 21775 8415
rect 22201 8381 22235 8415
rect 6653 8313 6687 8347
rect 7941 8313 7975 8347
rect 8861 8313 8895 8347
rect 9689 8313 9723 8347
rect 10333 8313 10367 8347
rect 13461 8313 13495 8347
rect 17417 8313 17451 8347
rect 18245 8313 18279 8347
rect 18981 8313 19015 8347
rect 29929 8517 29963 8551
rect 30205 8517 30239 8551
rect 40141 8517 40175 8551
rect 24317 8449 24351 8483
rect 24593 8449 24627 8483
rect 28825 8449 28859 8483
rect 29285 8449 29319 8483
rect 24501 8381 24535 8415
rect 25697 8381 25731 8415
rect 26065 8381 26099 8415
rect 26341 8381 26375 8415
rect 26617 8381 26651 8415
rect 27169 8381 27203 8415
rect 27629 8381 27663 8415
rect 27905 8381 27939 8415
rect 29377 8381 29411 8415
rect 22569 8313 22603 8347
rect 24133 8313 24167 8347
rect 29837 8313 29871 8347
rect 31769 8449 31803 8483
rect 32413 8449 32447 8483
rect 37105 8449 37139 8483
rect 37657 8449 37691 8483
rect 39037 8449 39071 8483
rect 39589 8449 39623 8483
rect 30665 8381 30699 8415
rect 31861 8381 31895 8415
rect 31953 8381 31987 8415
rect 33241 8381 33275 8415
rect 33793 8381 33827 8415
rect 34253 8381 34287 8415
rect 34529 8381 34563 8415
rect 34897 8381 34931 8415
rect 35265 8381 35299 8415
rect 35449 8381 35483 8415
rect 37197 8381 37231 8415
rect 37841 8381 37875 8415
rect 37933 8381 37967 8415
rect 39129 8381 39163 8415
rect 39865 8381 39899 8415
rect 35909 8313 35943 8347
rect 48513 8517 48547 8551
rect 51365 8517 51399 8551
rect 52009 8517 52043 8551
rect 52929 8517 52963 8551
rect 53205 8517 53239 8551
rect 61117 8517 61151 8551
rect 62221 8517 62255 8551
rect 41981 8449 42015 8483
rect 42717 8449 42751 8483
rect 44373 8449 44407 8483
rect 48697 8449 48731 8483
rect 50077 8449 50111 8483
rect 51089 8449 51123 8483
rect 51457 8449 51491 8483
rect 52101 8449 52135 8483
rect 40325 8381 40359 8415
rect 40509 8381 40543 8415
rect 40601 8381 40635 8415
rect 41061 8381 41095 8415
rect 42073 8381 42107 8415
rect 42809 8381 42843 8415
rect 43361 8381 43395 8415
rect 44511 8381 44545 8415
rect 44649 8381 44683 8415
rect 45937 8381 45971 8415
rect 46213 8381 46247 8415
rect 47041 8381 47075 8415
rect 47179 8381 47213 8415
rect 47501 8381 47535 8415
rect 47869 8381 47903 8415
rect 48830 8381 48864 8415
rect 49985 8381 50019 8415
rect 51365 8381 51399 8415
rect 51880 8381 51914 8415
rect 52929 8381 52963 8415
rect 54217 8381 54251 8415
rect 54953 8381 54987 8415
rect 55873 8381 55907 8415
rect 56195 8381 56229 8415
rect 56333 8381 56367 8415
rect 57529 8381 57563 8415
rect 58817 8381 58851 8415
rect 59093 8381 59127 8415
rect 60473 8381 60507 8415
rect 61301 8381 61335 8415
rect 38393 8313 38427 8347
rect 40141 8313 40175 8347
rect 41337 8313 41371 8347
rect 43821 8313 43855 8347
rect 45477 8313 45511 8347
rect 46305 8313 46339 8347
rect 50261 8313 50295 8347
rect 50445 8313 50479 8347
rect 50813 8313 50847 8347
rect 51733 8313 51767 8347
rect 52469 8313 52503 8347
rect 53849 8313 53883 8347
rect 54033 8313 54067 8347
rect 54585 8313 54619 8347
rect 55413 8313 55447 8347
rect 56701 8313 56735 8347
rect 57345 8313 57379 8347
rect 58173 8313 58207 8347
rect 5825 8245 5859 8279
rect 6285 8245 6319 8279
rect 10517 8245 10551 8279
rect 13277 8245 13311 8279
rect 16497 8245 16531 8279
rect 17785 8245 17819 8279
rect 19625 8245 19659 8279
rect 21373 8245 21407 8279
rect 23397 8245 23431 8279
rect 25053 8245 25087 8279
rect 27537 8245 27571 8279
rect 29929 8245 29963 8279
rect 30573 8245 30607 8279
rect 31309 8245 31343 8279
rect 32781 8245 32815 8279
rect 34529 8245 34563 8279
rect 36277 8245 36311 8279
rect 37841 8245 37875 8279
rect 41797 8245 41831 8279
rect 45109 8245 45143 8279
rect 49525 8245 49559 8279
rect 50353 8245 50387 8279
rect 57621 8245 57655 8279
rect 6377 8041 6411 8075
rect 6837 8041 6871 8075
rect 11529 8041 11563 8075
rect 17325 8041 17359 8075
rect 18981 8041 19015 8075
rect 20729 8041 20763 8075
rect 24777 8041 24811 8075
rect 30021 8041 30055 8075
rect 31861 8041 31895 8075
rect 32597 8041 32631 8075
rect 33425 8041 33459 8075
rect 34621 8041 34655 8075
rect 35265 8041 35299 8075
rect 43545 8041 43579 8075
rect 44097 8041 44131 8075
rect 45753 8041 45787 8075
rect 46949 8041 46983 8075
rect 48053 8041 48087 8075
rect 50997 8041 51031 8075
rect 51365 8041 51399 8075
rect 52837 8041 52871 8075
rect 53941 8041 53975 8075
rect 54309 8041 54343 8075
rect 55137 8041 55171 8075
rect 55505 8041 55539 8075
rect 57437 8041 57471 8075
rect 59001 8041 59035 8075
rect 59369 8041 59403 8075
rect 6101 7973 6135 8007
rect 8769 7973 8803 8007
rect 14105 7973 14139 8007
rect 21465 7973 21499 8007
rect 24593 7973 24627 8007
rect 4353 7905 4387 7939
rect 7205 7905 7239 7939
rect 7573 7905 7607 7939
rect 7757 7905 7791 7939
rect 9137 7905 9171 7939
rect 9965 7905 9999 7939
rect 10425 7905 10459 7939
rect 10517 7905 10551 7939
rect 11253 7905 11287 7939
rect 11437 7905 11471 7939
rect 12909 7905 12943 7939
rect 15025 7905 15059 7939
rect 15853 7905 15887 7939
rect 16129 7905 16163 7939
rect 20913 7905 20947 7939
rect 21097 7905 21131 7939
rect 22293 7905 22327 7939
rect 22937 7905 22971 7939
rect 4077 7837 4111 7871
rect 7021 7837 7055 7871
rect 8401 7837 8435 7871
rect 10057 7837 10091 7871
rect 11069 7837 11103 7871
rect 12081 7837 12115 7871
rect 12817 7837 12851 7871
rect 15301 7837 15335 7871
rect 16313 7837 16347 7871
rect 17601 7837 17635 7871
rect 17877 7837 17911 7871
rect 19717 7837 19751 7871
rect 22109 7837 22143 7871
rect 12541 7769 12575 7803
rect 19993 7769 20027 7803
rect 24133 7769 24167 7803
rect 29193 7973 29227 8007
rect 29377 7973 29411 8007
rect 32965 7973 32999 8007
rect 34345 7973 34379 8007
rect 37933 7973 37967 8007
rect 41889 7973 41923 8007
rect 44189 7973 44223 8007
rect 24869 7905 24903 7939
rect 25973 7905 26007 7939
rect 26801 7905 26835 7939
rect 28825 7905 28859 7939
rect 29285 7905 29319 7939
rect 30573 7905 30607 7939
rect 32413 7905 32447 7939
rect 33885 7905 33919 7939
rect 35173 7905 35207 7939
rect 36001 7905 36035 7939
rect 36369 7905 36403 7939
rect 39221 7905 39255 7939
rect 39589 7905 39623 7939
rect 41429 7905 41463 7939
rect 44833 7905 44867 7939
rect 45201 7905 45235 7939
rect 45385 7905 45419 7939
rect 47317 7905 47351 7939
rect 47685 7905 47719 7939
rect 47777 7905 47811 7939
rect 25237 7837 25271 7871
rect 26525 7837 26559 7871
rect 28181 7837 28215 7871
rect 29009 7837 29043 7871
rect 29745 7837 29779 7871
rect 33793 7837 33827 7871
rect 35081 7837 35115 7871
rect 35909 7837 35943 7871
rect 36921 7837 36955 7871
rect 37381 7837 37415 7871
rect 38485 7837 38519 7871
rect 39313 7837 39347 7871
rect 39681 7837 39715 7871
rect 41337 7837 41371 7871
rect 42257 7837 42291 7871
rect 44741 7837 44775 7871
rect 47133 7837 47167 7871
rect 26249 7769 26283 7803
rect 30389 7769 30423 7803
rect 36369 7769 36403 7803
rect 36645 7769 36679 7803
rect 38669 7769 38703 7803
rect 40141 7769 40175 7803
rect 57529 7973 57563 8007
rect 61209 7973 61243 8007
rect 48973 7905 49007 7939
rect 49157 7905 49191 7939
rect 50353 7905 50387 7939
rect 52009 7905 52043 7939
rect 53297 7905 53331 7939
rect 56149 7905 56183 7939
rect 56333 7905 56367 7939
rect 56517 7905 56551 7939
rect 58173 7905 58207 7939
rect 58265 7905 58299 7939
rect 58541 7905 58575 7939
rect 58725 7905 58759 7939
rect 60473 7905 60507 7939
rect 60933 7905 60967 7939
rect 48513 7837 48547 7871
rect 49525 7837 49559 7871
rect 50721 7837 50755 7871
rect 51733 7837 51767 7871
rect 51917 7837 51951 7871
rect 50491 7769 50525 7803
rect 53481 7769 53515 7803
rect 55965 7769 55999 7803
rect 60289 7769 60323 7803
rect 5641 7701 5675 7735
rect 8033 7701 8067 7735
rect 10517 7701 10551 7735
rect 10793 7701 10827 7735
rect 13093 7701 13127 7735
rect 13645 7701 13679 7735
rect 14473 7701 14507 7735
rect 16681 7701 16715 7735
rect 21833 7701 21867 7735
rect 22477 7701 22511 7735
rect 23305 7701 23339 7735
rect 23765 7701 23799 7735
rect 24777 7701 24811 7735
rect 25007 7701 25041 7735
rect 25145 7701 25179 7735
rect 25513 7701 25547 7735
rect 28457 7701 28491 7735
rect 30757 7701 30791 7735
rect 31217 7701 31251 7735
rect 31493 7701 31527 7735
rect 40509 7701 40543 7735
rect 40877 7701 40911 7735
rect 42625 7701 42659 7735
rect 43085 7701 43119 7735
rect 46213 7701 46247 7735
rect 48053 7701 48087 7735
rect 48237 7701 48271 7735
rect 49893 7701 49927 7735
rect 50629 7701 50663 7735
rect 52193 7701 52227 7735
rect 53205 7701 53239 7735
rect 54769 7701 54803 7735
rect 56977 7701 57011 7735
rect 59829 7701 59863 7735
rect 4353 7497 4387 7531
rect 7113 7497 7147 7531
rect 11437 7497 11471 7531
rect 12633 7497 12667 7531
rect 12909 7497 12943 7531
rect 16865 7497 16899 7531
rect 18245 7497 18279 7531
rect 19257 7497 19291 7531
rect 23489 7497 23523 7531
rect 25053 7497 25087 7531
rect 25881 7497 25915 7531
rect 27261 7497 27295 7531
rect 28457 7497 28491 7531
rect 28733 7497 28767 7531
rect 30665 7497 30699 7531
rect 31033 7497 31067 7531
rect 33885 7497 33919 7531
rect 35173 7497 35207 7531
rect 41705 7497 41739 7531
rect 42073 7497 42107 7531
rect 44741 7497 44775 7531
rect 45477 7497 45511 7531
rect 47225 7497 47259 7531
rect 47593 7497 47627 7531
rect 50629 7497 50663 7531
rect 52653 7497 52687 7531
rect 53757 7497 53791 7531
rect 55229 7497 55263 7531
rect 56701 7497 56735 7531
rect 57069 7497 57103 7531
rect 61025 7497 61059 7531
rect 8769 7429 8803 7463
rect 5457 7361 5491 7395
rect 6285 7361 6319 7395
rect 9045 7361 9079 7395
rect 9781 7361 9815 7395
rect 10149 7361 10183 7395
rect 5733 7293 5767 7327
rect 5917 7293 5951 7327
rect 7297 7293 7331 7327
rect 7481 7293 7515 7327
rect 7803 7293 7837 7327
rect 7941 7293 7975 7327
rect 9873 7293 9907 7327
rect 12449 7293 12483 7327
rect 13369 7429 13403 7463
rect 13093 7361 13127 7395
rect 14105 7361 14139 7395
rect 15761 7361 15795 7395
rect 24961 7361 24995 7395
rect 14013 7293 14047 7327
rect 14381 7293 14415 7327
rect 16589 7293 16623 7327
rect 16681 7293 16715 7327
rect 19441 7293 19475 7327
rect 19625 7293 19659 7327
rect 19993 7293 20027 7327
rect 20177 7293 20211 7327
rect 20453 7293 20487 7327
rect 21189 7293 21223 7327
rect 21833 7293 21867 7327
rect 22477 7293 22511 7327
rect 23029 7293 23063 7327
rect 24317 7293 24351 7327
rect 24409 7293 24443 7327
rect 24501 7293 24535 7327
rect 4905 7225 4939 7259
rect 8309 7225 8343 7259
rect 12909 7225 12943 7259
rect 17877 7225 17911 7259
rect 21005 7225 21039 7259
rect 22201 7225 22235 7259
rect 26525 7361 26559 7395
rect 26433 7293 26467 7327
rect 26801 7293 26835 7327
rect 26893 7293 26927 7327
rect 27629 7293 27663 7327
rect 27997 7293 28031 7327
rect 32781 7429 32815 7463
rect 38853 7429 38887 7463
rect 46489 7429 46523 7463
rect 34253 7361 34287 7395
rect 34713 7361 34747 7395
rect 35725 7361 35759 7395
rect 44005 7361 44039 7395
rect 44373 7361 44407 7395
rect 46360 7361 46394 7395
rect 46581 7361 46615 7395
rect 49893 7361 49927 7395
rect 53021 7429 53055 7463
rect 59737 7429 59771 7463
rect 52285 7361 52319 7395
rect 56057 7361 56091 7395
rect 57529 7361 57563 7395
rect 29469 7293 29503 7327
rect 30297 7293 30331 7327
rect 30849 7293 30883 7327
rect 31401 7293 31435 7327
rect 32597 7293 32631 7327
rect 33609 7293 33643 7327
rect 33701 7293 33735 7327
rect 34897 7293 34931 7327
rect 34989 7293 35023 7327
rect 36829 7293 36863 7327
rect 37013 7293 37047 7327
rect 37381 7293 37415 7327
rect 38485 7293 38519 7327
rect 39037 7293 39071 7327
rect 39221 7293 39255 7327
rect 39405 7293 39439 7327
rect 40233 7293 40267 7327
rect 40693 7293 40727 7327
rect 41337 7293 41371 7327
rect 42349 7293 42383 7327
rect 42625 7293 42659 7327
rect 44833 7293 44867 7327
rect 49985 7293 50019 7327
rect 50353 7293 50387 7327
rect 50537 7293 50571 7327
rect 50629 7293 50663 7327
rect 51733 7293 51767 7327
rect 52837 7293 52871 7327
rect 53389 7293 53423 7327
rect 53941 7293 53975 7327
rect 55597 7293 55631 7327
rect 55781 7293 55815 7327
rect 56241 7293 56275 7327
rect 57621 7293 57655 7327
rect 58081 7293 58115 7327
rect 58173 7293 58207 7327
rect 59461 7293 59495 7327
rect 59645 7293 59679 7327
rect 60197 7293 60231 7327
rect 60657 7293 60691 7327
rect 27813 7225 27847 7259
rect 28457 7225 28491 7259
rect 29285 7225 29319 7259
rect 29561 7225 29595 7259
rect 29653 7225 29687 7259
rect 30021 7225 30055 7259
rect 38025 7225 38059 7259
rect 40509 7225 40543 7259
rect 41061 7225 41095 7259
rect 45753 7225 45787 7259
rect 46213 7225 46247 7259
rect 46949 7225 46983 7259
rect 47777 7225 47811 7259
rect 47961 7225 47995 7259
rect 48145 7225 48179 7259
rect 48513 7225 48547 7259
rect 48789 7225 48823 7259
rect 49157 7225 49191 7259
rect 49341 7225 49375 7259
rect 50813 7225 50847 7259
rect 54493 7225 54527 7259
rect 58725 7225 58759 7259
rect 3709 7157 3743 7191
rect 3985 7157 4019 7191
rect 4721 7157 4755 7191
rect 6561 7157 6595 7191
rect 11897 7157 11931 7191
rect 12265 7157 12299 7191
rect 16221 7157 16255 7191
rect 17417 7157 17451 7191
rect 18797 7157 18831 7191
rect 20821 7157 20855 7191
rect 21281 7157 21315 7191
rect 22661 7157 22695 7191
rect 23949 7157 23983 7191
rect 25053 7157 25087 7191
rect 25329 7157 25363 7191
rect 25697 7157 25731 7191
rect 28089 7157 28123 7191
rect 29009 7157 29043 7191
rect 31769 7157 31803 7191
rect 32413 7157 32447 7191
rect 33241 7157 33275 7191
rect 36093 7157 36127 7191
rect 36645 7157 36679 7191
rect 39865 7157 39899 7191
rect 45017 7157 45051 7191
rect 48053 7157 48087 7191
rect 51273 7157 51307 7191
rect 51917 7157 51951 7191
rect 54125 7157 54159 7191
rect 59093 7157 59127 7191
rect 6469 6953 6503 6987
rect 6837 6953 6871 6987
rect 7941 6953 7975 6987
rect 9965 6953 9999 6987
rect 12357 6953 12391 6987
rect 12725 6953 12759 6987
rect 17601 6953 17635 6987
rect 17877 6953 17911 6987
rect 23213 6953 23247 6987
rect 23581 6953 23615 6987
rect 31217 6953 31251 6987
rect 32321 6953 32355 6987
rect 39681 6953 39715 6987
rect 46397 6953 46431 6987
rect 47501 6953 47535 6987
rect 51549 6953 51583 6987
rect 55137 6953 55171 6987
rect 5733 6885 5767 6919
rect 6101 6885 6135 6919
rect 6561 6885 6595 6919
rect 6745 6885 6779 6919
rect 6929 6885 6963 6919
rect 13185 6885 13219 6919
rect 16313 6885 16347 6919
rect 7297 6817 7331 6851
rect 8217 6817 8251 6851
rect 9505 6817 9539 6851
rect 13829 6817 13863 6851
rect 14197 6817 14231 6851
rect 14381 6817 14415 6851
rect 15025 6817 15059 6851
rect 16957 6817 16991 6851
rect 17325 6817 17359 6851
rect 17509 6817 17543 6851
rect 4077 6749 4111 6783
rect 4353 6749 4387 6783
rect 8125 6749 8159 6783
rect 8677 6749 8711 6783
rect 10057 6749 10091 6783
rect 10333 6749 10367 6783
rect 11713 6749 11747 6783
rect 13737 6749 13771 6783
rect 14749 6749 14783 6783
rect 15853 6749 15887 6783
rect 17049 6749 17083 6783
rect 18337 6885 18371 6919
rect 20913 6885 20947 6919
rect 36553 6885 36587 6919
rect 40785 6885 40819 6919
rect 43729 6885 43763 6919
rect 18981 6817 19015 6851
rect 19073 6817 19107 6851
rect 19315 6817 19349 6851
rect 19533 6817 19567 6851
rect 21097 6817 21131 6851
rect 22109 6817 22143 6851
rect 22569 6817 22603 6851
rect 22661 6817 22695 6851
rect 23765 6817 23799 6851
rect 25053 6817 25087 6851
rect 25145 6817 25179 6851
rect 26709 6817 26743 6851
rect 26801 6817 26835 6851
rect 27169 6817 27203 6851
rect 27349 6817 27383 6851
rect 28641 6817 28675 6851
rect 28825 6817 28859 6851
rect 29469 6817 29503 6851
rect 29745 6817 29779 6851
rect 30481 6817 30515 6851
rect 30665 6817 30699 6851
rect 32137 6817 32171 6851
rect 36134 6817 36168 6851
rect 36921 6817 36955 6851
rect 38393 6817 38427 6851
rect 38761 6817 38795 6851
rect 39957 6817 39991 6851
rect 40049 6817 40083 6851
rect 41153 6817 41187 6851
rect 41613 6817 41647 6851
rect 41705 6817 41739 6851
rect 42901 6817 42935 6851
rect 44281 6817 44315 6851
rect 45109 6817 45143 6851
rect 21465 6749 21499 6783
rect 21833 6749 21867 6783
rect 25605 6749 25639 6783
rect 25973 6749 26007 6783
rect 26341 6749 26375 6783
rect 33517 6749 33551 6783
rect 33793 6749 33827 6783
rect 34897 6749 34931 6783
rect 36001 6749 36035 6783
rect 37289 6749 37323 6783
rect 38025 6749 38059 6783
rect 38945 6749 38979 6783
rect 42165 6749 42199 6783
rect 44373 6749 44407 6783
rect 45201 6749 45235 6783
rect 45569 6749 45603 6783
rect 24777 6681 24811 6715
rect 27629 6681 27663 6715
rect 28917 6681 28951 6715
rect 30205 6681 30239 6715
rect 39221 6681 39255 6715
rect 47869 6885 47903 6919
rect 46489 6817 46523 6851
rect 48605 6817 48639 6851
rect 49801 6817 49835 6851
rect 50077 6817 50111 6851
rect 54861 6885 54895 6919
rect 60749 6885 60783 6919
rect 52285 6817 52319 6851
rect 52469 6817 52503 6851
rect 53665 6817 53699 6851
rect 54953 6817 54987 6851
rect 56149 6817 56183 6851
rect 56241 6817 56275 6851
rect 56333 6817 56367 6851
rect 56793 6817 56827 6851
rect 57529 6817 57563 6851
rect 58449 6817 58483 6851
rect 59277 6817 59311 6851
rect 59921 6817 59955 6851
rect 60289 6817 60323 6851
rect 61117 6817 61151 6851
rect 61669 6817 61703 6851
rect 46857 6749 46891 6783
rect 47225 6749 47259 6783
rect 48237 6749 48271 6783
rect 51457 6749 51491 6783
rect 51549 6749 51583 6783
rect 51733 6749 51767 6783
rect 52193 6749 52227 6783
rect 52837 6749 52871 6783
rect 55505 6749 55539 6783
rect 57069 6749 57103 6783
rect 57621 6749 57655 6783
rect 58173 6749 58207 6783
rect 58633 6749 58667 6783
rect 58909 6749 58943 6783
rect 60197 6749 60231 6783
rect 61393 6749 61427 6783
rect 61577 6749 61611 6783
rect 46765 6681 46799 6715
rect 3249 6613 3283 6647
rect 3525 6613 3559 6647
rect 8953 6613 8987 6647
rect 13093 6613 13127 6647
rect 16129 6613 16163 6647
rect 17601 6613 17635 6647
rect 18245 6613 18279 6647
rect 20177 6613 20211 6647
rect 20637 6613 20671 6647
rect 22845 6613 22879 6647
rect 23949 6613 23983 6647
rect 24317 6613 24351 6647
rect 24869 6613 24903 6647
rect 28273 6613 28307 6647
rect 30849 6613 30883 6647
rect 31953 6613 31987 6647
rect 32689 6613 32723 6647
rect 33057 6613 33091 6647
rect 35633 6613 35667 6647
rect 39773 6613 39807 6647
rect 40233 6613 40267 6647
rect 41429 6613 41463 6647
rect 42533 6613 42567 6647
rect 44097 6613 44131 6647
rect 46213 6613 46247 6647
rect 46397 6613 46431 6647
rect 46654 6613 46688 6647
rect 49157 6613 49191 6647
rect 49617 6613 49651 6647
rect 53297 6613 53331 6647
rect 54033 6613 54067 6647
rect 55873 6613 55907 6647
rect 61853 6613 61887 6647
rect 5181 6409 5215 6443
rect 6285 6409 6319 6443
rect 8493 6409 8527 6443
rect 11713 6409 11747 6443
rect 13185 6409 13219 6443
rect 33885 6409 33919 6443
rect 34437 6409 34471 6443
rect 34713 6409 34747 6443
rect 41981 6409 42015 6443
rect 43361 6409 43395 6443
rect 45017 6409 45051 6443
rect 45293 6409 45327 6443
rect 45569 6409 45603 6443
rect 47961 6409 47995 6443
rect 48881 6409 48915 6443
rect 50445 6409 50479 6443
rect 50997 6409 51031 6443
rect 54585 6409 54619 6443
rect 54953 6409 54987 6443
rect 55413 6409 55447 6443
rect 57161 6409 57195 6443
rect 59461 6409 59495 6443
rect 4813 6341 4847 6375
rect 9137 6341 9171 6375
rect 3525 6273 3559 6307
rect 5917 6273 5951 6307
rect 7757 6273 7791 6307
rect 8217 6273 8251 6307
rect 10149 6273 10183 6307
rect 10793 6273 10827 6307
rect 10977 6273 11011 6307
rect 3249 6205 3283 6239
rect 7021 6205 7055 6239
rect 8309 6205 8343 6239
rect 9597 6205 9631 6239
rect 9689 6205 9723 6239
rect 11069 6205 11103 6239
rect 11529 6205 11563 6239
rect 6561 6137 6595 6171
rect 6837 6137 6871 6171
rect 9413 6137 9447 6171
rect 10425 6137 10459 6171
rect 14473 6341 14507 6375
rect 17877 6341 17911 6375
rect 19165 6341 19199 6375
rect 19349 6341 19383 6375
rect 19993 6341 20027 6375
rect 23949 6341 23983 6375
rect 24409 6341 24443 6375
rect 11805 6273 11839 6307
rect 13553 6273 13587 6307
rect 16221 6273 16255 6307
rect 18613 6273 18647 6307
rect 34897 6341 34931 6375
rect 37933 6341 37967 6375
rect 39589 6341 39623 6375
rect 19809 6273 19843 6307
rect 22753 6273 22787 6307
rect 24501 6273 24535 6307
rect 25053 6273 25087 6307
rect 26341 6273 26375 6307
rect 28733 6273 28767 6307
rect 29561 6273 29595 6307
rect 32229 6273 32263 6307
rect 33241 6273 33275 6307
rect 34437 6273 34471 6307
rect 37105 6273 37139 6307
rect 39405 6273 39439 6307
rect 14657 6205 14691 6239
rect 15025 6205 15059 6239
rect 15117 6205 15151 6239
rect 15853 6205 15887 6239
rect 16129 6205 16163 6239
rect 16819 6205 16853 6239
rect 16957 6205 16991 6239
rect 18889 6205 18923 6239
rect 19073 6205 19107 6239
rect 19165 6205 19199 6239
rect 20085 6205 20119 6239
rect 20545 6205 20579 6239
rect 21097 6205 21131 6239
rect 21649 6205 21683 6239
rect 22293 6205 22327 6239
rect 23121 6205 23155 6239
rect 25329 6205 25363 6239
rect 25513 6205 25547 6239
rect 25789 6205 25823 6239
rect 26893 6205 26927 6239
rect 27169 6205 27203 6239
rect 27353 6205 27387 6239
rect 27445 6205 27479 6239
rect 28181 6205 28215 6239
rect 29285 6205 29319 6239
rect 31309 6205 31343 6239
rect 31769 6205 31803 6239
rect 31861 6205 31895 6239
rect 32045 6205 32079 6239
rect 33701 6205 33735 6239
rect 34253 6205 34287 6239
rect 35633 6205 35667 6239
rect 36001 6205 36035 6239
rect 36185 6205 36219 6239
rect 36553 6205 36587 6239
rect 37749 6205 37783 6239
rect 38301 6205 38335 6239
rect 38669 6205 38703 6239
rect 38853 6205 38887 6239
rect 39037 6205 39071 6239
rect 18061 6137 18095 6171
rect 21465 6137 21499 6171
rect 43913 6273 43947 6307
rect 44925 6273 44959 6307
rect 45017 6273 45051 6307
rect 47041 6341 47075 6375
rect 40693 6205 40727 6239
rect 41337 6205 41371 6239
rect 41797 6205 41831 6239
rect 42455 6205 42489 6239
rect 42625 6205 42659 6239
rect 42901 6205 42935 6239
rect 43085 6205 43119 6239
rect 44465 6205 44499 6239
rect 44741 6205 44775 6239
rect 46213 6205 46247 6239
rect 46489 6205 46523 6239
rect 47501 6341 47535 6375
rect 47593 6341 47627 6375
rect 51181 6341 51215 6375
rect 55229 6341 55263 6375
rect 55689 6341 55723 6375
rect 48329 6273 48363 6307
rect 49893 6273 49927 6307
rect 50997 6273 51031 6307
rect 53297 6273 53331 6307
rect 47501 6205 47535 6239
rect 47777 6205 47811 6239
rect 49065 6205 49099 6239
rect 49801 6205 49835 6239
rect 51917 6205 51951 6239
rect 53021 6205 53055 6239
rect 28273 6137 28307 6171
rect 29101 6137 29135 6171
rect 30941 6137 30975 6171
rect 35265 6137 35299 6171
rect 37473 6137 37507 6171
rect 39589 6137 39623 6171
rect 39681 6137 39715 6171
rect 40509 6137 40543 6171
rect 41061 6137 41095 6171
rect 43729 6137 43763 6171
rect 46397 6137 46431 6171
rect 46949 6137 46983 6171
rect 47041 6137 47075 6171
rect 52469 6137 52503 6171
rect 56425 6273 56459 6307
rect 60565 6273 60599 6307
rect 61117 6273 61151 6307
rect 56057 6205 56091 6239
rect 56701 6205 56735 6239
rect 58081 6205 58115 6239
rect 58357 6205 58391 6239
rect 60657 6205 60691 6239
rect 61945 6205 61979 6239
rect 55873 6137 55907 6171
rect 2605 6069 2639 6103
rect 2973 6069 3007 6103
rect 7113 6069 7147 6103
rect 8125 6069 8159 6103
rect 11713 6069 11747 6103
rect 12265 6069 12299 6103
rect 12817 6069 12851 6103
rect 13921 6069 13955 6103
rect 15577 6069 15611 6103
rect 17417 6069 17451 6103
rect 21741 6069 21775 6103
rect 23489 6069 23523 6103
rect 26249 6069 26283 6103
rect 27445 6069 27479 6103
rect 27629 6069 27663 6103
rect 27997 6069 28031 6103
rect 31585 6069 31619 6103
rect 32781 6069 32815 6103
rect 33517 6069 33551 6103
rect 40233 6069 40267 6103
rect 47225 6069 47259 6103
rect 49157 6069 49191 6103
rect 50813 6069 50847 6103
rect 52101 6069 52135 6103
rect 52837 6069 52871 6103
rect 55229 6069 55263 6103
rect 57529 6069 57563 6103
rect 57989 6069 58023 6103
rect 60013 6069 60047 6103
rect 60381 6069 60415 6103
rect 61577 6069 61611 6103
rect 5641 5865 5675 5899
rect 9413 5865 9447 5899
rect 16957 5865 16991 5899
rect 20729 5865 20763 5899
rect 22477 5865 22511 5899
rect 23121 5865 23155 5899
rect 23673 5865 23707 5899
rect 27261 5865 27295 5899
rect 31309 5865 31343 5899
rect 41613 5865 41647 5899
rect 42073 5865 42107 5899
rect 42625 5865 42659 5899
rect 42993 5865 43027 5899
rect 49157 5865 49191 5899
rect 49985 5865 50019 5899
rect 57069 5865 57103 5899
rect 58817 5865 58851 5899
rect 4261 5797 4295 5831
rect 6653 5797 6687 5831
rect 7849 5797 7883 5831
rect 12081 5797 12115 5831
rect 17509 5797 17543 5831
rect 18981 5797 19015 5831
rect 19165 5797 19199 5831
rect 19441 5797 19475 5831
rect 19993 5797 20027 5831
rect 21189 5797 21223 5831
rect 22753 5797 22787 5831
rect 25513 5797 25547 5831
rect 25881 5797 25915 5831
rect 26341 5797 26375 5831
rect 26617 5797 26651 5831
rect 28641 5797 28675 5831
rect 2697 5729 2731 5763
rect 3157 5729 3191 5763
rect 5089 5729 5123 5763
rect 5273 5729 5307 5763
rect 6101 5729 6135 5763
rect 7389 5729 7423 5763
rect 9781 5729 9815 5763
rect 10517 5729 10551 5763
rect 11621 5729 11655 5763
rect 13553 5729 13587 5763
rect 14105 5729 14139 5763
rect 15945 5729 15979 5763
rect 16313 5729 16347 5763
rect 16497 5729 16531 5763
rect 18245 5729 18279 5763
rect 18337 5729 18371 5763
rect 2605 5661 2639 5695
rect 4813 5661 4847 5695
rect 7297 5661 7331 5695
rect 9689 5661 9723 5695
rect 11529 5661 11563 5695
rect 14197 5661 14231 5695
rect 15577 5661 15611 5695
rect 17417 5661 17451 5695
rect 18521 5661 18555 5695
rect 6285 5593 6319 5627
rect 8309 5593 8343 5627
rect 11069 5593 11103 5627
rect 13093 5593 13127 5627
rect 14105 5593 14139 5627
rect 14749 5593 14783 5627
rect 19533 5729 19567 5763
rect 20269 5729 20303 5763
rect 21557 5729 21591 5763
rect 21649 5729 21683 5763
rect 22937 5729 22971 5763
rect 24133 5729 24167 5763
rect 24409 5729 24443 5763
rect 28549 5729 28583 5763
rect 28917 5729 28951 5763
rect 29469 5729 29503 5763
rect 29561 5729 29595 5763
rect 30021 5729 30055 5763
rect 31033 5729 31067 5763
rect 24869 5661 24903 5695
rect 25145 5661 25179 5695
rect 26764 5661 26798 5695
rect 26985 5661 27019 5695
rect 33057 5797 33091 5831
rect 33885 5797 33919 5831
rect 34345 5797 34379 5831
rect 38393 5797 38427 5831
rect 42809 5797 42843 5831
rect 43453 5797 43487 5831
rect 44005 5797 44039 5831
rect 53849 5797 53883 5831
rect 55045 5797 55079 5831
rect 56609 5797 56643 5831
rect 32137 5729 32171 5763
rect 33241 5729 33275 5763
rect 34897 5729 34931 5763
rect 34989 5729 35023 5763
rect 35173 5729 35207 5763
rect 35357 5729 35391 5763
rect 35633 5729 35667 5763
rect 36645 5729 36679 5763
rect 37473 5729 37507 5763
rect 37749 5729 37783 5763
rect 41797 5729 41831 5763
rect 41981 5729 42015 5763
rect 31493 5661 31527 5695
rect 39313 5661 39347 5695
rect 39589 5661 39623 5695
rect 40693 5661 40727 5695
rect 43637 5729 43671 5763
rect 44281 5729 44315 5763
rect 45017 5729 45051 5763
rect 45109 5729 45143 5763
rect 45845 5729 45879 5763
rect 46673 5729 46707 5763
rect 47133 5729 47167 5763
rect 48973 5729 49007 5763
rect 49525 5729 49559 5763
rect 50261 5729 50295 5763
rect 50905 5729 50939 5763
rect 53021 5729 53055 5763
rect 53389 5729 53423 5763
rect 54217 5729 54251 5763
rect 54585 5729 54619 5763
rect 55597 5729 55631 5763
rect 57713 5729 57747 5763
rect 57989 5729 58023 5763
rect 59001 5729 59035 5763
rect 60197 5729 60231 5763
rect 46765 5661 46799 5695
rect 48145 5661 48179 5695
rect 53481 5661 53515 5695
rect 55965 5661 55999 5695
rect 57161 5661 57195 5695
rect 58173 5661 58207 5695
rect 58449 5661 58483 5695
rect 60473 5661 60507 5695
rect 24225 5593 24259 5627
rect 30941 5593 30975 5627
rect 31309 5593 31343 5627
rect 32321 5593 32355 5627
rect 37105 5593 37139 5627
rect 42809 5593 42843 5627
rect 44649 5593 44683 5627
rect 44833 5593 44867 5627
rect 48789 5593 48823 5627
rect 52285 5593 52319 5627
rect 52837 5593 52871 5627
rect 55762 5593 55796 5627
rect 2421 5525 2455 5559
rect 3525 5525 3559 5559
rect 3801 5525 3835 5559
rect 5917 5525 5951 5559
rect 7021 5525 7055 5559
rect 8769 5525 8803 5559
rect 9965 5525 9999 5559
rect 12357 5525 12391 5559
rect 12817 5525 12851 5559
rect 15117 5525 15151 5559
rect 18521 5525 18555 5559
rect 18797 5525 18831 5559
rect 18981 5525 19015 5559
rect 19257 5525 19291 5559
rect 21373 5525 21407 5559
rect 21833 5525 21867 5559
rect 23949 5525 23983 5559
rect 26893 5525 26927 5559
rect 27813 5525 27847 5559
rect 30481 5525 30515 5559
rect 31125 5525 31159 5559
rect 31861 5525 31895 5559
rect 32689 5525 32723 5559
rect 33425 5525 33459 5559
rect 34253 5525 34287 5559
rect 36093 5525 36127 5559
rect 36461 5525 36495 5559
rect 36737 5525 36771 5559
rect 37933 5525 37967 5559
rect 38761 5525 38795 5559
rect 39221 5525 39255 5559
rect 41337 5525 41371 5559
rect 45293 5525 45327 5559
rect 46213 5525 46247 5559
rect 47501 5525 47535 5559
rect 47869 5525 47903 5559
rect 50353 5525 50387 5559
rect 51365 5525 51399 5559
rect 51733 5525 51767 5559
rect 54677 5525 54711 5559
rect 55505 5525 55539 5559
rect 55873 5525 55907 5559
rect 56241 5525 56275 5559
rect 59185 5525 59219 5559
rect 59553 5525 59587 5559
rect 59921 5525 59955 5559
rect 61761 5525 61795 5559
rect 2329 5321 2363 5355
rect 14473 5321 14507 5355
rect 16405 5321 16439 5355
rect 18061 5321 18095 5355
rect 18889 5321 18923 5355
rect 19073 5321 19107 5355
rect 24041 5321 24075 5355
rect 24225 5321 24259 5355
rect 32229 5321 32263 5355
rect 34437 5321 34471 5355
rect 35633 5321 35667 5355
rect 36001 5321 36035 5355
rect 39405 5321 39439 5355
rect 39589 5321 39623 5355
rect 39957 5321 39991 5355
rect 41429 5321 41463 5355
rect 41797 5321 41831 5355
rect 42717 5321 42751 5355
rect 43085 5321 43119 5355
rect 43545 5321 43579 5355
rect 44281 5321 44315 5355
rect 44925 5321 44959 5355
rect 45845 5321 45879 5355
rect 48973 5321 49007 5355
rect 51273 5321 51307 5355
rect 52377 5321 52411 5355
rect 54309 5321 54343 5355
rect 55965 5321 55999 5355
rect 58909 5321 58943 5355
rect 61485 5321 61519 5355
rect 4997 5253 5031 5287
rect 5273 5253 5307 5287
rect 6193 5253 6227 5287
rect 7849 5253 7883 5287
rect 8309 5253 8343 5287
rect 11897 5253 11931 5287
rect 14841 5253 14875 5287
rect 17417 5253 17451 5287
rect 7205 5185 7239 5219
rect 9413 5185 9447 5219
rect 10885 5185 10919 5219
rect 12449 5185 12483 5219
rect 12725 5185 12759 5219
rect 14933 5185 14967 5219
rect 15669 5185 15703 5219
rect 18797 5185 18831 5219
rect 18889 5185 18923 5219
rect 19441 5185 19475 5219
rect 21281 5185 21315 5219
rect 23121 5185 23155 5219
rect 2973 5117 3007 5151
rect 3249 5117 3283 5151
rect 5641 5117 5675 5151
rect 7021 5117 7055 5151
rect 7573 5117 7607 5151
rect 8493 5117 8527 5151
rect 9321 5117 9355 5151
rect 10333 5117 10367 5151
rect 10425 5117 10459 5151
rect 11621 5117 11655 5151
rect 15577 5117 15611 5151
rect 15945 5117 15979 5151
rect 16037 5117 16071 5151
rect 16773 5117 16807 5151
rect 18337 5117 18371 5151
rect 19625 5117 19659 5151
rect 20913 5117 20947 5151
rect 21465 5117 21499 5151
rect 21925 5117 21959 5151
rect 22477 5117 22511 5151
rect 23397 5117 23431 5151
rect 23673 5117 23707 5151
rect 8585 5049 8619 5083
rect 11161 5049 11195 5083
rect 14105 5049 14139 5083
rect 18245 5049 18279 5083
rect 24685 5253 24719 5287
rect 26893 5253 26927 5287
rect 28733 5253 28767 5287
rect 31217 5253 31251 5287
rect 2697 4981 2731 5015
rect 4537 4981 4571 5015
rect 5825 4981 5859 5015
rect 6653 4981 6687 5015
rect 9873 4981 9907 5015
rect 10241 4981 10275 5015
rect 17785 4981 17819 5015
rect 19809 4981 19843 5015
rect 20269 4981 20303 5015
rect 20821 4981 20855 5015
rect 22293 4981 22327 5015
rect 22661 4981 22695 5015
rect 23857 4981 23891 5015
rect 24041 4981 24075 5015
rect 24501 5185 24535 5219
rect 25053 5185 25087 5219
rect 26433 5185 26467 5219
rect 27261 5185 27295 5219
rect 24777 5117 24811 5151
rect 27813 5117 27847 5151
rect 28089 5117 28123 5151
rect 28273 5117 28307 5151
rect 29285 5117 29319 5151
rect 29837 5117 29871 5151
rect 29929 5117 29963 5151
rect 30113 5117 30147 5151
rect 30297 5117 30331 5151
rect 30665 5117 30699 5151
rect 29009 5049 29043 5083
rect 35265 5253 35299 5287
rect 35449 5253 35483 5287
rect 31401 5117 31435 5151
rect 31585 5117 31619 5151
rect 32689 5117 32723 5151
rect 32965 5117 32999 5151
rect 33701 5117 33735 5151
rect 34253 5117 34287 5151
rect 34437 5117 34471 5151
rect 34713 5117 34747 5151
rect 35081 5117 35115 5151
rect 32505 5049 32539 5083
rect 36185 5117 36219 5151
rect 36369 5117 36403 5151
rect 38025 5117 38059 5151
rect 38393 5117 38427 5151
rect 38761 5117 38795 5151
rect 38945 5117 38979 5151
rect 36737 5049 36771 5083
rect 40785 5253 40819 5287
rect 43913 5253 43947 5287
rect 46305 5253 46339 5287
rect 53389 5253 53423 5287
rect 41153 5185 41187 5219
rect 41429 5185 41463 5219
rect 45569 5185 45603 5219
rect 49157 5185 49191 5219
rect 49617 5185 49651 5219
rect 50537 5185 50571 5219
rect 57989 5185 58023 5219
rect 40601 5117 40635 5151
rect 41981 5117 42015 5151
rect 42441 5117 42475 5151
rect 43361 5117 43395 5151
rect 44465 5117 44499 5151
rect 44741 5117 44775 5151
rect 46489 5117 46523 5151
rect 47225 5117 47259 5151
rect 47501 5117 47535 5151
rect 48237 5117 48271 5151
rect 49341 5117 49375 5151
rect 49709 5117 49743 5151
rect 50905 5117 50939 5151
rect 52653 5117 52687 5151
rect 52929 5117 52963 5151
rect 53389 5117 53423 5151
rect 53941 5117 53975 5151
rect 55137 5117 55171 5151
rect 55413 5117 55447 5151
rect 55597 5117 55631 5151
rect 56793 5117 56827 5151
rect 57345 5117 57379 5151
rect 57437 5117 57471 5151
rect 57621 5117 57655 5151
rect 58357 5117 58391 5151
rect 59093 5117 59127 5151
rect 59277 5117 59311 5151
rect 59737 5117 59771 5151
rect 59829 5117 59863 5151
rect 44649 5049 44683 5083
rect 54585 5049 54619 5083
rect 24501 4981 24535 5015
rect 31033 4981 31067 5015
rect 31217 4981 31251 5015
rect 31769 4981 31803 5015
rect 32781 4981 32815 5015
rect 32965 4981 32999 5015
rect 33241 4981 33275 5015
rect 33609 4981 33643 5015
rect 33885 4981 33919 5015
rect 35449 4981 35483 5015
rect 37013 4981 37047 5015
rect 37381 4981 37415 5015
rect 39221 4981 39255 5015
rect 39405 4981 39439 5015
rect 41613 4981 41647 5015
rect 46581 4981 46615 5015
rect 47869 4981 47903 5015
rect 50169 4981 50203 5015
rect 51917 4981 51951 5015
rect 56333 4981 56367 5015
rect 57069 4981 57103 5015
rect 60289 4981 60323 5015
rect 60749 4981 60783 5015
rect 61117 4981 61151 5015
rect 6469 4777 6503 4811
rect 7665 4777 7699 4811
rect 8309 4777 8343 4811
rect 14933 4777 14967 4811
rect 15945 4777 15979 4811
rect 17877 4777 17911 4811
rect 19441 4777 19475 4811
rect 19625 4777 19659 4811
rect 24041 4777 24075 4811
rect 24409 4777 24443 4811
rect 24869 4777 24903 4811
rect 38853 4777 38887 4811
rect 2605 4709 2639 4743
rect 4077 4709 4111 4743
rect 8493 4709 8527 4743
rect 10793 4709 10827 4743
rect 2789 4641 2823 4675
rect 4537 4641 4571 4675
rect 4721 4641 4755 4675
rect 4905 4641 4939 4675
rect 5365 4641 5399 4675
rect 7021 4641 7055 4675
rect 7389 4641 7423 4675
rect 7665 4641 7699 4675
rect 8401 4641 8435 4675
rect 9873 4641 9907 4675
rect 10057 4641 10091 4675
rect 11621 4641 11655 4675
rect 11805 4641 11839 4675
rect 12817 4641 12851 4675
rect 13277 4641 13311 4675
rect 13737 4641 13771 4675
rect 15301 4641 15335 4675
rect 16589 4641 16623 4675
rect 17049 4641 17083 4675
rect 18245 4641 18279 4675
rect 18429 4641 18463 4675
rect 18613 4641 18647 4675
rect 18705 4641 18739 4675
rect 3157 4573 3191 4607
rect 7113 4573 7147 4607
rect 7297 4573 7331 4607
rect 8953 4573 8987 4607
rect 9505 4573 9539 4607
rect 10425 4573 10459 4607
rect 14013 4573 14047 4607
rect 17417 4573 17451 4607
rect 19165 4573 19199 4607
rect 10222 4505 10256 4539
rect 13093 4505 13127 4539
rect 16773 4505 16807 4539
rect 29837 4709 29871 4743
rect 31585 4709 31619 4743
rect 31769 4709 31803 4743
rect 34161 4709 34195 4743
rect 20913 4641 20947 4675
rect 21189 4641 21223 4675
rect 22385 4641 22419 4675
rect 22477 4641 22511 4675
rect 22661 4641 22695 4675
rect 23857 4641 23891 4675
rect 25145 4641 25179 4675
rect 25329 4641 25363 4675
rect 25881 4641 25915 4675
rect 26893 4641 26927 4675
rect 27169 4641 27203 4675
rect 27445 4641 27479 4675
rect 27997 4641 28031 4675
rect 28457 4641 28491 4675
rect 29377 4641 29411 4675
rect 29929 4641 29963 4675
rect 21005 4573 21039 4607
rect 21373 4573 21407 4607
rect 32965 4641 32999 4675
rect 33701 4641 33735 4675
rect 34621 4641 34655 4675
rect 34805 4641 34839 4675
rect 34989 4641 35023 4675
rect 35265 4641 35299 4675
rect 35449 4641 35483 4675
rect 36461 4641 36495 4675
rect 37933 4641 37967 4675
rect 38761 4641 38795 4675
rect 28825 4573 28859 4607
rect 31401 4573 31435 4607
rect 31585 4573 31619 4607
rect 35909 4573 35943 4607
rect 37013 4573 37047 4607
rect 26525 4505 26559 4539
rect 32413 4505 32447 4539
rect 32873 4505 32907 4539
rect 33149 4505 33183 4539
rect 36277 4505 36311 4539
rect 36645 4505 36679 4539
rect 38117 4505 38151 4539
rect 38945 4777 38979 4811
rect 48697 4777 48731 4811
rect 49801 4777 49835 4811
rect 57345 4777 57379 4811
rect 58081 4777 58115 4811
rect 39221 4709 39255 4743
rect 42533 4709 42567 4743
rect 43177 4709 43211 4743
rect 47133 4709 47167 4743
rect 47501 4709 47535 4743
rect 50169 4709 50203 4743
rect 50997 4709 51031 4743
rect 51549 4709 51583 4743
rect 52285 4709 52319 4743
rect 53941 4709 53975 4743
rect 55413 4709 55447 4743
rect 58265 4709 58299 4743
rect 39865 4641 39899 4675
rect 40233 4641 40267 4675
rect 40417 4641 40451 4675
rect 41245 4641 41279 4675
rect 41705 4641 41739 4675
rect 41889 4641 41923 4675
rect 42073 4641 42107 4675
rect 44005 4641 44039 4675
rect 44741 4641 44775 4675
rect 45753 4641 45787 4675
rect 46121 4641 46155 4675
rect 46305 4641 46339 4675
rect 47317 4641 47351 4675
rect 47409 4641 47443 4675
rect 50261 4641 50295 4675
rect 50721 4641 50755 4675
rect 53113 4641 53147 4675
rect 53297 4641 53331 4675
rect 54585 4641 54619 4675
rect 59093 4641 59127 4675
rect 59921 4641 59955 4675
rect 61025 4641 61059 4675
rect 61209 4641 61243 4675
rect 38945 4573 38979 4607
rect 39957 4573 39991 4607
rect 41061 4573 41095 4607
rect 45661 4573 45695 4607
rect 46949 4573 46983 4607
rect 47869 4573 47903 4607
rect 49985 4573 50019 4607
rect 51917 4573 51951 4607
rect 53665 4573 53699 4607
rect 55781 4573 55815 4607
rect 56057 4573 56091 4607
rect 58817 4573 58851 4607
rect 59277 4573 59311 4607
rect 60197 4573 60231 4607
rect 60749 4573 60783 4607
rect 39037 4505 39071 4539
rect 51714 4505 51748 4539
rect 54309 4505 54343 4539
rect 54769 4505 54803 4539
rect 3525 4437 3559 4471
rect 5825 4437 5859 4471
rect 6285 4437 6319 4471
rect 7941 4437 7975 4471
rect 10333 4437 10367 4471
rect 11253 4437 11287 4471
rect 11897 4437 11931 4471
rect 12541 4437 12575 4471
rect 14657 4437 14691 4471
rect 15485 4437 15519 4471
rect 16313 4437 16347 4471
rect 19625 4437 19659 4471
rect 19809 4437 19843 4471
rect 20269 4437 20303 4471
rect 20729 4437 20763 4471
rect 22201 4437 22235 4471
rect 22385 4437 22419 4471
rect 22753 4437 22787 4471
rect 23305 4437 23339 4471
rect 23673 4437 23707 4471
rect 25513 4437 25547 4471
rect 26341 4437 26375 4471
rect 29653 4437 29687 4471
rect 30113 4437 30147 4471
rect 30665 4437 30699 4471
rect 31125 4437 31159 4471
rect 33977 4437 34011 4471
rect 37381 4437 37415 4471
rect 38853 4437 38887 4471
rect 40785 4437 40819 4471
rect 43637 4437 43671 4471
rect 44189 4437 44223 4471
rect 45201 4437 45235 4471
rect 46673 4437 46707 4471
rect 48421 4437 48455 4471
rect 49157 4437 49191 4471
rect 51365 4437 51399 4471
rect 51825 4437 51859 4471
rect 52561 4437 52595 4471
rect 52929 4437 52963 4471
rect 59553 4437 59587 4471
rect 61485 4437 61519 4471
rect 2513 4233 2547 4267
rect 3617 4233 3651 4267
rect 4721 4233 4755 4267
rect 7297 4233 7331 4267
rect 8769 4233 8803 4267
rect 9965 4233 9999 4267
rect 12265 4233 12299 4267
rect 12587 4233 12621 4267
rect 12725 4233 12759 4267
rect 13921 4233 13955 4267
rect 16221 4233 16255 4267
rect 17325 4233 17359 4267
rect 22109 4233 22143 4267
rect 23857 4233 23891 4267
rect 27445 4233 27479 4267
rect 31125 4233 31159 4267
rect 32413 4233 32447 4267
rect 34253 4233 34287 4267
rect 34621 4233 34655 4267
rect 37105 4233 37139 4267
rect 38853 4233 38887 4267
rect 40325 4233 40359 4267
rect 40601 4233 40635 4267
rect 47317 4233 47351 4267
rect 47869 4233 47903 4267
rect 58357 4233 58391 4267
rect 58725 4233 58759 4267
rect 61117 4233 61151 4267
rect 5181 4165 5215 4199
rect 8493 4165 8527 4199
rect 11437 4165 11471 4199
rect 11897 4165 11931 4199
rect 14841 4165 14875 4199
rect 17693 4165 17727 4199
rect 26157 4165 26191 4199
rect 28825 4165 28859 4199
rect 31493 4165 31527 4199
rect 2145 4097 2179 4131
rect 3709 4097 3743 4131
rect 5825 4097 5859 4131
rect 6653 4097 6687 4131
rect 8125 4097 8159 4131
rect 10057 4097 10091 4131
rect 12909 4097 12943 4131
rect 13461 4097 13495 4131
rect 15025 4097 15059 4131
rect 17049 4097 17083 4131
rect 19441 4097 19475 4131
rect 19993 4097 20027 4131
rect 21005 4097 21039 4131
rect 21373 4097 21407 4131
rect 24225 4097 24259 4131
rect 25881 4097 25915 4131
rect 3488 4029 3522 4063
rect 4077 4029 4111 4063
rect 5365 4029 5399 4063
rect 5733 4029 5767 4063
rect 6285 4029 6319 4063
rect 9229 4029 9263 4063
rect 9836 4029 9870 4063
rect 11253 4029 11287 4063
rect 12788 4029 12822 4063
rect 14381 4029 14415 4063
rect 14933 4029 14967 4063
rect 18797 4029 18831 4063
rect 20545 4029 20579 4063
rect 20821 4029 20855 4063
rect 21649 4029 21683 4063
rect 22385 4029 22419 4063
rect 22753 4029 22787 4063
rect 24685 4029 24719 4063
rect 24869 4029 24903 4063
rect 26341 4029 26375 4063
rect 26801 4029 26835 4063
rect 27721 4029 27755 4063
rect 27905 4029 27939 4063
rect 29009 4097 29043 4131
rect 29745 4097 29779 4131
rect 30205 4097 30239 4131
rect 32229 4097 32263 4131
rect 30113 4029 30147 4063
rect 30297 4029 30331 4063
rect 30757 4029 30791 4063
rect 31610 4029 31644 4063
rect 3249 3961 3283 3995
rect 3341 3961 3375 3995
rect 4353 3961 4387 3995
rect 7389 3961 7423 3995
rect 7757 3961 7791 3995
rect 9597 3961 9631 3995
rect 9689 3961 9723 3995
rect 10425 3961 10459 3995
rect 12449 3961 12483 3995
rect 15485 3961 15519 3995
rect 16313 3961 16347 3995
rect 16681 3961 16715 3995
rect 18521 3961 18555 3995
rect 18613 3961 18647 3995
rect 19165 3961 19199 3995
rect 19901 3961 19935 3995
rect 22201 3961 22235 3995
rect 27813 3961 27847 3995
rect 28365 3961 28399 3995
rect 28825 3961 28859 3995
rect 32597 4165 32631 4199
rect 34897 4165 34931 4199
rect 39957 4165 39991 4199
rect 42257 4165 42291 4199
rect 44005 4165 44039 4199
rect 49157 4165 49191 4199
rect 53021 4165 53055 4199
rect 54493 4165 54527 4199
rect 61485 4165 61519 4199
rect 33241 4097 33275 4131
rect 37473 4097 37507 4131
rect 38301 4097 38335 4131
rect 38669 4097 38703 4131
rect 39589 4097 39623 4131
rect 43729 4097 43763 4131
rect 47317 4097 47351 4131
rect 48053 4097 48087 4131
rect 52285 4097 52319 4131
rect 54217 4097 54251 4131
rect 55413 4097 55447 4131
rect 57437 4097 57471 4131
rect 59093 4097 59127 4131
rect 62221 4097 62255 4131
rect 32689 4029 32723 4063
rect 33517 4029 33551 4063
rect 33701 4029 33735 4063
rect 35357 4029 35391 4063
rect 36001 4029 36035 4063
rect 36277 4029 36311 4063
rect 36553 4029 36587 4063
rect 37657 4029 37691 4063
rect 39129 4029 39163 4063
rect 40785 4029 40819 4063
rect 41245 4029 41279 4063
rect 42073 4029 42107 4063
rect 42625 4029 42659 4063
rect 44741 4029 44775 4063
rect 45017 4029 45051 4063
rect 45201 4029 45235 4063
rect 46213 4029 46247 4063
rect 47041 4029 47075 4063
rect 47179 4029 47213 4063
rect 47501 4029 47535 4063
rect 48605 4029 48639 4063
rect 48881 4029 48915 4063
rect 49065 4029 49099 4063
rect 49157 4029 49191 4063
rect 50077 4029 50111 4063
rect 50721 4029 50755 4063
rect 50905 4029 50939 4063
rect 51733 4029 51767 4063
rect 51825 4029 51859 4063
rect 53389 4029 53423 4063
rect 53481 4029 53515 4063
rect 53665 4029 53699 4063
rect 54861 4029 54895 4063
rect 54953 4029 54987 4063
rect 55689 4029 55723 4063
rect 56425 4029 56459 4063
rect 57529 4029 57563 4063
rect 58817 4029 58851 4063
rect 61301 4029 61335 4063
rect 61853 4029 61887 4063
rect 35265 3961 35299 3995
rect 39037 3961 39071 3995
rect 44189 3961 44223 3995
rect 45477 3961 45511 3995
rect 46305 3961 46339 3995
rect 49709 3961 49743 3995
rect 49893 3961 49927 3995
rect 51549 3961 51583 3995
rect 52653 3961 52687 3995
rect 54677 3961 54711 3995
rect 55045 3961 55079 3995
rect 57069 3961 57103 3995
rect 57989 3961 58023 3995
rect 2881 3893 2915 3927
rect 7573 3893 7607 3927
rect 7665 3893 7699 3927
rect 10701 3893 10735 3927
rect 11161 3893 11195 3927
rect 16497 3893 16531 3927
rect 16589 3893 16623 3927
rect 23029 3893 23063 3927
rect 23397 3893 23431 3927
rect 24961 3893 24995 3927
rect 25513 3893 25547 3927
rect 27169 3893 27203 3927
rect 28641 3893 28675 3927
rect 31769 3893 31803 3927
rect 32413 3893 32447 3927
rect 32781 3893 32815 3927
rect 33885 3893 33919 3927
rect 37841 3893 37875 3927
rect 41613 3893 41647 3927
rect 41981 3893 42015 3927
rect 43361 3893 43395 3927
rect 45937 3893 45971 3927
rect 49341 3893 49375 3927
rect 50169 3893 50203 3927
rect 50905 3893 50939 3927
rect 51089 3893 51123 3927
rect 56057 3893 56091 3927
rect 60197 3893 60231 3927
rect 4169 3689 4203 3723
rect 4905 3689 4939 3723
rect 9413 3689 9447 3723
rect 14105 3689 14139 3723
rect 14749 3689 14783 3723
rect 18153 3689 18187 3723
rect 23213 3689 23247 3723
rect 25513 3689 25547 3723
rect 25973 3689 26007 3723
rect 31953 3689 31987 3723
rect 32413 3689 32447 3723
rect 36553 3689 36587 3723
rect 37933 3689 37967 3723
rect 39865 3689 39899 3723
rect 41981 3689 42015 3723
rect 42257 3689 42291 3723
rect 44373 3689 44407 3723
rect 47593 3689 47627 3723
rect 47961 3689 47995 3723
rect 48789 3689 48823 3723
rect 49157 3689 49191 3723
rect 49893 3689 49927 3723
rect 51825 3689 51859 3723
rect 54217 3689 54251 3723
rect 54769 3689 54803 3723
rect 56241 3689 56275 3723
rect 56793 3689 56827 3723
rect 57897 3689 57931 3723
rect 58081 3689 58115 3723
rect 8677 3621 8711 3655
rect 11989 3621 12023 3655
rect 17233 3621 17267 3655
rect 22569 3621 22603 3655
rect 29377 3621 29411 3655
rect 32505 3621 32539 3655
rect 35081 3621 35115 3655
rect 36829 3621 36863 3655
rect 41613 3621 41647 3655
rect 47225 3621 47259 3655
rect 52745 3621 52779 3655
rect 55689 3621 55723 3655
rect 57345 3621 57379 3655
rect 59277 3621 59311 3655
rect 2697 3553 2731 3587
rect 3525 3553 3559 3587
rect 4077 3553 4111 3587
rect 4537 3553 4571 3587
rect 5917 3553 5951 3587
rect 6285 3553 6319 3587
rect 7573 3553 7607 3587
rect 8033 3553 8067 3587
rect 10149 3553 10183 3587
rect 11069 3553 11103 3587
rect 12265 3553 12299 3587
rect 12817 3553 12851 3587
rect 13001 3553 13035 3587
rect 15669 3553 15703 3587
rect 16221 3553 16255 3587
rect 17417 3553 17451 3587
rect 17785 3553 17819 3587
rect 19257 3553 19291 3587
rect 19993 3553 20027 3587
rect 20637 3553 20671 3587
rect 21189 3553 21223 3587
rect 24225 3553 24259 3587
rect 25329 3553 25363 3587
rect 26525 3553 26559 3587
rect 28089 3553 28123 3587
rect 28273 3553 28307 3587
rect 28549 3553 28583 3587
rect 28733 3553 28767 3587
rect 29009 3553 29043 3587
rect 29745 3553 29779 3587
rect 30205 3553 30239 3587
rect 30573 3553 30607 3587
rect 32321 3553 32355 3587
rect 34253 3553 34287 3587
rect 34621 3553 34655 3587
rect 34713 3553 34747 3587
rect 35725 3553 35759 3587
rect 38669 3553 38703 3587
rect 38853 3553 38887 3587
rect 40693 3553 40727 3587
rect 41061 3553 41095 3587
rect 42073 3553 42107 3587
rect 43729 3553 43763 3587
rect 45569 3553 45603 3587
rect 47501 3553 47535 3587
rect 47777 3553 47811 3587
rect 48973 3553 49007 3587
rect 50077 3553 50111 3587
rect 50905 3553 50939 3587
rect 51089 3553 51123 3587
rect 52009 3553 52043 3587
rect 52101 3553 52135 3587
rect 52285 3553 52319 3587
rect 53389 3553 53423 3587
rect 54953 3553 54987 3587
rect 55045 3553 55079 3587
rect 55229 3553 55263 3587
rect 56517 3553 56551 3587
rect 56701 3553 56735 3587
rect 57897 3553 57931 3587
rect 58357 3553 58391 3587
rect 58541 3553 58575 3587
rect 58817 3553 58851 3587
rect 59553 3553 59587 3587
rect 59921 3553 59955 3587
rect 60197 3553 60231 3587
rect 60381 3553 60415 3587
rect 2605 3485 2639 3519
rect 3157 3485 3191 3519
rect 5825 3485 5859 3519
rect 6377 3485 6411 3519
rect 9137 3485 9171 3519
rect 10241 3485 10275 3519
rect 10793 3485 10827 3519
rect 11253 3485 11287 3519
rect 12081 3485 12115 3519
rect 15025 3485 15059 3519
rect 15485 3485 15519 3519
rect 16405 3485 16439 3519
rect 18429 3485 18463 3519
rect 19625 3485 19659 3519
rect 20913 3485 20947 3519
rect 23397 3485 23431 3519
rect 23949 3485 23983 3519
rect 24409 3485 24443 3519
rect 27629 3485 27663 3519
rect 31585 3485 31619 3519
rect 32137 3485 32171 3519
rect 32873 3485 32907 3519
rect 35357 3485 35391 3519
rect 35633 3485 35667 3519
rect 36185 3485 36219 3519
rect 38577 3485 38611 3519
rect 39221 3485 39255 3519
rect 40601 3485 40635 3519
rect 41153 3485 41187 3519
rect 43637 3485 43671 3519
rect 44097 3485 44131 3519
rect 45293 3485 45327 3519
rect 3893 3417 3927 3451
rect 7389 3417 7423 3451
rect 8309 3417 8343 3451
rect 11621 3417 11655 3451
rect 20361 3417 20395 3451
rect 26709 3417 26743 3451
rect 30021 3417 30055 3451
rect 31125 3417 31159 3451
rect 34069 3417 34103 3451
rect 42717 3417 42751 3451
rect 43894 3417 43928 3451
rect 44833 3417 44867 3451
rect 45109 3417 45143 3451
rect 46673 3417 46707 3451
rect 58633 3485 58667 3519
rect 50813 3417 50847 3451
rect 53849 3417 53883 3451
rect 5365 3349 5399 3383
rect 6837 3349 6871 3383
rect 7205 3349 7239 3383
rect 13277 3349 13311 3383
rect 13829 3349 13863 3383
rect 16681 3349 16715 3383
rect 17141 3349 17175 3383
rect 19165 3349 19199 3383
rect 22845 3349 22879 3383
rect 24685 3349 24719 3383
rect 25053 3349 25087 3383
rect 26341 3349 26375 3383
rect 27169 3349 27203 3383
rect 27445 3349 27479 3383
rect 33241 3349 33275 3383
rect 33517 3349 33551 3383
rect 35357 3349 35391 3383
rect 35449 3349 35483 3383
rect 37197 3349 37231 3383
rect 39497 3349 39531 3383
rect 40141 3349 40175 3383
rect 42993 3349 43027 3383
rect 44005 3349 44039 3383
rect 47501 3349 47535 3383
rect 48421 3349 48455 3383
rect 49525 3349 49559 3383
rect 51549 3349 51583 3383
rect 53021 3349 53055 3383
rect 60473 3349 60507 3383
rect 61117 3349 61151 3383
rect 61577 3349 61611 3383
rect 2697 3145 2731 3179
rect 2973 3145 3007 3179
rect 5089 3145 5123 3179
rect 5917 3145 5951 3179
rect 6377 3145 6411 3179
rect 8309 3145 8343 3179
rect 10241 3145 10275 3179
rect 10885 3145 10919 3179
rect 11621 3145 11655 3179
rect 11897 3145 11931 3179
rect 14473 3145 14507 3179
rect 16773 3145 16807 3179
rect 17785 3145 17819 3179
rect 18061 3145 18095 3179
rect 21281 3145 21315 3179
rect 21465 3145 21499 3179
rect 25329 3145 25363 3179
rect 28365 3145 28399 3179
rect 32229 3145 32263 3179
rect 34713 3145 34747 3179
rect 35633 3145 35667 3179
rect 38117 3145 38151 3179
rect 42073 3145 42107 3179
rect 42717 3145 42751 3179
rect 45477 3145 45511 3179
rect 48789 3145 48823 3179
rect 49249 3145 49283 3179
rect 51549 3145 51583 3179
rect 52561 3145 52595 3179
rect 53849 3145 53883 3179
rect 55965 3145 55999 3179
rect 56333 3145 56367 3179
rect 56701 3145 56735 3179
rect 57161 3145 57195 3179
rect 57621 3145 57655 3179
rect 57989 3145 58023 3179
rect 58633 3145 58667 3179
rect 58909 3145 58943 3179
rect 61117 3145 61151 3179
rect 61301 3145 61335 3179
rect 62313 3145 62347 3179
rect 3709 3009 3743 3043
rect 3985 3009 4019 3043
rect 7389 3009 7423 3043
rect 7941 3009 7975 3043
rect 8677 3009 8711 3043
rect 9505 3009 9539 3043
rect 9965 3009 9999 3043
rect 10425 3009 10459 3043
rect 11529 3009 11563 3043
rect 2329 2941 2363 2975
rect 3617 2941 3651 2975
rect 7481 2941 7515 2975
rect 7849 2941 7883 2975
rect 9427 2941 9461 2975
rect 9873 2941 9907 2975
rect 10241 2941 10275 2975
rect 11161 2941 11195 2975
rect 16405 3077 16439 3111
rect 12725 3009 12759 3043
rect 13737 3009 13771 3043
rect 14013 3009 14047 3043
rect 14841 3009 14875 3043
rect 15669 3009 15703 3043
rect 18797 3009 18831 3043
rect 20637 3009 20671 3043
rect 21649 3077 21683 3111
rect 25605 3077 25639 3111
rect 31493 3077 31527 3111
rect 35081 3077 35115 3111
rect 22293 3009 22327 3043
rect 23489 3009 23523 3043
rect 23765 3009 23799 3043
rect 12265 2941 12299 2975
rect 13277 2941 13311 2975
rect 13553 2941 13587 2975
rect 15577 2941 15611 2975
rect 15945 2941 15979 2975
rect 16129 2941 16163 2975
rect 18337 2941 18371 2975
rect 19901 2941 19935 2975
rect 20085 2941 20119 2975
rect 20177 2941 20211 2975
rect 21465 2941 21499 2975
rect 22201 2941 22235 2975
rect 22569 2941 22603 2975
rect 22753 2941 22787 2975
rect 24593 2941 24627 2975
rect 24731 2941 24765 2975
rect 6837 2873 6871 2907
rect 8861 2873 8895 2907
rect 10977 2873 11011 2907
rect 11621 2873 11655 2907
rect 14933 2873 14967 2907
rect 17417 2873 17451 2907
rect 18245 2873 18279 2907
rect 19073 2873 19107 2907
rect 23857 2873 23891 2907
rect 37841 3077 37875 3111
rect 39957 3077 39991 3111
rect 40325 3077 40359 3111
rect 42809 3077 42843 3111
rect 47593 3077 47627 3111
rect 52745 3077 52779 3111
rect 61006 3077 61040 3111
rect 25697 3009 25731 3043
rect 26525 3009 26559 3043
rect 27353 3009 27387 3043
rect 29745 3009 29779 3043
rect 30849 3009 30883 3043
rect 32597 3009 32631 3043
rect 33977 3009 34011 3043
rect 34069 3009 34103 3043
rect 34345 3009 34379 3043
rect 35633 3009 35667 3043
rect 36093 3009 36127 3043
rect 39589 3009 39623 3043
rect 40785 3009 40819 3043
rect 42717 3009 42751 3043
rect 50813 3009 50847 3043
rect 52653 3009 52687 3043
rect 53297 3009 53331 3043
rect 54585 3009 54619 3043
rect 55597 3009 55631 3043
rect 59369 3009 59403 3043
rect 61206 3009 61240 3043
rect 27261 2941 27295 2975
rect 27629 2941 27663 2975
rect 27721 2941 27755 2975
rect 29285 2941 29319 2975
rect 29469 2941 29503 2975
rect 30297 2941 30331 2975
rect 31033 2941 31067 2975
rect 31493 2941 31527 2975
rect 33333 2941 33367 2975
rect 33517 2941 33551 2975
rect 26065 2873 26099 2907
rect 26617 2873 26651 2907
rect 28825 2873 28859 2907
rect 30481 2873 30515 2907
rect 33425 2873 33459 2907
rect 34897 2941 34931 2975
rect 36277 2941 36311 2975
rect 36369 2941 36403 2975
rect 36829 2941 36863 2975
rect 37933 2941 37967 2975
rect 39221 2941 39255 2975
rect 40509 2941 40543 2975
rect 42993 2941 43027 2975
rect 44649 2941 44683 2975
rect 44741 2941 44775 2975
rect 45017 2941 45051 2975
rect 45201 2941 45235 2975
rect 46213 2941 46247 2975
rect 46305 2941 46339 2975
rect 47041 2941 47075 2975
rect 47133 2941 47167 2975
rect 47961 2941 47995 2975
rect 49341 2941 49375 2975
rect 49893 2941 49927 2975
rect 50353 2941 50387 2975
rect 50721 2941 50755 2975
rect 52193 2941 52227 2975
rect 52432 2941 52466 2975
rect 54125 2941 54159 2975
rect 54861 2941 54895 2975
rect 55321 2941 55355 2975
rect 56149 2941 56183 2975
rect 59461 2941 59495 2975
rect 59829 2941 59863 2975
rect 60013 2941 60047 2975
rect 36461 2873 36495 2907
rect 38485 2873 38519 2907
rect 39037 2873 39071 2907
rect 42533 2873 42567 2907
rect 44005 2873 44039 2907
rect 45845 2873 45879 2907
rect 51181 2873 51215 2907
rect 52285 2873 52319 2907
rect 54033 2873 54067 2907
rect 58265 2873 58299 2907
rect 60289 2873 60323 2907
rect 60749 2873 60783 2907
rect 60841 2873 60875 2907
rect 1961 2805 1995 2839
rect 19441 2805 19475 2839
rect 23029 2805 23063 2839
rect 25605 2805 25639 2839
rect 30113 2805 30147 2839
rect 30297 2805 30331 2839
rect 32965 2805 32999 2839
rect 34069 2805 34103 2839
rect 35817 2805 35851 2839
rect 37105 2805 37139 2839
rect 38853 2805 38887 2839
rect 43085 2805 43119 2839
rect 43821 2805 43855 2839
rect 48421 2805 48455 2839
rect 53757 2805 53791 2839
rect 61853 2805 61887 2839
rect 3065 2601 3099 2635
rect 5733 2601 5767 2635
rect 6285 2601 6319 2635
rect 9505 2601 9539 2635
rect 10701 2601 10735 2635
rect 10793 2601 10827 2635
rect 12173 2601 12207 2635
rect 12357 2601 12391 2635
rect 12909 2601 12943 2635
rect 13461 2601 13495 2635
rect 14749 2601 14783 2635
rect 15209 2601 15243 2635
rect 17785 2601 17819 2635
rect 19625 2601 19659 2635
rect 25145 2601 25179 2635
rect 26617 2601 26651 2635
rect 28273 2601 28307 2635
rect 29193 2601 29227 2635
rect 32321 2601 32355 2635
rect 34897 2601 34931 2635
rect 36093 2601 36127 2635
rect 38577 2601 38611 2635
rect 39313 2601 39347 2635
rect 40785 2601 40819 2635
rect 43821 2601 43855 2635
rect 46213 2601 46247 2635
rect 47041 2601 47075 2635
rect 49893 2601 49927 2635
rect 51917 2601 51951 2635
rect 53849 2601 53883 2635
rect 54677 2601 54711 2635
rect 54953 2601 54987 2635
rect 55689 2601 55723 2635
rect 58541 2601 58575 2635
rect 62221 2601 62255 2635
rect 8861 2533 8895 2567
rect 9229 2533 9263 2567
rect 10149 2533 10183 2567
rect 2973 2465 3007 2499
rect 3433 2465 3467 2499
rect 3893 2465 3927 2499
rect 4629 2465 4663 2499
rect 6745 2465 6779 2499
rect 7481 2465 7515 2499
rect 10701 2465 10735 2499
rect 10977 2465 11011 2499
rect 11161 2465 11195 2499
rect 11253 2465 11287 2499
rect 2513 2397 2547 2431
rect 2881 2397 2915 2431
rect 4353 2397 4387 2431
rect 7205 2397 7239 2431
rect 10517 2397 10551 2431
rect 14013 2465 14047 2499
rect 14381 2465 14415 2499
rect 14473 2465 14507 2499
rect 17141 2533 17175 2567
rect 18889 2533 18923 2567
rect 20269 2533 20303 2567
rect 23121 2533 23155 2567
rect 23489 2533 23523 2567
rect 24225 2533 24259 2567
rect 25421 2533 25455 2567
rect 28825 2533 28859 2567
rect 39681 2533 39715 2567
rect 40233 2533 40267 2567
rect 45937 2533 45971 2567
rect 48789 2533 48823 2567
rect 50077 2533 50111 2567
rect 50813 2533 50847 2567
rect 52377 2533 52411 2567
rect 53205 2533 53239 2567
rect 59001 2533 59035 2567
rect 59461 2533 59495 2567
rect 15485 2465 15519 2499
rect 15761 2465 15795 2499
rect 18153 2465 18187 2499
rect 18337 2465 18371 2499
rect 18521 2465 18555 2499
rect 19165 2465 19199 2499
rect 19717 2465 19751 2499
rect 19901 2465 19935 2499
rect 20545 2465 20579 2499
rect 21005 2465 21039 2499
rect 21741 2465 21775 2499
rect 24317 2465 24351 2499
rect 25605 2465 25639 2499
rect 26157 2465 26191 2499
rect 27169 2465 27203 2499
rect 30113 2465 30147 2499
rect 30757 2465 30791 2499
rect 31125 2465 31159 2499
rect 31953 2465 31987 2499
rect 32597 2465 32631 2499
rect 35909 2465 35943 2499
rect 36001 2465 36035 2499
rect 36645 2465 36679 2499
rect 36829 2465 36863 2499
rect 38393 2465 38427 2499
rect 39497 2465 39531 2499
rect 39773 2465 39807 2499
rect 41797 2465 41831 2499
rect 44557 2465 44591 2499
rect 46857 2465 46891 2499
rect 47961 2465 47995 2499
rect 48053 2465 48087 2499
rect 50905 2465 50939 2499
rect 53352 2465 53386 2499
rect 59608 2465 59642 2499
rect 60841 2465 60875 2499
rect 61117 2465 61151 2499
rect 62129 2465 62163 2499
rect 14657 2397 14691 2431
rect 14749 2397 14783 2431
rect 21465 2397 21499 2431
rect 24777 2397 24811 2431
rect 26893 2397 26927 2431
rect 30481 2397 30515 2431
rect 31401 2397 31435 2431
rect 32873 2397 32907 2431
rect 37381 2397 37415 2431
rect 39037 2397 39071 2431
rect 41705 2397 41739 2431
rect 42165 2397 42199 2431
rect 42809 2397 42843 2431
rect 44281 2397 44315 2431
rect 48421 2397 48455 2431
rect 50445 2397 50479 2431
rect 13829 2329 13863 2363
rect 2145 2261 2179 2295
rect 11437 2261 11471 2295
rect 12173 2261 12207 2295
rect 25789 2329 25823 2363
rect 30849 2329 30883 2363
rect 42073 2329 42107 2363
rect 43177 2329 43211 2363
rect 50353 2329 50387 2363
rect 53573 2397 53607 2431
rect 54217 2397 54251 2431
rect 56793 2397 56827 2431
rect 57989 2397 58023 2431
rect 59829 2397 59863 2431
rect 60473 2397 60507 2431
rect 61209 2397 61243 2431
rect 51089 2329 51123 2363
rect 53113 2329 53147 2363
rect 59369 2329 59403 2363
rect 14657 2261 14691 2295
rect 14933 2261 14967 2295
rect 23857 2261 23891 2295
rect 24041 2261 24075 2295
rect 33977 2261 34011 2295
rect 34529 2261 34563 2295
rect 37841 2261 37875 2295
rect 41962 2261 41996 2295
rect 42441 2261 42475 2295
rect 46581 2261 46615 2295
rect 47593 2261 47627 2295
rect 48218 2261 48252 2295
rect 48329 2261 48363 2295
rect 49065 2261 49099 2295
rect 49525 2261 49559 2295
rect 50215 2261 50249 2295
rect 50905 2261 50939 2295
rect 51549 2261 51583 2295
rect 53481 2261 53515 2295
rect 55965 2261 55999 2295
rect 56333 2261 56367 2295
rect 59737 2261 59771 2295
rect 59921 2261 59955 2295
rect 61577 2261 61611 2295
rect 62589 2261 62623 2295
rect 9597 2057 9631 2091
rect 9597 1921 9631 1955
<< metal1 >>
rect 1104 17434 63480 17456
rect 1104 17382 11378 17434
rect 11430 17382 11442 17434
rect 11494 17382 11506 17434
rect 11558 17382 11570 17434
rect 11622 17382 32170 17434
rect 32222 17382 32234 17434
rect 32286 17382 32298 17434
rect 32350 17382 32362 17434
rect 32414 17382 52962 17434
rect 53014 17382 53026 17434
rect 53078 17382 53090 17434
rect 53142 17382 53154 17434
rect 53206 17382 63480 17434
rect 1104 17360 63480 17382
rect 14369 17323 14427 17329
rect 14369 17289 14381 17323
rect 14415 17320 14427 17323
rect 14642 17320 14648 17332
rect 14415 17292 14648 17320
rect 14415 17289 14427 17292
rect 14369 17283 14427 17289
rect 14642 17280 14648 17292
rect 14700 17280 14706 17332
rect 23477 17323 23535 17329
rect 23477 17289 23489 17323
rect 23523 17320 23535 17323
rect 24394 17320 24400 17332
rect 23523 17292 24400 17320
rect 23523 17289 23535 17292
rect 23477 17283 23535 17289
rect 19150 17212 19156 17264
rect 19208 17252 19214 17264
rect 20441 17255 20499 17261
rect 20441 17252 20453 17255
rect 19208 17224 20453 17252
rect 19208 17212 19214 17224
rect 12250 17144 12256 17196
rect 12308 17184 12314 17196
rect 12437 17187 12495 17193
rect 12437 17184 12449 17187
rect 12308 17156 12449 17184
rect 12308 17144 12314 17156
rect 12437 17153 12449 17156
rect 12483 17184 12495 17187
rect 12805 17187 12863 17193
rect 12805 17184 12817 17187
rect 12483 17156 12817 17184
rect 12483 17153 12495 17156
rect 12437 17147 12495 17153
rect 12805 17153 12817 17156
rect 12851 17184 12863 17187
rect 15746 17184 15752 17196
rect 12851 17156 15752 17184
rect 12851 17153 12863 17156
rect 12805 17147 12863 17153
rect 15746 17144 15752 17156
rect 15804 17144 15810 17196
rect 19260 17193 19288 17224
rect 20441 17221 20453 17224
rect 20487 17252 20499 17255
rect 22738 17252 22744 17264
rect 20487 17224 22744 17252
rect 20487 17221 20499 17224
rect 20441 17215 20499 17221
rect 22738 17212 22744 17224
rect 22796 17212 22802 17264
rect 19245 17187 19303 17193
rect 19245 17153 19257 17187
rect 19291 17153 19303 17187
rect 23492 17184 23520 17283
rect 24394 17280 24400 17292
rect 24452 17280 24458 17332
rect 28350 17280 28356 17332
rect 28408 17320 28414 17332
rect 28537 17323 28595 17329
rect 28537 17320 28549 17323
rect 28408 17292 28549 17320
rect 28408 17280 28414 17292
rect 28537 17289 28549 17292
rect 28583 17320 28595 17323
rect 28902 17320 28908 17332
rect 28583 17292 28908 17320
rect 28583 17289 28595 17292
rect 28537 17283 28595 17289
rect 28902 17280 28908 17292
rect 28960 17280 28966 17332
rect 42058 17280 42064 17332
rect 42116 17320 42122 17332
rect 42521 17323 42579 17329
rect 42521 17320 42533 17323
rect 42116 17292 42533 17320
rect 42116 17280 42122 17292
rect 42521 17289 42533 17292
rect 42567 17289 42579 17323
rect 42521 17283 42579 17289
rect 45922 17280 45928 17332
rect 45980 17320 45986 17332
rect 48130 17320 48136 17332
rect 45980 17292 48136 17320
rect 45980 17280 45986 17292
rect 48130 17280 48136 17292
rect 48188 17320 48194 17332
rect 48409 17323 48467 17329
rect 48409 17320 48421 17323
rect 48188 17292 48421 17320
rect 48188 17280 48194 17292
rect 48409 17289 48421 17292
rect 48455 17289 48467 17323
rect 48409 17283 48467 17289
rect 53834 17280 53840 17332
rect 53892 17320 53898 17332
rect 53929 17323 53987 17329
rect 53929 17320 53941 17323
rect 53892 17292 53941 17320
rect 53892 17280 53898 17292
rect 53929 17289 53941 17292
rect 53975 17289 53987 17323
rect 53929 17283 53987 17289
rect 33778 17252 33784 17264
rect 33739 17224 33784 17252
rect 33778 17212 33784 17224
rect 33836 17212 33842 17264
rect 49970 17252 49976 17264
rect 49931 17224 49976 17252
rect 49970 17212 49976 17224
rect 50028 17212 50034 17264
rect 19245 17147 19303 17153
rect 22572 17156 23520 17184
rect 26697 17187 26755 17193
rect 13081 17119 13139 17125
rect 13081 17085 13093 17119
rect 13127 17116 13139 17119
rect 13906 17116 13912 17128
rect 13127 17088 13912 17116
rect 13127 17085 13139 17088
rect 13081 17079 13139 17085
rect 13906 17076 13912 17088
rect 13964 17076 13970 17128
rect 18506 17076 18512 17128
rect 18564 17116 18570 17128
rect 22572 17125 22600 17156
rect 26697 17153 26709 17187
rect 26743 17184 26755 17187
rect 26743 17156 27476 17184
rect 26743 17153 26755 17156
rect 26697 17147 26755 17153
rect 18785 17119 18843 17125
rect 18785 17116 18797 17119
rect 18564 17088 18797 17116
rect 18564 17076 18570 17088
rect 18785 17085 18797 17088
rect 18831 17085 18843 17119
rect 18785 17079 18843 17085
rect 19153 17119 19211 17125
rect 19153 17085 19165 17119
rect 19199 17116 19211 17119
rect 22557 17119 22615 17125
rect 19199 17088 20116 17116
rect 19199 17085 19211 17088
rect 19153 17079 19211 17085
rect 18322 17048 18328 17060
rect 18283 17020 18328 17048
rect 18322 17008 18328 17020
rect 18380 17008 18386 17060
rect 18800 17048 18828 17079
rect 19242 17048 19248 17060
rect 18800 17020 19248 17048
rect 19242 17008 19248 17020
rect 19300 17048 19306 17060
rect 19613 17051 19671 17057
rect 19613 17048 19625 17051
rect 19300 17020 19625 17048
rect 19300 17008 19306 17020
rect 19613 17017 19625 17020
rect 19659 17017 19671 17051
rect 19613 17011 19671 17017
rect 20088 16989 20116 17088
rect 22557 17085 22569 17119
rect 22603 17085 22615 17119
rect 22738 17116 22744 17128
rect 22699 17088 22744 17116
rect 22557 17079 22615 17085
rect 22738 17076 22744 17088
rect 22796 17076 22802 17128
rect 22925 17119 22983 17125
rect 22925 17085 22937 17119
rect 22971 17116 22983 17119
rect 23106 17116 23112 17128
rect 22971 17088 23112 17116
rect 22971 17085 22983 17088
rect 22925 17079 22983 17085
rect 23106 17076 23112 17088
rect 23164 17116 23170 17128
rect 27448 17125 27476 17156
rect 27522 17144 27528 17196
rect 27580 17184 27586 17196
rect 29733 17187 29791 17193
rect 29733 17184 29745 17187
rect 27580 17156 29745 17184
rect 27580 17144 27586 17156
rect 29733 17153 29745 17156
rect 29779 17153 29791 17187
rect 31021 17187 31079 17193
rect 31021 17184 31033 17187
rect 29733 17147 29791 17153
rect 30208 17156 31033 17184
rect 23753 17119 23811 17125
rect 23753 17116 23765 17119
rect 23164 17088 23765 17116
rect 23164 17076 23170 17088
rect 23753 17085 23765 17088
rect 23799 17085 23811 17119
rect 23753 17079 23811 17085
rect 27157 17119 27215 17125
rect 27157 17085 27169 17119
rect 27203 17085 27215 17119
rect 27157 17079 27215 17085
rect 27433 17119 27491 17125
rect 27433 17085 27445 17119
rect 27479 17116 27491 17119
rect 28350 17116 28356 17128
rect 27479 17088 28356 17116
rect 27479 17085 27491 17088
rect 27433 17079 27491 17085
rect 22097 17051 22155 17057
rect 22097 17017 22109 17051
rect 22143 17048 22155 17051
rect 23566 17048 23572 17060
rect 22143 17020 23572 17048
rect 22143 17017 22155 17020
rect 22097 17011 22155 17017
rect 23566 17008 23572 17020
rect 23624 17008 23630 17060
rect 20073 16983 20131 16989
rect 20073 16949 20085 16983
rect 20119 16980 20131 16983
rect 20438 16980 20444 16992
rect 20119 16952 20444 16980
rect 20119 16949 20131 16952
rect 20073 16943 20131 16949
rect 20438 16940 20444 16952
rect 20496 16940 20502 16992
rect 20714 16980 20720 16992
rect 20675 16952 20720 16980
rect 20714 16940 20720 16952
rect 20772 16980 20778 16992
rect 21361 16983 21419 16989
rect 21361 16980 21373 16983
rect 20772 16952 21373 16980
rect 20772 16940 20778 16952
rect 21361 16949 21373 16952
rect 21407 16980 21419 16983
rect 21729 16983 21787 16989
rect 21729 16980 21741 16983
rect 21407 16952 21741 16980
rect 21407 16949 21419 16952
rect 21361 16943 21419 16949
rect 21729 16949 21741 16952
rect 21775 16949 21787 16983
rect 27172 16980 27200 17079
rect 28350 17076 28356 17088
rect 28408 17076 28414 17128
rect 28718 17076 28724 17128
rect 28776 17116 28782 17128
rect 30208 17125 30236 17156
rect 31021 17153 31033 17156
rect 31067 17153 31079 17187
rect 34238 17184 34244 17196
rect 31021 17147 31079 17153
rect 33980 17156 34244 17184
rect 30193 17119 30251 17125
rect 30193 17116 30205 17119
rect 28776 17088 30205 17116
rect 28776 17076 28782 17088
rect 30193 17085 30205 17088
rect 30239 17085 30251 17119
rect 30558 17116 30564 17128
rect 30519 17088 30564 17116
rect 30193 17079 30251 17085
rect 30558 17076 30564 17088
rect 30616 17076 30622 17128
rect 30653 17119 30711 17125
rect 30653 17085 30665 17119
rect 30699 17116 30711 17119
rect 30742 17116 30748 17128
rect 30699 17088 30748 17116
rect 30699 17085 30711 17088
rect 30653 17079 30711 17085
rect 30742 17076 30748 17088
rect 30800 17076 30806 17128
rect 33980 17125 34008 17156
rect 34238 17144 34244 17156
rect 34296 17184 34302 17196
rect 34793 17187 34851 17193
rect 34793 17184 34805 17187
rect 34296 17156 34805 17184
rect 34296 17144 34302 17156
rect 34793 17153 34805 17156
rect 34839 17153 34851 17187
rect 40313 17187 40371 17193
rect 40313 17184 40325 17187
rect 34793 17147 34851 17153
rect 39500 17156 40325 17184
rect 39500 17128 39528 17156
rect 40313 17153 40325 17156
rect 40359 17153 40371 17187
rect 40313 17147 40371 17153
rect 40957 17187 41015 17193
rect 40957 17153 40969 17187
rect 41003 17184 41015 17187
rect 46661 17187 46719 17193
rect 41003 17156 41460 17184
rect 41003 17153 41015 17156
rect 40957 17147 41015 17153
rect 33965 17119 34023 17125
rect 33965 17085 33977 17119
rect 34011 17085 34023 17119
rect 34146 17116 34152 17128
rect 34107 17088 34152 17116
rect 33965 17079 34023 17085
rect 34146 17076 34152 17088
rect 34204 17076 34210 17128
rect 34330 17116 34336 17128
rect 34291 17088 34336 17116
rect 34330 17076 34336 17088
rect 34388 17116 34394 17128
rect 35161 17119 35219 17125
rect 35161 17116 35173 17119
rect 34388 17088 35173 17116
rect 34388 17076 34394 17088
rect 35161 17085 35173 17088
rect 35207 17085 35219 17119
rect 39482 17116 39488 17128
rect 39443 17088 39488 17116
rect 35161 17079 35219 17085
rect 39482 17076 39488 17088
rect 39540 17076 39546 17128
rect 39669 17119 39727 17125
rect 39669 17116 39681 17119
rect 39592 17088 39681 17116
rect 30576 17048 30604 17076
rect 31389 17051 31447 17057
rect 31389 17048 31401 17051
rect 30576 17020 31401 17048
rect 31389 17017 31401 17020
rect 31435 17017 31447 17051
rect 39022 17048 39028 17060
rect 38983 17020 39028 17048
rect 31389 17011 31447 17017
rect 39022 17008 39028 17020
rect 39080 17008 39086 17060
rect 29362 16980 29368 16992
rect 27172 16952 29368 16980
rect 21729 16943 21787 16949
rect 29362 16940 29368 16952
rect 29420 16940 29426 16992
rect 38933 16983 38991 16989
rect 38933 16949 38945 16983
rect 38979 16980 38991 16983
rect 39206 16980 39212 16992
rect 38979 16952 39212 16980
rect 38979 16949 38991 16952
rect 38933 16943 38991 16949
rect 39206 16940 39212 16952
rect 39264 16980 39270 16992
rect 39592 16980 39620 17088
rect 39669 17085 39681 17088
rect 39715 17085 39727 17119
rect 39850 17116 39856 17128
rect 39811 17088 39856 17116
rect 39669 17079 39727 17085
rect 39850 17076 39856 17088
rect 39908 17076 39914 17128
rect 40218 17076 40224 17128
rect 40276 17116 40282 17128
rect 41432 17125 41460 17156
rect 46661 17153 46673 17187
rect 46707 17184 46719 17187
rect 50985 17187 51043 17193
rect 50985 17184 50997 17187
rect 46707 17156 47164 17184
rect 46707 17153 46719 17156
rect 46661 17147 46719 17153
rect 47136 17128 47164 17156
rect 50172 17156 50997 17184
rect 41141 17119 41199 17125
rect 41141 17116 41153 17119
rect 40276 17088 41153 17116
rect 40276 17076 40282 17088
rect 41141 17085 41153 17088
rect 41187 17085 41199 17119
rect 41141 17079 41199 17085
rect 41417 17119 41475 17125
rect 41417 17085 41429 17119
rect 41463 17116 41475 17119
rect 43622 17116 43628 17128
rect 41463 17088 43628 17116
rect 41463 17085 41475 17088
rect 41417 17079 41475 17085
rect 43622 17076 43628 17088
rect 43680 17076 43686 17128
rect 46845 17119 46903 17125
rect 46845 17085 46857 17119
rect 46891 17116 46903 17119
rect 46934 17116 46940 17128
rect 46891 17088 46940 17116
rect 46891 17085 46903 17088
rect 46845 17079 46903 17085
rect 46934 17076 46940 17088
rect 46992 17076 46998 17128
rect 47118 17116 47124 17128
rect 47079 17088 47124 17116
rect 47118 17076 47124 17088
rect 47176 17076 47182 17128
rect 49878 17076 49884 17128
rect 49936 17116 49942 17128
rect 50172 17125 50200 17156
rect 50985 17153 50997 17156
rect 51031 17153 51043 17187
rect 53852 17184 53880 17280
rect 50985 17147 51043 17153
rect 53116 17156 53880 17184
rect 50157 17119 50215 17125
rect 50157 17116 50169 17119
rect 49936 17088 50169 17116
rect 49936 17076 49942 17088
rect 50157 17085 50169 17088
rect 50203 17085 50215 17119
rect 50338 17116 50344 17128
rect 50299 17088 50344 17116
rect 50157 17079 50215 17085
rect 50338 17076 50344 17088
rect 50396 17076 50402 17128
rect 53116 17125 53144 17156
rect 50525 17119 50583 17125
rect 50525 17085 50537 17119
rect 50571 17085 50583 17119
rect 50525 17079 50583 17085
rect 53101 17119 53159 17125
rect 53101 17085 53113 17119
rect 53147 17085 53159 17119
rect 53101 17079 53159 17085
rect 53469 17119 53527 17125
rect 53469 17085 53481 17119
rect 53515 17085 53527 17119
rect 53469 17079 53527 17085
rect 53561 17119 53619 17125
rect 53561 17085 53573 17119
rect 53607 17116 53619 17119
rect 53926 17116 53932 17128
rect 53607 17088 53932 17116
rect 53607 17085 53619 17088
rect 53561 17079 53619 17085
rect 48774 17008 48780 17060
rect 48832 17048 48838 17060
rect 50540 17048 50568 17079
rect 52641 17051 52699 17057
rect 48832 17020 51488 17048
rect 48832 17008 48838 17020
rect 43070 16980 43076 16992
rect 39264 16952 39620 16980
rect 43031 16952 43076 16980
rect 39264 16940 39270 16952
rect 43070 16940 43076 16952
rect 43128 16940 43134 16992
rect 51460 16989 51488 17020
rect 52641 17017 52653 17051
rect 52687 17048 52699 17051
rect 52822 17048 52828 17060
rect 52687 17020 52828 17048
rect 52687 17017 52699 17020
rect 52641 17011 52699 17017
rect 52822 17008 52828 17020
rect 52880 17008 52886 17060
rect 53484 16992 53512 17079
rect 53926 17076 53932 17088
rect 53984 17076 53990 17128
rect 51445 16983 51503 16989
rect 51445 16949 51457 16983
rect 51491 16980 51503 16983
rect 53466 16980 53472 16992
rect 51491 16952 53472 16980
rect 51491 16949 51503 16952
rect 51445 16943 51503 16949
rect 53466 16940 53472 16952
rect 53524 16980 53530 16992
rect 54297 16983 54355 16989
rect 54297 16980 54309 16983
rect 53524 16952 54309 16980
rect 53524 16940 53530 16952
rect 54297 16949 54309 16952
rect 54343 16949 54355 16983
rect 54297 16943 54355 16949
rect 1104 16890 63480 16912
rect 1104 16838 21774 16890
rect 21826 16838 21838 16890
rect 21890 16838 21902 16890
rect 21954 16838 21966 16890
rect 22018 16838 42566 16890
rect 42618 16838 42630 16890
rect 42682 16838 42694 16890
rect 42746 16838 42758 16890
rect 42810 16838 63480 16890
rect 1104 16816 63480 16838
rect 12618 16776 12624 16788
rect 12579 16748 12624 16776
rect 12618 16736 12624 16748
rect 12676 16736 12682 16788
rect 16666 16736 16672 16788
rect 16724 16776 16730 16788
rect 17126 16776 17132 16788
rect 16724 16748 17132 16776
rect 16724 16736 16730 16748
rect 17126 16736 17132 16748
rect 17184 16736 17190 16788
rect 19242 16736 19248 16788
rect 19300 16776 19306 16788
rect 19613 16779 19671 16785
rect 19613 16776 19625 16779
rect 19300 16748 19625 16776
rect 19300 16736 19306 16748
rect 19613 16745 19625 16748
rect 19659 16745 19671 16779
rect 22462 16776 22468 16788
rect 22423 16748 22468 16776
rect 19613 16739 19671 16745
rect 22462 16736 22468 16748
rect 22520 16736 22526 16788
rect 24486 16736 24492 16788
rect 24544 16776 24550 16788
rect 24949 16779 25007 16785
rect 24949 16776 24961 16779
rect 24544 16748 24961 16776
rect 24544 16736 24550 16748
rect 24949 16745 24961 16748
rect 24995 16745 25007 16779
rect 24949 16739 25007 16745
rect 34238 16736 34244 16788
rect 34296 16776 34302 16788
rect 35989 16779 36047 16785
rect 35989 16776 36001 16779
rect 34296 16748 36001 16776
rect 34296 16736 34302 16748
rect 35989 16745 36001 16748
rect 36035 16745 36047 16779
rect 35989 16739 36047 16745
rect 40126 16736 40132 16788
rect 40184 16776 40190 16788
rect 41601 16779 41659 16785
rect 41601 16776 41613 16779
rect 40184 16748 41613 16776
rect 40184 16736 40190 16748
rect 41601 16745 41613 16748
rect 41647 16745 41659 16779
rect 48774 16776 48780 16788
rect 48735 16748 48780 16776
rect 41601 16739 41659 16745
rect 48774 16736 48780 16748
rect 48832 16736 48838 16788
rect 49878 16736 49884 16788
rect 49936 16776 49942 16788
rect 50341 16779 50399 16785
rect 50341 16776 50353 16779
rect 49936 16748 50353 16776
rect 49936 16736 49942 16748
rect 50341 16745 50353 16748
rect 50387 16745 50399 16779
rect 50341 16739 50399 16745
rect 50801 16779 50859 16785
rect 50801 16745 50813 16779
rect 50847 16776 50859 16779
rect 53926 16776 53932 16788
rect 50847 16748 53932 16776
rect 50847 16745 50859 16748
rect 50801 16739 50859 16745
rect 53926 16736 53932 16748
rect 53984 16776 53990 16788
rect 54113 16779 54171 16785
rect 54113 16776 54125 16779
rect 53984 16748 54125 16776
rect 53984 16736 53990 16748
rect 54113 16745 54125 16748
rect 54159 16745 54171 16779
rect 54113 16739 54171 16745
rect 47946 16708 47952 16720
rect 47504 16680 47952 16708
rect 8110 16600 8116 16652
rect 8168 16640 8174 16652
rect 8205 16643 8263 16649
rect 8205 16640 8217 16643
rect 8168 16612 8217 16640
rect 8168 16600 8174 16612
rect 8205 16609 8217 16612
rect 8251 16609 8263 16643
rect 8205 16603 8263 16609
rect 8389 16643 8447 16649
rect 8389 16609 8401 16643
rect 8435 16609 8447 16643
rect 8389 16603 8447 16609
rect 8573 16643 8631 16649
rect 8573 16609 8585 16643
rect 8619 16640 8631 16643
rect 9490 16640 9496 16652
rect 8619 16612 9496 16640
rect 8619 16609 8631 16612
rect 8573 16603 8631 16609
rect 7926 16532 7932 16584
rect 7984 16572 7990 16584
rect 8404 16572 8432 16603
rect 9490 16600 9496 16612
rect 9548 16600 9554 16652
rect 11057 16643 11115 16649
rect 11057 16609 11069 16643
rect 11103 16640 11115 16643
rect 12250 16640 12256 16652
rect 11103 16612 12256 16640
rect 11103 16609 11115 16612
rect 11057 16603 11115 16609
rect 12250 16600 12256 16612
rect 12308 16600 12314 16652
rect 13173 16643 13231 16649
rect 13173 16609 13185 16643
rect 13219 16640 13231 16643
rect 13906 16640 13912 16652
rect 13219 16612 13912 16640
rect 13219 16609 13231 16612
rect 13173 16603 13231 16609
rect 13906 16600 13912 16612
rect 13964 16600 13970 16652
rect 18046 16640 18052 16652
rect 18007 16612 18052 16640
rect 18046 16600 18052 16612
rect 18104 16640 18110 16652
rect 18233 16643 18291 16649
rect 18233 16640 18245 16643
rect 18104 16612 18245 16640
rect 18104 16600 18110 16612
rect 18233 16609 18245 16612
rect 18279 16609 18291 16643
rect 18233 16603 18291 16609
rect 21361 16643 21419 16649
rect 21361 16609 21373 16643
rect 21407 16640 21419 16643
rect 22094 16640 22100 16652
rect 21407 16612 22100 16640
rect 21407 16609 21419 16612
rect 21361 16603 21419 16609
rect 22094 16600 22100 16612
rect 22152 16600 22158 16652
rect 23569 16643 23627 16649
rect 23569 16640 23581 16643
rect 22204 16612 23581 16640
rect 7984 16544 8432 16572
rect 7984 16532 7990 16544
rect 11238 16532 11244 16584
rect 11296 16572 11302 16584
rect 11333 16575 11391 16581
rect 11333 16572 11345 16575
rect 11296 16544 11345 16572
rect 11296 16532 11302 16544
rect 11333 16541 11345 16544
rect 11379 16541 11391 16575
rect 15746 16572 15752 16584
rect 15707 16544 15752 16572
rect 11333 16535 11391 16541
rect 15746 16532 15752 16544
rect 15804 16532 15810 16584
rect 16022 16572 16028 16584
rect 15983 16544 16028 16572
rect 16022 16532 16028 16544
rect 16080 16532 16086 16584
rect 18506 16572 18512 16584
rect 18467 16544 18512 16572
rect 18506 16532 18512 16544
rect 18564 16532 18570 16584
rect 19978 16532 19984 16584
rect 20036 16572 20042 16584
rect 20714 16572 20720 16584
rect 20036 16544 20720 16572
rect 20036 16532 20042 16544
rect 20714 16532 20720 16544
rect 20772 16572 20778 16584
rect 21085 16575 21143 16581
rect 21085 16572 21097 16575
rect 20772 16544 21097 16572
rect 20772 16532 20778 16544
rect 21085 16541 21097 16544
rect 21131 16572 21143 16575
rect 21450 16572 21456 16584
rect 21131 16544 21456 16572
rect 21131 16541 21143 16544
rect 21085 16535 21143 16541
rect 21450 16532 21456 16544
rect 21508 16572 21514 16584
rect 22204 16572 22232 16612
rect 23569 16609 23581 16612
rect 23615 16640 23627 16643
rect 25038 16640 25044 16652
rect 23615 16612 25044 16640
rect 23615 16609 23627 16612
rect 23569 16603 23627 16609
rect 25038 16600 25044 16612
rect 25096 16600 25102 16652
rect 30282 16640 30288 16652
rect 30243 16612 30288 16640
rect 30282 16600 30288 16612
rect 30340 16600 30346 16652
rect 30650 16640 30656 16652
rect 30611 16612 30656 16640
rect 30650 16600 30656 16612
rect 30708 16600 30714 16652
rect 33318 16640 33324 16652
rect 30760 16612 33324 16640
rect 30760 16584 30788 16612
rect 33318 16600 33324 16612
rect 33376 16640 33382 16652
rect 34057 16643 34115 16649
rect 34057 16640 34069 16643
rect 33376 16612 34069 16640
rect 33376 16600 33382 16612
rect 34057 16609 34069 16612
rect 34103 16640 34115 16643
rect 34146 16640 34152 16652
rect 34103 16612 34152 16640
rect 34103 16609 34115 16612
rect 34057 16603 34115 16609
rect 34146 16600 34152 16612
rect 34204 16640 34210 16652
rect 34425 16643 34483 16649
rect 34425 16640 34437 16643
rect 34204 16612 34437 16640
rect 34204 16600 34210 16612
rect 34425 16609 34437 16612
rect 34471 16609 34483 16643
rect 34425 16603 34483 16609
rect 47302 16600 47308 16652
rect 47360 16640 47366 16652
rect 47504 16649 47532 16680
rect 47946 16668 47952 16680
rect 48004 16668 48010 16720
rect 47489 16643 47547 16649
rect 47489 16640 47501 16643
rect 47360 16612 47501 16640
rect 47360 16600 47366 16612
rect 47489 16609 47501 16612
rect 47535 16609 47547 16643
rect 47489 16603 47547 16609
rect 47673 16643 47731 16649
rect 47673 16609 47685 16643
rect 47719 16609 47731 16643
rect 47673 16603 47731 16609
rect 47857 16643 47915 16649
rect 47857 16609 47869 16643
rect 47903 16640 47915 16643
rect 48792 16640 48820 16736
rect 47903 16612 48820 16640
rect 48961 16643 49019 16649
rect 47903 16609 47915 16612
rect 47857 16603 47915 16609
rect 48961 16609 48973 16643
rect 49007 16640 49019 16643
rect 49007 16612 50660 16640
rect 49007 16609 49019 16612
rect 48961 16603 49019 16609
rect 23842 16572 23848 16584
rect 21508 16544 22232 16572
rect 23803 16544 23848 16572
rect 21508 16532 21514 16544
rect 23842 16532 23848 16544
rect 23900 16532 23906 16584
rect 27065 16575 27123 16581
rect 27065 16541 27077 16575
rect 27111 16572 27123 16575
rect 27341 16575 27399 16581
rect 27341 16572 27353 16575
rect 27111 16544 27353 16572
rect 27111 16541 27123 16544
rect 27065 16535 27123 16541
rect 27341 16541 27353 16544
rect 27387 16541 27399 16575
rect 27614 16572 27620 16584
rect 27575 16544 27620 16572
rect 27341 16535 27399 16541
rect 27614 16532 27620 16544
rect 27672 16532 27678 16584
rect 30742 16572 30748 16584
rect 30655 16544 30748 16572
rect 30742 16532 30748 16544
rect 30800 16532 30806 16584
rect 31938 16532 31944 16584
rect 31996 16572 32002 16584
rect 32125 16575 32183 16581
rect 32125 16572 32137 16575
rect 31996 16544 32137 16572
rect 31996 16532 32002 16544
rect 32125 16541 32137 16544
rect 32171 16541 32183 16575
rect 32125 16535 32183 16541
rect 32401 16575 32459 16581
rect 32401 16541 32413 16575
rect 32447 16572 32459 16575
rect 32582 16572 32588 16584
rect 32447 16544 32588 16572
rect 32447 16541 32459 16544
rect 32401 16535 32459 16541
rect 32582 16532 32588 16544
rect 32640 16532 32646 16584
rect 34606 16572 34612 16584
rect 34567 16544 34612 16572
rect 34606 16532 34612 16544
rect 34664 16532 34670 16584
rect 34885 16575 34943 16581
rect 34885 16541 34897 16575
rect 34931 16572 34943 16575
rect 35066 16572 35072 16584
rect 34931 16544 35072 16572
rect 34931 16541 34943 16544
rect 34885 16535 34943 16541
rect 35066 16532 35072 16544
rect 35124 16532 35130 16584
rect 37737 16575 37795 16581
rect 37737 16541 37749 16575
rect 37783 16541 37795 16575
rect 37737 16535 37795 16541
rect 38013 16575 38071 16581
rect 38013 16541 38025 16575
rect 38059 16572 38071 16575
rect 38102 16572 38108 16584
rect 38059 16544 38108 16572
rect 38059 16541 38071 16544
rect 38013 16535 38071 16541
rect 8021 16507 8079 16513
rect 8021 16473 8033 16507
rect 8067 16504 8079 16507
rect 8202 16504 8208 16516
rect 8067 16476 8208 16504
rect 8067 16473 8079 16476
rect 8021 16467 8079 16473
rect 8202 16464 8208 16476
rect 8260 16464 8266 16516
rect 8864 16476 11100 16504
rect 4798 16396 4804 16448
rect 4856 16436 4862 16448
rect 8864 16436 8892 16476
rect 9030 16436 9036 16448
rect 4856 16408 8892 16436
rect 8991 16408 9036 16436
rect 4856 16396 4862 16408
rect 9030 16396 9036 16408
rect 9088 16396 9094 16448
rect 9490 16436 9496 16448
rect 9451 16408 9496 16436
rect 9490 16396 9496 16408
rect 9548 16396 9554 16448
rect 10870 16436 10876 16448
rect 10831 16408 10876 16436
rect 10870 16396 10876 16408
rect 10928 16396 10934 16448
rect 11072 16436 11100 16476
rect 26326 16464 26332 16516
rect 26384 16504 26390 16516
rect 30098 16504 30104 16516
rect 26384 16476 27384 16504
rect 30059 16476 30104 16504
rect 26384 16464 26390 16476
rect 11974 16436 11980 16448
rect 11072 16408 11980 16436
rect 11974 16396 11980 16408
rect 12032 16396 12038 16448
rect 14274 16436 14280 16448
rect 14235 16408 14280 16436
rect 14274 16396 14280 16408
rect 14332 16396 14338 16448
rect 20346 16436 20352 16448
rect 20307 16408 20352 16436
rect 20346 16396 20352 16408
rect 20404 16396 20410 16448
rect 22554 16396 22560 16448
rect 22612 16436 22618 16448
rect 22738 16436 22744 16448
rect 22612 16408 22744 16436
rect 22612 16396 22618 16408
rect 22738 16396 22744 16408
rect 22796 16436 22802 16448
rect 23109 16439 23167 16445
rect 23109 16436 23121 16439
rect 22796 16408 23121 16436
rect 22796 16396 22802 16408
rect 23109 16405 23121 16408
rect 23155 16436 23167 16439
rect 25406 16436 25412 16448
rect 23155 16408 25412 16436
rect 23155 16405 23167 16408
rect 23109 16399 23167 16405
rect 25406 16396 25412 16408
rect 25464 16396 25470 16448
rect 26142 16396 26148 16448
rect 26200 16436 26206 16448
rect 27065 16439 27123 16445
rect 27065 16436 27077 16439
rect 26200 16408 27077 16436
rect 26200 16396 26206 16408
rect 27065 16405 27077 16408
rect 27111 16436 27123 16439
rect 27157 16439 27215 16445
rect 27157 16436 27169 16439
rect 27111 16408 27169 16436
rect 27111 16405 27123 16408
rect 27065 16399 27123 16405
rect 27157 16405 27169 16408
rect 27203 16405 27215 16439
rect 27356 16436 27384 16476
rect 30098 16464 30104 16476
rect 30156 16464 30162 16516
rect 28718 16436 28724 16448
rect 27356 16408 28724 16436
rect 27157 16399 27215 16405
rect 28718 16396 28724 16408
rect 28776 16396 28782 16448
rect 29546 16436 29552 16448
rect 29507 16408 29552 16436
rect 29546 16396 29552 16408
rect 29604 16396 29610 16448
rect 30760 16436 30788 16532
rect 31110 16436 31116 16448
rect 30760 16408 31116 16436
rect 31110 16396 31116 16408
rect 31168 16396 31174 16448
rect 32490 16396 32496 16448
rect 32548 16436 32554 16448
rect 32858 16436 32864 16448
rect 32548 16408 32864 16436
rect 32548 16396 32554 16408
rect 32858 16396 32864 16408
rect 32916 16436 32922 16448
rect 33505 16439 33563 16445
rect 33505 16436 33517 16439
rect 32916 16408 33517 16436
rect 32916 16396 32922 16408
rect 33505 16405 33517 16408
rect 33551 16436 33563 16439
rect 33686 16436 33692 16448
rect 33551 16408 33692 16436
rect 33551 16405 33563 16408
rect 33505 16399 33563 16405
rect 33686 16396 33692 16408
rect 33744 16396 33750 16448
rect 37366 16436 37372 16448
rect 37327 16408 37372 16436
rect 37366 16396 37372 16408
rect 37424 16396 37430 16448
rect 37752 16436 37780 16535
rect 38102 16532 38108 16544
rect 38160 16532 38166 16584
rect 38194 16532 38200 16584
rect 38252 16572 38258 16584
rect 39117 16575 39175 16581
rect 39117 16572 39129 16575
rect 38252 16544 39129 16572
rect 38252 16532 38258 16544
rect 39117 16541 39129 16544
rect 39163 16572 39175 16575
rect 39482 16572 39488 16584
rect 39163 16544 39488 16572
rect 39163 16541 39175 16544
rect 39117 16535 39175 16541
rect 39482 16532 39488 16544
rect 39540 16532 39546 16584
rect 40218 16572 40224 16584
rect 39776 16544 40224 16572
rect 38470 16436 38476 16448
rect 37752 16408 38476 16436
rect 38470 16396 38476 16408
rect 38528 16436 38534 16448
rect 39776 16436 39804 16544
rect 40218 16532 40224 16544
rect 40276 16532 40282 16584
rect 40497 16575 40555 16581
rect 40497 16541 40509 16575
rect 40543 16572 40555 16575
rect 40954 16572 40960 16584
rect 40543 16544 40960 16572
rect 40543 16541 40555 16544
rect 40497 16535 40555 16541
rect 40954 16532 40960 16544
rect 41012 16532 41018 16584
rect 47026 16532 47032 16584
rect 47084 16572 47090 16584
rect 47688 16572 47716 16603
rect 48222 16572 48228 16584
rect 47084 16544 48228 16572
rect 47084 16532 47090 16544
rect 48222 16532 48228 16544
rect 48280 16532 48286 16584
rect 49237 16575 49295 16581
rect 49237 16541 49249 16575
rect 49283 16572 49295 16575
rect 49418 16572 49424 16584
rect 49283 16544 49424 16572
rect 49283 16541 49295 16544
rect 49237 16535 49295 16541
rect 49418 16532 49424 16544
rect 49476 16532 49482 16584
rect 41598 16464 41604 16516
rect 41656 16504 41662 16516
rect 42521 16507 42579 16513
rect 42521 16504 42533 16507
rect 41656 16476 42533 16504
rect 41656 16464 41662 16476
rect 42521 16473 42533 16476
rect 42567 16504 42579 16507
rect 42889 16507 42947 16513
rect 42889 16504 42901 16507
rect 42567 16476 42901 16504
rect 42567 16473 42579 16476
rect 42521 16467 42579 16473
rect 42889 16473 42901 16476
rect 42935 16504 42947 16507
rect 43070 16504 43076 16516
rect 42935 16476 43076 16504
rect 42935 16473 42947 16476
rect 42889 16467 42947 16473
rect 43070 16464 43076 16476
rect 43128 16464 43134 16516
rect 47210 16464 47216 16516
rect 47268 16504 47274 16516
rect 47305 16507 47363 16513
rect 47305 16504 47317 16507
rect 47268 16476 47317 16504
rect 47268 16464 47274 16476
rect 47305 16473 47317 16476
rect 47351 16473 47363 16507
rect 48240 16504 48268 16532
rect 50632 16516 50660 16612
rect 53374 16600 53380 16652
rect 53432 16640 53438 16652
rect 54757 16643 54815 16649
rect 54757 16640 54769 16643
rect 53432 16612 54769 16640
rect 53432 16600 53438 16612
rect 54757 16609 54769 16612
rect 54803 16609 54815 16643
rect 54757 16603 54815 16609
rect 51813 16575 51871 16581
rect 51813 16541 51825 16575
rect 51859 16541 51871 16575
rect 52086 16572 52092 16584
rect 52047 16544 52092 16572
rect 51813 16535 51871 16541
rect 48240 16476 49004 16504
rect 47305 16467 47363 16473
rect 38528 16408 39804 16436
rect 38528 16396 38534 16408
rect 39850 16396 39856 16448
rect 39908 16436 39914 16448
rect 39945 16439 40003 16445
rect 39945 16436 39957 16439
rect 39908 16408 39957 16436
rect 39908 16396 39914 16408
rect 39945 16405 39957 16408
rect 39991 16436 40003 16439
rect 40678 16436 40684 16448
rect 39991 16408 40684 16436
rect 39991 16405 40003 16408
rect 39945 16399 40003 16405
rect 40678 16396 40684 16408
rect 40736 16396 40742 16448
rect 42150 16436 42156 16448
rect 42111 16408 42156 16436
rect 42150 16396 42156 16408
rect 42208 16396 42214 16448
rect 46569 16439 46627 16445
rect 46569 16405 46581 16439
rect 46615 16436 46627 16439
rect 46934 16436 46940 16448
rect 46615 16408 46940 16436
rect 46615 16405 46627 16408
rect 46569 16399 46627 16405
rect 46934 16396 46940 16408
rect 46992 16436 46998 16448
rect 47394 16436 47400 16448
rect 46992 16408 47400 16436
rect 46992 16396 46998 16408
rect 47394 16396 47400 16408
rect 47452 16396 47458 16448
rect 48314 16436 48320 16448
rect 48275 16408 48320 16436
rect 48314 16396 48320 16408
rect 48372 16396 48378 16448
rect 48976 16436 49004 16476
rect 50614 16464 50620 16516
rect 50672 16504 50678 16516
rect 51828 16504 51856 16535
rect 52086 16532 52092 16544
rect 52144 16532 52150 16584
rect 50672 16476 51856 16504
rect 50672 16464 50678 16476
rect 49694 16436 49700 16448
rect 48976 16408 49700 16436
rect 49694 16396 49700 16408
rect 49752 16436 49758 16448
rect 50338 16436 50344 16448
rect 49752 16408 50344 16436
rect 49752 16396 49758 16408
rect 50338 16396 50344 16408
rect 50396 16436 50402 16448
rect 50801 16439 50859 16445
rect 50801 16436 50813 16439
rect 50396 16408 50813 16436
rect 50396 16396 50402 16408
rect 50801 16405 50813 16408
rect 50847 16436 50859 16439
rect 50893 16439 50951 16445
rect 50893 16436 50905 16439
rect 50847 16408 50905 16436
rect 50847 16405 50859 16408
rect 50801 16399 50859 16405
rect 50893 16405 50905 16408
rect 50939 16405 50951 16439
rect 50893 16399 50951 16405
rect 51810 16396 51816 16448
rect 51868 16436 51874 16448
rect 53193 16439 53251 16445
rect 53193 16436 53205 16439
rect 51868 16408 53205 16436
rect 51868 16396 51874 16408
rect 53193 16405 53205 16408
rect 53239 16436 53251 16439
rect 53282 16436 53288 16448
rect 53239 16408 53288 16436
rect 53239 16405 53251 16408
rect 53193 16399 53251 16405
rect 53282 16396 53288 16408
rect 53340 16396 53346 16448
rect 53742 16436 53748 16448
rect 53703 16408 53748 16436
rect 53742 16396 53748 16408
rect 53800 16396 53806 16448
rect 1104 16346 63480 16368
rect 1104 16294 11378 16346
rect 11430 16294 11442 16346
rect 11494 16294 11506 16346
rect 11558 16294 11570 16346
rect 11622 16294 32170 16346
rect 32222 16294 32234 16346
rect 32286 16294 32298 16346
rect 32350 16294 32362 16346
rect 32414 16294 52962 16346
rect 53014 16294 53026 16346
rect 53078 16294 53090 16346
rect 53142 16294 53154 16346
rect 53206 16294 63480 16346
rect 1104 16272 63480 16294
rect 8110 16192 8116 16244
rect 8168 16232 8174 16244
rect 8205 16235 8263 16241
rect 8205 16232 8217 16235
rect 8168 16204 8217 16232
rect 8168 16192 8174 16204
rect 8205 16201 8217 16204
rect 8251 16232 8263 16235
rect 9861 16235 9919 16241
rect 9861 16232 9873 16235
rect 8251 16204 9873 16232
rect 8251 16201 8263 16204
rect 8205 16195 8263 16201
rect 9861 16201 9873 16204
rect 9907 16232 9919 16235
rect 10686 16232 10692 16244
rect 9907 16204 10692 16232
rect 9907 16201 9919 16204
rect 9861 16195 9919 16201
rect 10686 16192 10692 16204
rect 10744 16192 10750 16244
rect 11238 16232 11244 16244
rect 11199 16204 11244 16232
rect 11238 16192 11244 16204
rect 11296 16232 11302 16244
rect 11793 16235 11851 16241
rect 11793 16232 11805 16235
rect 11296 16204 11805 16232
rect 11296 16192 11302 16204
rect 11793 16201 11805 16204
rect 11839 16201 11851 16235
rect 12250 16232 12256 16244
rect 12211 16204 12256 16232
rect 11793 16195 11851 16201
rect 12250 16192 12256 16204
rect 12308 16192 12314 16244
rect 14642 16232 14648 16244
rect 14603 16204 14648 16232
rect 14642 16192 14648 16204
rect 14700 16192 14706 16244
rect 16022 16192 16028 16244
rect 16080 16232 16086 16244
rect 16117 16235 16175 16241
rect 16117 16232 16129 16235
rect 16080 16204 16129 16232
rect 16080 16192 16086 16204
rect 16117 16201 16129 16204
rect 16163 16232 16175 16235
rect 16761 16235 16819 16241
rect 16761 16232 16773 16235
rect 16163 16204 16773 16232
rect 16163 16201 16175 16204
rect 16117 16195 16175 16201
rect 16761 16201 16773 16204
rect 16807 16201 16819 16235
rect 16761 16195 16819 16201
rect 18046 16192 18052 16244
rect 18104 16232 18110 16244
rect 19978 16232 19984 16244
rect 18104 16204 19984 16232
rect 18104 16192 18110 16204
rect 19978 16192 19984 16204
rect 20036 16192 20042 16244
rect 20530 16192 20536 16244
rect 20588 16232 20594 16244
rect 20990 16232 20996 16244
rect 20588 16204 20996 16232
rect 20588 16192 20594 16204
rect 20990 16192 20996 16204
rect 21048 16232 21054 16244
rect 21453 16235 21511 16241
rect 21453 16232 21465 16235
rect 21048 16204 21465 16232
rect 21048 16192 21054 16204
rect 21453 16201 21465 16204
rect 21499 16201 21511 16235
rect 49694 16232 49700 16244
rect 21453 16195 21511 16201
rect 21560 16204 49556 16232
rect 49655 16204 49700 16232
rect 19794 16164 19800 16176
rect 9232 16136 19800 16164
rect 8573 16099 8631 16105
rect 6288 16068 8432 16096
rect 934 15852 940 15904
rect 992 15892 998 15904
rect 3602 15892 3608 15904
rect 992 15864 3608 15892
rect 992 15852 998 15864
rect 3602 15852 3608 15864
rect 3660 15892 3666 15904
rect 6288 15892 6316 16068
rect 8297 16031 8355 16037
rect 8297 16028 8309 16031
rect 7392 16000 8309 16028
rect 3660 15864 6316 15892
rect 3660 15852 3666 15864
rect 7282 15852 7288 15904
rect 7340 15892 7346 15904
rect 7392 15901 7420 16000
rect 8297 15997 8309 16000
rect 8343 15997 8355 16031
rect 8404 16028 8432 16068
rect 8573 16065 8585 16099
rect 8619 16096 8631 16099
rect 9030 16096 9036 16108
rect 8619 16068 9036 16096
rect 8619 16065 8631 16068
rect 8573 16059 8631 16065
rect 9030 16056 9036 16068
rect 9088 16056 9094 16108
rect 9232 16028 9260 16136
rect 19794 16124 19800 16136
rect 19852 16124 19858 16176
rect 21082 16124 21088 16176
rect 21140 16164 21146 16176
rect 21560 16164 21588 16204
rect 21140 16136 21588 16164
rect 21140 16124 21146 16136
rect 22370 16124 22376 16176
rect 22428 16164 22434 16176
rect 22465 16167 22523 16173
rect 22465 16164 22477 16167
rect 22428 16136 22477 16164
rect 22428 16124 22434 16136
rect 22465 16133 22477 16136
rect 22511 16164 22523 16167
rect 22554 16164 22560 16176
rect 22511 16136 22560 16164
rect 22511 16133 22523 16136
rect 22465 16127 22523 16133
rect 22554 16124 22560 16136
rect 22612 16124 22618 16176
rect 25406 16164 25412 16176
rect 25367 16136 25412 16164
rect 25406 16124 25412 16136
rect 25464 16124 25470 16176
rect 27525 16167 27583 16173
rect 27525 16133 27537 16167
rect 27571 16164 27583 16167
rect 27614 16164 27620 16176
rect 27571 16136 27620 16164
rect 27571 16133 27583 16136
rect 27525 16127 27583 16133
rect 27614 16124 27620 16136
rect 27672 16124 27678 16176
rect 29270 16164 29276 16176
rect 27724 16136 29276 16164
rect 10321 16099 10379 16105
rect 10321 16065 10333 16099
rect 10367 16096 10379 16099
rect 14642 16096 14648 16108
rect 10367 16068 11100 16096
rect 10367 16065 10379 16068
rect 10321 16059 10379 16065
rect 10870 16028 10876 16040
rect 8404 16000 9260 16028
rect 10831 16000 10876 16028
rect 8297 15991 8355 15997
rect 10870 15988 10876 16000
rect 10928 15988 10934 16040
rect 11072 16037 11100 16068
rect 13832 16068 14648 16096
rect 11057 16031 11115 16037
rect 11057 15997 11069 16031
rect 11103 16028 11115 16031
rect 12250 16028 12256 16040
rect 11103 16000 12256 16028
rect 11103 15997 11115 16000
rect 11057 15991 11115 15997
rect 12250 15988 12256 16000
rect 12308 15988 12314 16040
rect 13832 16037 13860 16068
rect 14642 16056 14648 16068
rect 14700 16056 14706 16108
rect 16301 16099 16359 16105
rect 16301 16065 16313 16099
rect 16347 16096 16359 16099
rect 16758 16096 16764 16108
rect 16347 16068 16764 16096
rect 16347 16065 16359 16068
rect 16301 16059 16359 16065
rect 16758 16056 16764 16068
rect 16816 16056 16822 16108
rect 17034 16056 17040 16108
rect 17092 16096 17098 16108
rect 17773 16099 17831 16105
rect 17773 16096 17785 16099
rect 17092 16068 17785 16096
rect 17092 16056 17098 16068
rect 17773 16065 17785 16068
rect 17819 16096 17831 16099
rect 18046 16096 18052 16108
rect 17819 16068 18052 16096
rect 17819 16065 17831 16068
rect 17773 16059 17831 16065
rect 18046 16056 18052 16068
rect 18104 16056 18110 16108
rect 19337 16099 19395 16105
rect 19337 16096 19349 16099
rect 18524 16068 19349 16096
rect 13817 16031 13875 16037
rect 13817 15997 13829 16031
rect 13863 15997 13875 16031
rect 13817 15991 13875 15997
rect 14185 16031 14243 16037
rect 14185 15997 14197 16031
rect 14231 15997 14243 16031
rect 14185 15991 14243 15997
rect 10689 15963 10747 15969
rect 10689 15929 10701 15963
rect 10735 15960 10747 15963
rect 10965 15963 11023 15969
rect 10965 15960 10977 15963
rect 10735 15932 10977 15960
rect 10735 15929 10747 15932
rect 10689 15923 10747 15929
rect 10965 15929 10977 15932
rect 11011 15960 11023 15963
rect 11146 15960 11152 15972
rect 11011 15932 11152 15960
rect 11011 15929 11023 15932
rect 10965 15923 11023 15929
rect 11146 15920 11152 15932
rect 11204 15920 11210 15972
rect 13354 15960 13360 15972
rect 13315 15932 13360 15960
rect 13354 15920 13360 15932
rect 13412 15920 13418 15972
rect 7377 15895 7435 15901
rect 7377 15892 7389 15895
rect 7340 15864 7389 15892
rect 7340 15852 7346 15864
rect 7377 15861 7389 15864
rect 7423 15861 7435 15895
rect 7377 15855 7435 15861
rect 7837 15895 7895 15901
rect 7837 15861 7849 15895
rect 7883 15892 7895 15895
rect 7926 15892 7932 15904
rect 7883 15864 7932 15892
rect 7883 15861 7895 15864
rect 7837 15855 7895 15861
rect 7926 15852 7932 15864
rect 7984 15852 7990 15904
rect 13262 15852 13268 15904
rect 13320 15892 13326 15904
rect 14200 15892 14228 15991
rect 14274 15988 14280 16040
rect 14332 16028 14338 16040
rect 14332 16000 14377 16028
rect 14332 15988 14338 16000
rect 16390 15988 16396 16040
rect 16448 16028 16454 16040
rect 16577 16031 16635 16037
rect 16577 16028 16589 16031
rect 16448 16000 16589 16028
rect 16448 15988 16454 16000
rect 16577 15997 16589 16000
rect 16623 15997 16635 16031
rect 16577 15991 16635 15997
rect 17126 15988 17132 16040
rect 17184 16028 17190 16040
rect 18524 16037 18552 16068
rect 19337 16065 19349 16068
rect 19383 16065 19395 16099
rect 19337 16059 19395 16065
rect 23109 16099 23167 16105
rect 23109 16065 23121 16099
rect 23155 16096 23167 16099
rect 23155 16068 23796 16096
rect 23155 16065 23167 16068
rect 23109 16059 23167 16065
rect 18509 16031 18567 16037
rect 18509 16028 18521 16031
rect 17184 16000 18521 16028
rect 17184 15988 17190 16000
rect 18509 15997 18521 16000
rect 18555 15997 18567 16031
rect 18509 15991 18567 15997
rect 18877 16031 18935 16037
rect 18877 15997 18889 16031
rect 18923 15997 18935 16031
rect 18877 15991 18935 15997
rect 18969 16031 19027 16037
rect 18969 15997 18981 16031
rect 19015 16028 19027 16031
rect 19150 16028 19156 16040
rect 19015 16000 19156 16028
rect 19015 15997 19027 16000
rect 18969 15991 19027 15997
rect 16485 15963 16543 15969
rect 16485 15929 16497 15963
rect 16531 15929 16543 15963
rect 16485 15923 16543 15929
rect 17405 15963 17463 15969
rect 17405 15929 17417 15963
rect 17451 15960 17463 15963
rect 18049 15963 18107 15969
rect 18049 15960 18061 15963
rect 17451 15932 18061 15960
rect 17451 15929 17463 15932
rect 17405 15923 17463 15929
rect 18049 15929 18061 15932
rect 18095 15929 18107 15963
rect 18892 15960 18920 15991
rect 19150 15988 19156 16000
rect 19208 15988 19214 16040
rect 19981 16031 20039 16037
rect 19981 15997 19993 16031
rect 20027 16028 20039 16031
rect 20073 16031 20131 16037
rect 20073 16028 20085 16031
rect 20027 16000 20085 16028
rect 20027 15997 20039 16000
rect 19981 15991 20039 15997
rect 20073 15997 20085 16000
rect 20119 15997 20131 16031
rect 20346 16028 20352 16040
rect 20307 16000 20352 16028
rect 20073 15991 20131 15997
rect 20346 15988 20352 16000
rect 20404 15988 20410 16040
rect 23658 16028 23664 16040
rect 23619 16000 23664 16028
rect 23658 15988 23664 16000
rect 23716 15988 23722 16040
rect 23768 16028 23796 16068
rect 23842 16056 23848 16108
rect 23900 16096 23906 16108
rect 24397 16099 24455 16105
rect 24397 16096 24409 16099
rect 23900 16068 24409 16096
rect 23900 16056 23906 16068
rect 24397 16065 24409 16068
rect 24443 16096 24455 16099
rect 24673 16099 24731 16105
rect 24673 16096 24685 16099
rect 24443 16068 24685 16096
rect 24443 16065 24455 16068
rect 24397 16059 24455 16065
rect 24673 16065 24685 16068
rect 24719 16065 24731 16099
rect 25038 16096 25044 16108
rect 24999 16068 25044 16096
rect 24673 16059 24731 16065
rect 25038 16056 25044 16068
rect 25096 16096 25102 16108
rect 26142 16096 26148 16108
rect 25096 16068 26148 16096
rect 25096 16056 25102 16068
rect 26142 16056 26148 16068
rect 26200 16096 26206 16108
rect 26697 16099 26755 16105
rect 26697 16096 26709 16099
rect 26200 16068 26709 16096
rect 26200 16056 26206 16068
rect 26697 16065 26709 16068
rect 26743 16065 26755 16099
rect 26697 16059 26755 16065
rect 23937 16031 23995 16037
rect 23937 16028 23949 16031
rect 23768 16000 23949 16028
rect 23937 15997 23949 16000
rect 23983 15997 23995 16031
rect 23937 15991 23995 15997
rect 18892 15932 19840 15960
rect 18049 15923 18107 15929
rect 15013 15895 15071 15901
rect 15013 15892 15025 15895
rect 13320 15864 15025 15892
rect 13320 15852 13326 15864
rect 15013 15861 15025 15864
rect 15059 15892 15071 15895
rect 15562 15892 15568 15904
rect 15059 15864 15568 15892
rect 15059 15861 15071 15864
rect 15013 15855 15071 15861
rect 15562 15852 15568 15864
rect 15620 15852 15626 15904
rect 15746 15892 15752 15904
rect 15707 15864 15752 15892
rect 15746 15852 15752 15864
rect 15804 15852 15810 15904
rect 16500 15892 16528 15923
rect 17420 15892 17448 15923
rect 19812 15901 19840 15932
rect 22094 15920 22100 15972
rect 22152 15960 22158 15972
rect 22554 15960 22560 15972
rect 22152 15932 22560 15960
rect 22152 15920 22158 15932
rect 22554 15920 22560 15932
rect 22612 15920 22618 15972
rect 23566 15920 23572 15972
rect 23624 15960 23630 15972
rect 23845 15963 23903 15969
rect 23845 15960 23857 15963
rect 23624 15932 23857 15960
rect 23624 15920 23630 15932
rect 23845 15929 23857 15932
rect 23891 15929 23903 15963
rect 23952 15960 23980 15991
rect 24118 15988 24124 16040
rect 24176 16028 24182 16040
rect 25225 16031 25283 16037
rect 25225 16028 25237 16031
rect 24176 16000 25237 16028
rect 24176 15988 24182 16000
rect 25225 15997 25237 16000
rect 25271 16028 25283 16031
rect 25777 16031 25835 16037
rect 25777 16028 25789 16031
rect 25271 16000 25789 16028
rect 25271 15997 25283 16000
rect 25225 15991 25283 15997
rect 25777 15997 25789 16000
rect 25823 16028 25835 16031
rect 26970 16028 26976 16040
rect 25823 16000 26976 16028
rect 25823 15997 25835 16000
rect 25777 15991 25835 15997
rect 26970 15988 26976 16000
rect 27028 15988 27034 16040
rect 27062 15988 27068 16040
rect 27120 16028 27126 16040
rect 27724 16037 27752 16136
rect 29270 16124 29276 16136
rect 29328 16124 29334 16176
rect 30282 16124 30288 16176
rect 30340 16164 30346 16176
rect 30653 16167 30711 16173
rect 30653 16164 30665 16167
rect 30340 16136 30665 16164
rect 30340 16124 30346 16136
rect 30653 16133 30665 16136
rect 30699 16133 30711 16167
rect 30653 16127 30711 16133
rect 30742 16124 30748 16176
rect 30800 16164 30806 16176
rect 32674 16164 32680 16176
rect 30800 16136 32680 16164
rect 30800 16124 30806 16136
rect 32674 16124 32680 16136
rect 32732 16164 32738 16176
rect 33686 16164 33692 16176
rect 32732 16136 33456 16164
rect 33647 16136 33692 16164
rect 32732 16124 32738 16136
rect 28350 16096 28356 16108
rect 28311 16068 28356 16096
rect 28350 16056 28356 16068
rect 28408 16056 28414 16108
rect 33318 16096 33324 16108
rect 31220 16068 32996 16096
rect 33279 16068 33324 16096
rect 27157 16031 27215 16037
rect 27157 16028 27169 16031
rect 27120 16000 27169 16028
rect 27120 15988 27126 16000
rect 27157 15997 27169 16000
rect 27203 16028 27215 16031
rect 27709 16031 27767 16037
rect 27709 16028 27721 16031
rect 27203 16000 27721 16028
rect 27203 15997 27215 16000
rect 27157 15991 27215 15997
rect 27709 15997 27721 16000
rect 27755 15997 27767 16031
rect 27709 15991 27767 15997
rect 27893 16031 27951 16037
rect 27893 15997 27905 16031
rect 27939 16028 27951 16031
rect 28258 16028 28264 16040
rect 27939 16000 28264 16028
rect 27939 15997 27951 16000
rect 27893 15991 27951 15997
rect 28258 15988 28264 16000
rect 28316 16028 28322 16040
rect 28997 16031 29055 16037
rect 28997 16028 29009 16031
rect 28316 16000 29009 16028
rect 28316 15988 28322 16000
rect 28997 15997 29009 16000
rect 29043 15997 29055 16031
rect 28997 15991 29055 15997
rect 29273 16031 29331 16037
rect 29273 15997 29285 16031
rect 29319 16028 29331 16031
rect 29362 16028 29368 16040
rect 29319 16000 29368 16028
rect 29319 15997 29331 16000
rect 29273 15991 29331 15997
rect 29362 15988 29368 16000
rect 29420 15988 29426 16040
rect 29546 16028 29552 16040
rect 29507 16000 29552 16028
rect 29546 15988 29552 16000
rect 29604 15988 29610 16040
rect 27801 15963 27859 15969
rect 23952 15932 27752 15960
rect 23845 15923 23903 15929
rect 27724 15904 27752 15932
rect 27801 15929 27813 15963
rect 27847 15929 27859 15963
rect 27801 15923 27859 15929
rect 16500 15864 17448 15892
rect 19797 15895 19855 15901
rect 19797 15861 19809 15895
rect 19843 15892 19855 15895
rect 20438 15892 20444 15904
rect 19843 15864 20444 15892
rect 19843 15861 19855 15864
rect 19797 15855 19855 15861
rect 20438 15852 20444 15864
rect 20496 15852 20502 15904
rect 23477 15895 23535 15901
rect 23477 15861 23489 15895
rect 23523 15892 23535 15895
rect 23658 15892 23664 15904
rect 23523 15864 23664 15892
rect 23523 15861 23535 15864
rect 23477 15855 23535 15861
rect 23658 15852 23664 15864
rect 23716 15852 23722 15904
rect 27706 15852 27712 15904
rect 27764 15852 27770 15904
rect 27816 15892 27844 15923
rect 28534 15892 28540 15904
rect 27816 15864 28540 15892
rect 28534 15852 28540 15864
rect 28592 15892 28598 15904
rect 28629 15895 28687 15901
rect 28629 15892 28641 15895
rect 28592 15864 28641 15892
rect 28592 15852 28598 15864
rect 28629 15861 28641 15864
rect 28675 15861 28687 15895
rect 28629 15855 28687 15861
rect 29362 15852 29368 15904
rect 29420 15892 29426 15904
rect 30650 15892 30656 15904
rect 29420 15864 30656 15892
rect 29420 15852 29426 15864
rect 30650 15852 30656 15864
rect 30708 15892 30714 15904
rect 31220 15901 31248 16068
rect 32858 16028 32864 16040
rect 32819 16000 32864 16028
rect 32858 15988 32864 16000
rect 32916 15988 32922 16040
rect 32968 16028 32996 16068
rect 33318 16056 33324 16068
rect 33376 16056 33382 16108
rect 33428 16096 33456 16136
rect 33686 16124 33692 16136
rect 33744 16124 33750 16176
rect 35710 16124 35716 16176
rect 35768 16164 35774 16176
rect 39761 16167 39819 16173
rect 39761 16164 39773 16167
rect 35768 16136 39773 16164
rect 35768 16124 35774 16136
rect 39761 16133 39773 16136
rect 39807 16133 39819 16167
rect 39761 16127 39819 16133
rect 39945 16167 40003 16173
rect 39945 16133 39957 16167
rect 39991 16164 40003 16167
rect 40126 16164 40132 16176
rect 39991 16136 40132 16164
rect 39991 16133 40003 16136
rect 39945 16127 40003 16133
rect 39960 16096 39988 16127
rect 40126 16124 40132 16136
rect 40184 16124 40190 16176
rect 43438 16164 43444 16176
rect 43351 16136 43444 16164
rect 43438 16124 43444 16136
rect 43496 16164 43502 16176
rect 43990 16164 43996 16176
rect 43496 16136 43996 16164
rect 43496 16124 43502 16136
rect 43990 16124 43996 16136
rect 44048 16124 44054 16176
rect 46385 16167 46443 16173
rect 46385 16133 46397 16167
rect 46431 16164 46443 16167
rect 47026 16164 47032 16176
rect 46431 16136 47032 16164
rect 46431 16133 46443 16136
rect 46385 16127 46443 16133
rect 47026 16124 47032 16136
rect 47084 16124 47090 16176
rect 47213 16167 47271 16173
rect 47213 16133 47225 16167
rect 47259 16164 47271 16167
rect 47302 16164 47308 16176
rect 47259 16136 47308 16164
rect 47259 16133 47271 16136
rect 47213 16127 47271 16133
rect 47302 16124 47308 16136
rect 47360 16124 47366 16176
rect 33428 16068 37412 16096
rect 37384 16040 37412 16068
rect 39040 16068 39988 16096
rect 33229 16031 33287 16037
rect 33229 16028 33241 16031
rect 32968 16000 33241 16028
rect 33229 15997 33241 16000
rect 33275 16028 33287 16031
rect 34057 16031 34115 16037
rect 34057 16028 34069 16031
rect 33275 16000 34069 16028
rect 33275 15997 33287 16000
rect 33229 15991 33287 15997
rect 34057 15997 34069 16000
rect 34103 16028 34115 16031
rect 34330 16028 34336 16040
rect 34103 16000 34336 16028
rect 34103 15997 34115 16000
rect 34057 15991 34115 15997
rect 34330 15988 34336 16000
rect 34388 15988 34394 16040
rect 34885 16031 34943 16037
rect 34885 15997 34897 16031
rect 34931 16028 34943 16031
rect 36449 16031 36507 16037
rect 36449 16028 36461 16031
rect 34931 16000 36461 16028
rect 34931 15997 34943 16000
rect 34885 15991 34943 15997
rect 36449 15997 36461 16000
rect 36495 16028 36507 16031
rect 37185 16031 37243 16037
rect 37185 16028 37197 16031
rect 36495 16000 37197 16028
rect 36495 15997 36507 16000
rect 36449 15991 36507 15997
rect 37185 15997 37197 16000
rect 37231 15997 37243 16031
rect 37366 16028 37372 16040
rect 37327 16000 37372 16028
rect 37185 15991 37243 15997
rect 37366 15988 37372 16000
rect 37424 15988 37430 16040
rect 38930 16028 38936 16040
rect 37476 16000 38936 16028
rect 32306 15920 32312 15972
rect 32364 15960 32370 15972
rect 32401 15963 32459 15969
rect 32401 15960 32413 15963
rect 32364 15932 32413 15960
rect 32364 15920 32370 15932
rect 32401 15929 32413 15932
rect 32447 15929 32459 15963
rect 32401 15923 32459 15929
rect 33686 15920 33692 15972
rect 33744 15960 33750 15972
rect 37476 15960 37504 16000
rect 38930 15988 38936 16000
rect 38988 15988 38994 16040
rect 39040 16037 39068 16068
rect 41598 16056 41604 16108
rect 41656 16096 41662 16108
rect 41877 16099 41935 16105
rect 41877 16096 41889 16099
rect 41656 16068 41889 16096
rect 41656 16056 41662 16068
rect 41877 16065 41889 16068
rect 41923 16065 41935 16099
rect 47581 16099 47639 16105
rect 41877 16059 41935 16065
rect 41984 16068 47532 16096
rect 39025 16031 39083 16037
rect 39025 15997 39037 16031
rect 39071 15997 39083 16031
rect 39206 16028 39212 16040
rect 39167 16000 39212 16028
rect 39025 15991 39083 15997
rect 39206 15988 39212 16000
rect 39264 15988 39270 16040
rect 39393 16031 39451 16037
rect 39393 15997 39405 16031
rect 39439 15997 39451 16031
rect 39393 15991 39451 15997
rect 39761 16031 39819 16037
rect 39761 15997 39773 16031
rect 39807 16028 39819 16031
rect 40313 16031 40371 16037
rect 40313 16028 40325 16031
rect 39807 16000 40325 16028
rect 39807 15997 39819 16000
rect 39761 15991 39819 15997
rect 40313 15997 40325 16000
rect 40359 16028 40371 16031
rect 40497 16031 40555 16037
rect 40497 16028 40509 16031
rect 40359 16000 40509 16028
rect 40359 15997 40371 16000
rect 40313 15991 40371 15997
rect 40497 15997 40509 16000
rect 40543 16028 40555 16031
rect 41984 16028 42012 16068
rect 42150 16028 42156 16040
rect 40543 16000 42012 16028
rect 42111 16000 42156 16028
rect 40543 15997 40555 16000
rect 40497 15991 40555 15997
rect 33744 15932 37504 15960
rect 38565 15963 38623 15969
rect 33744 15920 33750 15932
rect 38565 15929 38577 15963
rect 38611 15960 38623 15963
rect 38654 15960 38660 15972
rect 38611 15932 38660 15960
rect 38611 15929 38623 15932
rect 38565 15923 38623 15929
rect 38654 15920 38660 15932
rect 38712 15920 38718 15972
rect 39408 15960 39436 15991
rect 42150 15988 42156 16000
rect 42208 15988 42214 16040
rect 46198 16028 46204 16040
rect 46159 16000 46204 16028
rect 46198 15988 46204 16000
rect 46256 16028 46262 16040
rect 46750 16028 46756 16040
rect 46256 16000 46756 16028
rect 46256 15988 46262 16000
rect 46750 15988 46756 16000
rect 46808 15988 46814 16040
rect 47305 16031 47363 16037
rect 47305 15997 47317 16031
rect 47351 16028 47363 16031
rect 47394 16028 47400 16040
rect 47351 16000 47400 16028
rect 47351 15997 47363 16000
rect 47305 15991 47363 15997
rect 47394 15988 47400 16000
rect 47452 15988 47458 16040
rect 47504 16028 47532 16068
rect 47581 16065 47593 16099
rect 47627 16096 47639 16099
rect 48314 16096 48320 16108
rect 47627 16068 48320 16096
rect 47627 16065 47639 16068
rect 47581 16059 47639 16065
rect 48314 16056 48320 16068
rect 48372 16056 48378 16108
rect 49528 16096 49556 16204
rect 49694 16192 49700 16204
rect 49752 16192 49758 16244
rect 52086 16192 52092 16244
rect 52144 16232 52150 16244
rect 52181 16235 52239 16241
rect 52181 16232 52193 16235
rect 52144 16204 52193 16232
rect 52144 16192 52150 16204
rect 52181 16201 52193 16204
rect 52227 16232 52239 16235
rect 52733 16235 52791 16241
rect 52733 16232 52745 16235
rect 52227 16204 52745 16232
rect 52227 16201 52239 16204
rect 52181 16195 52239 16201
rect 52733 16201 52745 16204
rect 52779 16201 52791 16235
rect 52733 16195 52791 16201
rect 53926 16192 53932 16244
rect 53984 16232 53990 16244
rect 54665 16235 54723 16241
rect 54665 16232 54677 16235
rect 53984 16204 54677 16232
rect 53984 16192 53990 16204
rect 54665 16201 54677 16204
rect 54711 16201 54723 16235
rect 54665 16195 54723 16201
rect 49973 16167 50031 16173
rect 49973 16133 49985 16167
rect 50019 16164 50031 16167
rect 51626 16164 51632 16176
rect 50019 16136 51632 16164
rect 50019 16133 50031 16136
rect 49973 16127 50031 16133
rect 51626 16124 51632 16136
rect 51684 16124 51690 16176
rect 53561 16099 53619 16105
rect 49528 16068 53420 16096
rect 49789 16031 49847 16037
rect 49789 16028 49801 16031
rect 47504 16000 49801 16028
rect 49789 15997 49801 16000
rect 49835 16028 49847 16031
rect 50341 16031 50399 16037
rect 50341 16028 50353 16031
rect 49835 16000 50353 16028
rect 49835 15997 49847 16000
rect 49789 15991 49847 15997
rect 50341 15997 50353 16000
rect 50387 16028 50399 16031
rect 51442 16028 51448 16040
rect 50387 16000 51448 16028
rect 50387 15997 50399 16000
rect 50341 15991 50399 15997
rect 51442 15988 51448 16000
rect 51500 15988 51506 16040
rect 51534 15988 51540 16040
rect 51592 16028 51598 16040
rect 51721 16031 51779 16037
rect 51721 16028 51733 16031
rect 51592 16000 51733 16028
rect 51592 15988 51598 16000
rect 51721 15997 51733 16000
rect 51767 15997 51779 16031
rect 51721 15991 51779 15997
rect 51997 16031 52055 16037
rect 51997 15997 52009 16031
rect 52043 16028 52055 16031
rect 52454 16028 52460 16040
rect 52043 16000 52460 16028
rect 52043 15997 52055 16000
rect 51997 15991 52055 15997
rect 52454 15988 52460 16000
rect 52512 15988 52518 16040
rect 53285 16031 53343 16037
rect 53285 15997 53297 16031
rect 53331 15997 53343 16031
rect 53392 16028 53420 16068
rect 53561 16065 53573 16099
rect 53607 16096 53619 16099
rect 53742 16096 53748 16108
rect 53607 16068 53748 16096
rect 53607 16065 53619 16068
rect 53561 16059 53619 16065
rect 53742 16056 53748 16068
rect 53800 16056 53806 16108
rect 57146 16028 57152 16040
rect 53392 16000 57152 16028
rect 53285 15991 53343 15997
rect 51905 15963 51963 15969
rect 39408 15932 40724 15960
rect 31205 15895 31263 15901
rect 31205 15892 31217 15895
rect 30708 15864 31217 15892
rect 30708 15852 30714 15864
rect 31205 15861 31217 15864
rect 31251 15861 31263 15895
rect 31938 15892 31944 15904
rect 31899 15864 31944 15892
rect 31205 15855 31263 15861
rect 31938 15852 31944 15864
rect 31996 15852 32002 15904
rect 32217 15895 32275 15901
rect 32217 15861 32229 15895
rect 32263 15892 32275 15895
rect 32582 15892 32588 15904
rect 32263 15864 32588 15892
rect 32263 15861 32275 15864
rect 32217 15855 32275 15861
rect 32582 15852 32588 15864
rect 32640 15852 32646 15904
rect 32766 15852 32772 15904
rect 32824 15892 32830 15904
rect 34606 15892 34612 15904
rect 32824 15864 34612 15892
rect 32824 15852 32830 15864
rect 34606 15852 34612 15864
rect 34664 15892 34670 15904
rect 34885 15895 34943 15901
rect 34885 15892 34897 15895
rect 34664 15864 34897 15892
rect 34664 15852 34670 15864
rect 34885 15861 34897 15864
rect 34931 15861 34943 15895
rect 35066 15892 35072 15904
rect 35027 15864 35072 15892
rect 34885 15855 34943 15861
rect 35066 15852 35072 15864
rect 35124 15852 35130 15904
rect 35529 15895 35587 15901
rect 35529 15861 35541 15895
rect 35575 15892 35587 15895
rect 35618 15892 35624 15904
rect 35575 15864 35624 15892
rect 35575 15861 35587 15864
rect 35529 15855 35587 15861
rect 35618 15852 35624 15864
rect 35676 15852 35682 15904
rect 35894 15852 35900 15904
rect 35952 15892 35958 15904
rect 35989 15895 36047 15901
rect 35989 15892 36001 15895
rect 35952 15864 36001 15892
rect 35952 15852 35958 15864
rect 35989 15861 36001 15864
rect 36035 15861 36047 15895
rect 35989 15855 36047 15861
rect 37553 15895 37611 15901
rect 37553 15861 37565 15895
rect 37599 15892 37611 15895
rect 37918 15892 37924 15904
rect 37599 15864 37924 15892
rect 37599 15861 37611 15864
rect 37553 15855 37611 15861
rect 37918 15852 37924 15864
rect 37976 15852 37982 15904
rect 38102 15892 38108 15904
rect 38063 15864 38108 15892
rect 38102 15852 38108 15864
rect 38160 15852 38166 15904
rect 38473 15895 38531 15901
rect 38473 15861 38485 15895
rect 38519 15892 38531 15895
rect 39408 15892 39436 15932
rect 40696 15901 40724 15932
rect 51905 15929 51917 15963
rect 51951 15929 51963 15963
rect 51905 15923 51963 15929
rect 38519 15864 39436 15892
rect 40681 15895 40739 15901
rect 38519 15861 38531 15864
rect 38473 15855 38531 15861
rect 40681 15861 40693 15895
rect 40727 15892 40739 15895
rect 40770 15892 40776 15904
rect 40727 15864 40776 15892
rect 40727 15861 40739 15864
rect 40681 15855 40739 15861
rect 40770 15852 40776 15864
rect 40828 15852 40834 15904
rect 41046 15892 41052 15904
rect 41007 15864 41052 15892
rect 41046 15852 41052 15864
rect 41104 15852 41110 15904
rect 41598 15892 41604 15904
rect 41559 15864 41604 15892
rect 41598 15852 41604 15864
rect 41656 15852 41662 15904
rect 47946 15852 47952 15904
rect 48004 15892 48010 15904
rect 48685 15895 48743 15901
rect 48685 15892 48697 15895
rect 48004 15864 48697 15892
rect 48004 15852 48010 15864
rect 48685 15861 48697 15864
rect 48731 15861 48743 15895
rect 48685 15855 48743 15861
rect 49329 15895 49387 15901
rect 49329 15861 49341 15895
rect 49375 15892 49387 15895
rect 49418 15892 49424 15904
rect 49375 15864 49424 15892
rect 49375 15861 49387 15864
rect 49329 15855 49387 15861
rect 49418 15852 49424 15864
rect 49476 15852 49482 15904
rect 50614 15852 50620 15904
rect 50672 15892 50678 15904
rect 50709 15895 50767 15901
rect 50709 15892 50721 15895
rect 50672 15864 50721 15892
rect 50672 15852 50678 15864
rect 50709 15861 50721 15864
rect 50755 15861 50767 15895
rect 50709 15855 50767 15861
rect 50982 15852 50988 15904
rect 51040 15892 51046 15904
rect 51074 15892 51080 15904
rect 51040 15864 51080 15892
rect 51040 15852 51046 15864
rect 51074 15852 51080 15864
rect 51132 15852 51138 15904
rect 51169 15895 51227 15901
rect 51169 15861 51181 15895
rect 51215 15892 51227 15895
rect 51920 15892 51948 15923
rect 52638 15892 52644 15904
rect 51215 15864 52644 15892
rect 51215 15861 51227 15864
rect 51169 15855 51227 15861
rect 52638 15852 52644 15864
rect 52696 15852 52702 15904
rect 53193 15895 53251 15901
rect 53193 15861 53205 15895
rect 53239 15892 53251 15895
rect 53300 15892 53328 15991
rect 57146 15988 57152 16000
rect 57204 15988 57210 16040
rect 53374 15892 53380 15904
rect 53239 15864 53380 15892
rect 53239 15861 53251 15864
rect 53193 15855 53251 15861
rect 53374 15852 53380 15864
rect 53432 15852 53438 15904
rect 56962 15852 56968 15904
rect 57020 15892 57026 15904
rect 57517 15895 57575 15901
rect 57517 15892 57529 15895
rect 57020 15864 57529 15892
rect 57020 15852 57026 15864
rect 57517 15861 57529 15864
rect 57563 15861 57575 15895
rect 57517 15855 57575 15861
rect 1104 15802 63480 15824
rect 1104 15750 21774 15802
rect 21826 15750 21838 15802
rect 21890 15750 21902 15802
rect 21954 15750 21966 15802
rect 22018 15750 42566 15802
rect 42618 15750 42630 15802
rect 42682 15750 42694 15802
rect 42746 15750 42758 15802
rect 42810 15750 63480 15802
rect 1104 15728 63480 15750
rect 6730 15648 6736 15700
rect 6788 15688 6794 15700
rect 6917 15691 6975 15697
rect 6917 15688 6929 15691
rect 6788 15660 6929 15688
rect 6788 15648 6794 15660
rect 6917 15657 6929 15660
rect 6963 15688 6975 15691
rect 7834 15688 7840 15700
rect 6963 15660 7840 15688
rect 6963 15657 6975 15660
rect 6917 15651 6975 15657
rect 7834 15648 7840 15660
rect 7892 15648 7898 15700
rect 9125 15691 9183 15697
rect 9125 15688 9137 15691
rect 8220 15660 9137 15688
rect 8220 15632 8248 15660
rect 9125 15657 9137 15660
rect 9171 15657 9183 15691
rect 9125 15651 9183 15657
rect 10870 15648 10876 15700
rect 10928 15688 10934 15700
rect 10928 15660 13308 15688
rect 10928 15648 10934 15660
rect 8202 15620 8208 15632
rect 8163 15592 8208 15620
rect 8202 15580 8208 15592
rect 8260 15580 8266 15632
rect 8757 15623 8815 15629
rect 8757 15589 8769 15623
rect 8803 15620 8815 15623
rect 9030 15620 9036 15632
rect 8803 15592 9036 15620
rect 8803 15589 8815 15592
rect 8757 15583 8815 15589
rect 9030 15580 9036 15592
rect 9088 15580 9094 15632
rect 8294 15552 8300 15564
rect 8255 15524 8300 15552
rect 8294 15512 8300 15524
rect 8352 15512 8358 15564
rect 10321 15555 10379 15561
rect 10321 15521 10333 15555
rect 10367 15552 10379 15555
rect 10965 15555 11023 15561
rect 10965 15552 10977 15555
rect 10367 15524 10977 15552
rect 10367 15521 10379 15524
rect 10321 15515 10379 15521
rect 10965 15521 10977 15524
rect 11011 15552 11023 15555
rect 12158 15552 12164 15564
rect 11011 15524 12164 15552
rect 11011 15521 11023 15524
rect 10965 15515 11023 15521
rect 5350 15484 5356 15496
rect 5311 15456 5356 15484
rect 5350 15444 5356 15456
rect 5408 15444 5414 15496
rect 5626 15484 5632 15496
rect 5587 15456 5632 15484
rect 5626 15444 5632 15456
rect 5684 15444 5690 15496
rect 7282 15444 7288 15496
rect 7340 15484 7346 15496
rect 10336 15484 10364 15515
rect 12158 15512 12164 15524
rect 12216 15512 12222 15564
rect 13280 15552 13308 15660
rect 14274 15648 14280 15700
rect 14332 15688 14338 15700
rect 15473 15691 15531 15697
rect 15473 15688 15485 15691
rect 14332 15660 15485 15688
rect 14332 15648 14338 15660
rect 15473 15657 15485 15660
rect 15519 15657 15531 15691
rect 19150 15688 19156 15700
rect 19111 15660 19156 15688
rect 15473 15651 15531 15657
rect 19150 15648 19156 15660
rect 19208 15648 19214 15700
rect 23477 15691 23535 15697
rect 23477 15688 23489 15691
rect 19628 15660 23489 15688
rect 13354 15580 13360 15632
rect 13412 15620 13418 15632
rect 13633 15623 13691 15629
rect 13633 15620 13645 15623
rect 13412 15592 13645 15620
rect 13412 15580 13418 15592
rect 13633 15589 13645 15592
rect 13679 15620 13691 15623
rect 14461 15623 14519 15629
rect 14461 15620 14473 15623
rect 13679 15592 14473 15620
rect 13679 15589 13691 15592
rect 13633 15583 13691 15589
rect 14461 15589 14473 15592
rect 14507 15589 14519 15623
rect 17589 15623 17647 15629
rect 14461 15583 14519 15589
rect 15580 15592 17172 15620
rect 13449 15555 13507 15561
rect 13449 15552 13461 15555
rect 13280 15524 13461 15552
rect 13449 15521 13461 15524
rect 13495 15521 13507 15555
rect 13449 15515 13507 15521
rect 13725 15555 13783 15561
rect 13725 15521 13737 15555
rect 13771 15552 13783 15555
rect 13998 15552 14004 15564
rect 13771 15524 14004 15552
rect 13771 15521 13783 15524
rect 13725 15515 13783 15521
rect 11238 15484 11244 15496
rect 7340 15456 10364 15484
rect 11199 15456 11244 15484
rect 7340 15444 7346 15456
rect 11238 15444 11244 15456
rect 11296 15444 11302 15496
rect 13464 15484 13492 15515
rect 13998 15512 14004 15524
rect 14056 15512 14062 15564
rect 15194 15512 15200 15564
rect 15252 15552 15258 15564
rect 15289 15555 15347 15561
rect 15289 15552 15301 15555
rect 15252 15524 15301 15552
rect 15252 15512 15258 15524
rect 15289 15521 15301 15524
rect 15335 15552 15347 15555
rect 15580 15552 15608 15592
rect 15335 15524 15608 15552
rect 15335 15521 15347 15524
rect 15289 15515 15347 15521
rect 14090 15484 14096 15496
rect 13464 15456 14096 15484
rect 14090 15444 14096 15456
rect 14148 15444 14154 15496
rect 15746 15444 15752 15496
rect 15804 15484 15810 15496
rect 17144 15484 17172 15592
rect 17589 15589 17601 15623
rect 17635 15620 17647 15623
rect 17865 15623 17923 15629
rect 17865 15620 17877 15623
rect 17635 15592 17877 15620
rect 17635 15589 17647 15592
rect 17589 15583 17647 15589
rect 17865 15589 17877 15592
rect 17911 15620 17923 15623
rect 18322 15620 18328 15632
rect 17911 15592 18328 15620
rect 17911 15589 17923 15592
rect 17865 15583 17923 15589
rect 18322 15580 18328 15592
rect 18380 15580 18386 15632
rect 18417 15623 18475 15629
rect 18417 15589 18429 15623
rect 18463 15620 18475 15623
rect 18506 15620 18512 15632
rect 18463 15592 18512 15620
rect 18463 15589 18475 15592
rect 18417 15583 18475 15589
rect 18506 15580 18512 15592
rect 18564 15620 18570 15632
rect 18693 15623 18751 15629
rect 18693 15620 18705 15623
rect 18564 15592 18705 15620
rect 18564 15580 18570 15592
rect 18693 15589 18705 15592
rect 18739 15589 18751 15623
rect 18693 15583 18751 15589
rect 17221 15555 17279 15561
rect 17221 15521 17233 15555
rect 17267 15552 17279 15555
rect 17957 15555 18015 15561
rect 17957 15552 17969 15555
rect 17267 15524 17969 15552
rect 17267 15521 17279 15524
rect 17221 15515 17279 15521
rect 17957 15521 17969 15524
rect 18003 15552 18015 15555
rect 19334 15552 19340 15564
rect 18003 15524 19340 15552
rect 18003 15521 18015 15524
rect 17957 15515 18015 15521
rect 19334 15512 19340 15524
rect 19392 15512 19398 15564
rect 19518 15552 19524 15564
rect 19479 15524 19524 15552
rect 19518 15512 19524 15524
rect 19576 15512 19582 15564
rect 19628 15484 19656 15660
rect 23477 15657 23489 15660
rect 23523 15657 23535 15691
rect 23477 15651 23535 15657
rect 23566 15648 23572 15700
rect 23624 15688 23630 15700
rect 24029 15691 24087 15697
rect 24029 15688 24041 15691
rect 23624 15660 24041 15688
rect 23624 15648 23630 15660
rect 24029 15657 24041 15660
rect 24075 15657 24087 15691
rect 24029 15651 24087 15657
rect 24397 15691 24455 15697
rect 24397 15657 24409 15691
rect 24443 15657 24455 15691
rect 24397 15651 24455 15657
rect 20349 15623 20407 15629
rect 20349 15589 20361 15623
rect 20395 15620 20407 15623
rect 21082 15620 21088 15632
rect 20395 15592 21088 15620
rect 20395 15589 20407 15592
rect 20349 15583 20407 15589
rect 19794 15552 19800 15564
rect 19707 15524 19800 15552
rect 19794 15512 19800 15524
rect 19852 15552 19858 15564
rect 20364 15552 20392 15583
rect 21082 15580 21088 15592
rect 21140 15580 21146 15632
rect 21450 15620 21456 15632
rect 21411 15592 21456 15620
rect 21450 15580 21456 15592
rect 21508 15620 21514 15632
rect 21637 15623 21695 15629
rect 21637 15620 21649 15623
rect 21508 15592 21649 15620
rect 21508 15580 21514 15592
rect 21637 15589 21649 15592
rect 21683 15589 21695 15623
rect 21637 15583 21695 15589
rect 23106 15580 23112 15632
rect 23164 15620 23170 15632
rect 24412 15620 24440 15651
rect 26970 15648 26976 15700
rect 27028 15688 27034 15700
rect 29733 15691 29791 15697
rect 29733 15688 29745 15691
rect 27028 15660 29745 15688
rect 27028 15648 27034 15660
rect 29733 15657 29745 15660
rect 29779 15657 29791 15691
rect 29733 15651 29791 15657
rect 30282 15648 30288 15700
rect 30340 15688 30346 15700
rect 30377 15691 30435 15697
rect 30377 15688 30389 15691
rect 30340 15660 30389 15688
rect 30340 15648 30346 15660
rect 30377 15657 30389 15660
rect 30423 15657 30435 15691
rect 31110 15688 31116 15700
rect 31023 15660 31116 15688
rect 30377 15651 30435 15657
rect 31110 15648 31116 15660
rect 31168 15648 31174 15700
rect 31573 15691 31631 15697
rect 31573 15657 31585 15691
rect 31619 15688 31631 15691
rect 31938 15688 31944 15700
rect 31619 15660 31944 15688
rect 31619 15657 31631 15660
rect 31573 15651 31631 15657
rect 31938 15648 31944 15660
rect 31996 15688 32002 15700
rect 32766 15688 32772 15700
rect 31996 15660 32772 15688
rect 31996 15648 32002 15660
rect 32766 15648 32772 15660
rect 32824 15648 32830 15700
rect 33686 15688 33692 15700
rect 33647 15660 33692 15688
rect 33686 15648 33692 15660
rect 33744 15648 33750 15700
rect 34793 15691 34851 15697
rect 34793 15688 34805 15691
rect 33980 15660 34805 15688
rect 26050 15620 26056 15632
rect 23164 15592 24440 15620
rect 26011 15592 26056 15620
rect 23164 15580 23170 15592
rect 26050 15580 26056 15592
rect 26108 15580 26114 15632
rect 27154 15620 27160 15632
rect 27067 15592 27160 15620
rect 27154 15580 27160 15592
rect 27212 15620 27218 15632
rect 27522 15620 27528 15632
rect 27212 15592 27528 15620
rect 27212 15580 27218 15592
rect 27522 15580 27528 15592
rect 27580 15580 27586 15632
rect 27614 15580 27620 15632
rect 27672 15620 27678 15632
rect 27709 15623 27767 15629
rect 27709 15620 27721 15623
rect 27672 15592 27721 15620
rect 27672 15580 27678 15592
rect 27709 15589 27721 15592
rect 27755 15589 27767 15623
rect 27709 15583 27767 15589
rect 27985 15623 28043 15629
rect 27985 15589 27997 15623
rect 28031 15620 28043 15623
rect 28166 15620 28172 15632
rect 28031 15592 28172 15620
rect 28031 15589 28043 15592
rect 27985 15583 28043 15589
rect 28166 15580 28172 15592
rect 28224 15580 28230 15632
rect 28534 15620 28540 15632
rect 28495 15592 28540 15620
rect 28534 15580 28540 15592
rect 28592 15580 28598 15632
rect 30653 15623 30711 15629
rect 30653 15620 30665 15623
rect 29196 15592 30665 15620
rect 19852 15524 20392 15552
rect 19852 15512 19858 15524
rect 20438 15512 20444 15564
rect 20496 15552 20502 15564
rect 20717 15555 20775 15561
rect 20717 15552 20729 15555
rect 20496 15524 20729 15552
rect 20496 15512 20502 15524
rect 20717 15521 20729 15524
rect 20763 15552 20775 15555
rect 23124 15552 23152 15580
rect 29196 15564 29224 15592
rect 30653 15589 30665 15592
rect 30699 15620 30711 15623
rect 31128 15620 31156 15648
rect 32306 15620 32312 15632
rect 30699 15592 31156 15620
rect 32267 15592 32312 15620
rect 30699 15589 30711 15592
rect 30653 15583 30711 15589
rect 32306 15580 32312 15592
rect 32364 15580 32370 15632
rect 33778 15580 33784 15632
rect 33836 15620 33842 15632
rect 33980 15629 34008 15660
rect 34793 15657 34805 15660
rect 34839 15657 34851 15691
rect 34793 15651 34851 15657
rect 36170 15648 36176 15700
rect 36228 15688 36234 15700
rect 40034 15688 40040 15700
rect 36228 15660 40040 15688
rect 36228 15648 36234 15660
rect 40034 15648 40040 15660
rect 40092 15688 40098 15700
rect 40129 15691 40187 15697
rect 40129 15688 40141 15691
rect 40092 15660 40141 15688
rect 40092 15648 40098 15660
rect 40129 15657 40141 15660
rect 40175 15657 40187 15691
rect 40129 15651 40187 15657
rect 40218 15648 40224 15700
rect 40276 15688 40282 15700
rect 40865 15691 40923 15697
rect 40865 15688 40877 15691
rect 40276 15660 40877 15688
rect 40276 15648 40282 15660
rect 40865 15657 40877 15660
rect 40911 15688 40923 15691
rect 41598 15688 41604 15700
rect 40911 15660 41604 15688
rect 40911 15657 40923 15660
rect 40865 15651 40923 15657
rect 41598 15648 41604 15660
rect 41656 15648 41662 15700
rect 47210 15688 47216 15700
rect 47171 15660 47216 15688
rect 47210 15648 47216 15660
rect 47268 15688 47274 15700
rect 48593 15691 48651 15697
rect 47268 15660 47532 15688
rect 47268 15648 47274 15660
rect 33965 15623 34023 15629
rect 33965 15620 33977 15623
rect 33836 15592 33977 15620
rect 33836 15580 33842 15592
rect 33965 15589 33977 15592
rect 34011 15589 34023 15623
rect 33965 15583 34023 15589
rect 34517 15623 34575 15629
rect 34517 15589 34529 15623
rect 34563 15620 34575 15623
rect 35066 15620 35072 15632
rect 34563 15592 35072 15620
rect 34563 15589 34575 15592
rect 34517 15583 34575 15589
rect 35066 15580 35072 15592
rect 35124 15580 35130 15632
rect 43438 15620 43444 15632
rect 41892 15592 43444 15620
rect 20763 15524 23152 15552
rect 23477 15555 23535 15561
rect 20763 15521 20775 15524
rect 20717 15515 20775 15521
rect 23477 15521 23489 15555
rect 23523 15552 23535 15555
rect 24118 15552 24124 15564
rect 23523 15524 24124 15552
rect 23523 15521 23535 15524
rect 23477 15515 23535 15521
rect 24118 15512 24124 15524
rect 24176 15512 24182 15564
rect 24213 15555 24271 15561
rect 24213 15521 24225 15555
rect 24259 15552 24271 15555
rect 24670 15552 24676 15564
rect 24259 15524 24676 15552
rect 24259 15521 24271 15524
rect 24213 15515 24271 15521
rect 24670 15512 24676 15524
rect 24728 15512 24734 15564
rect 25869 15555 25927 15561
rect 25869 15521 25881 15555
rect 25915 15552 25927 15555
rect 27062 15552 27068 15564
rect 25915 15524 26280 15552
rect 27023 15524 27068 15552
rect 25915 15521 25927 15524
rect 25869 15515 25927 15521
rect 15804 15456 16896 15484
rect 17144 15456 19656 15484
rect 19981 15487 20039 15493
rect 15804 15444 15810 15456
rect 16868 15428 16896 15456
rect 19981 15453 19993 15487
rect 20027 15484 20039 15487
rect 20027 15456 21220 15484
rect 20027 15453 20039 15456
rect 19981 15447 20039 15453
rect 7190 15376 7196 15428
rect 7248 15416 7254 15428
rect 7466 15416 7472 15428
rect 7248 15388 7472 15416
rect 7248 15376 7254 15388
rect 7466 15376 7472 15388
rect 7524 15416 7530 15428
rect 8021 15419 8079 15425
rect 8021 15416 8033 15419
rect 7524 15388 8033 15416
rect 7524 15376 7530 15388
rect 8021 15385 8033 15388
rect 8067 15416 8079 15419
rect 10870 15416 10876 15428
rect 8067 15388 10876 15416
rect 8067 15385 8079 15388
rect 8021 15379 8079 15385
rect 10870 15376 10876 15388
rect 10928 15376 10934 15428
rect 12989 15419 13047 15425
rect 11900 15388 12940 15416
rect 7650 15348 7656 15360
rect 7611 15320 7656 15348
rect 7650 15308 7656 15320
rect 7708 15308 7714 15360
rect 8938 15308 8944 15360
rect 8996 15348 9002 15360
rect 9490 15348 9496 15360
rect 8996 15320 9496 15348
rect 8996 15308 9002 15320
rect 9490 15308 9496 15320
rect 9548 15348 9554 15360
rect 10502 15348 10508 15360
rect 9548 15320 10508 15348
rect 9548 15308 9554 15320
rect 10502 15308 10508 15320
rect 10560 15348 10566 15360
rect 10597 15351 10655 15357
rect 10597 15348 10609 15351
rect 10560 15320 10609 15348
rect 10560 15308 10566 15320
rect 10597 15317 10609 15320
rect 10643 15348 10655 15351
rect 11900 15348 11928 15388
rect 10643 15320 11928 15348
rect 10643 15317 10655 15320
rect 10597 15311 10655 15317
rect 11974 15308 11980 15360
rect 12032 15348 12038 15360
rect 12529 15351 12587 15357
rect 12529 15348 12541 15351
rect 12032 15320 12541 15348
rect 12032 15308 12038 15320
rect 12529 15317 12541 15320
rect 12575 15317 12587 15351
rect 12912 15348 12940 15388
rect 12989 15385 13001 15419
rect 13035 15416 13047 15419
rect 13814 15416 13820 15428
rect 13035 15388 13820 15416
rect 13035 15385 13047 15388
rect 12989 15379 13047 15385
rect 13814 15376 13820 15388
rect 13872 15376 13878 15428
rect 16114 15376 16120 15428
rect 16172 15416 16178 15428
rect 16390 15416 16396 15428
rect 16172 15388 16396 15416
rect 16172 15376 16178 15388
rect 16390 15376 16396 15388
rect 16448 15416 16454 15428
rect 16669 15419 16727 15425
rect 16669 15416 16681 15419
rect 16448 15388 16681 15416
rect 16448 15376 16454 15388
rect 16669 15385 16681 15388
rect 16715 15385 16727 15419
rect 16669 15379 16727 15385
rect 16850 15376 16856 15428
rect 16908 15416 16914 15428
rect 16908 15388 18092 15416
rect 16908 15376 16914 15388
rect 13262 15348 13268 15360
rect 12912 15320 13268 15348
rect 12529 15311 12587 15317
rect 13262 15308 13268 15320
rect 13320 15308 13326 15360
rect 13906 15348 13912 15360
rect 13867 15320 13912 15348
rect 13906 15308 13912 15320
rect 13964 15308 13970 15360
rect 16301 15351 16359 15357
rect 16301 15317 16313 15351
rect 16347 15348 16359 15351
rect 16758 15348 16764 15360
rect 16347 15320 16764 15348
rect 16347 15317 16359 15320
rect 16301 15311 16359 15317
rect 16758 15308 16764 15320
rect 16816 15348 16822 15360
rect 17681 15351 17739 15357
rect 17681 15348 17693 15351
rect 16816 15320 17693 15348
rect 16816 15308 16822 15320
rect 17681 15317 17693 15320
rect 17727 15348 17739 15351
rect 17862 15348 17868 15360
rect 17727 15320 17868 15348
rect 17727 15317 17739 15320
rect 17681 15311 17739 15317
rect 17862 15308 17868 15320
rect 17920 15308 17926 15360
rect 18064 15348 18092 15388
rect 18138 15376 18144 15428
rect 18196 15416 18202 15428
rect 19996 15416 20024 15447
rect 18196 15388 20024 15416
rect 18196 15376 18202 15388
rect 19794 15348 19800 15360
rect 18064 15320 19800 15348
rect 19794 15308 19800 15320
rect 19852 15348 19858 15360
rect 21085 15351 21143 15357
rect 21085 15348 21097 15351
rect 19852 15320 21097 15348
rect 19852 15308 19858 15320
rect 21085 15317 21097 15320
rect 21131 15317 21143 15351
rect 21192 15348 21220 15456
rect 21634 15444 21640 15496
rect 21692 15484 21698 15496
rect 21729 15487 21787 15493
rect 21729 15484 21741 15487
rect 21692 15456 21741 15484
rect 21692 15444 21698 15456
rect 21729 15453 21741 15456
rect 21775 15453 21787 15487
rect 22002 15484 22008 15496
rect 21963 15456 22008 15484
rect 21729 15447 21787 15453
rect 22002 15444 22008 15456
rect 22060 15444 22066 15496
rect 24688 15484 24716 15512
rect 24688 15456 26096 15484
rect 25869 15419 25927 15425
rect 25869 15416 25881 15419
rect 23124 15388 25881 15416
rect 23124 15348 23152 15388
rect 25869 15385 25881 15388
rect 25915 15385 25927 15419
rect 25869 15379 25927 15385
rect 23290 15348 23296 15360
rect 21192 15320 23152 15348
rect 23251 15320 23296 15348
rect 21085 15311 21143 15317
rect 23290 15308 23296 15320
rect 23348 15308 23354 15360
rect 23658 15348 23664 15360
rect 23619 15320 23664 15348
rect 23658 15308 23664 15320
rect 23716 15308 23722 15360
rect 25038 15308 25044 15360
rect 25096 15348 25102 15360
rect 25593 15351 25651 15357
rect 25593 15348 25605 15351
rect 25096 15320 25605 15348
rect 25096 15308 25102 15320
rect 25593 15317 25605 15320
rect 25639 15348 25651 15351
rect 25958 15348 25964 15360
rect 25639 15320 25964 15348
rect 25639 15317 25651 15320
rect 25593 15311 25651 15317
rect 25958 15308 25964 15320
rect 26016 15308 26022 15360
rect 26068 15348 26096 15456
rect 26252 15416 26280 15524
rect 27062 15512 27068 15524
rect 27120 15512 27126 15564
rect 27249 15555 27307 15561
rect 27249 15521 27261 15555
rect 27295 15552 27307 15555
rect 28074 15552 28080 15564
rect 27295 15524 28080 15552
rect 27295 15521 27307 15524
rect 27249 15515 27307 15521
rect 26881 15487 26939 15493
rect 26881 15453 26893 15487
rect 26927 15484 26939 15487
rect 27264 15484 27292 15515
rect 28074 15512 28080 15524
rect 28132 15512 28138 15564
rect 28902 15512 28908 15564
rect 28960 15552 28966 15564
rect 28997 15555 29055 15561
rect 28997 15552 29009 15555
rect 28960 15524 29009 15552
rect 28960 15512 28966 15524
rect 28997 15521 29009 15524
rect 29043 15521 29055 15555
rect 29178 15552 29184 15564
rect 29139 15524 29184 15552
rect 28997 15515 29055 15521
rect 29178 15512 29184 15524
rect 29236 15512 29242 15564
rect 29362 15552 29368 15564
rect 29323 15524 29368 15552
rect 29362 15512 29368 15524
rect 29420 15512 29426 15564
rect 29733 15555 29791 15561
rect 29733 15521 29745 15555
rect 29779 15552 29791 15555
rect 30929 15555 30987 15561
rect 30929 15552 30941 15555
rect 29779 15524 30941 15552
rect 29779 15521 29791 15524
rect 29733 15515 29791 15521
rect 30929 15521 30941 15524
rect 30975 15552 30987 15555
rect 31294 15552 31300 15564
rect 30975 15524 31300 15552
rect 30975 15521 30987 15524
rect 30929 15515 30987 15521
rect 31294 15512 31300 15524
rect 31352 15512 31358 15564
rect 31754 15512 31760 15564
rect 31812 15552 31818 15564
rect 32401 15555 32459 15561
rect 32401 15552 32413 15555
rect 31812 15524 32413 15552
rect 31812 15512 31818 15524
rect 32401 15521 32413 15524
rect 32447 15521 32459 15555
rect 32401 15515 32459 15521
rect 34057 15555 34115 15561
rect 34057 15521 34069 15555
rect 34103 15552 34115 15555
rect 34790 15552 34796 15564
rect 34103 15524 34796 15552
rect 34103 15521 34115 15524
rect 34057 15515 34115 15521
rect 34790 15512 34796 15524
rect 34848 15512 34854 15564
rect 35345 15555 35403 15561
rect 35345 15521 35357 15555
rect 35391 15521 35403 15555
rect 36538 15552 36544 15564
rect 36499 15524 36544 15552
rect 35345 15515 35403 15521
rect 26927 15456 27292 15484
rect 26927 15453 26939 15456
rect 26881 15447 26939 15453
rect 27430 15444 27436 15496
rect 27488 15484 27494 15496
rect 28353 15487 28411 15493
rect 28353 15484 28365 15487
rect 27488 15456 28365 15484
rect 27488 15444 27494 15456
rect 28353 15453 28365 15456
rect 28399 15453 28411 15487
rect 28353 15447 28411 15453
rect 29270 15444 29276 15496
rect 29328 15484 29334 15496
rect 29917 15487 29975 15493
rect 29917 15484 29929 15487
rect 29328 15456 29929 15484
rect 29328 15444 29334 15456
rect 29917 15453 29929 15456
rect 29963 15484 29975 15487
rect 32030 15484 32036 15496
rect 29963 15456 32036 15484
rect 29963 15453 29975 15456
rect 29917 15447 29975 15453
rect 32030 15444 32036 15456
rect 32088 15484 32094 15496
rect 32125 15487 32183 15493
rect 32125 15484 32137 15487
rect 32088 15456 32137 15484
rect 32088 15444 32094 15456
rect 32125 15453 32137 15456
rect 32171 15453 32183 15487
rect 35360 15484 35388 15515
rect 36538 15512 36544 15524
rect 36596 15512 36602 15564
rect 41892 15561 41920 15592
rect 43438 15580 43444 15592
rect 43496 15580 43502 15632
rect 47504 15629 47532 15660
rect 48593 15657 48605 15691
rect 48639 15688 48651 15691
rect 48774 15688 48780 15700
rect 48639 15660 48780 15688
rect 48639 15657 48651 15660
rect 48593 15651 48651 15657
rect 48774 15648 48780 15660
rect 48832 15648 48838 15700
rect 49970 15688 49976 15700
rect 49160 15660 49976 15688
rect 47489 15623 47547 15629
rect 47489 15589 47501 15623
rect 47535 15589 47547 15623
rect 47489 15583 47547 15589
rect 48041 15623 48099 15629
rect 48041 15589 48053 15623
rect 48087 15620 48099 15623
rect 48314 15620 48320 15632
rect 48087 15592 48320 15620
rect 48087 15589 48099 15592
rect 48041 15583 48099 15589
rect 48314 15580 48320 15592
rect 48372 15580 48378 15632
rect 49160 15629 49188 15660
rect 49970 15648 49976 15660
rect 50028 15648 50034 15700
rect 52454 15688 52460 15700
rect 52415 15660 52460 15688
rect 52454 15648 52460 15660
rect 52512 15648 52518 15700
rect 54018 15688 54024 15700
rect 53979 15660 54024 15688
rect 54018 15648 54024 15660
rect 54076 15648 54082 15700
rect 61654 15688 61660 15700
rect 54128 15660 61660 15688
rect 49145 15623 49203 15629
rect 49145 15589 49157 15623
rect 49191 15589 49203 15623
rect 49145 15583 49203 15589
rect 50706 15580 50712 15632
rect 50764 15620 50770 15632
rect 52472 15620 52500 15648
rect 52638 15620 52644 15632
rect 50764 15592 52500 15620
rect 52599 15592 52644 15620
rect 50764 15580 50770 15592
rect 52638 15580 52644 15592
rect 52696 15580 52702 15632
rect 41877 15555 41935 15561
rect 41877 15521 41889 15555
rect 41923 15521 41935 15555
rect 41877 15515 41935 15521
rect 42061 15555 42119 15561
rect 42061 15521 42073 15555
rect 42107 15521 42119 15555
rect 42242 15552 42248 15564
rect 42203 15524 42248 15552
rect 42061 15515 42119 15521
rect 35710 15484 35716 15496
rect 32125 15447 32183 15453
rect 34440 15456 35716 15484
rect 30742 15416 30748 15428
rect 26252 15388 30748 15416
rect 30742 15376 30748 15388
rect 30800 15376 30806 15428
rect 34440 15416 34468 15456
rect 35710 15444 35716 15456
rect 35768 15444 35774 15496
rect 38289 15487 38347 15493
rect 38289 15453 38301 15487
rect 38335 15484 38347 15487
rect 38470 15484 38476 15496
rect 38335 15456 38476 15484
rect 38335 15453 38347 15456
rect 38289 15447 38347 15453
rect 38470 15444 38476 15456
rect 38528 15484 38534 15496
rect 38565 15487 38623 15493
rect 38565 15484 38577 15487
rect 38528 15456 38577 15484
rect 38528 15444 38534 15456
rect 38565 15453 38577 15456
rect 38611 15453 38623 15487
rect 38565 15447 38623 15453
rect 38841 15487 38899 15493
rect 38841 15453 38853 15487
rect 38887 15484 38899 15487
rect 40126 15484 40132 15496
rect 38887 15456 40132 15484
rect 38887 15453 38899 15456
rect 38841 15447 38899 15453
rect 40126 15444 40132 15456
rect 40184 15444 40190 15496
rect 42076 15484 42104 15515
rect 42242 15512 42248 15524
rect 42300 15512 42306 15564
rect 46198 15552 46204 15564
rect 46159 15524 46204 15552
rect 46198 15512 46204 15524
rect 46256 15512 46262 15564
rect 46845 15555 46903 15561
rect 46845 15521 46857 15555
rect 46891 15552 46903 15555
rect 47578 15552 47584 15564
rect 46891 15524 47584 15552
rect 46891 15521 46903 15524
rect 46845 15515 46903 15521
rect 47578 15512 47584 15524
rect 47636 15512 47642 15564
rect 49237 15555 49295 15561
rect 49237 15521 49249 15555
rect 49283 15552 49295 15555
rect 49602 15552 49608 15564
rect 49283 15524 49608 15552
rect 49283 15521 49295 15524
rect 49237 15515 49295 15521
rect 49602 15512 49608 15524
rect 49660 15512 49666 15564
rect 51261 15555 51319 15561
rect 51261 15521 51273 15555
rect 51307 15521 51319 15555
rect 51626 15552 51632 15564
rect 51587 15524 51632 15552
rect 51261 15515 51319 15521
rect 42334 15484 42340 15496
rect 41248 15456 42340 15484
rect 35529 15419 35587 15425
rect 35529 15416 35541 15419
rect 30852 15388 34468 15416
rect 34532 15388 35541 15416
rect 30852 15348 30880 15388
rect 32582 15348 32588 15360
rect 26068 15320 30880 15348
rect 32543 15320 32588 15348
rect 32582 15308 32588 15320
rect 32640 15308 32646 15360
rect 32858 15308 32864 15360
rect 32916 15348 32922 15360
rect 33321 15351 33379 15357
rect 33321 15348 33333 15351
rect 32916 15320 33333 15348
rect 32916 15308 32922 15320
rect 33321 15317 33333 15320
rect 33367 15348 33379 15351
rect 33781 15351 33839 15357
rect 33781 15348 33793 15351
rect 33367 15320 33793 15348
rect 33367 15317 33379 15320
rect 33321 15311 33379 15317
rect 33781 15317 33793 15320
rect 33827 15317 33839 15351
rect 33781 15311 33839 15317
rect 34330 15308 34336 15360
rect 34388 15348 34394 15360
rect 34532 15348 34560 15388
rect 35529 15385 35541 15388
rect 35575 15385 35587 15419
rect 35529 15379 35587 15385
rect 36725 15419 36783 15425
rect 36725 15385 36737 15419
rect 36771 15416 36783 15419
rect 36771 15388 38608 15416
rect 36771 15385 36783 15388
rect 36725 15379 36783 15385
rect 35158 15348 35164 15360
rect 34388 15320 34560 15348
rect 35119 15320 35164 15348
rect 34388 15308 34394 15320
rect 35158 15308 35164 15320
rect 35216 15308 35222 15360
rect 36170 15348 36176 15360
rect 36131 15320 36176 15348
rect 36170 15308 36176 15320
rect 36228 15308 36234 15360
rect 37182 15348 37188 15360
rect 37143 15320 37188 15348
rect 37182 15308 37188 15320
rect 37240 15308 37246 15360
rect 37458 15348 37464 15360
rect 37419 15320 37464 15348
rect 37458 15308 37464 15320
rect 37516 15308 37522 15360
rect 38010 15308 38016 15360
rect 38068 15348 38074 15360
rect 38289 15351 38347 15357
rect 38289 15348 38301 15351
rect 38068 15320 38301 15348
rect 38068 15308 38074 15320
rect 38289 15317 38301 15320
rect 38335 15348 38347 15351
rect 38381 15351 38439 15357
rect 38381 15348 38393 15351
rect 38335 15320 38393 15348
rect 38335 15317 38347 15320
rect 38289 15311 38347 15317
rect 38381 15317 38393 15320
rect 38427 15317 38439 15351
rect 38580 15348 38608 15388
rect 39850 15376 39856 15428
rect 39908 15416 39914 15428
rect 41248 15425 41276 15456
rect 42334 15444 42340 15456
rect 42392 15444 42398 15496
rect 50246 15444 50252 15496
rect 50304 15484 50310 15496
rect 50801 15487 50859 15493
rect 50801 15484 50813 15487
rect 50304 15456 50813 15484
rect 50304 15444 50310 15456
rect 50801 15453 50813 15456
rect 50847 15453 50859 15487
rect 50801 15447 50859 15453
rect 41233 15419 41291 15425
rect 41233 15416 41245 15419
rect 39908 15388 41245 15416
rect 39908 15376 39914 15388
rect 41233 15385 41245 15388
rect 41279 15385 41291 15419
rect 41690 15416 41696 15428
rect 41651 15388 41696 15416
rect 41233 15379 41291 15385
rect 41690 15376 41696 15388
rect 41748 15376 41754 15428
rect 46385 15419 46443 15425
rect 46385 15385 46397 15419
rect 46431 15416 46443 15419
rect 48774 15416 48780 15428
rect 46431 15388 48780 15416
rect 46431 15385 46443 15388
rect 46385 15379 46443 15385
rect 48774 15376 48780 15388
rect 48832 15376 48838 15428
rect 51276 15416 51304 15515
rect 51626 15512 51632 15524
rect 51684 15512 51690 15564
rect 53101 15555 53159 15561
rect 53101 15521 53113 15555
rect 53147 15552 53159 15555
rect 53282 15552 53288 15564
rect 53147 15524 53288 15552
rect 53147 15521 53159 15524
rect 53101 15515 53159 15521
rect 53282 15512 53288 15524
rect 53340 15512 53346 15564
rect 53466 15552 53472 15564
rect 53427 15524 53472 15552
rect 53466 15512 53472 15524
rect 53524 15512 53530 15564
rect 53561 15555 53619 15561
rect 53561 15521 53573 15555
rect 53607 15552 53619 15555
rect 54036 15552 54064 15648
rect 53607 15524 54064 15552
rect 53607 15521 53619 15524
rect 53561 15515 53619 15521
rect 51718 15484 51724 15496
rect 51679 15456 51724 15484
rect 51718 15444 51724 15456
rect 51776 15444 51782 15496
rect 51350 15416 51356 15428
rect 51263 15388 51356 15416
rect 51350 15376 51356 15388
rect 51408 15416 51414 15428
rect 54128 15416 54156 15660
rect 61654 15648 61660 15660
rect 61712 15648 61718 15700
rect 57698 15620 57704 15632
rect 56888 15592 57704 15620
rect 56888 15564 56916 15592
rect 57698 15580 57704 15592
rect 57756 15580 57762 15632
rect 56870 15552 56876 15564
rect 56783 15524 56876 15552
rect 56870 15512 56876 15524
rect 56928 15512 56934 15564
rect 56962 15512 56968 15564
rect 57020 15552 57026 15564
rect 57057 15555 57115 15561
rect 57057 15552 57069 15555
rect 57020 15524 57069 15552
rect 57020 15512 57026 15524
rect 57057 15521 57069 15524
rect 57103 15521 57115 15555
rect 57057 15515 57115 15521
rect 57241 15555 57299 15561
rect 57241 15521 57253 15555
rect 57287 15521 57299 15555
rect 57241 15515 57299 15521
rect 55858 15444 55864 15496
rect 55916 15484 55922 15496
rect 56137 15487 56195 15493
rect 56137 15484 56149 15487
rect 55916 15456 56149 15484
rect 55916 15444 55922 15456
rect 56137 15453 56149 15456
rect 56183 15484 56195 15487
rect 56413 15487 56471 15493
rect 56413 15484 56425 15487
rect 56183 15456 56425 15484
rect 56183 15453 56195 15456
rect 56137 15447 56195 15453
rect 56413 15453 56425 15456
rect 56459 15453 56471 15487
rect 56413 15447 56471 15453
rect 56778 15444 56784 15496
rect 56836 15484 56842 15496
rect 57256 15484 57284 15515
rect 58069 15487 58127 15493
rect 58069 15484 58081 15487
rect 56836 15456 58081 15484
rect 56836 15444 56842 15456
rect 58069 15453 58081 15456
rect 58115 15484 58127 15487
rect 58158 15484 58164 15496
rect 58115 15456 58164 15484
rect 58115 15453 58127 15456
rect 58069 15447 58127 15453
rect 58158 15444 58164 15456
rect 58216 15444 58222 15496
rect 51408 15388 54156 15416
rect 51408 15376 51414 15388
rect 58894 15376 58900 15428
rect 58952 15416 58958 15428
rect 59722 15416 59728 15428
rect 58952 15388 59728 15416
rect 58952 15376 58958 15388
rect 59722 15376 59728 15388
rect 59780 15376 59786 15428
rect 38930 15348 38936 15360
rect 38580 15320 38936 15348
rect 38381 15311 38439 15317
rect 38930 15308 38936 15320
rect 38988 15308 38994 15360
rect 40494 15348 40500 15360
rect 40455 15320 40500 15348
rect 40494 15308 40500 15320
rect 40552 15308 40558 15360
rect 42886 15348 42892 15360
rect 42847 15320 42892 15348
rect 42886 15308 42892 15320
rect 42944 15308 42950 15360
rect 43070 15308 43076 15360
rect 43128 15348 43134 15360
rect 43533 15351 43591 15357
rect 43533 15348 43545 15351
rect 43128 15320 43545 15348
rect 43128 15308 43134 15320
rect 43533 15317 43545 15320
rect 43579 15317 43591 15351
rect 43898 15348 43904 15360
rect 43859 15320 43904 15348
rect 43533 15311 43591 15317
rect 43898 15308 43904 15320
rect 43956 15308 43962 15360
rect 47302 15348 47308 15360
rect 47263 15320 47308 15348
rect 47302 15308 47308 15320
rect 47360 15308 47366 15360
rect 48961 15351 49019 15357
rect 48961 15317 48973 15351
rect 49007 15348 49019 15351
rect 49142 15348 49148 15360
rect 49007 15320 49148 15348
rect 49007 15317 49019 15320
rect 48961 15311 49019 15317
rect 49142 15308 49148 15320
rect 49200 15308 49206 15360
rect 49418 15348 49424 15360
rect 49379 15320 49424 15348
rect 49418 15308 49424 15320
rect 49476 15308 49482 15360
rect 50338 15348 50344 15360
rect 50299 15320 50344 15348
rect 50338 15308 50344 15320
rect 50396 15308 50402 15360
rect 52181 15351 52239 15357
rect 52181 15317 52193 15351
rect 52227 15348 52239 15351
rect 52270 15348 52276 15360
rect 52227 15320 52276 15348
rect 52227 15317 52239 15320
rect 52181 15311 52239 15317
rect 52270 15308 52276 15320
rect 52328 15308 52334 15360
rect 55674 15348 55680 15360
rect 55635 15320 55680 15348
rect 55674 15308 55680 15320
rect 55732 15308 55738 15360
rect 57793 15351 57851 15357
rect 57793 15317 57805 15351
rect 57839 15348 57851 15351
rect 57974 15348 57980 15360
rect 57839 15320 57980 15348
rect 57839 15317 57851 15320
rect 57793 15311 57851 15317
rect 57974 15308 57980 15320
rect 58032 15308 58038 15360
rect 1104 15258 63480 15280
rect 1104 15206 11378 15258
rect 11430 15206 11442 15258
rect 11494 15206 11506 15258
rect 11558 15206 11570 15258
rect 11622 15206 32170 15258
rect 32222 15206 32234 15258
rect 32286 15206 32298 15258
rect 32350 15206 32362 15258
rect 32414 15206 52962 15258
rect 53014 15206 53026 15258
rect 53078 15206 53090 15258
rect 53142 15206 53154 15258
rect 53206 15206 63480 15258
rect 1104 15184 63480 15206
rect 4525 15147 4583 15153
rect 4525 15113 4537 15147
rect 4571 15144 4583 15147
rect 5350 15144 5356 15156
rect 4571 15116 5356 15144
rect 4571 15113 4583 15116
rect 4525 15107 4583 15113
rect 5350 15104 5356 15116
rect 5408 15104 5414 15156
rect 5626 15104 5632 15156
rect 5684 15144 5690 15156
rect 6181 15147 6239 15153
rect 6181 15144 6193 15147
rect 5684 15116 6193 15144
rect 5684 15104 5690 15116
rect 6181 15113 6193 15116
rect 6227 15144 6239 15147
rect 6270 15144 6276 15156
rect 6227 15116 6276 15144
rect 6227 15113 6239 15116
rect 6181 15107 6239 15113
rect 6270 15104 6276 15116
rect 6328 15104 6334 15156
rect 7190 15144 7196 15156
rect 7151 15116 7196 15144
rect 7190 15104 7196 15116
rect 7248 15104 7254 15156
rect 7300 15116 22416 15144
rect 2866 15036 2872 15088
rect 2924 15076 2930 15088
rect 7300 15076 7328 15116
rect 2924 15048 7328 15076
rect 2924 15036 2930 15048
rect 8754 15036 8760 15088
rect 8812 15076 8818 15088
rect 8849 15079 8907 15085
rect 8849 15076 8861 15079
rect 8812 15048 8861 15076
rect 8812 15036 8818 15048
rect 8849 15045 8861 15048
rect 8895 15076 8907 15079
rect 11057 15079 11115 15085
rect 11057 15076 11069 15079
rect 8895 15048 11069 15076
rect 8895 15045 8907 15048
rect 8849 15039 8907 15045
rect 4062 14968 4068 15020
rect 4120 15008 4126 15020
rect 4120 14980 7236 15008
rect 4120 14968 4126 14980
rect 5261 14943 5319 14949
rect 5261 14909 5273 14943
rect 5307 14940 5319 14943
rect 5350 14940 5356 14952
rect 5307 14912 5356 14940
rect 5307 14909 5319 14912
rect 5261 14903 5319 14909
rect 5350 14900 5356 14912
rect 5408 14900 5414 14952
rect 5445 14943 5503 14949
rect 5445 14909 5457 14943
rect 5491 14940 5503 14943
rect 5534 14940 5540 14952
rect 5491 14912 5540 14940
rect 5491 14909 5503 14912
rect 5445 14903 5503 14909
rect 4893 14875 4951 14881
rect 4893 14841 4905 14875
rect 4939 14872 4951 14875
rect 5460 14872 5488 14903
rect 5534 14900 5540 14912
rect 5592 14900 5598 14952
rect 5902 14872 5908 14884
rect 4939 14844 5488 14872
rect 5863 14844 5908 14872
rect 4939 14841 4951 14844
rect 4893 14835 4951 14841
rect 5902 14832 5908 14844
rect 5960 14832 5966 14884
rect 5442 14764 5448 14816
rect 5500 14804 5506 14816
rect 6549 14807 6607 14813
rect 6549 14804 6561 14807
rect 5500 14776 6561 14804
rect 5500 14764 5506 14776
rect 6549 14773 6561 14776
rect 6595 14804 6607 14807
rect 7098 14804 7104 14816
rect 6595 14776 7104 14804
rect 6595 14773 6607 14776
rect 6549 14767 6607 14773
rect 7098 14764 7104 14776
rect 7156 14764 7162 14816
rect 7208 14804 7236 14980
rect 7742 14968 7748 15020
rect 7800 15008 7806 15020
rect 9769 15011 9827 15017
rect 9769 15008 9781 15011
rect 7800 14980 9781 15008
rect 7800 14968 7806 14980
rect 9769 14977 9781 14980
rect 9815 14977 9827 15011
rect 9769 14971 9827 14977
rect 7282 14900 7288 14952
rect 7340 14940 7346 14952
rect 7561 14943 7619 14949
rect 7340 14912 7385 14940
rect 7340 14900 7346 14912
rect 7561 14909 7573 14943
rect 7607 14940 7619 14943
rect 7650 14940 7656 14952
rect 7607 14912 7656 14940
rect 7607 14909 7619 14912
rect 7561 14903 7619 14909
rect 7650 14900 7656 14912
rect 7708 14940 7714 14952
rect 8018 14940 8024 14952
rect 7708 14912 8024 14940
rect 7708 14900 7714 14912
rect 8018 14900 8024 14912
rect 8076 14900 8082 14952
rect 10244 14949 10272 15048
rect 11057 15045 11069 15048
rect 11103 15045 11115 15079
rect 14090 15076 14096 15088
rect 14051 15048 14096 15076
rect 11057 15039 11115 15045
rect 14090 15036 14096 15048
rect 14148 15076 14154 15088
rect 14461 15079 14519 15085
rect 14461 15076 14473 15079
rect 14148 15048 14473 15076
rect 14148 15036 14154 15048
rect 14461 15045 14473 15048
rect 14507 15045 14519 15079
rect 15562 15076 15568 15088
rect 15523 15048 15568 15076
rect 14461 15039 14519 15045
rect 15562 15036 15568 15048
rect 15620 15036 15626 15088
rect 16393 15079 16451 15085
rect 16393 15045 16405 15079
rect 16439 15076 16451 15079
rect 17034 15076 17040 15088
rect 16439 15048 17040 15076
rect 16439 15045 16451 15048
rect 16393 15039 16451 15045
rect 17034 15036 17040 15048
rect 17092 15036 17098 15088
rect 17497 15079 17555 15085
rect 17497 15045 17509 15079
rect 17543 15076 17555 15079
rect 18138 15076 18144 15088
rect 17543 15048 18144 15076
rect 17543 15045 17555 15048
rect 17497 15039 17555 15045
rect 13725 15011 13783 15017
rect 13725 15008 13737 15011
rect 11072 14980 12572 15008
rect 10229 14943 10287 14949
rect 10229 14909 10241 14943
rect 10275 14909 10287 14943
rect 10410 14940 10416 14952
rect 10371 14912 10416 14940
rect 10229 14903 10287 14909
rect 10410 14900 10416 14912
rect 10468 14900 10474 14952
rect 10502 14900 10508 14952
rect 10560 14949 10566 14952
rect 10560 14943 10609 14949
rect 10560 14909 10563 14943
rect 10597 14909 10609 14943
rect 10560 14903 10609 14909
rect 10560 14900 10566 14903
rect 8294 14832 8300 14884
rect 8352 14872 8358 14884
rect 9217 14875 9275 14881
rect 9217 14872 9229 14875
rect 8352 14844 9229 14872
rect 8352 14832 8358 14844
rect 9217 14841 9229 14844
rect 9263 14841 9275 14875
rect 9217 14835 9275 14841
rect 11072 14804 11100 14980
rect 11146 14900 11152 14952
rect 11204 14940 11210 14952
rect 12437 14943 12495 14949
rect 12437 14940 12449 14943
rect 11204 14912 12449 14940
rect 11204 14900 11210 14912
rect 12437 14909 12449 14912
rect 12483 14909 12495 14943
rect 12437 14903 12495 14909
rect 11514 14832 11520 14884
rect 11572 14872 11578 14884
rect 11885 14875 11943 14881
rect 11885 14872 11897 14875
rect 11572 14844 11897 14872
rect 11572 14832 11578 14844
rect 11885 14841 11897 14844
rect 11931 14872 11943 14875
rect 12158 14872 12164 14884
rect 11931 14844 12164 14872
rect 11931 14841 11943 14844
rect 11885 14835 11943 14841
rect 12158 14832 12164 14844
rect 12216 14832 12222 14884
rect 12544 14872 12572 14980
rect 12912 14980 13737 15008
rect 12618 14900 12624 14952
rect 12676 14940 12682 14952
rect 12912 14949 12940 14980
rect 13725 14977 13737 14980
rect 13771 14977 13783 15011
rect 14182 15008 14188 15020
rect 13725 14971 13783 14977
rect 13813 14980 14188 15008
rect 12897 14943 12955 14949
rect 12897 14940 12909 14943
rect 12676 14912 12909 14940
rect 12676 14900 12682 14912
rect 12897 14909 12909 14912
rect 12943 14909 12955 14943
rect 13262 14940 13268 14952
rect 13223 14912 13268 14940
rect 12897 14903 12955 14909
rect 13262 14900 13268 14912
rect 13320 14900 13326 14952
rect 13357 14943 13415 14949
rect 13357 14909 13369 14943
rect 13403 14940 13415 14943
rect 13446 14940 13452 14952
rect 13403 14912 13452 14940
rect 13403 14909 13415 14912
rect 13357 14903 13415 14909
rect 13446 14900 13452 14912
rect 13504 14940 13510 14952
rect 13813 14940 13841 14980
rect 14182 14968 14188 14980
rect 14240 14968 14246 15020
rect 15194 15008 15200 15020
rect 15155 14980 15200 15008
rect 15194 14968 15200 14980
rect 15252 14968 15258 15020
rect 15304 14980 16896 15008
rect 14274 14940 14280 14952
rect 13504 14912 13841 14940
rect 14187 14912 14280 14940
rect 13504 14900 13510 14912
rect 14274 14900 14280 14912
rect 14332 14940 14338 14952
rect 14921 14943 14979 14949
rect 14921 14940 14933 14943
rect 14332 14912 14933 14940
rect 14332 14900 14338 14912
rect 14921 14909 14933 14912
rect 14967 14940 14979 14943
rect 15304 14940 15332 14980
rect 14967 14912 15332 14940
rect 15381 14943 15439 14949
rect 14967 14909 14979 14912
rect 14921 14903 14979 14909
rect 15381 14909 15393 14943
rect 15427 14940 15439 14943
rect 16022 14940 16028 14952
rect 15427 14912 16028 14940
rect 15427 14909 15439 14912
rect 15381 14903 15439 14909
rect 16022 14900 16028 14912
rect 16080 14900 16086 14952
rect 16868 14949 16896 14980
rect 16853 14943 16911 14949
rect 16853 14909 16865 14943
rect 16899 14940 16911 14943
rect 17512 14940 17540 15039
rect 18138 15036 18144 15048
rect 18196 15036 18202 15088
rect 20806 15076 20812 15088
rect 18248 15048 20812 15076
rect 18248 15008 18276 15048
rect 20806 15036 20812 15048
rect 20864 15036 20870 15088
rect 20990 15076 20996 15088
rect 20951 15048 20996 15076
rect 20990 15036 20996 15048
rect 21048 15036 21054 15088
rect 21082 15036 21088 15088
rect 21140 15076 21146 15088
rect 21361 15079 21419 15085
rect 21361 15076 21373 15079
rect 21140 15048 21373 15076
rect 21140 15036 21146 15048
rect 21361 15045 21373 15048
rect 21407 15076 21419 15079
rect 22002 15076 22008 15088
rect 21407 15048 22008 15076
rect 21407 15045 21419 15048
rect 21361 15039 21419 15045
rect 22002 15036 22008 15048
rect 22060 15036 22066 15088
rect 22388 15076 22416 15116
rect 22462 15104 22468 15156
rect 22520 15144 22526 15156
rect 22741 15147 22799 15153
rect 22741 15144 22753 15147
rect 22520 15116 22753 15144
rect 22520 15104 22526 15116
rect 22741 15113 22753 15116
rect 22787 15113 22799 15147
rect 28258 15144 28264 15156
rect 22741 15107 22799 15113
rect 22848 15116 28028 15144
rect 28219 15116 28264 15144
rect 22848 15076 22876 15116
rect 23106 15076 23112 15088
rect 22388 15048 22876 15076
rect 23067 15048 23112 15076
rect 23106 15036 23112 15048
rect 23164 15036 23170 15088
rect 23290 15036 23296 15088
rect 23348 15076 23354 15088
rect 25593 15079 25651 15085
rect 25593 15076 25605 15079
rect 23348 15048 25605 15076
rect 23348 15036 23354 15048
rect 25593 15045 25605 15048
rect 25639 15076 25651 15079
rect 25685 15079 25743 15085
rect 25685 15076 25697 15079
rect 25639 15048 25697 15076
rect 25639 15045 25651 15048
rect 25593 15039 25651 15045
rect 25685 15045 25697 15048
rect 25731 15045 25743 15079
rect 27062 15076 27068 15088
rect 27023 15048 27068 15076
rect 25685 15039 25743 15045
rect 27062 15036 27068 15048
rect 27120 15036 27126 15088
rect 27430 15036 27436 15088
rect 27488 15076 27494 15088
rect 27893 15079 27951 15085
rect 27893 15076 27905 15079
rect 27488 15048 27905 15076
rect 27488 15036 27494 15048
rect 27893 15045 27905 15048
rect 27939 15045 27951 15079
rect 28000 15076 28028 15116
rect 28258 15104 28264 15116
rect 28316 15104 28322 15156
rect 28994 15144 29000 15156
rect 28955 15116 29000 15144
rect 28994 15104 29000 15116
rect 29052 15104 29058 15156
rect 29270 15144 29276 15156
rect 29231 15116 29276 15144
rect 29270 15104 29276 15116
rect 29328 15104 29334 15156
rect 29546 15104 29552 15156
rect 29604 15144 29610 15156
rect 29733 15147 29791 15153
rect 29733 15144 29745 15147
rect 29604 15116 29745 15144
rect 29604 15104 29610 15116
rect 29733 15113 29745 15116
rect 29779 15113 29791 15147
rect 29733 15107 29791 15113
rect 30098 15104 30104 15156
rect 30156 15144 30162 15156
rect 30285 15147 30343 15153
rect 30285 15144 30297 15147
rect 30156 15116 30297 15144
rect 30156 15104 30162 15116
rect 30285 15113 30297 15116
rect 30331 15113 30343 15147
rect 31294 15144 31300 15156
rect 31255 15116 31300 15144
rect 30285 15107 30343 15113
rect 31294 15104 31300 15116
rect 31352 15104 31358 15156
rect 31754 15104 31760 15156
rect 31812 15144 31818 15156
rect 32030 15144 32036 15156
rect 31812 15116 31857 15144
rect 31943 15116 32036 15144
rect 31812 15104 31818 15116
rect 32030 15104 32036 15116
rect 32088 15144 32094 15156
rect 32858 15144 32864 15156
rect 32088 15116 32864 15144
rect 32088 15104 32094 15116
rect 32858 15104 32864 15116
rect 32916 15104 32922 15156
rect 34057 15147 34115 15153
rect 34057 15144 34069 15147
rect 33152 15116 34069 15144
rect 31113 15079 31171 15085
rect 31113 15076 31125 15079
rect 28000 15048 31125 15076
rect 27893 15039 27951 15045
rect 31113 15045 31125 15048
rect 31159 15045 31171 15079
rect 31312 15076 31340 15104
rect 32398 15076 32404 15088
rect 31312 15048 32404 15076
rect 31113 15039 31171 15045
rect 32398 15036 32404 15048
rect 32456 15036 32462 15088
rect 32493 15079 32551 15085
rect 32493 15045 32505 15079
rect 32539 15076 32551 15079
rect 32674 15076 32680 15088
rect 32539 15048 32680 15076
rect 32539 15045 32551 15048
rect 32493 15039 32551 15045
rect 32674 15036 32680 15048
rect 32732 15036 32738 15088
rect 16899 14912 17540 14940
rect 17604 14980 18276 15008
rect 18785 15011 18843 15017
rect 16899 14909 16911 14912
rect 16853 14903 16911 14909
rect 17604 14872 17632 14980
rect 18785 14977 18797 15011
rect 18831 15008 18843 15011
rect 20346 15008 20352 15020
rect 18831 14980 20352 15008
rect 18831 14977 18843 14980
rect 18785 14971 18843 14977
rect 20346 14968 20352 14980
rect 20404 14968 20410 15020
rect 20530 14968 20536 15020
rect 20588 15008 20594 15020
rect 22370 15008 22376 15020
rect 20588 14980 22376 15008
rect 20588 14968 20594 14980
rect 22370 14968 22376 14980
rect 22428 14968 22434 15020
rect 22554 14968 22560 15020
rect 22612 15008 22618 15020
rect 24397 15011 24455 15017
rect 24397 15008 24409 15011
rect 22612 14980 24409 15008
rect 22612 14968 22618 14980
rect 24397 14977 24409 14980
rect 24443 14977 24455 15011
rect 25038 15008 25044 15020
rect 24999 14980 25044 15008
rect 24397 14971 24455 14977
rect 25038 14968 25044 14980
rect 25096 14968 25102 15020
rect 25222 14968 25228 15020
rect 25280 15008 25286 15020
rect 27985 15011 28043 15017
rect 25280 14980 27936 15008
rect 25280 14968 25286 14980
rect 17862 14900 17868 14952
rect 17920 14940 17926 14952
rect 18049 14943 18107 14949
rect 18049 14940 18061 14943
rect 17920 14912 18061 14940
rect 17920 14900 17926 14912
rect 18049 14909 18061 14912
rect 18095 14909 18107 14943
rect 18322 14940 18328 14952
rect 18283 14912 18328 14940
rect 18049 14903 18107 14909
rect 18322 14900 18328 14912
rect 18380 14900 18386 14952
rect 19337 14943 19395 14949
rect 19337 14909 19349 14943
rect 19383 14940 19395 14943
rect 19978 14940 19984 14952
rect 19383 14912 19984 14940
rect 19383 14909 19395 14912
rect 19337 14903 19395 14909
rect 19978 14900 19984 14912
rect 20036 14900 20042 14952
rect 20073 14943 20131 14949
rect 20073 14909 20085 14943
rect 20119 14909 20131 14943
rect 20438 14940 20444 14952
rect 20399 14912 20444 14940
rect 20073 14903 20131 14909
rect 12544 14844 17632 14872
rect 18233 14875 18291 14881
rect 18233 14841 18245 14875
rect 18279 14872 18291 14875
rect 18874 14872 18880 14884
rect 18279 14844 18880 14872
rect 18279 14841 18291 14844
rect 18233 14835 18291 14841
rect 18874 14832 18880 14844
rect 18932 14872 18938 14884
rect 19613 14875 19671 14881
rect 19613 14872 19625 14875
rect 18932 14844 19625 14872
rect 18932 14832 18938 14844
rect 19613 14841 19625 14844
rect 19659 14841 19671 14875
rect 20088 14872 20116 14903
rect 20438 14900 20444 14912
rect 20496 14900 20502 14952
rect 21910 14940 21916 14952
rect 21871 14912 21916 14940
rect 21910 14900 21916 14912
rect 21968 14900 21974 14952
rect 22281 14943 22339 14949
rect 22281 14909 22293 14943
rect 22327 14940 22339 14943
rect 23106 14940 23112 14952
rect 22327 14912 23112 14940
rect 22327 14909 22339 14912
rect 22281 14903 22339 14909
rect 23106 14900 23112 14912
rect 23164 14900 23170 14952
rect 23658 14940 23664 14952
rect 23619 14912 23664 14940
rect 23658 14900 23664 14912
rect 23716 14900 23722 14952
rect 23934 14940 23940 14952
rect 23895 14912 23940 14940
rect 23934 14900 23940 14912
rect 23992 14900 23998 14952
rect 25593 14943 25651 14949
rect 25593 14909 25605 14943
rect 25639 14940 25651 14943
rect 25869 14943 25927 14949
rect 25869 14940 25881 14943
rect 25639 14912 25881 14940
rect 25639 14909 25651 14912
rect 25593 14903 25651 14909
rect 25869 14909 25881 14912
rect 25915 14909 25927 14943
rect 25869 14903 25927 14909
rect 25961 14943 26019 14949
rect 25961 14909 25973 14943
rect 26007 14940 26019 14943
rect 26050 14940 26056 14952
rect 26007 14912 26056 14940
rect 26007 14909 26019 14912
rect 25961 14903 26019 14909
rect 20990 14872 20996 14884
rect 20088 14844 20996 14872
rect 19613 14835 19671 14841
rect 20990 14832 20996 14844
rect 21048 14832 21054 14884
rect 21453 14875 21511 14881
rect 21453 14841 21465 14875
rect 21499 14872 21511 14875
rect 23842 14872 23848 14884
rect 21499 14844 23848 14872
rect 21499 14841 21511 14844
rect 21453 14835 21511 14841
rect 23842 14832 23848 14844
rect 23900 14832 23906 14884
rect 24670 14872 24676 14884
rect 24631 14844 24676 14872
rect 24670 14832 24676 14844
rect 24728 14832 24734 14884
rect 25130 14832 25136 14884
rect 25188 14872 25194 14884
rect 25976 14872 26004 14903
rect 26050 14900 26056 14912
rect 26108 14900 26114 14952
rect 27338 14900 27344 14952
rect 27396 14940 27402 14952
rect 27798 14949 27804 14952
rect 27617 14943 27675 14949
rect 27617 14940 27629 14943
rect 27396 14912 27629 14940
rect 27396 14900 27402 14912
rect 27617 14909 27629 14912
rect 27663 14909 27675 14943
rect 27617 14903 27675 14909
rect 27764 14943 27804 14949
rect 27764 14909 27776 14943
rect 27764 14903 27804 14909
rect 27798 14900 27804 14903
rect 27856 14900 27862 14952
rect 27908 14940 27936 14980
rect 27985 14977 27997 15011
rect 28031 15008 28043 15011
rect 28166 15008 28172 15020
rect 28031 14980 28172 15008
rect 28031 14977 28043 14980
rect 27985 14971 28043 14977
rect 28166 14968 28172 14980
rect 28224 14968 28230 15020
rect 28721 15011 28779 15017
rect 28721 14977 28733 15011
rect 28767 15008 28779 15011
rect 29178 15008 29184 15020
rect 28767 14980 29184 15008
rect 28767 14977 28779 14980
rect 28721 14971 28779 14977
rect 29178 14968 29184 14980
rect 29236 14968 29242 15020
rect 30374 15008 30380 15020
rect 29288 14980 30380 15008
rect 29288 14940 29316 14980
rect 30374 14968 30380 14980
rect 30432 14968 30438 15020
rect 33152 15008 33180 15116
rect 34057 15113 34069 15116
rect 34103 15113 34115 15147
rect 34057 15107 34115 15113
rect 34238 15104 34244 15156
rect 34296 15144 34302 15156
rect 36817 15147 36875 15153
rect 36817 15144 36829 15147
rect 34296 15116 36829 15144
rect 34296 15104 34302 15116
rect 36817 15113 36829 15116
rect 36863 15113 36875 15147
rect 36817 15107 36875 15113
rect 38381 15147 38439 15153
rect 38381 15113 38393 15147
rect 38427 15144 38439 15147
rect 38654 15144 38660 15156
rect 38427 15116 38660 15144
rect 38427 15113 38439 15116
rect 38381 15107 38439 15113
rect 38654 15104 38660 15116
rect 38712 15104 38718 15156
rect 39206 15104 39212 15156
rect 39264 15144 39270 15156
rect 39850 15144 39856 15156
rect 39264 15116 39856 15144
rect 39264 15104 39270 15116
rect 39850 15104 39856 15116
rect 39908 15104 39914 15156
rect 41782 15144 41788 15156
rect 39960 15116 41788 15144
rect 33229 15079 33287 15085
rect 33229 15045 33241 15079
rect 33275 15076 33287 15079
rect 35342 15076 35348 15088
rect 33275 15048 35348 15076
rect 33275 15045 33287 15048
rect 33229 15039 33287 15045
rect 35342 15036 35348 15048
rect 35400 15036 35406 15088
rect 35710 15076 35716 15088
rect 35671 15048 35716 15076
rect 35710 15036 35716 15048
rect 35768 15036 35774 15088
rect 36078 15036 36084 15088
rect 36136 15076 36142 15088
rect 39960 15076 39988 15116
rect 41782 15104 41788 15116
rect 41840 15104 41846 15156
rect 42058 15104 42064 15156
rect 42116 15144 42122 15156
rect 42337 15147 42395 15153
rect 42337 15144 42349 15147
rect 42116 15116 42349 15144
rect 42116 15104 42122 15116
rect 42337 15113 42349 15116
rect 42383 15113 42395 15147
rect 42337 15107 42395 15113
rect 42426 15104 42432 15156
rect 42484 15144 42490 15156
rect 43901 15147 43959 15153
rect 43901 15144 43913 15147
rect 42484 15116 43913 15144
rect 42484 15104 42490 15116
rect 43901 15113 43913 15116
rect 43947 15113 43959 15147
rect 43901 15107 43959 15113
rect 47118 15104 47124 15156
rect 47176 15144 47182 15156
rect 49973 15147 50031 15153
rect 49973 15144 49985 15147
rect 47176 15116 49985 15144
rect 47176 15104 47182 15116
rect 49973 15113 49985 15116
rect 50019 15113 50031 15147
rect 51350 15144 51356 15156
rect 51311 15116 51356 15144
rect 49973 15107 50031 15113
rect 51350 15104 51356 15116
rect 51408 15104 51414 15156
rect 51537 15147 51595 15153
rect 51537 15113 51549 15147
rect 51583 15144 51595 15147
rect 51718 15144 51724 15156
rect 51583 15116 51724 15144
rect 51583 15113 51595 15116
rect 51537 15107 51595 15113
rect 51718 15104 51724 15116
rect 51776 15144 51782 15156
rect 51905 15147 51963 15153
rect 51905 15144 51917 15147
rect 51776 15116 51917 15144
rect 51776 15104 51782 15116
rect 51905 15113 51917 15116
rect 51951 15113 51963 15147
rect 51905 15107 51963 15113
rect 53282 15104 53288 15156
rect 53340 15144 53346 15156
rect 53837 15147 53895 15153
rect 53837 15144 53849 15147
rect 53340 15116 53849 15144
rect 53340 15104 53346 15116
rect 53837 15113 53849 15116
rect 53883 15113 53895 15147
rect 56870 15144 56876 15156
rect 56831 15116 56876 15144
rect 53837 15107 53895 15113
rect 56870 15104 56876 15116
rect 56928 15104 56934 15156
rect 58894 15144 58900 15156
rect 58855 15116 58900 15144
rect 58894 15104 58900 15116
rect 58952 15104 58958 15156
rect 36136 15048 39988 15076
rect 41325 15079 41383 15085
rect 36136 15036 36142 15048
rect 41325 15045 41337 15079
rect 41371 15076 41383 15079
rect 43070 15076 43076 15088
rect 41371 15048 43076 15076
rect 41371 15045 41383 15048
rect 41325 15039 41383 15045
rect 43070 15036 43076 15048
rect 43128 15036 43134 15088
rect 46753 15079 46811 15085
rect 46753 15045 46765 15079
rect 46799 15076 46811 15079
rect 47302 15076 47308 15088
rect 46799 15048 47308 15076
rect 46799 15045 46811 15048
rect 46753 15039 46811 15045
rect 47302 15036 47308 15048
rect 47360 15076 47366 15088
rect 47581 15079 47639 15085
rect 47581 15076 47593 15079
rect 47360 15048 47593 15076
rect 47360 15036 47366 15048
rect 47581 15045 47593 15048
rect 47627 15076 47639 15079
rect 49142 15076 49148 15088
rect 47627 15048 49148 15076
rect 47627 15045 47639 15048
rect 47581 15039 47639 15045
rect 49142 15036 49148 15048
rect 49200 15076 49206 15088
rect 49421 15079 49479 15085
rect 49421 15076 49433 15079
rect 49200 15048 49433 15076
rect 49200 15036 49206 15048
rect 49421 15045 49433 15048
rect 49467 15076 49479 15079
rect 49513 15079 49571 15085
rect 49513 15076 49525 15079
rect 49467 15048 49525 15076
rect 49467 15045 49479 15048
rect 49421 15039 49479 15045
rect 49513 15045 49525 15048
rect 49559 15076 49571 15079
rect 50982 15076 50988 15088
rect 49559 15048 50988 15076
rect 49559 15045 49571 15048
rect 49513 15039 49571 15045
rect 50982 15036 50988 15048
rect 51040 15076 51046 15088
rect 52641 15079 52699 15085
rect 52641 15076 52653 15079
rect 51040 15048 52653 15076
rect 51040 15036 51046 15048
rect 52641 15045 52653 15048
rect 52687 15076 52699 15079
rect 52825 15079 52883 15085
rect 52825 15076 52837 15079
rect 52687 15048 52837 15076
rect 52687 15045 52699 15048
rect 52641 15039 52699 15045
rect 52825 15045 52837 15048
rect 52871 15045 52883 15079
rect 52825 15039 52883 15045
rect 53466 15036 53472 15088
rect 53524 15076 53530 15088
rect 54205 15079 54263 15085
rect 54205 15076 54217 15079
rect 53524 15048 54217 15076
rect 53524 15036 53530 15048
rect 54205 15045 54217 15048
rect 54251 15045 54263 15079
rect 54205 15039 54263 15045
rect 33686 15008 33692 15020
rect 30484 14980 33180 15008
rect 33612 14980 33692 15008
rect 29546 14940 29552 14952
rect 27908 14912 29316 14940
rect 29507 14912 29552 14940
rect 29546 14900 29552 14912
rect 29604 14900 29610 14952
rect 29822 14900 29828 14952
rect 29880 14940 29886 14952
rect 30484 14940 30512 14980
rect 29880 14912 30512 14940
rect 30561 14943 30619 14949
rect 29880 14900 29886 14912
rect 30561 14909 30573 14943
rect 30607 14940 30619 14943
rect 30837 14943 30895 14949
rect 30837 14940 30849 14943
rect 30607 14912 30849 14940
rect 30607 14909 30619 14912
rect 30561 14903 30619 14909
rect 30837 14909 30849 14912
rect 30883 14909 30895 14943
rect 30837 14903 30895 14909
rect 31849 14943 31907 14949
rect 31849 14909 31861 14943
rect 31895 14940 31907 14943
rect 32674 14940 32680 14952
rect 31895 14912 32680 14940
rect 31895 14909 31907 14912
rect 31849 14903 31907 14909
rect 32674 14900 32680 14912
rect 32732 14900 32738 14952
rect 33612 14949 33640 14980
rect 33686 14968 33692 14980
rect 33744 14968 33750 15020
rect 34701 15011 34759 15017
rect 34701 15008 34713 15011
rect 33796 14980 34713 15008
rect 33796 14952 33824 14980
rect 34701 14977 34713 14980
rect 34747 15008 34759 15011
rect 36446 15008 36452 15020
rect 34747 14980 36452 15008
rect 34747 14977 34759 14980
rect 34701 14971 34759 14977
rect 36446 14968 36452 14980
rect 36504 14968 36510 15020
rect 36538 14968 36544 15020
rect 36596 15008 36602 15020
rect 37369 15011 37427 15017
rect 37369 15008 37381 15011
rect 36596 14980 37381 15008
rect 36596 14968 36602 14980
rect 37369 14977 37381 14980
rect 37415 14977 37427 15011
rect 37369 14971 37427 14977
rect 38654 14968 38660 15020
rect 38712 15008 38718 15020
rect 39577 15011 39635 15017
rect 38712 14980 39068 15008
rect 38712 14968 38718 14980
rect 33413 14943 33471 14949
rect 33413 14940 33425 14943
rect 32876 14912 33425 14940
rect 26418 14872 26424 14884
rect 25188 14844 26004 14872
rect 26379 14844 26424 14872
rect 25188 14832 25194 14844
rect 26418 14832 26424 14844
rect 26476 14832 26482 14884
rect 27525 14875 27583 14881
rect 27525 14841 27537 14875
rect 27571 14872 27583 14875
rect 27890 14872 27896 14884
rect 27571 14844 27896 14872
rect 27571 14841 27583 14844
rect 27525 14835 27583 14841
rect 27890 14832 27896 14844
rect 27948 14832 27954 14884
rect 29457 14875 29515 14881
rect 29457 14841 29469 14875
rect 29503 14872 29515 14875
rect 30098 14872 30104 14884
rect 29503 14844 30104 14872
rect 29503 14841 29515 14844
rect 29457 14835 29515 14841
rect 30098 14832 30104 14844
rect 30156 14832 30162 14884
rect 30929 14875 30987 14881
rect 30929 14872 30941 14875
rect 30208 14844 30941 14872
rect 7208 14776 11100 14804
rect 11238 14764 11244 14816
rect 11296 14804 11302 14816
rect 11425 14807 11483 14813
rect 11425 14804 11437 14807
rect 11296 14776 11437 14804
rect 11296 14764 11302 14776
rect 11425 14773 11437 14776
rect 11471 14773 11483 14807
rect 11425 14767 11483 14773
rect 12253 14807 12311 14813
rect 12253 14773 12265 14807
rect 12299 14804 12311 14807
rect 12894 14804 12900 14816
rect 12299 14776 12900 14804
rect 12299 14773 12311 14776
rect 12253 14767 12311 14773
rect 12894 14764 12900 14776
rect 12952 14764 12958 14816
rect 16022 14804 16028 14816
rect 15983 14776 16028 14804
rect 16022 14764 16028 14776
rect 16080 14764 16086 14816
rect 16761 14807 16819 14813
rect 16761 14773 16773 14807
rect 16807 14804 16819 14807
rect 16850 14804 16856 14816
rect 16807 14776 16856 14804
rect 16807 14773 16819 14776
rect 16761 14767 16819 14773
rect 16850 14764 16856 14776
rect 16908 14764 16914 14816
rect 17037 14807 17095 14813
rect 17037 14773 17049 14807
rect 17083 14804 17095 14807
rect 17862 14804 17868 14816
rect 17083 14776 17868 14804
rect 17083 14773 17095 14776
rect 17037 14767 17095 14773
rect 17862 14764 17868 14776
rect 17920 14804 17926 14816
rect 19153 14807 19211 14813
rect 19153 14804 19165 14807
rect 17920 14776 19165 14804
rect 17920 14764 17926 14776
rect 19153 14773 19165 14776
rect 19199 14804 19211 14807
rect 19337 14807 19395 14813
rect 19337 14804 19349 14807
rect 19199 14776 19349 14804
rect 19199 14773 19211 14776
rect 19153 14767 19211 14773
rect 19337 14773 19349 14776
rect 19383 14773 19395 14807
rect 19518 14804 19524 14816
rect 19431 14776 19524 14804
rect 19337 14767 19395 14773
rect 19518 14764 19524 14776
rect 19576 14804 19582 14816
rect 20162 14804 20168 14816
rect 19576 14776 20168 14804
rect 19576 14764 19582 14776
rect 20162 14764 20168 14776
rect 20220 14764 20226 14816
rect 22370 14764 22376 14816
rect 22428 14804 22434 14816
rect 30208 14804 30236 14844
rect 30929 14841 30941 14844
rect 30975 14841 30987 14875
rect 30929 14835 30987 14841
rect 31113 14875 31171 14881
rect 31113 14841 31125 14875
rect 31159 14872 31171 14875
rect 32876 14872 32904 14912
rect 33413 14909 33425 14912
rect 33459 14909 33471 14943
rect 33413 14903 33471 14909
rect 33597 14943 33655 14949
rect 33597 14909 33609 14943
rect 33643 14909 33655 14943
rect 33778 14940 33784 14952
rect 33691 14912 33784 14940
rect 33597 14903 33655 14909
rect 31159 14844 32904 14872
rect 33428 14872 33456 14903
rect 33778 14900 33784 14912
rect 33836 14900 33842 14952
rect 34057 14943 34115 14949
rect 34057 14909 34069 14943
rect 34103 14940 34115 14943
rect 35069 14943 35127 14949
rect 34103 14912 34468 14940
rect 34103 14909 34115 14912
rect 34057 14903 34115 14909
rect 34146 14872 34152 14884
rect 33428 14844 34152 14872
rect 31159 14841 31171 14844
rect 31113 14835 31171 14841
rect 22428 14776 30236 14804
rect 22428 14764 22434 14776
rect 30282 14764 30288 14816
rect 30340 14804 30346 14816
rect 30561 14807 30619 14813
rect 30561 14804 30573 14807
rect 30340 14776 30573 14804
rect 30340 14764 30346 14776
rect 30561 14773 30573 14776
rect 30607 14804 30619 14807
rect 30653 14807 30711 14813
rect 30653 14804 30665 14807
rect 30607 14776 30665 14804
rect 30607 14773 30619 14776
rect 30561 14767 30619 14773
rect 30653 14773 30665 14776
rect 30699 14773 30711 14807
rect 30944 14804 30972 14835
rect 34146 14832 34152 14844
rect 34204 14872 34210 14884
rect 34241 14875 34299 14881
rect 34241 14872 34253 14875
rect 34204 14844 34253 14872
rect 34204 14832 34210 14844
rect 34241 14841 34253 14844
rect 34287 14841 34299 14875
rect 34241 14835 34299 14841
rect 34330 14804 34336 14816
rect 30944 14776 34336 14804
rect 30653 14767 30711 14773
rect 34330 14764 34336 14776
rect 34388 14764 34394 14816
rect 34440 14804 34468 14912
rect 35069 14909 35081 14943
rect 35115 14940 35127 14943
rect 35158 14940 35164 14952
rect 35115 14912 35164 14940
rect 35115 14909 35127 14912
rect 35069 14903 35127 14909
rect 35158 14900 35164 14912
rect 35216 14900 35222 14952
rect 35434 14940 35440 14952
rect 35395 14912 35440 14940
rect 35434 14900 35440 14912
rect 35492 14900 35498 14952
rect 36725 14943 36783 14949
rect 36725 14940 36737 14943
rect 36372 14912 36737 14940
rect 34885 14875 34943 14881
rect 34885 14841 34897 14875
rect 34931 14872 34943 14875
rect 35618 14872 35624 14884
rect 34931 14844 35624 14872
rect 34931 14841 34943 14844
rect 34885 14835 34943 14841
rect 35618 14832 35624 14844
rect 35676 14832 35682 14884
rect 36372 14813 36400 14912
rect 36725 14909 36737 14912
rect 36771 14940 36783 14943
rect 37826 14940 37832 14952
rect 36771 14912 37832 14940
rect 36771 14909 36783 14912
rect 36725 14903 36783 14909
rect 37826 14900 37832 14912
rect 37884 14900 37890 14952
rect 37918 14900 37924 14952
rect 37976 14940 37982 14952
rect 39040 14949 39068 14980
rect 39577 14977 39589 15011
rect 39623 15008 39635 15011
rect 41046 15008 41052 15020
rect 39623 14980 41052 15008
rect 39623 14977 39635 14980
rect 39577 14971 39635 14977
rect 41046 14968 41052 14980
rect 41104 14968 41110 15020
rect 42058 15008 42064 15020
rect 41524 14980 42064 15008
rect 41524 14949 41552 14980
rect 42058 14968 42064 14980
rect 42116 14968 42122 15020
rect 42797 15011 42855 15017
rect 42797 14977 42809 15011
rect 42843 15008 42855 15011
rect 43438 15008 43444 15020
rect 42843 14980 43444 15008
rect 42843 14977 42855 14980
rect 42797 14971 42855 14977
rect 43438 14968 43444 14980
rect 43496 14968 43502 15020
rect 43622 15008 43628 15020
rect 43583 14980 43628 15008
rect 43622 14968 43628 14980
rect 43680 14968 43686 15020
rect 48961 15011 49019 15017
rect 48961 15008 48973 15011
rect 48148 14980 48973 15008
rect 48148 14952 48176 14980
rect 48961 14977 48973 14980
rect 49007 14977 49019 15011
rect 48961 14971 49019 14977
rect 51626 14968 51632 15020
rect 51684 15008 51690 15020
rect 52362 15008 52368 15020
rect 51684 14980 52368 15008
rect 51684 14968 51690 14980
rect 52362 14968 52368 14980
rect 52420 14968 52426 15020
rect 53561 15011 53619 15017
rect 53561 14977 53573 15011
rect 53607 15008 53619 15011
rect 53742 15008 53748 15020
rect 53607 14980 53748 15008
rect 53607 14977 53619 14980
rect 53561 14971 53619 14977
rect 53742 14968 53748 14980
rect 53800 14968 53806 15020
rect 63586 15008 63592 15020
rect 53944 14980 63592 15008
rect 38841 14943 38899 14949
rect 38841 14940 38853 14943
rect 37976 14912 38853 14940
rect 37976 14900 37982 14912
rect 36541 14875 36599 14881
rect 36541 14841 36553 14875
rect 36587 14872 36599 14875
rect 37182 14872 37188 14884
rect 36587 14844 37188 14872
rect 36587 14841 36599 14844
rect 36541 14835 36599 14841
rect 37182 14832 37188 14844
rect 37240 14832 37246 14884
rect 38378 14872 38384 14884
rect 37292 14844 38384 14872
rect 36357 14807 36415 14813
rect 36357 14804 36369 14807
rect 34440 14776 36369 14804
rect 36357 14773 36369 14776
rect 36403 14773 36415 14807
rect 36357 14767 36415 14773
rect 36446 14764 36452 14816
rect 36504 14804 36510 14816
rect 37292 14804 37320 14844
rect 38378 14832 38384 14844
rect 38436 14832 38442 14884
rect 37734 14804 37740 14816
rect 36504 14776 37320 14804
rect 37695 14776 37740 14804
rect 36504 14764 36510 14776
rect 37734 14764 37740 14776
rect 37792 14764 37798 14816
rect 38672 14804 38700 14912
rect 38841 14909 38853 14912
rect 38887 14909 38899 14943
rect 38841 14903 38899 14909
rect 39025 14943 39083 14949
rect 39025 14909 39037 14943
rect 39071 14909 39083 14943
rect 39025 14903 39083 14909
rect 39117 14943 39175 14949
rect 39117 14909 39129 14943
rect 39163 14940 39175 14943
rect 41509 14943 41567 14949
rect 39163 14912 40356 14940
rect 39163 14909 39175 14912
rect 39117 14903 39175 14909
rect 38749 14875 38807 14881
rect 38749 14841 38761 14875
rect 38795 14872 38807 14875
rect 40126 14872 40132 14884
rect 38795 14844 40132 14872
rect 38795 14841 38807 14844
rect 38749 14835 38807 14841
rect 40126 14832 40132 14844
rect 40184 14832 40190 14884
rect 40328 14881 40356 14912
rect 41509 14909 41521 14943
rect 41555 14909 41567 14943
rect 41509 14903 41567 14909
rect 41598 14900 41604 14952
rect 41656 14940 41662 14952
rect 41874 14940 41880 14952
rect 41656 14912 41880 14940
rect 41656 14900 41662 14912
rect 41874 14900 41880 14912
rect 41932 14900 41938 14952
rect 41969 14943 42027 14949
rect 41969 14909 41981 14943
rect 42015 14940 42027 14943
rect 42334 14940 42340 14952
rect 42015 14912 42340 14940
rect 42015 14909 42027 14912
rect 41969 14903 42027 14909
rect 42334 14900 42340 14912
rect 42392 14900 42398 14952
rect 42886 14940 42892 14952
rect 42847 14912 42892 14940
rect 42886 14900 42892 14912
rect 42944 14900 42950 14952
rect 43070 14940 43076 14952
rect 43031 14912 43076 14940
rect 43070 14900 43076 14912
rect 43128 14900 43134 14952
rect 43162 14900 43168 14952
rect 43220 14940 43226 14952
rect 43898 14940 43904 14952
rect 43220 14912 43904 14940
rect 43220 14900 43226 14912
rect 43898 14900 43904 14912
rect 43956 14900 43962 14952
rect 46477 14943 46535 14949
rect 46477 14909 46489 14943
rect 46523 14940 46535 14943
rect 46569 14943 46627 14949
rect 46569 14940 46581 14943
rect 46523 14912 46581 14940
rect 46523 14909 46535 14912
rect 46477 14903 46535 14909
rect 46569 14909 46581 14912
rect 46615 14940 46627 14943
rect 47121 14943 47179 14949
rect 47121 14940 47133 14943
rect 46615 14912 47133 14940
rect 46615 14909 46627 14912
rect 46569 14903 46627 14909
rect 47121 14909 47133 14912
rect 47167 14909 47179 14943
rect 48130 14940 48136 14952
rect 48091 14912 48136 14940
rect 47121 14903 47179 14909
rect 40313 14875 40371 14881
rect 40313 14841 40325 14875
rect 40359 14872 40371 14875
rect 41138 14872 41144 14884
rect 40359 14844 41144 14872
rect 40359 14841 40371 14844
rect 40313 14835 40371 14841
rect 41138 14832 41144 14844
rect 41196 14832 41202 14884
rect 41230 14832 41236 14884
rect 41288 14872 41294 14884
rect 46198 14872 46204 14884
rect 41288 14844 46204 14872
rect 41288 14832 41294 14844
rect 46198 14832 46204 14844
rect 46256 14872 46262 14884
rect 46293 14875 46351 14881
rect 46293 14872 46305 14875
rect 46256 14844 46305 14872
rect 46256 14832 46262 14844
rect 46293 14841 46305 14844
rect 46339 14872 46351 14875
rect 46842 14872 46848 14884
rect 46339 14844 46848 14872
rect 46339 14841 46351 14844
rect 46293 14835 46351 14841
rect 46842 14832 46848 14844
rect 46900 14832 46906 14884
rect 40586 14804 40592 14816
rect 38672 14776 40592 14804
rect 40586 14764 40592 14776
rect 40644 14764 40650 14816
rect 40678 14764 40684 14816
rect 40736 14804 40742 14816
rect 40736 14776 40781 14804
rect 40736 14764 40742 14776
rect 41782 14764 41788 14816
rect 41840 14804 41846 14816
rect 45186 14804 45192 14816
rect 41840 14776 45192 14804
rect 41840 14764 41846 14776
rect 45186 14764 45192 14776
rect 45244 14804 45250 14816
rect 46477 14807 46535 14813
rect 46477 14804 46489 14807
rect 45244 14776 46489 14804
rect 45244 14764 45250 14776
rect 46477 14773 46489 14776
rect 46523 14773 46535 14807
rect 47136 14804 47164 14903
rect 48130 14900 48136 14912
rect 48188 14900 48194 14952
rect 48222 14900 48228 14952
rect 48280 14940 48286 14952
rect 48317 14943 48375 14949
rect 48317 14940 48329 14943
rect 48280 14912 48329 14940
rect 48280 14900 48286 14912
rect 48317 14909 48329 14912
rect 48363 14909 48375 14943
rect 48317 14903 48375 14909
rect 48501 14943 48559 14949
rect 48501 14909 48513 14943
rect 48547 14940 48559 14943
rect 48774 14940 48780 14952
rect 48547 14912 48780 14940
rect 48547 14909 48559 14912
rect 48501 14903 48559 14909
rect 48774 14900 48780 14912
rect 48832 14900 48838 14952
rect 49786 14940 49792 14952
rect 49699 14912 49792 14940
rect 49786 14900 49792 14912
rect 49844 14940 49850 14952
rect 50338 14940 50344 14952
rect 49844 14912 50344 14940
rect 49844 14900 49850 14912
rect 50338 14900 50344 14912
rect 50396 14900 50402 14952
rect 51721 14943 51779 14949
rect 51721 14909 51733 14943
rect 51767 14940 51779 14943
rect 52270 14940 52276 14952
rect 51767 14912 52276 14940
rect 51767 14909 51779 14912
rect 51721 14903 51779 14909
rect 52270 14900 52276 14912
rect 52328 14900 52334 14952
rect 52822 14900 52828 14952
rect 52880 14940 52886 14952
rect 53009 14943 53067 14949
rect 53009 14940 53021 14943
rect 52880 14912 53021 14940
rect 52880 14900 52886 14912
rect 53009 14909 53021 14912
rect 53055 14909 53067 14943
rect 53009 14903 53067 14909
rect 53101 14943 53159 14949
rect 53101 14909 53113 14943
rect 53147 14940 53159 14943
rect 53834 14940 53840 14952
rect 53147 14912 53840 14940
rect 53147 14909 53159 14912
rect 53101 14903 53159 14909
rect 53834 14900 53840 14912
rect 53892 14900 53898 14952
rect 47673 14875 47731 14881
rect 47673 14841 47685 14875
rect 47719 14872 47731 14875
rect 49697 14875 49755 14881
rect 49697 14872 49709 14875
rect 47719 14844 49709 14872
rect 47719 14841 47731 14844
rect 47673 14835 47731 14841
rect 49697 14841 49709 14844
rect 49743 14841 49755 14875
rect 49697 14835 49755 14841
rect 50985 14875 51043 14881
rect 50985 14841 50997 14875
rect 51031 14872 51043 14875
rect 51537 14875 51595 14881
rect 51537 14872 51549 14875
rect 51031 14844 51549 14872
rect 51031 14841 51043 14844
rect 50985 14835 51043 14841
rect 51537 14841 51549 14844
rect 51583 14872 51595 14875
rect 51583 14844 52684 14872
rect 51583 14841 51595 14844
rect 51537 14835 51595 14841
rect 48958 14804 48964 14816
rect 47136 14776 48964 14804
rect 46477 14767 46535 14773
rect 48958 14764 48964 14776
rect 49016 14764 49022 14816
rect 49712 14804 49740 14835
rect 50525 14807 50583 14813
rect 50525 14804 50537 14807
rect 49712 14776 50537 14804
rect 50525 14773 50537 14776
rect 50571 14773 50583 14807
rect 52656 14804 52684 14844
rect 52730 14832 52736 14884
rect 52788 14872 52794 14884
rect 53944 14872 53972 14980
rect 63586 14968 63592 14980
rect 63644 14968 63650 15020
rect 55674 14940 55680 14952
rect 55635 14912 55680 14940
rect 55674 14900 55680 14912
rect 55732 14900 55738 14952
rect 55858 14940 55864 14952
rect 55819 14912 55864 14940
rect 55858 14900 55864 14912
rect 55916 14900 55922 14952
rect 55953 14943 56011 14949
rect 55953 14909 55965 14943
rect 55999 14940 56011 14943
rect 56226 14940 56232 14952
rect 55999 14912 56232 14940
rect 55999 14909 56011 14912
rect 55953 14903 56011 14909
rect 52788 14844 53972 14872
rect 55585 14875 55643 14881
rect 52788 14832 52794 14844
rect 55585 14841 55597 14875
rect 55631 14872 55643 14875
rect 55968 14872 55996 14903
rect 56226 14900 56232 14912
rect 56284 14900 56290 14952
rect 57238 14900 57244 14952
rect 57296 14940 57302 14952
rect 57333 14943 57391 14949
rect 57333 14940 57345 14943
rect 57296 14912 57345 14940
rect 57296 14900 57302 14912
rect 57333 14909 57345 14912
rect 57379 14909 57391 14943
rect 57333 14903 57391 14909
rect 57609 14943 57667 14949
rect 57609 14909 57621 14943
rect 57655 14940 57667 14943
rect 57974 14940 57980 14952
rect 57655 14912 57980 14940
rect 57655 14909 57667 14912
rect 57609 14903 57667 14909
rect 57974 14900 57980 14912
rect 58032 14940 58038 14952
rect 58710 14940 58716 14952
rect 58032 14912 58716 14940
rect 58032 14900 58038 14912
rect 58710 14900 58716 14912
rect 58768 14900 58774 14952
rect 56410 14872 56416 14884
rect 55631 14844 55996 14872
rect 56371 14844 56416 14872
rect 55631 14841 55643 14844
rect 55585 14835 55643 14841
rect 56410 14832 56416 14844
rect 56468 14832 56474 14884
rect 55490 14804 55496 14816
rect 52656 14776 55496 14804
rect 50525 14767 50583 14773
rect 55490 14764 55496 14776
rect 55548 14764 55554 14816
rect 1104 14714 63480 14736
rect 1104 14662 21774 14714
rect 21826 14662 21838 14714
rect 21890 14662 21902 14714
rect 21954 14662 21966 14714
rect 22018 14662 42566 14714
rect 42618 14662 42630 14714
rect 42682 14662 42694 14714
rect 42746 14662 42758 14714
rect 42810 14662 63480 14714
rect 1104 14640 63480 14662
rect 4890 14560 4896 14612
rect 4948 14600 4954 14612
rect 10689 14603 10747 14609
rect 10689 14600 10701 14603
rect 4948 14572 10701 14600
rect 4948 14560 4954 14572
rect 10689 14569 10701 14572
rect 10735 14569 10747 14603
rect 10689 14563 10747 14569
rect 10778 14560 10784 14612
rect 10836 14600 10842 14612
rect 10873 14603 10931 14609
rect 10873 14600 10885 14603
rect 10836 14572 10885 14600
rect 10836 14560 10842 14572
rect 10873 14569 10885 14572
rect 10919 14600 10931 14603
rect 14185 14603 14243 14609
rect 14185 14600 14197 14603
rect 10919 14572 14197 14600
rect 10919 14569 10931 14572
rect 10873 14563 10931 14569
rect 14185 14569 14197 14572
rect 14231 14600 14243 14603
rect 18874 14600 18880 14612
rect 14231 14572 17816 14600
rect 18835 14572 18880 14600
rect 14231 14569 14243 14572
rect 14185 14563 14243 14569
rect 7466 14532 7472 14544
rect 5828 14504 7472 14532
rect 5828 14473 5856 14504
rect 7466 14492 7472 14504
rect 7524 14492 7530 14544
rect 7926 14492 7932 14544
rect 7984 14532 7990 14544
rect 8757 14535 8815 14541
rect 8757 14532 8769 14535
rect 7984 14504 8769 14532
rect 7984 14492 7990 14504
rect 5813 14467 5871 14473
rect 5813 14433 5825 14467
rect 5859 14433 5871 14467
rect 5994 14464 6000 14476
rect 5955 14436 6000 14464
rect 5813 14427 5871 14433
rect 5994 14424 6000 14436
rect 6052 14424 6058 14476
rect 6089 14467 6147 14473
rect 6089 14433 6101 14467
rect 6135 14464 6147 14467
rect 6641 14467 6699 14473
rect 6641 14464 6653 14467
rect 6135 14436 6653 14464
rect 6135 14433 6147 14436
rect 6089 14427 6147 14433
rect 6641 14433 6653 14436
rect 6687 14433 6699 14467
rect 7834 14464 7840 14476
rect 7795 14436 7840 14464
rect 6641 14427 6699 14433
rect 7834 14424 7840 14436
rect 7892 14464 7898 14476
rect 8110 14464 8116 14476
rect 7892 14436 8116 14464
rect 7892 14424 7898 14436
rect 8110 14424 8116 14436
rect 8168 14424 8174 14476
rect 8312 14473 8340 14504
rect 8757 14501 8769 14504
rect 8803 14532 8815 14535
rect 13173 14535 13231 14541
rect 8803 14504 10456 14532
rect 8803 14501 8815 14504
rect 8757 14495 8815 14501
rect 10428 14476 10456 14504
rect 13173 14501 13185 14535
rect 13219 14532 13231 14535
rect 14090 14532 14096 14544
rect 13219 14504 14096 14532
rect 13219 14501 13231 14504
rect 13173 14495 13231 14501
rect 14090 14492 14096 14504
rect 14148 14492 14154 14544
rect 17788 14532 17816 14572
rect 18874 14560 18880 14572
rect 18932 14560 18938 14612
rect 20530 14600 20536 14612
rect 20491 14572 20536 14600
rect 20530 14560 20536 14572
rect 20588 14560 20594 14612
rect 20640 14572 30328 14600
rect 20640 14532 20668 14572
rect 17788 14504 20668 14532
rect 20714 14492 20720 14544
rect 20772 14532 20778 14544
rect 21634 14532 21640 14544
rect 20772 14504 21640 14532
rect 20772 14492 20778 14504
rect 21634 14492 21640 14504
rect 21692 14492 21698 14544
rect 23842 14532 23848 14544
rect 23803 14504 23848 14532
rect 23842 14492 23848 14504
rect 23900 14492 23906 14544
rect 26418 14492 26424 14544
rect 26476 14532 26482 14544
rect 27709 14535 27767 14541
rect 27709 14532 27721 14535
rect 26476 14504 27721 14532
rect 26476 14492 26482 14504
rect 27709 14501 27721 14504
rect 27755 14532 27767 14535
rect 28258 14532 28264 14544
rect 27755 14504 28264 14532
rect 27755 14501 27767 14504
rect 27709 14495 27767 14501
rect 28258 14492 28264 14504
rect 28316 14492 28322 14544
rect 29362 14532 29368 14544
rect 29323 14504 29368 14532
rect 29362 14492 29368 14504
rect 29420 14492 29426 14544
rect 8205 14467 8263 14473
rect 8205 14433 8217 14467
rect 8251 14433 8263 14467
rect 8205 14427 8263 14433
rect 8297 14467 8355 14473
rect 8297 14433 8309 14467
rect 8343 14464 8355 14467
rect 9674 14464 9680 14476
rect 8343 14436 8377 14464
rect 9635 14436 9680 14464
rect 8343 14433 8355 14436
rect 8297 14427 8355 14433
rect 6012 14396 6040 14424
rect 7377 14399 7435 14405
rect 7377 14396 7389 14399
rect 6012 14368 7389 14396
rect 7377 14365 7389 14368
rect 7423 14365 7435 14399
rect 8220 14396 8248 14427
rect 9674 14424 9680 14436
rect 9732 14424 9738 14476
rect 9858 14464 9864 14476
rect 9819 14436 9864 14464
rect 9858 14424 9864 14436
rect 9916 14424 9922 14476
rect 10410 14424 10416 14476
rect 10468 14464 10474 14476
rect 11241 14467 11299 14473
rect 11241 14464 11253 14467
rect 10468 14436 11253 14464
rect 10468 14424 10474 14436
rect 11241 14433 11253 14436
rect 11287 14464 11299 14467
rect 13446 14464 13452 14476
rect 11287 14436 13452 14464
rect 11287 14433 11299 14436
rect 11241 14427 11299 14433
rect 13446 14424 13452 14436
rect 13504 14424 13510 14476
rect 14001 14467 14059 14473
rect 14001 14433 14013 14467
rect 14047 14464 14059 14467
rect 14274 14464 14280 14476
rect 14047 14436 14280 14464
rect 14047 14433 14059 14436
rect 14001 14427 14059 14433
rect 14274 14424 14280 14436
rect 14332 14424 14338 14476
rect 15289 14467 15347 14473
rect 15289 14433 15301 14467
rect 15335 14464 15347 14467
rect 15930 14464 15936 14476
rect 15335 14436 15936 14464
rect 15335 14433 15347 14436
rect 15289 14427 15347 14433
rect 15930 14424 15936 14436
rect 15988 14424 15994 14476
rect 16022 14424 16028 14476
rect 16080 14464 16086 14476
rect 18509 14467 18567 14473
rect 16080 14436 17264 14464
rect 16080 14424 16086 14436
rect 8938 14396 8944 14408
rect 8220 14368 8944 14396
rect 7377 14359 7435 14365
rect 8938 14356 8944 14368
rect 8996 14356 9002 14408
rect 10229 14399 10287 14405
rect 10229 14365 10241 14399
rect 10275 14396 10287 14399
rect 10318 14396 10324 14408
rect 10275 14368 10324 14396
rect 10275 14365 10287 14368
rect 10229 14359 10287 14365
rect 10318 14356 10324 14368
rect 10376 14356 10382 14408
rect 11514 14396 11520 14408
rect 11475 14368 11520 14396
rect 11514 14356 11520 14368
rect 11572 14356 11578 14408
rect 11793 14399 11851 14405
rect 11793 14365 11805 14399
rect 11839 14396 11851 14399
rect 12434 14396 12440 14408
rect 11839 14368 12440 14396
rect 11839 14365 11851 14368
rect 11793 14359 11851 14365
rect 12434 14356 12440 14368
rect 12492 14356 12498 14408
rect 16850 14396 16856 14408
rect 16811 14368 16856 14396
rect 16850 14356 16856 14368
rect 16908 14356 16914 14408
rect 17126 14396 17132 14408
rect 17087 14368 17132 14396
rect 17126 14356 17132 14368
rect 17184 14356 17190 14408
rect 17236 14396 17264 14436
rect 18509 14433 18521 14467
rect 18555 14464 18567 14467
rect 19613 14467 19671 14473
rect 19613 14464 19625 14467
rect 18555 14436 19625 14464
rect 18555 14433 18567 14436
rect 18509 14427 18567 14433
rect 19613 14433 19625 14436
rect 19659 14464 19671 14467
rect 19886 14464 19892 14476
rect 19659 14436 19892 14464
rect 19659 14433 19671 14436
rect 19613 14427 19671 14433
rect 19886 14424 19892 14436
rect 19944 14464 19950 14476
rect 19981 14467 20039 14473
rect 19981 14464 19993 14467
rect 19944 14436 19993 14464
rect 19944 14424 19950 14436
rect 19981 14433 19993 14436
rect 20027 14464 20039 14467
rect 24854 14464 24860 14476
rect 20027 14436 24860 14464
rect 20027 14433 20039 14436
rect 19981 14427 20039 14433
rect 24854 14424 24860 14436
rect 24912 14424 24918 14476
rect 25130 14464 25136 14476
rect 25091 14436 25136 14464
rect 25130 14424 25136 14436
rect 25188 14424 25194 14476
rect 25774 14424 25780 14476
rect 25832 14464 25838 14476
rect 26605 14467 26663 14473
rect 26605 14464 26617 14467
rect 25832 14436 26617 14464
rect 25832 14424 25838 14436
rect 26605 14433 26617 14436
rect 26651 14433 26663 14467
rect 27154 14464 27160 14476
rect 27115 14436 27160 14464
rect 26605 14427 26663 14433
rect 27154 14424 27160 14436
rect 27212 14424 27218 14476
rect 28445 14467 28503 14473
rect 28445 14433 28457 14467
rect 28491 14464 28503 14467
rect 29546 14464 29552 14476
rect 28491 14436 29552 14464
rect 28491 14433 28503 14436
rect 28445 14427 28503 14433
rect 29546 14424 29552 14436
rect 29604 14464 29610 14476
rect 29733 14467 29791 14473
rect 29733 14464 29745 14467
rect 29604 14436 29745 14464
rect 29604 14424 29610 14436
rect 29733 14433 29745 14436
rect 29779 14433 29791 14467
rect 30190 14464 30196 14476
rect 30151 14436 30196 14464
rect 29733 14427 29791 14433
rect 30190 14424 30196 14436
rect 30248 14424 30254 14476
rect 30300 14464 30328 14572
rect 30374 14560 30380 14612
rect 30432 14600 30438 14612
rect 32306 14600 32312 14612
rect 30432 14572 32312 14600
rect 30432 14560 30438 14572
rect 32306 14560 32312 14572
rect 32364 14560 32370 14612
rect 32401 14603 32459 14609
rect 32401 14569 32413 14603
rect 32447 14600 32459 14603
rect 32490 14600 32496 14612
rect 32447 14572 32496 14600
rect 32447 14569 32459 14572
rect 32401 14563 32459 14569
rect 32490 14560 32496 14572
rect 32548 14560 32554 14612
rect 34146 14600 34152 14612
rect 32600 14572 33732 14600
rect 34107 14572 34152 14600
rect 30929 14535 30987 14541
rect 30929 14501 30941 14535
rect 30975 14532 30987 14535
rect 31754 14532 31760 14544
rect 30975 14504 31760 14532
rect 30975 14501 30987 14504
rect 30929 14495 30987 14501
rect 31754 14492 31760 14504
rect 31812 14492 31818 14544
rect 32600 14532 32628 14572
rect 32324 14504 32628 14532
rect 33704 14532 33732 14572
rect 34146 14560 34152 14572
rect 34204 14560 34210 14612
rect 34330 14560 34336 14612
rect 34388 14600 34394 14612
rect 34698 14600 34704 14612
rect 34388 14572 34704 14600
rect 34388 14560 34394 14572
rect 34698 14560 34704 14572
rect 34756 14560 34762 14612
rect 37182 14560 37188 14612
rect 37240 14600 37246 14612
rect 40310 14600 40316 14612
rect 37240 14572 40316 14600
rect 37240 14560 37246 14572
rect 40310 14560 40316 14572
rect 40368 14560 40374 14612
rect 42242 14560 42248 14612
rect 42300 14600 42306 14612
rect 42705 14603 42763 14609
rect 42705 14600 42717 14603
rect 42300 14572 42717 14600
rect 42300 14560 42306 14572
rect 42705 14569 42717 14572
rect 42751 14600 42763 14603
rect 42981 14603 43039 14609
rect 42981 14600 42993 14603
rect 42751 14572 42993 14600
rect 42751 14569 42763 14572
rect 42705 14563 42763 14569
rect 42981 14569 42993 14572
rect 43027 14569 43039 14603
rect 47121 14603 47179 14609
rect 42981 14563 43039 14569
rect 43088 14572 46520 14600
rect 33704 14504 34284 14532
rect 32324 14464 32352 14504
rect 30300 14436 32352 14464
rect 32490 14424 32496 14476
rect 32548 14464 32554 14476
rect 33318 14464 33324 14476
rect 32548 14436 33324 14464
rect 32548 14424 32554 14436
rect 33318 14424 33324 14436
rect 33376 14464 33382 14476
rect 34146 14464 34152 14476
rect 33376 14436 34152 14464
rect 33376 14424 33382 14436
rect 34146 14424 34152 14436
rect 34204 14424 34210 14476
rect 21542 14396 21548 14408
rect 17236 14368 21548 14396
rect 21542 14356 21548 14368
rect 21600 14356 21606 14408
rect 21634 14356 21640 14408
rect 21692 14396 21698 14408
rect 21821 14399 21879 14405
rect 21821 14396 21833 14399
rect 21692 14368 21833 14396
rect 21692 14356 21698 14368
rect 21821 14365 21833 14368
rect 21867 14365 21879 14399
rect 21821 14359 21879 14365
rect 22097 14399 22155 14405
rect 22097 14365 22109 14399
rect 22143 14396 22155 14399
rect 22554 14396 22560 14408
rect 22143 14368 22560 14396
rect 22143 14365 22155 14368
rect 22097 14359 22155 14365
rect 22554 14356 22560 14368
rect 22612 14356 22618 14408
rect 25038 14396 25044 14408
rect 24999 14368 25044 14396
rect 25038 14356 25044 14368
rect 25096 14356 25102 14408
rect 25593 14399 25651 14405
rect 25593 14365 25605 14399
rect 25639 14396 25651 14399
rect 27522 14396 27528 14408
rect 25639 14368 27528 14396
rect 25639 14365 25651 14368
rect 25593 14359 25651 14365
rect 27522 14356 27528 14368
rect 27580 14356 27586 14408
rect 27856 14399 27914 14405
rect 27856 14365 27868 14399
rect 27902 14396 27914 14399
rect 27982 14396 27988 14408
rect 27902 14368 27988 14396
rect 27902 14365 27914 14368
rect 27856 14359 27914 14365
rect 27982 14356 27988 14368
rect 28040 14356 28046 14408
rect 28077 14399 28135 14405
rect 28077 14365 28089 14399
rect 28123 14396 28135 14399
rect 28166 14396 28172 14408
rect 28123 14368 28172 14396
rect 28123 14365 28135 14368
rect 28077 14359 28135 14365
rect 28166 14356 28172 14368
rect 28224 14356 28230 14408
rect 28350 14356 28356 14408
rect 28408 14396 28414 14408
rect 30098 14396 30104 14408
rect 28408 14368 30104 14396
rect 28408 14356 28414 14368
rect 30098 14356 30104 14368
rect 30156 14356 30162 14408
rect 30561 14399 30619 14405
rect 30561 14365 30573 14399
rect 30607 14396 30619 14399
rect 31202 14396 31208 14408
rect 30607 14368 31208 14396
rect 30607 14365 30619 14368
rect 30561 14359 30619 14365
rect 5350 14288 5356 14340
rect 5408 14328 5414 14340
rect 11146 14328 11152 14340
rect 5408 14300 11152 14328
rect 5408 14288 5414 14300
rect 11146 14288 11152 14300
rect 11204 14288 11210 14340
rect 16390 14328 16396 14340
rect 13832 14300 16396 14328
rect 5629 14263 5687 14269
rect 5629 14229 5641 14263
rect 5675 14260 5687 14263
rect 5718 14260 5724 14272
rect 5675 14232 5724 14260
rect 5675 14229 5687 14232
rect 5629 14223 5687 14229
rect 5718 14220 5724 14232
rect 5776 14220 5782 14272
rect 6270 14260 6276 14272
rect 6231 14232 6276 14260
rect 6270 14220 6276 14232
rect 6328 14220 6334 14272
rect 6641 14263 6699 14269
rect 6641 14229 6653 14263
rect 6687 14260 6699 14263
rect 6917 14263 6975 14269
rect 6917 14260 6929 14263
rect 6687 14232 6929 14260
rect 6687 14229 6699 14232
rect 6641 14223 6699 14229
rect 6917 14229 6929 14232
rect 6963 14260 6975 14263
rect 7098 14260 7104 14272
rect 6963 14232 7104 14260
rect 6963 14229 6975 14232
rect 6917 14223 6975 14229
rect 7098 14220 7104 14232
rect 7156 14220 7162 14272
rect 9309 14263 9367 14269
rect 9309 14229 9321 14263
rect 9355 14260 9367 14263
rect 9490 14260 9496 14272
rect 9355 14232 9496 14260
rect 9355 14229 9367 14232
rect 9309 14223 9367 14229
rect 9490 14220 9496 14232
rect 9548 14220 9554 14272
rect 10689 14263 10747 14269
rect 10689 14229 10701 14263
rect 10735 14260 10747 14263
rect 13832 14260 13860 14300
rect 16390 14288 16396 14300
rect 16448 14288 16454 14340
rect 27540 14328 27568 14356
rect 29270 14328 29276 14340
rect 27540 14300 29276 14328
rect 29270 14288 29276 14300
rect 29328 14288 29334 14340
rect 30576 14328 30604 14359
rect 31202 14356 31208 14368
rect 31260 14356 31266 14408
rect 32766 14396 32772 14408
rect 32727 14368 32772 14396
rect 32766 14356 32772 14368
rect 32824 14356 32830 14408
rect 33042 14396 33048 14408
rect 33003 14368 33048 14396
rect 33042 14356 33048 14368
rect 33100 14356 33106 14408
rect 34256 14396 34284 14504
rect 35342 14492 35348 14544
rect 35400 14532 35406 14544
rect 35437 14535 35495 14541
rect 35437 14532 35449 14535
rect 35400 14504 35449 14532
rect 35400 14492 35406 14504
rect 35437 14501 35449 14504
rect 35483 14532 35495 14535
rect 36354 14532 36360 14544
rect 35483 14504 36360 14532
rect 35483 14501 35495 14504
rect 35437 14495 35495 14501
rect 36354 14492 36360 14504
rect 36412 14492 36418 14544
rect 37553 14535 37611 14541
rect 37553 14501 37565 14535
rect 37599 14532 37611 14535
rect 38105 14535 38163 14541
rect 38105 14532 38117 14535
rect 37599 14504 38117 14532
rect 37599 14501 37611 14504
rect 37553 14495 37611 14501
rect 38105 14501 38117 14504
rect 38151 14532 38163 14535
rect 39022 14532 39028 14544
rect 38151 14504 39028 14532
rect 38151 14501 38163 14504
rect 38105 14495 38163 14501
rect 39022 14492 39028 14504
rect 39080 14492 39086 14544
rect 39850 14492 39856 14544
rect 39908 14532 39914 14544
rect 40770 14532 40776 14544
rect 39908 14504 40172 14532
rect 39908 14492 39914 14504
rect 35529 14467 35587 14473
rect 35529 14433 35541 14467
rect 35575 14464 35587 14467
rect 36262 14464 36268 14476
rect 35575 14436 36268 14464
rect 35575 14433 35587 14436
rect 35529 14427 35587 14433
rect 36262 14424 36268 14436
rect 36320 14424 36326 14476
rect 37918 14464 37924 14476
rect 37879 14436 37924 14464
rect 37918 14424 37924 14436
rect 37976 14424 37982 14476
rect 38194 14424 38200 14476
rect 38252 14464 38258 14476
rect 38252 14436 38297 14464
rect 38252 14424 38258 14436
rect 38378 14424 38384 14476
rect 38436 14464 38442 14476
rect 39945 14467 40003 14473
rect 38436 14436 39160 14464
rect 38436 14424 38442 14436
rect 35253 14399 35311 14405
rect 35253 14396 35265 14399
rect 34256 14368 35265 14396
rect 35253 14365 35265 14368
rect 35299 14396 35311 14399
rect 36078 14396 36084 14408
rect 35299 14368 36084 14396
rect 35299 14365 35311 14368
rect 35253 14359 35311 14365
rect 36078 14356 36084 14368
rect 36136 14356 36142 14408
rect 37936 14396 37964 14424
rect 38933 14399 38991 14405
rect 38933 14396 38945 14399
rect 37936 14368 38945 14396
rect 38933 14365 38945 14368
rect 38979 14365 38991 14399
rect 38933 14359 38991 14365
rect 29380 14300 30604 14328
rect 31573 14331 31631 14337
rect 10735 14232 13860 14260
rect 13909 14263 13967 14269
rect 10735 14229 10747 14232
rect 10689 14223 10747 14229
rect 13909 14229 13921 14263
rect 13955 14260 13967 14263
rect 13998 14260 14004 14272
rect 13955 14232 14004 14260
rect 13955 14229 13967 14232
rect 13909 14223 13967 14229
rect 13998 14220 14004 14232
rect 14056 14220 14062 14272
rect 14734 14260 14740 14272
rect 14695 14232 14740 14260
rect 14734 14220 14740 14232
rect 14792 14220 14798 14272
rect 14826 14220 14832 14272
rect 14884 14260 14890 14272
rect 15473 14263 15531 14269
rect 15473 14260 15485 14263
rect 14884 14232 15485 14260
rect 14884 14220 14890 14232
rect 15473 14229 15485 14232
rect 15519 14229 15531 14263
rect 15930 14260 15936 14272
rect 15891 14232 15936 14260
rect 15473 14223 15531 14229
rect 15930 14220 15936 14232
rect 15988 14220 15994 14272
rect 16301 14263 16359 14269
rect 16301 14229 16313 14263
rect 16347 14260 16359 14263
rect 16574 14260 16580 14272
rect 16347 14232 16580 14260
rect 16347 14229 16359 14232
rect 16301 14223 16359 14229
rect 16574 14220 16580 14232
rect 16632 14220 16638 14272
rect 16758 14260 16764 14272
rect 16719 14232 16764 14260
rect 16758 14220 16764 14232
rect 16816 14220 16822 14272
rect 18322 14220 18328 14272
rect 18380 14260 18386 14272
rect 19245 14263 19303 14269
rect 19245 14260 19257 14263
rect 18380 14232 19257 14260
rect 18380 14220 18386 14232
rect 19245 14229 19257 14232
rect 19291 14260 19303 14263
rect 19978 14260 19984 14272
rect 19291 14232 19984 14260
rect 19291 14229 19303 14232
rect 19245 14223 19303 14229
rect 19978 14220 19984 14232
rect 20036 14220 20042 14272
rect 20714 14220 20720 14272
rect 20772 14260 20778 14272
rect 21085 14263 21143 14269
rect 21085 14260 21097 14263
rect 20772 14232 21097 14260
rect 20772 14220 20778 14232
rect 21085 14229 21097 14232
rect 21131 14229 21143 14263
rect 21085 14223 21143 14229
rect 21358 14220 21364 14272
rect 21416 14260 21422 14272
rect 21453 14263 21511 14269
rect 21453 14260 21465 14263
rect 21416 14232 21465 14260
rect 21416 14220 21422 14232
rect 21453 14229 21465 14232
rect 21499 14229 21511 14263
rect 23382 14260 23388 14272
rect 23343 14232 23388 14260
rect 21453 14223 21511 14229
rect 23382 14220 23388 14232
rect 23440 14220 23446 14272
rect 23566 14220 23572 14272
rect 23624 14260 23630 14272
rect 23934 14260 23940 14272
rect 23624 14232 23940 14260
rect 23624 14220 23630 14232
rect 23934 14220 23940 14232
rect 23992 14260 23998 14272
rect 24213 14263 24271 14269
rect 24213 14260 24225 14263
rect 23992 14232 24225 14260
rect 23992 14220 23998 14232
rect 24213 14229 24225 14232
rect 24259 14229 24271 14263
rect 24213 14223 24271 14229
rect 25774 14220 25780 14272
rect 25832 14260 25838 14272
rect 25869 14263 25927 14269
rect 25869 14260 25881 14263
rect 25832 14232 25881 14260
rect 25832 14220 25838 14232
rect 25869 14229 25881 14232
rect 25915 14229 25927 14263
rect 26234 14260 26240 14272
rect 26195 14232 26240 14260
rect 25869 14223 25927 14229
rect 26234 14220 26240 14232
rect 26292 14220 26298 14272
rect 26786 14260 26792 14272
rect 26747 14232 26792 14260
rect 26786 14220 26792 14232
rect 26844 14220 26850 14272
rect 27338 14220 27344 14272
rect 27396 14260 27402 14272
rect 27525 14263 27583 14269
rect 27525 14260 27537 14263
rect 27396 14232 27537 14260
rect 27396 14220 27402 14232
rect 27525 14229 27537 14232
rect 27571 14229 27583 14263
rect 27525 14223 27583 14229
rect 27985 14263 28043 14269
rect 27985 14229 27997 14263
rect 28031 14260 28043 14263
rect 28810 14260 28816 14272
rect 28031 14232 28816 14260
rect 28031 14229 28043 14232
rect 27985 14223 28043 14229
rect 28810 14220 28816 14232
rect 28868 14220 28874 14272
rect 28902 14220 28908 14272
rect 28960 14260 28966 14272
rect 29380 14260 29408 14300
rect 31573 14297 31585 14331
rect 31619 14328 31631 14331
rect 34790 14328 34796 14340
rect 31619 14300 32812 14328
rect 34703 14300 34796 14328
rect 31619 14297 31631 14300
rect 31573 14291 31631 14297
rect 30374 14269 30380 14272
rect 28960 14232 29408 14260
rect 30358 14263 30380 14269
rect 28960 14220 28966 14232
rect 30358 14229 30370 14263
rect 30358 14223 30380 14229
rect 30374 14220 30380 14223
rect 30432 14220 30438 14272
rect 30466 14220 30472 14272
rect 30524 14260 30530 14272
rect 31938 14260 31944 14272
rect 30524 14232 30569 14260
rect 31899 14232 31944 14260
rect 30524 14220 30530 14232
rect 31938 14220 31944 14232
rect 31996 14220 32002 14272
rect 32784 14260 32812 14300
rect 34790 14288 34796 14300
rect 34848 14328 34854 14340
rect 39022 14328 39028 14340
rect 34848 14300 39028 14328
rect 34848 14288 34854 14300
rect 39022 14288 39028 14300
rect 39080 14288 39086 14340
rect 39132 14328 39160 14436
rect 39945 14433 39957 14467
rect 39991 14464 40003 14467
rect 40034 14464 40040 14476
rect 39991 14436 40040 14464
rect 39991 14433 40003 14436
rect 39945 14427 40003 14433
rect 40034 14424 40040 14436
rect 40092 14424 40098 14476
rect 40144 14473 40172 14504
rect 40328 14504 40776 14532
rect 40328 14473 40356 14504
rect 40770 14492 40776 14504
rect 40828 14532 40834 14544
rect 40865 14535 40923 14541
rect 40865 14532 40877 14535
rect 40828 14504 40877 14532
rect 40828 14492 40834 14504
rect 40865 14501 40877 14504
rect 40911 14532 40923 14535
rect 41598 14532 41604 14544
rect 40911 14504 41604 14532
rect 40911 14501 40923 14504
rect 40865 14495 40923 14501
rect 41598 14492 41604 14504
rect 41656 14492 41662 14544
rect 41690 14492 41696 14544
rect 41748 14532 41754 14544
rect 41785 14535 41843 14541
rect 41785 14532 41797 14535
rect 41748 14504 41797 14532
rect 41748 14492 41754 14504
rect 41785 14501 41797 14504
rect 41831 14501 41843 14535
rect 42058 14532 42064 14544
rect 41785 14495 41843 14501
rect 41892 14504 42064 14532
rect 40129 14467 40187 14473
rect 40129 14433 40141 14467
rect 40175 14433 40187 14467
rect 40129 14427 40187 14433
rect 40313 14467 40371 14473
rect 40313 14433 40325 14467
rect 40359 14433 40371 14467
rect 40313 14427 40371 14433
rect 39298 14396 39304 14408
rect 39259 14368 39304 14396
rect 39298 14356 39304 14368
rect 39356 14356 39362 14408
rect 39482 14396 39488 14408
rect 39443 14368 39488 14396
rect 39482 14356 39488 14368
rect 39540 14356 39546 14408
rect 40144 14396 40172 14427
rect 40586 14424 40592 14476
rect 40644 14464 40650 14476
rect 41892 14473 41920 14504
rect 42058 14492 42064 14504
rect 42116 14492 42122 14544
rect 42150 14492 42156 14544
rect 42208 14532 42214 14544
rect 42337 14535 42395 14541
rect 42337 14532 42349 14535
rect 42208 14504 42349 14532
rect 42208 14492 42214 14504
rect 42337 14501 42349 14504
rect 42383 14501 42395 14535
rect 42337 14495 42395 14501
rect 41877 14467 41935 14473
rect 40644 14436 41644 14464
rect 40644 14424 40650 14436
rect 40402 14396 40408 14408
rect 40144 14368 40408 14396
rect 40402 14356 40408 14368
rect 40460 14356 40466 14408
rect 41616 14405 41644 14436
rect 41877 14433 41889 14467
rect 41923 14433 41935 14467
rect 41877 14427 41935 14433
rect 41966 14424 41972 14476
rect 42024 14464 42030 14476
rect 43088 14464 43116 14572
rect 46492 14532 46520 14572
rect 47121 14569 47133 14603
rect 47167 14600 47179 14603
rect 47486 14600 47492 14612
rect 47167 14572 47492 14600
rect 47167 14569 47179 14572
rect 47121 14563 47179 14569
rect 47486 14560 47492 14572
rect 47544 14600 47550 14612
rect 52730 14600 52736 14612
rect 47544 14572 52736 14600
rect 47544 14560 47550 14572
rect 52730 14560 52736 14572
rect 52788 14560 52794 14612
rect 52822 14560 52828 14612
rect 52880 14600 52886 14612
rect 53193 14603 53251 14609
rect 53193 14600 53205 14603
rect 52880 14572 53205 14600
rect 52880 14560 52886 14572
rect 53193 14569 53205 14572
rect 53239 14569 53251 14603
rect 53193 14563 53251 14569
rect 55766 14560 55772 14612
rect 55824 14600 55830 14612
rect 55953 14603 56011 14609
rect 55953 14600 55965 14603
rect 55824 14572 55965 14600
rect 55824 14560 55830 14572
rect 55953 14569 55965 14572
rect 55999 14569 56011 14603
rect 55953 14563 56011 14569
rect 57698 14560 57704 14612
rect 57756 14600 57762 14612
rect 58437 14603 58495 14609
rect 58437 14600 58449 14603
rect 57756 14572 58449 14600
rect 57756 14560 57762 14572
rect 58437 14569 58449 14572
rect 58483 14569 58495 14603
rect 58437 14563 58495 14569
rect 46492 14504 49096 14532
rect 42024 14436 43116 14464
rect 43349 14467 43407 14473
rect 42024 14424 42030 14436
rect 43349 14433 43361 14467
rect 43395 14464 43407 14467
rect 43438 14464 43444 14476
rect 43395 14436 43444 14464
rect 43395 14433 43407 14436
rect 43349 14427 43407 14433
rect 43438 14424 43444 14436
rect 43496 14424 43502 14476
rect 45465 14467 45523 14473
rect 45465 14433 45477 14467
rect 45511 14464 45523 14467
rect 45557 14467 45615 14473
rect 45557 14464 45569 14467
rect 45511 14436 45569 14464
rect 45511 14433 45523 14436
rect 45465 14427 45523 14433
rect 45557 14433 45569 14436
rect 45603 14464 45615 14467
rect 47394 14464 47400 14476
rect 45603 14436 47400 14464
rect 45603 14433 45615 14436
rect 45557 14427 45615 14433
rect 47394 14424 47400 14436
rect 47452 14424 47458 14476
rect 48222 14424 48228 14476
rect 48280 14464 48286 14476
rect 48501 14467 48559 14473
rect 48501 14464 48513 14467
rect 48280 14436 48513 14464
rect 48280 14424 48286 14436
rect 48501 14433 48513 14436
rect 48547 14433 48559 14467
rect 48958 14464 48964 14476
rect 48919 14436 48964 14464
rect 48501 14427 48559 14433
rect 48958 14424 48964 14436
rect 49016 14424 49022 14476
rect 49068 14464 49096 14504
rect 49142 14492 49148 14544
rect 49200 14532 49206 14544
rect 49513 14535 49571 14541
rect 49513 14532 49525 14535
rect 49200 14504 49525 14532
rect 49200 14492 49206 14504
rect 49513 14501 49525 14504
rect 49559 14501 49571 14535
rect 52270 14532 52276 14544
rect 49513 14495 49571 14501
rect 52012 14504 52276 14532
rect 52012 14464 52040 14504
rect 52270 14492 52276 14504
rect 52328 14492 52334 14544
rect 52362 14492 52368 14544
rect 52420 14532 52426 14544
rect 56778 14532 56784 14544
rect 52420 14504 54708 14532
rect 52420 14492 52426 14504
rect 52638 14464 52644 14476
rect 49068 14436 52040 14464
rect 52599 14436 52644 14464
rect 52638 14424 52644 14436
rect 52696 14424 52702 14476
rect 54680 14464 54708 14504
rect 55876 14504 56784 14532
rect 55876 14476 55904 14504
rect 56778 14492 56784 14504
rect 56836 14492 56842 14544
rect 55858 14464 55864 14476
rect 54680 14436 55864 14464
rect 55858 14424 55864 14436
rect 55916 14424 55922 14476
rect 56410 14424 56416 14476
rect 56468 14464 56474 14476
rect 57333 14467 57391 14473
rect 57333 14464 57345 14467
rect 56468 14436 57345 14464
rect 56468 14424 56474 14436
rect 57333 14433 57345 14436
rect 57379 14433 57391 14467
rect 57333 14427 57391 14433
rect 41601 14399 41659 14405
rect 41601 14365 41613 14399
rect 41647 14396 41659 14399
rect 41647 14368 41736 14396
rect 41647 14365 41659 14368
rect 41601 14359 41659 14365
rect 41230 14328 41236 14340
rect 39132 14300 41236 14328
rect 41230 14288 41236 14300
rect 41288 14288 41294 14340
rect 41708 14328 41736 14368
rect 42978 14356 42984 14408
rect 43036 14396 43042 14408
rect 44637 14399 44695 14405
rect 44637 14396 44649 14399
rect 43036 14368 44649 14396
rect 43036 14356 43042 14368
rect 44637 14365 44649 14368
rect 44683 14396 44695 14399
rect 45005 14399 45063 14405
rect 45005 14396 45017 14399
rect 44683 14368 45017 14396
rect 44683 14365 44695 14368
rect 44637 14359 44695 14365
rect 45005 14365 45017 14368
rect 45051 14365 45063 14399
rect 45830 14396 45836 14408
rect 45791 14368 45836 14396
rect 45005 14359 45063 14365
rect 45830 14356 45836 14368
rect 45888 14356 45894 14408
rect 46750 14356 46756 14408
rect 46808 14396 46814 14408
rect 47489 14399 47547 14405
rect 47489 14396 47501 14399
rect 46808 14368 47501 14396
rect 46808 14356 46814 14368
rect 47489 14365 47501 14368
rect 47535 14396 47547 14399
rect 47762 14396 47768 14408
rect 47535 14368 47768 14396
rect 47535 14365 47547 14368
rect 47489 14359 47547 14365
rect 47762 14356 47768 14368
rect 47820 14356 47826 14408
rect 50157 14399 50215 14405
rect 50157 14365 50169 14399
rect 50203 14365 50215 14399
rect 50157 14359 50215 14365
rect 50433 14399 50491 14405
rect 50433 14365 50445 14399
rect 50479 14396 50491 14399
rect 50522 14396 50528 14408
rect 50479 14368 50528 14396
rect 50479 14365 50491 14368
rect 50433 14359 50491 14365
rect 41782 14328 41788 14340
rect 41695 14300 41788 14328
rect 41782 14288 41788 14300
rect 41840 14328 41846 14340
rect 42886 14328 42892 14340
rect 41840 14300 42892 14328
rect 41840 14288 41846 14300
rect 42886 14288 42892 14300
rect 42944 14288 42950 14340
rect 43622 14288 43628 14340
rect 43680 14328 43686 14340
rect 44269 14331 44327 14337
rect 44269 14328 44281 14331
rect 43680 14300 44281 14328
rect 43680 14288 43686 14300
rect 44269 14297 44281 14300
rect 44315 14297 44327 14331
rect 44269 14291 44327 14297
rect 47394 14288 47400 14340
rect 47452 14328 47458 14340
rect 48038 14328 48044 14340
rect 47452 14300 48044 14328
rect 47452 14288 47458 14300
rect 48038 14288 48044 14300
rect 48096 14328 48102 14340
rect 50172 14328 50200 14359
rect 50522 14356 50528 14368
rect 50580 14356 50586 14408
rect 50614 14356 50620 14408
rect 50672 14396 50678 14408
rect 50672 14368 51304 14396
rect 50672 14356 50678 14368
rect 48096 14300 50200 14328
rect 51276 14328 51304 14368
rect 51350 14356 51356 14408
rect 51408 14396 51414 14408
rect 51537 14399 51595 14405
rect 51537 14396 51549 14399
rect 51408 14368 51549 14396
rect 51408 14356 51414 14368
rect 51537 14365 51549 14368
rect 51583 14365 51595 14399
rect 53374 14396 53380 14408
rect 51537 14359 51595 14365
rect 52104 14368 53380 14396
rect 52104 14337 52132 14368
rect 53374 14356 53380 14368
rect 53432 14396 53438 14408
rect 53742 14396 53748 14408
rect 53432 14368 53748 14396
rect 53432 14356 53438 14368
rect 53742 14356 53748 14368
rect 53800 14396 53806 14408
rect 54573 14399 54631 14405
rect 54573 14396 54585 14399
rect 53800 14368 54585 14396
rect 53800 14356 53806 14368
rect 54573 14365 54585 14368
rect 54619 14365 54631 14399
rect 54573 14359 54631 14365
rect 54849 14399 54907 14405
rect 54849 14365 54861 14399
rect 54895 14396 54907 14399
rect 55214 14396 55220 14408
rect 54895 14368 55220 14396
rect 54895 14365 54907 14368
rect 54849 14359 54907 14365
rect 55214 14356 55220 14368
rect 55272 14356 55278 14408
rect 55490 14356 55496 14408
rect 55548 14396 55554 14408
rect 56505 14399 56563 14405
rect 56505 14396 56517 14399
rect 55548 14368 56517 14396
rect 55548 14356 55554 14368
rect 56505 14365 56517 14368
rect 56551 14396 56563 14399
rect 56962 14396 56968 14408
rect 56551 14368 56968 14396
rect 56551 14365 56563 14368
rect 56505 14359 56563 14365
rect 56962 14356 56968 14368
rect 57020 14356 57026 14408
rect 57057 14399 57115 14405
rect 57057 14365 57069 14399
rect 57103 14396 57115 14399
rect 57238 14396 57244 14408
rect 57103 14368 57244 14396
rect 57103 14365 57115 14368
rect 57057 14359 57115 14365
rect 52089 14331 52147 14337
rect 52089 14328 52101 14331
rect 51276 14300 52101 14328
rect 48096 14288 48102 14300
rect 32950 14260 32956 14272
rect 32784 14232 32956 14260
rect 32950 14220 32956 14232
rect 33008 14220 33014 14272
rect 34882 14220 34888 14272
rect 34940 14260 34946 14272
rect 35069 14263 35127 14269
rect 35069 14260 35081 14263
rect 34940 14232 35081 14260
rect 34940 14220 34946 14232
rect 35069 14229 35081 14232
rect 35115 14229 35127 14263
rect 35710 14260 35716 14272
rect 35671 14232 35716 14260
rect 35069 14223 35127 14229
rect 35710 14220 35716 14232
rect 35768 14220 35774 14272
rect 36262 14260 36268 14272
rect 36223 14232 36268 14260
rect 36262 14220 36268 14232
rect 36320 14220 36326 14272
rect 36722 14260 36728 14272
rect 36683 14232 36728 14260
rect 36722 14220 36728 14232
rect 36780 14220 36786 14272
rect 36998 14260 37004 14272
rect 36959 14232 37004 14260
rect 36998 14220 37004 14232
rect 37056 14220 37062 14272
rect 38102 14220 38108 14272
rect 38160 14260 38166 14272
rect 38381 14263 38439 14269
rect 38381 14260 38393 14263
rect 38160 14232 38393 14260
rect 38160 14220 38166 14232
rect 38381 14229 38393 14232
rect 38427 14229 38439 14263
rect 41414 14260 41420 14272
rect 41375 14232 41420 14260
rect 38381 14223 38439 14229
rect 41414 14220 41420 14232
rect 41472 14220 41478 14272
rect 43530 14260 43536 14272
rect 43491 14232 43536 14260
rect 43530 14220 43536 14232
rect 43588 14220 43594 14272
rect 43806 14220 43812 14272
rect 43864 14260 43870 14272
rect 43901 14263 43959 14269
rect 43901 14260 43913 14263
rect 43864 14232 43913 14260
rect 43864 14220 43870 14232
rect 43901 14229 43913 14232
rect 43947 14229 43959 14263
rect 43901 14223 43959 14229
rect 48225 14263 48283 14269
rect 48225 14229 48237 14263
rect 48271 14260 48283 14263
rect 48314 14260 48320 14272
rect 48271 14232 48320 14260
rect 48271 14229 48283 14232
rect 48225 14223 48283 14229
rect 48314 14220 48320 14232
rect 48372 14220 48378 14272
rect 49142 14260 49148 14272
rect 49103 14232 49148 14260
rect 49142 14220 49148 14232
rect 49200 14220 49206 14272
rect 49602 14220 49608 14272
rect 49660 14260 49666 14272
rect 49881 14263 49939 14269
rect 49881 14260 49893 14263
rect 49660 14232 49893 14260
rect 49660 14220 49666 14232
rect 49881 14229 49893 14232
rect 49927 14229 49939 14263
rect 50172 14260 50200 14300
rect 52089 14297 52101 14300
rect 52135 14297 52147 14331
rect 57072 14328 57100 14359
rect 57238 14356 57244 14368
rect 57296 14356 57302 14408
rect 52089 14291 52147 14297
rect 56888 14300 57100 14328
rect 50614 14260 50620 14272
rect 50172 14232 50620 14260
rect 49881 14223 49939 14229
rect 50614 14220 50620 14232
rect 50672 14220 50678 14272
rect 52822 14260 52828 14272
rect 52783 14232 52828 14260
rect 52822 14220 52828 14232
rect 52880 14220 52886 14272
rect 53653 14263 53711 14269
rect 53653 14229 53665 14263
rect 53699 14260 53711 14263
rect 53834 14260 53840 14272
rect 53699 14232 53840 14260
rect 53699 14229 53711 14232
rect 53653 14223 53711 14229
rect 53834 14220 53840 14232
rect 53892 14260 53898 14272
rect 54570 14260 54576 14272
rect 53892 14232 54576 14260
rect 53892 14220 53898 14232
rect 54570 14220 54576 14232
rect 54628 14220 54634 14272
rect 55582 14220 55588 14272
rect 55640 14260 55646 14272
rect 56778 14260 56784 14272
rect 55640 14232 56784 14260
rect 55640 14220 55646 14232
rect 56778 14220 56784 14232
rect 56836 14260 56842 14272
rect 56888 14269 56916 14300
rect 56873 14263 56931 14269
rect 56873 14260 56885 14263
rect 56836 14232 56885 14260
rect 56836 14220 56842 14232
rect 56873 14229 56885 14232
rect 56919 14229 56931 14263
rect 56873 14223 56931 14229
rect 56962 14220 56968 14272
rect 57020 14260 57026 14272
rect 58989 14263 59047 14269
rect 58989 14260 59001 14263
rect 57020 14232 59001 14260
rect 57020 14220 57026 14232
rect 58989 14229 59001 14232
rect 59035 14229 59047 14263
rect 58989 14223 59047 14229
rect 1104 14170 63480 14192
rect 1104 14118 11378 14170
rect 11430 14118 11442 14170
rect 11494 14118 11506 14170
rect 11558 14118 11570 14170
rect 11622 14118 32170 14170
rect 32222 14118 32234 14170
rect 32286 14118 32298 14170
rect 32350 14118 32362 14170
rect 32414 14118 52962 14170
rect 53014 14118 53026 14170
rect 53078 14118 53090 14170
rect 53142 14118 53154 14170
rect 53206 14118 63480 14170
rect 1104 14096 63480 14118
rect 4890 14056 4896 14068
rect 4851 14028 4896 14056
rect 4890 14016 4896 14028
rect 4948 14016 4954 14068
rect 5994 14016 6000 14068
rect 6052 14056 6058 14068
rect 6549 14059 6607 14065
rect 6549 14056 6561 14059
rect 6052 14028 6561 14056
rect 6052 14016 6058 14028
rect 6549 14025 6561 14028
rect 6595 14025 6607 14059
rect 6549 14019 6607 14025
rect 6825 14059 6883 14065
rect 6825 14025 6837 14059
rect 6871 14056 6883 14059
rect 7466 14056 7472 14068
rect 6871 14028 7472 14056
rect 6871 14025 6883 14028
rect 6825 14019 6883 14025
rect 7466 14016 7472 14028
rect 7524 14056 7530 14068
rect 7561 14059 7619 14065
rect 7561 14056 7573 14059
rect 7524 14028 7573 14056
rect 7524 14016 7530 14028
rect 7561 14025 7573 14028
rect 7607 14025 7619 14059
rect 8018 14056 8024 14068
rect 7979 14028 8024 14056
rect 7561 14019 7619 14025
rect 8018 14016 8024 14028
rect 8076 14016 8082 14068
rect 8110 14016 8116 14068
rect 8168 14056 8174 14068
rect 8573 14059 8631 14065
rect 8573 14056 8585 14059
rect 8168 14028 8585 14056
rect 8168 14016 8174 14028
rect 8573 14025 8585 14028
rect 8619 14025 8631 14059
rect 8938 14056 8944 14068
rect 8899 14028 8944 14056
rect 8573 14019 8631 14025
rect 8938 14016 8944 14028
rect 8996 14016 9002 14068
rect 10778 14056 10784 14068
rect 10739 14028 10784 14056
rect 10778 14016 10784 14028
rect 10836 14016 10842 14068
rect 11238 14056 11244 14068
rect 11199 14028 11244 14056
rect 11238 14016 11244 14028
rect 11296 14016 11302 14068
rect 12069 14059 12127 14065
rect 12069 14025 12081 14059
rect 12115 14056 12127 14059
rect 12621 14059 12679 14065
rect 12621 14056 12633 14059
rect 12115 14028 12633 14056
rect 12115 14025 12127 14028
rect 12069 14019 12127 14025
rect 12621 14025 12633 14028
rect 12667 14056 12679 14059
rect 14366 14056 14372 14068
rect 12667 14028 14372 14056
rect 12667 14025 12679 14028
rect 12621 14019 12679 14025
rect 14366 14016 14372 14028
rect 14424 14016 14430 14068
rect 14734 14016 14740 14068
rect 14792 14056 14798 14068
rect 15286 14056 15292 14068
rect 14792 14028 15292 14056
rect 14792 14016 14798 14028
rect 15286 14016 15292 14028
rect 15344 14016 15350 14068
rect 16390 14056 16396 14068
rect 16303 14028 16396 14056
rect 16390 14016 16396 14028
rect 16448 14056 16454 14068
rect 20165 14059 20223 14065
rect 16448 14028 18184 14056
rect 16448 14016 16454 14028
rect 3142 13948 3148 14000
rect 3200 13988 3206 14000
rect 14093 13991 14151 13997
rect 3200 13960 13400 13988
rect 3200 13948 3206 13960
rect 4890 13920 4896 13932
rect 4172 13892 4896 13920
rect 4172 13864 4200 13892
rect 4890 13880 4896 13892
rect 4948 13880 4954 13932
rect 5626 13920 5632 13932
rect 5368 13892 5632 13920
rect 3881 13855 3939 13861
rect 3881 13821 3893 13855
rect 3927 13852 3939 13855
rect 3973 13855 4031 13861
rect 3973 13852 3985 13855
rect 3927 13824 3985 13852
rect 3927 13821 3939 13824
rect 3881 13815 3939 13821
rect 3973 13821 3985 13824
rect 4019 13852 4031 13855
rect 4019 13824 4108 13852
rect 4019 13821 4031 13824
rect 3973 13815 4031 13821
rect 4080 13784 4108 13824
rect 4154 13812 4160 13864
rect 4212 13852 4218 13864
rect 4522 13852 4528 13864
rect 4212 13824 4305 13852
rect 4483 13824 4528 13852
rect 4212 13812 4218 13824
rect 4522 13812 4528 13824
rect 4580 13812 4586 13864
rect 5368 13861 5396 13892
rect 5626 13880 5632 13892
rect 5684 13880 5690 13932
rect 5905 13923 5963 13929
rect 5905 13889 5917 13923
rect 5951 13920 5963 13923
rect 8754 13920 8760 13932
rect 5951 13892 8760 13920
rect 5951 13889 5963 13892
rect 5905 13883 5963 13889
rect 8754 13880 8760 13892
rect 8812 13880 8818 13932
rect 9125 13923 9183 13929
rect 9125 13889 9137 13923
rect 9171 13920 9183 13923
rect 9950 13920 9956 13932
rect 9171 13892 9956 13920
rect 9171 13889 9183 13892
rect 9125 13883 9183 13889
rect 9950 13880 9956 13892
rect 10008 13880 10014 13932
rect 10689 13923 10747 13929
rect 10689 13889 10701 13923
rect 10735 13920 10747 13923
rect 10735 13892 11008 13920
rect 10735 13889 10747 13892
rect 10689 13883 10747 13889
rect 5261 13855 5319 13861
rect 5261 13821 5273 13855
rect 5307 13852 5319 13855
rect 5353 13855 5411 13861
rect 5353 13852 5365 13855
rect 5307 13824 5365 13852
rect 5307 13821 5319 13824
rect 5261 13815 5319 13821
rect 5353 13821 5365 13824
rect 5399 13821 5411 13855
rect 5353 13815 5411 13821
rect 5537 13855 5595 13861
rect 5537 13821 5549 13855
rect 5583 13821 5595 13855
rect 5537 13815 5595 13821
rect 6273 13855 6331 13861
rect 6273 13821 6285 13855
rect 6319 13852 6331 13855
rect 6825 13855 6883 13861
rect 6825 13852 6837 13855
rect 6319 13824 6837 13852
rect 6319 13821 6331 13824
rect 6273 13815 6331 13821
rect 6825 13821 6837 13824
rect 6871 13821 6883 13855
rect 6825 13815 6883 13821
rect 4706 13784 4712 13796
rect 4080 13756 4712 13784
rect 4706 13744 4712 13756
rect 4764 13744 4770 13796
rect 5552 13716 5580 13815
rect 6914 13812 6920 13864
rect 6972 13852 6978 13864
rect 7009 13855 7067 13861
rect 7009 13852 7021 13855
rect 6972 13824 7021 13852
rect 6972 13812 6978 13824
rect 7009 13821 7021 13824
rect 7055 13821 7067 13855
rect 7742 13852 7748 13864
rect 7703 13824 7748 13852
rect 7009 13815 7067 13821
rect 7742 13812 7748 13824
rect 7800 13812 7806 13864
rect 7837 13855 7895 13861
rect 7837 13821 7849 13855
rect 7883 13852 7895 13855
rect 8018 13852 8024 13864
rect 7883 13824 8024 13852
rect 7883 13821 7895 13824
rect 7837 13815 7895 13821
rect 8018 13812 8024 13824
rect 8076 13812 8082 13864
rect 9217 13855 9275 13861
rect 9217 13821 9229 13855
rect 9263 13852 9275 13855
rect 9490 13852 9496 13864
rect 9263 13824 9496 13852
rect 9263 13821 9275 13824
rect 9217 13815 9275 13821
rect 9490 13812 9496 13824
rect 9548 13812 9554 13864
rect 10980 13861 11008 13892
rect 11238 13880 11244 13932
rect 11296 13920 11302 13932
rect 12069 13923 12127 13929
rect 12069 13920 12081 13923
rect 11296 13892 12081 13920
rect 11296 13880 11302 13892
rect 12069 13889 12081 13892
rect 12115 13920 12127 13923
rect 12161 13923 12219 13929
rect 12161 13920 12173 13923
rect 12115 13892 12173 13920
rect 12115 13889 12127 13892
rect 12069 13883 12127 13889
rect 12161 13889 12173 13892
rect 12207 13889 12219 13923
rect 13262 13920 13268 13932
rect 12161 13883 12219 13889
rect 12820 13892 13268 13920
rect 10965 13855 11023 13861
rect 10965 13821 10977 13855
rect 11011 13821 11023 13855
rect 10965 13815 11023 13821
rect 11057 13855 11115 13861
rect 11057 13821 11069 13855
rect 11103 13852 11115 13855
rect 11146 13852 11152 13864
rect 11103 13824 11152 13852
rect 11103 13821 11115 13824
rect 11057 13815 11115 13821
rect 9582 13744 9588 13796
rect 9640 13784 9646 13796
rect 9677 13787 9735 13793
rect 9677 13784 9689 13787
rect 9640 13756 9689 13784
rect 9640 13744 9646 13756
rect 9677 13753 9689 13756
rect 9723 13753 9735 13787
rect 10980 13784 11008 13815
rect 11146 13812 11152 13824
rect 11204 13812 11210 13864
rect 11885 13855 11943 13861
rect 11885 13821 11897 13855
rect 11931 13852 11943 13855
rect 12434 13852 12440 13864
rect 11931 13824 12440 13852
rect 11931 13821 11943 13824
rect 11885 13815 11943 13821
rect 11698 13784 11704 13796
rect 10980 13756 11704 13784
rect 9677 13747 9735 13753
rect 11698 13744 11704 13756
rect 11756 13744 11762 13796
rect 12360 13784 12388 13824
rect 12434 13812 12440 13824
rect 12492 13812 12498 13864
rect 12820 13861 12848 13892
rect 13262 13880 13268 13892
rect 13320 13880 13326 13932
rect 13372 13929 13400 13960
rect 14093 13957 14105 13991
rect 14139 13988 14151 13991
rect 14274 13988 14280 14000
rect 14139 13960 14280 13988
rect 14139 13957 14151 13960
rect 14093 13951 14151 13957
rect 14274 13948 14280 13960
rect 14332 13948 14338 14000
rect 14918 13988 14924 14000
rect 14384 13960 14924 13988
rect 13357 13923 13415 13929
rect 13357 13889 13369 13923
rect 13403 13889 13415 13923
rect 13357 13883 13415 13889
rect 13446 13880 13452 13932
rect 13504 13920 13510 13932
rect 13725 13923 13783 13929
rect 13725 13920 13737 13923
rect 13504 13892 13737 13920
rect 13504 13880 13510 13892
rect 13725 13889 13737 13892
rect 13771 13920 13783 13923
rect 13906 13920 13912 13932
rect 13771 13892 13912 13920
rect 13771 13889 13783 13892
rect 13725 13883 13783 13889
rect 13906 13880 13912 13892
rect 13964 13880 13970 13932
rect 14182 13880 14188 13932
rect 14240 13920 14246 13932
rect 14384 13920 14412 13960
rect 14918 13948 14924 13960
rect 14976 13948 14982 14000
rect 16117 13991 16175 13997
rect 16117 13988 16129 13991
rect 15212 13960 16129 13988
rect 14734 13920 14740 13932
rect 14240 13892 14412 13920
rect 14695 13892 14740 13920
rect 14240 13880 14246 13892
rect 14734 13880 14740 13892
rect 14792 13880 14798 13932
rect 12805 13855 12863 13861
rect 12805 13821 12817 13855
rect 12851 13821 12863 13855
rect 12805 13815 12863 13821
rect 12897 13855 12955 13861
rect 12897 13821 12909 13855
rect 12943 13852 12955 13855
rect 13814 13852 13820 13864
rect 12943 13824 13820 13852
rect 12943 13821 12955 13824
rect 12897 13815 12955 13821
rect 13814 13812 13820 13824
rect 13872 13852 13878 13864
rect 15212 13861 15240 13960
rect 16117 13957 16129 13960
rect 16163 13988 16175 13991
rect 17678 13988 17684 14000
rect 16163 13960 17684 13988
rect 16163 13957 16175 13960
rect 16117 13951 16175 13957
rect 17678 13948 17684 13960
rect 17736 13948 17742 14000
rect 15930 13880 15936 13932
rect 15988 13920 15994 13932
rect 16853 13923 16911 13929
rect 16853 13920 16865 13923
rect 15988 13892 16865 13920
rect 15988 13880 15994 13892
rect 16224 13864 16252 13892
rect 16853 13889 16865 13892
rect 16899 13920 16911 13923
rect 17034 13920 17040 13932
rect 16899 13892 17040 13920
rect 16899 13889 16911 13892
rect 16853 13883 16911 13889
rect 17034 13880 17040 13892
rect 17092 13880 17098 13932
rect 17126 13880 17132 13932
rect 17184 13920 17190 13932
rect 17221 13923 17279 13929
rect 17221 13920 17233 13923
rect 17184 13892 17233 13920
rect 17184 13880 17190 13892
rect 17221 13889 17233 13892
rect 17267 13920 17279 13923
rect 18049 13923 18107 13929
rect 18049 13920 18061 13923
rect 17267 13892 18061 13920
rect 17267 13889 17279 13892
rect 17221 13883 17279 13889
rect 18049 13889 18061 13892
rect 18095 13889 18107 13923
rect 18156 13920 18184 14028
rect 20165 14025 20177 14059
rect 20211 14056 20223 14059
rect 21082 14056 21088 14068
rect 20211 14028 21088 14056
rect 20211 14025 20223 14028
rect 20165 14019 20223 14025
rect 21082 14016 21088 14028
rect 21140 14016 21146 14068
rect 21174 14016 21180 14068
rect 21232 14056 21238 14068
rect 22370 14056 22376 14068
rect 21232 14028 22376 14056
rect 21232 14016 21238 14028
rect 22370 14016 22376 14028
rect 22428 14016 22434 14068
rect 22554 14056 22560 14068
rect 22515 14028 22560 14056
rect 22554 14016 22560 14028
rect 22612 14016 22618 14068
rect 24118 14016 24124 14068
rect 24176 14056 24182 14068
rect 26050 14056 26056 14068
rect 24176 14028 26056 14056
rect 24176 14016 24182 14028
rect 26050 14016 26056 14028
rect 26108 14056 26114 14068
rect 27157 14059 27215 14065
rect 26108 14028 26464 14056
rect 26108 14016 26114 14028
rect 18690 13948 18696 14000
rect 18748 13988 18754 14000
rect 19337 13991 19395 13997
rect 19337 13988 19349 13991
rect 18748 13960 19349 13988
rect 18748 13948 18754 13960
rect 19337 13957 19349 13960
rect 19383 13988 19395 13991
rect 21818 13988 21824 14000
rect 19383 13960 21824 13988
rect 19383 13957 19395 13960
rect 19337 13951 19395 13957
rect 21818 13948 21824 13960
rect 21876 13948 21882 14000
rect 22094 13988 22100 14000
rect 21928 13960 22100 13988
rect 21928 13920 21956 13960
rect 22094 13948 22100 13960
rect 22152 13948 22158 14000
rect 23845 13991 23903 13997
rect 23845 13957 23857 13991
rect 23891 13988 23903 13991
rect 24486 13988 24492 14000
rect 23891 13960 24492 13988
rect 23891 13957 23903 13960
rect 23845 13951 23903 13957
rect 24486 13948 24492 13960
rect 24544 13988 24550 14000
rect 25222 13988 25228 14000
rect 24544 13960 25228 13988
rect 24544 13948 24550 13960
rect 25222 13948 25228 13960
rect 25280 13948 25286 14000
rect 23290 13920 23296 13932
rect 18156 13892 21956 13920
rect 22112 13892 23296 13920
rect 18049 13883 18107 13889
rect 22112 13864 22140 13892
rect 23290 13880 23296 13892
rect 23348 13880 23354 13932
rect 24854 13920 24860 13932
rect 24815 13892 24860 13920
rect 24854 13880 24860 13892
rect 24912 13880 24918 13932
rect 25961 13923 26019 13929
rect 25961 13889 25973 13923
rect 26007 13920 26019 13923
rect 26053 13923 26111 13929
rect 26053 13920 26065 13923
rect 26007 13892 26065 13920
rect 26007 13889 26019 13892
rect 25961 13883 26019 13889
rect 26053 13889 26065 13892
rect 26099 13920 26111 13923
rect 26099 13892 26188 13920
rect 26099 13889 26111 13892
rect 26053 13883 26111 13889
rect 14829 13855 14887 13861
rect 13872 13824 14228 13852
rect 13872 13812 13878 13824
rect 13630 13784 13636 13796
rect 11808 13756 12296 13784
rect 12360 13756 13636 13784
rect 5718 13716 5724 13728
rect 5552 13688 5724 13716
rect 5718 13676 5724 13688
rect 5776 13716 5782 13728
rect 9306 13716 9312 13728
rect 5776 13688 9312 13716
rect 5776 13676 5782 13688
rect 9306 13676 9312 13688
rect 9364 13676 9370 13728
rect 9950 13676 9956 13728
rect 10008 13716 10014 13728
rect 10045 13719 10103 13725
rect 10045 13716 10057 13719
rect 10008 13688 10057 13716
rect 10008 13676 10014 13688
rect 10045 13685 10057 13688
rect 10091 13716 10103 13719
rect 10594 13716 10600 13728
rect 10091 13688 10600 13716
rect 10091 13685 10103 13688
rect 10045 13679 10103 13685
rect 10594 13676 10600 13688
rect 10652 13716 10658 13728
rect 11808 13716 11836 13756
rect 10652 13688 11836 13716
rect 12268 13716 12296 13756
rect 13630 13744 13636 13756
rect 13688 13744 13694 13796
rect 14200 13793 14228 13824
rect 14829 13821 14841 13855
rect 14875 13821 14887 13855
rect 14829 13815 14887 13821
rect 15197 13855 15255 13861
rect 15197 13821 15209 13855
rect 15243 13821 15255 13855
rect 15197 13815 15255 13821
rect 15289 13855 15347 13861
rect 15289 13821 15301 13855
rect 15335 13852 15347 13855
rect 15562 13852 15568 13864
rect 15335 13824 15568 13852
rect 15335 13821 15347 13824
rect 15289 13815 15347 13821
rect 14185 13787 14243 13793
rect 14185 13753 14197 13787
rect 14231 13753 14243 13787
rect 14185 13747 14243 13753
rect 14734 13744 14740 13796
rect 14792 13784 14798 13796
rect 14844 13784 14872 13815
rect 15562 13812 15568 13824
rect 15620 13812 15626 13864
rect 15749 13855 15807 13861
rect 15749 13821 15761 13855
rect 15795 13821 15807 13855
rect 16206 13852 16212 13864
rect 16119 13824 16212 13852
rect 15749 13815 15807 13821
rect 15764 13784 15792 13815
rect 16206 13812 16212 13824
rect 16264 13812 16270 13864
rect 16758 13812 16764 13864
rect 16816 13852 16822 13864
rect 18230 13852 18236 13864
rect 16816 13824 18236 13852
rect 16816 13812 16822 13824
rect 18230 13812 18236 13824
rect 18288 13812 18294 13864
rect 18509 13855 18567 13861
rect 18509 13821 18521 13855
rect 18555 13852 18567 13855
rect 18598 13852 18604 13864
rect 18555 13824 18604 13852
rect 18555 13821 18567 13824
rect 18509 13815 18567 13821
rect 18598 13812 18604 13824
rect 18656 13812 18662 13864
rect 18690 13812 18696 13864
rect 18748 13852 18754 13864
rect 18877 13855 18935 13861
rect 18748 13824 18793 13852
rect 18748 13812 18754 13824
rect 18877 13821 18889 13855
rect 18923 13852 18935 13855
rect 19886 13852 19892 13864
rect 18923 13824 19892 13852
rect 18923 13821 18935 13824
rect 18877 13815 18935 13821
rect 19886 13812 19892 13824
rect 19944 13812 19950 13864
rect 20073 13855 20131 13861
rect 20073 13821 20085 13855
rect 20119 13852 20131 13855
rect 20714 13852 20720 13864
rect 20119 13824 20720 13852
rect 20119 13821 20131 13824
rect 20073 13815 20131 13821
rect 20714 13812 20720 13824
rect 20772 13812 20778 13864
rect 20990 13812 20996 13864
rect 21048 13852 21054 13864
rect 21269 13855 21327 13861
rect 21269 13852 21281 13855
rect 21048 13824 21281 13852
rect 21048 13812 21054 13824
rect 21269 13821 21281 13824
rect 21315 13821 21327 13855
rect 21634 13852 21640 13864
rect 21269 13815 21327 13821
rect 21376 13824 21640 13852
rect 20438 13784 20444 13796
rect 14792 13756 20444 13784
rect 14792 13744 14798 13756
rect 20438 13744 20444 13756
rect 20496 13744 20502 13796
rect 21177 13787 21235 13793
rect 21177 13753 21189 13787
rect 21223 13784 21235 13787
rect 21376 13784 21404 13824
rect 21634 13812 21640 13824
rect 21692 13852 21698 13864
rect 21729 13855 21787 13861
rect 21729 13852 21741 13855
rect 21692 13824 21741 13852
rect 21692 13812 21698 13824
rect 21729 13821 21741 13824
rect 21775 13821 21787 13855
rect 21729 13815 21787 13821
rect 21818 13812 21824 13864
rect 21876 13852 21882 13864
rect 21913 13855 21971 13861
rect 21913 13852 21925 13855
rect 21876 13824 21925 13852
rect 21876 13812 21882 13824
rect 21913 13821 21925 13824
rect 21959 13821 21971 13855
rect 22094 13852 22100 13864
rect 22055 13824 22100 13852
rect 21913 13815 21971 13821
rect 21223 13756 21404 13784
rect 21928 13784 21956 13815
rect 22094 13812 22100 13824
rect 22152 13812 22158 13864
rect 23474 13812 23480 13864
rect 23532 13852 23538 13864
rect 23661 13855 23719 13861
rect 23661 13852 23673 13855
rect 23532 13824 23673 13852
rect 23532 13812 23538 13824
rect 23661 13821 23673 13824
rect 23707 13852 23719 13855
rect 24213 13855 24271 13861
rect 24213 13852 24225 13855
rect 23707 13824 24225 13852
rect 23707 13821 23719 13824
rect 23661 13815 23719 13821
rect 24213 13821 24225 13824
rect 24259 13821 24271 13855
rect 24213 13815 24271 13821
rect 24949 13855 25007 13861
rect 24949 13821 24961 13855
rect 24995 13821 25007 13855
rect 24949 13815 25007 13821
rect 25409 13855 25467 13861
rect 25409 13821 25421 13855
rect 25455 13852 25467 13855
rect 26160 13852 26188 13892
rect 26234 13880 26240 13932
rect 26292 13920 26298 13932
rect 26292 13892 26337 13920
rect 26292 13880 26298 13892
rect 26329 13855 26387 13861
rect 26329 13852 26341 13855
rect 25455 13824 26096 13852
rect 26160 13824 26341 13852
rect 25455 13821 25467 13824
rect 25409 13815 25467 13821
rect 22186 13784 22192 13796
rect 21928 13756 22192 13784
rect 21223 13753 21235 13756
rect 21177 13747 21235 13753
rect 22186 13744 22192 13756
rect 22244 13784 22250 13796
rect 22922 13784 22928 13796
rect 22244 13756 22928 13784
rect 22244 13744 22250 13756
rect 22922 13744 22928 13756
rect 22980 13744 22986 13796
rect 23014 13744 23020 13796
rect 23072 13784 23078 13796
rect 24673 13787 24731 13793
rect 24673 13784 24685 13787
rect 23072 13756 24685 13784
rect 23072 13744 23078 13756
rect 24673 13753 24685 13756
rect 24719 13784 24731 13787
rect 24964 13784 24992 13815
rect 25130 13784 25136 13796
rect 24719 13756 25136 13784
rect 24719 13753 24731 13756
rect 24673 13747 24731 13753
rect 25130 13744 25136 13756
rect 25188 13784 25194 13796
rect 25685 13787 25743 13793
rect 25685 13784 25697 13787
rect 25188 13756 25697 13784
rect 25188 13744 25194 13756
rect 25685 13753 25697 13756
rect 25731 13784 25743 13787
rect 25961 13787 26019 13793
rect 25961 13784 25973 13787
rect 25731 13756 25973 13784
rect 25731 13753 25743 13756
rect 25685 13747 25743 13753
rect 25961 13753 25973 13756
rect 26007 13753 26019 13787
rect 26068 13784 26096 13824
rect 26329 13821 26341 13824
rect 26375 13821 26387 13855
rect 26436 13852 26464 14028
rect 27157 14025 27169 14059
rect 27203 14056 27215 14059
rect 27982 14056 27988 14068
rect 27203 14028 27988 14056
rect 27203 14025 27215 14028
rect 27157 14019 27215 14025
rect 27982 14016 27988 14028
rect 28040 14016 28046 14068
rect 28074 14016 28080 14068
rect 28132 14056 28138 14068
rect 28132 14028 28177 14056
rect 28132 14016 28138 14028
rect 28258 14016 28264 14068
rect 28316 14056 28322 14068
rect 28997 14059 29055 14065
rect 28997 14056 29009 14059
rect 28316 14028 29009 14056
rect 28316 14016 28322 14028
rect 28997 14025 29009 14028
rect 29043 14025 29055 14059
rect 28997 14019 29055 14025
rect 29825 14059 29883 14065
rect 29825 14025 29837 14059
rect 29871 14056 29883 14059
rect 30374 14056 30380 14068
rect 29871 14028 30380 14056
rect 29871 14025 29883 14028
rect 29825 14019 29883 14025
rect 30374 14016 30380 14028
rect 30432 14016 30438 14068
rect 33042 14016 33048 14068
rect 33100 14056 33106 14068
rect 33597 14059 33655 14065
rect 33597 14056 33609 14059
rect 33100 14028 33609 14056
rect 33100 14016 33106 14028
rect 33597 14025 33609 14028
rect 33643 14056 33655 14059
rect 35710 14056 35716 14068
rect 33643 14028 35716 14056
rect 33643 14025 33655 14028
rect 33597 14019 33655 14025
rect 35710 14016 35716 14028
rect 35768 14016 35774 14068
rect 35989 14059 36047 14065
rect 35989 14025 36001 14059
rect 36035 14056 36047 14059
rect 36078 14056 36084 14068
rect 36035 14028 36084 14056
rect 36035 14025 36047 14028
rect 35989 14019 36047 14025
rect 36078 14016 36084 14028
rect 36136 14016 36142 14068
rect 36354 14056 36360 14068
rect 36315 14028 36360 14056
rect 36354 14016 36360 14028
rect 36412 14016 36418 14068
rect 38194 14016 38200 14068
rect 38252 14056 38258 14068
rect 39301 14059 39359 14065
rect 39301 14056 39313 14059
rect 38252 14028 39313 14056
rect 38252 14016 38258 14028
rect 39301 14025 39313 14028
rect 39347 14025 39359 14059
rect 41693 14059 41751 14065
rect 39301 14019 39359 14025
rect 40236 14028 41276 14056
rect 27430 13948 27436 14000
rect 27488 13988 27494 14000
rect 27525 13991 27583 13997
rect 27525 13988 27537 13991
rect 27488 13960 27537 13988
rect 27488 13948 27494 13960
rect 27525 13957 27537 13960
rect 27571 13988 27583 13991
rect 27893 13991 27951 13997
rect 27893 13988 27905 13991
rect 27571 13960 27905 13988
rect 27571 13957 27583 13960
rect 27525 13951 27583 13957
rect 27893 13957 27905 13960
rect 27939 13988 27951 13991
rect 28810 13988 28816 14000
rect 27939 13960 28816 13988
rect 27939 13957 27951 13960
rect 27893 13951 27951 13957
rect 28810 13948 28816 13960
rect 28868 13948 28874 14000
rect 31021 13991 31079 13997
rect 31021 13957 31033 13991
rect 31067 13988 31079 13991
rect 35342 13988 35348 14000
rect 31067 13960 35348 13988
rect 31067 13957 31079 13960
rect 31021 13951 31079 13957
rect 35342 13948 35348 13960
rect 35400 13948 35406 14000
rect 35434 13948 35440 14000
rect 35492 13988 35498 14000
rect 36633 13991 36691 13997
rect 36633 13988 36645 13991
rect 35492 13960 36645 13988
rect 35492 13948 35498 13960
rect 36633 13957 36645 13960
rect 36679 13957 36691 13991
rect 36633 13951 36691 13957
rect 37918 13948 37924 14000
rect 37976 13988 37982 14000
rect 38286 13988 38292 14000
rect 37976 13960 38292 13988
rect 37976 13948 37982 13960
rect 38286 13948 38292 13960
rect 38344 13948 38350 14000
rect 38749 13991 38807 13997
rect 38749 13957 38761 13991
rect 38795 13988 38807 13991
rect 39117 13991 39175 13997
rect 39117 13988 39129 13991
rect 38795 13960 39129 13988
rect 38795 13957 38807 13960
rect 38749 13951 38807 13957
rect 39117 13957 39129 13960
rect 39163 13988 39175 13991
rect 40236 13988 40264 14028
rect 41248 14000 41276 14028
rect 41693 14025 41705 14059
rect 41739 14056 41751 14059
rect 41782 14056 41788 14068
rect 41739 14028 41788 14056
rect 41739 14025 41751 14028
rect 41693 14019 41751 14025
rect 41782 14016 41788 14028
rect 41840 14016 41846 14068
rect 42058 14016 42064 14068
rect 42116 14056 42122 14068
rect 42518 14056 42524 14068
rect 42116 14028 42524 14056
rect 42116 14016 42122 14028
rect 42518 14016 42524 14028
rect 42576 14016 42582 14068
rect 42613 14059 42671 14065
rect 42613 14025 42625 14059
rect 42659 14056 42671 14059
rect 43162 14056 43168 14068
rect 42659 14028 43168 14056
rect 42659 14025 42671 14028
rect 42613 14019 42671 14025
rect 43162 14016 43168 14028
rect 43220 14016 43226 14068
rect 43257 14059 43315 14065
rect 43257 14025 43269 14059
rect 43303 14056 43315 14059
rect 43530 14056 43536 14068
rect 43303 14028 43536 14056
rect 43303 14025 43315 14028
rect 43257 14019 43315 14025
rect 43530 14016 43536 14028
rect 43588 14016 43594 14068
rect 43990 14056 43996 14068
rect 43951 14028 43996 14056
rect 43990 14016 43996 14028
rect 44048 14016 44054 14068
rect 45830 14056 45836 14068
rect 45791 14028 45836 14056
rect 45830 14016 45836 14028
rect 45888 14016 45894 14068
rect 47486 14056 47492 14068
rect 46584 14028 47492 14056
rect 39163 13960 40264 13988
rect 40328 13960 40632 13988
rect 39163 13957 39175 13960
rect 39117 13951 39175 13957
rect 26789 13923 26847 13929
rect 26789 13889 26801 13923
rect 26835 13920 26847 13923
rect 27338 13920 27344 13932
rect 26835 13892 27344 13920
rect 26835 13889 26847 13892
rect 26789 13883 26847 13889
rect 27338 13880 27344 13892
rect 27396 13880 27402 13932
rect 27985 13923 28043 13929
rect 27985 13889 27997 13923
rect 28031 13920 28043 13923
rect 28166 13920 28172 13932
rect 28031 13892 28172 13920
rect 28031 13889 28043 13892
rect 27985 13883 28043 13889
rect 28166 13880 28172 13892
rect 28224 13920 28230 13932
rect 28721 13923 28779 13929
rect 28721 13920 28733 13923
rect 28224 13892 28733 13920
rect 28224 13880 28230 13892
rect 28721 13889 28733 13892
rect 28767 13920 28779 13923
rect 28902 13920 28908 13932
rect 28767 13892 28908 13920
rect 28767 13889 28779 13892
rect 28721 13883 28779 13889
rect 28902 13880 28908 13892
rect 28960 13880 28966 13932
rect 29822 13920 29828 13932
rect 29012 13892 29828 13920
rect 26436 13824 27476 13852
rect 26329 13815 26387 13821
rect 26234 13784 26240 13796
rect 26068 13756 26240 13784
rect 25961 13747 26019 13753
rect 26234 13744 26240 13756
rect 26292 13744 26298 13796
rect 27448 13784 27476 13824
rect 27522 13812 27528 13864
rect 27580 13852 27586 13864
rect 27617 13855 27675 13861
rect 27617 13852 27629 13855
rect 27580 13824 27629 13852
rect 27580 13812 27586 13824
rect 27617 13821 27629 13824
rect 27663 13821 27675 13855
rect 27617 13815 27675 13821
rect 27764 13855 27822 13861
rect 27764 13821 27776 13855
rect 27810 13852 27822 13855
rect 28534 13852 28540 13864
rect 27810 13824 28540 13852
rect 27810 13821 27822 13824
rect 27764 13815 27822 13821
rect 28534 13812 28540 13824
rect 28592 13812 28598 13864
rect 29012 13852 29040 13892
rect 29822 13880 29828 13892
rect 29880 13880 29886 13932
rect 30190 13880 30196 13932
rect 30248 13920 30254 13932
rect 30469 13923 30527 13929
rect 30469 13920 30481 13923
rect 30248 13892 30481 13920
rect 30248 13880 30254 13892
rect 30469 13889 30481 13892
rect 30515 13920 30527 13923
rect 31481 13923 31539 13929
rect 31481 13920 31493 13923
rect 30515 13892 31493 13920
rect 30515 13889 30527 13892
rect 30469 13883 30527 13889
rect 31481 13889 31493 13892
rect 31527 13889 31539 13923
rect 31481 13883 31539 13889
rect 31938 13880 31944 13932
rect 31996 13920 32002 13932
rect 33229 13923 33287 13929
rect 33229 13920 33241 13923
rect 31996 13892 33241 13920
rect 31996 13880 32002 13892
rect 33229 13889 33241 13892
rect 33275 13920 33287 13923
rect 35621 13923 35679 13929
rect 35621 13920 35633 13923
rect 33275 13892 35633 13920
rect 33275 13889 33287 13892
rect 33229 13883 33287 13889
rect 35621 13889 35633 13892
rect 35667 13889 35679 13923
rect 35621 13883 35679 13889
rect 35710 13880 35716 13932
rect 35768 13920 35774 13932
rect 37458 13920 37464 13932
rect 35768 13892 37464 13920
rect 35768 13880 35774 13892
rect 37458 13880 37464 13892
rect 37516 13880 37522 13932
rect 38013 13923 38071 13929
rect 38013 13889 38025 13923
rect 38059 13920 38071 13923
rect 39209 13923 39267 13929
rect 38059 13892 39160 13920
rect 38059 13889 38071 13892
rect 38013 13883 38071 13889
rect 28644 13824 29040 13852
rect 28644 13784 28672 13824
rect 29730 13812 29736 13864
rect 29788 13852 29794 13864
rect 29917 13855 29975 13861
rect 29917 13852 29929 13855
rect 29788 13824 29929 13852
rect 29788 13812 29794 13824
rect 29917 13821 29929 13824
rect 29963 13821 29975 13855
rect 29917 13815 29975 13821
rect 30009 13855 30067 13861
rect 30009 13821 30021 13855
rect 30055 13821 30067 13855
rect 30009 13815 30067 13821
rect 27448 13756 28672 13784
rect 30024 13784 30052 13815
rect 30098 13812 30104 13864
rect 30156 13852 30162 13864
rect 32217 13855 32275 13861
rect 32217 13852 32229 13855
rect 30156 13824 32229 13852
rect 30156 13812 30162 13824
rect 32217 13821 32229 13824
rect 32263 13821 32275 13855
rect 32217 13815 32275 13821
rect 32769 13855 32827 13861
rect 32769 13821 32781 13855
rect 32815 13821 32827 13855
rect 33042 13852 33048 13864
rect 33003 13824 33048 13852
rect 32769 13815 32827 13821
rect 30745 13787 30803 13793
rect 30745 13784 30757 13787
rect 30024 13756 30757 13784
rect 30745 13753 30757 13756
rect 30791 13784 30803 13787
rect 31021 13787 31079 13793
rect 31021 13784 31033 13787
rect 30791 13756 31033 13784
rect 30791 13753 30803 13756
rect 30745 13747 30803 13753
rect 31021 13753 31033 13756
rect 31067 13753 31079 13787
rect 31202 13784 31208 13796
rect 31163 13756 31208 13784
rect 31021 13747 31079 13753
rect 31202 13744 31208 13756
rect 31260 13744 31266 13796
rect 32122 13784 32128 13796
rect 32083 13756 32128 13784
rect 32122 13744 32128 13756
rect 32180 13784 32186 13796
rect 32784 13784 32812 13815
rect 33042 13812 33048 13824
rect 33100 13812 33106 13864
rect 33134 13812 33140 13864
rect 33192 13852 33198 13864
rect 33870 13852 33876 13864
rect 33192 13824 33876 13852
rect 33192 13812 33198 13824
rect 33870 13812 33876 13824
rect 33928 13812 33934 13864
rect 34146 13812 34152 13864
rect 34204 13852 34210 13864
rect 34333 13855 34391 13861
rect 34204 13824 34284 13852
rect 34204 13812 34210 13824
rect 32180 13756 32812 13784
rect 34256 13784 34284 13824
rect 34333 13821 34345 13855
rect 34379 13852 34391 13855
rect 34379 13824 35204 13852
rect 34379 13821 34391 13824
rect 34333 13815 34391 13821
rect 34609 13787 34667 13793
rect 34609 13784 34621 13787
rect 34256 13756 34621 13784
rect 32180 13744 32186 13756
rect 34609 13753 34621 13756
rect 34655 13753 34667 13787
rect 34882 13784 34888 13796
rect 34843 13756 34888 13784
rect 34609 13747 34667 13753
rect 17402 13716 17408 13728
rect 12268 13688 17408 13716
rect 10652 13676 10658 13688
rect 17402 13676 17408 13688
rect 17460 13676 17466 13728
rect 17862 13716 17868 13728
rect 17823 13688 17868 13716
rect 17862 13676 17868 13688
rect 17920 13676 17926 13728
rect 19518 13676 19524 13728
rect 19576 13716 19582 13728
rect 19705 13719 19763 13725
rect 19705 13716 19717 13719
rect 19576 13688 19717 13716
rect 19576 13676 19582 13688
rect 19705 13685 19717 13688
rect 19751 13685 19763 13719
rect 19705 13679 19763 13685
rect 22738 13676 22744 13728
rect 22796 13716 22802 13728
rect 29822 13716 29828 13728
rect 22796 13688 29828 13716
rect 22796 13676 22802 13688
rect 29822 13676 29828 13688
rect 29880 13676 29886 13728
rect 30006 13676 30012 13728
rect 30064 13716 30070 13728
rect 33502 13716 33508 13728
rect 30064 13688 33508 13716
rect 30064 13676 30070 13688
rect 33502 13676 33508 13688
rect 33560 13716 33566 13728
rect 33962 13716 33968 13728
rect 33560 13688 33968 13716
rect 33560 13676 33566 13688
rect 33962 13676 33968 13688
rect 34020 13676 34026 13728
rect 34624 13716 34652 13747
rect 34882 13744 34888 13756
rect 34940 13744 34946 13796
rect 35176 13725 35204 13824
rect 35342 13812 35348 13864
rect 35400 13852 35406 13864
rect 37277 13855 37335 13861
rect 37277 13852 37289 13855
rect 35400 13824 37289 13852
rect 35400 13812 35406 13824
rect 37277 13821 37289 13824
rect 37323 13852 37335 13855
rect 37553 13855 37611 13861
rect 37553 13852 37565 13855
rect 37323 13824 37565 13852
rect 37323 13821 37335 13824
rect 37277 13815 37335 13821
rect 37553 13821 37565 13824
rect 37599 13852 37611 13855
rect 38102 13852 38108 13864
rect 37599 13824 38108 13852
rect 37599 13821 37611 13824
rect 37553 13815 37611 13821
rect 38102 13812 38108 13824
rect 38160 13812 38166 13864
rect 39022 13861 39028 13864
rect 38988 13855 39028 13861
rect 38988 13821 39000 13855
rect 38988 13815 39028 13821
rect 39022 13812 39028 13815
rect 39080 13812 39086 13864
rect 39132 13852 39160 13892
rect 39209 13889 39221 13923
rect 39255 13920 39267 13923
rect 39298 13920 39304 13932
rect 39255 13892 39304 13920
rect 39255 13889 39267 13892
rect 39209 13883 39267 13889
rect 39298 13880 39304 13892
rect 39356 13880 39362 13932
rect 40034 13920 40040 13932
rect 39995 13892 40040 13920
rect 40034 13880 40040 13892
rect 40092 13880 40098 13932
rect 40328 13852 40356 13960
rect 40494 13920 40500 13932
rect 40455 13892 40500 13920
rect 40494 13880 40500 13892
rect 40552 13880 40558 13932
rect 40604 13920 40632 13960
rect 41230 13948 41236 14000
rect 41288 13988 41294 14000
rect 42245 13991 42303 13997
rect 42245 13988 42257 13991
rect 41288 13960 42257 13988
rect 41288 13948 41294 13960
rect 42245 13957 42257 13960
rect 42291 13988 42303 13991
rect 43806 13988 43812 14000
rect 42291 13960 43812 13988
rect 42291 13957 42303 13960
rect 42245 13951 42303 13957
rect 43806 13948 43812 13960
rect 43864 13988 43870 14000
rect 44913 13991 44971 13997
rect 44913 13988 44925 13991
rect 43864 13960 44925 13988
rect 43864 13948 43870 13960
rect 44913 13957 44925 13960
rect 44959 13957 44971 13991
rect 44913 13951 44971 13957
rect 40604 13892 42472 13920
rect 40586 13852 40592 13864
rect 39132 13824 40356 13852
rect 40547 13824 40592 13852
rect 40586 13812 40592 13824
rect 40644 13812 40650 13864
rect 40678 13812 40684 13864
rect 40736 13852 40742 13864
rect 41049 13855 41107 13861
rect 41049 13852 41061 13855
rect 40736 13824 41061 13852
rect 40736 13812 40742 13824
rect 41049 13821 41061 13824
rect 41095 13821 41107 13855
rect 41966 13852 41972 13864
rect 41927 13824 41972 13852
rect 41049 13815 41107 13821
rect 41966 13812 41972 13824
rect 42024 13812 42030 13864
rect 42150 13861 42156 13864
rect 42116 13855 42156 13861
rect 42116 13821 42128 13855
rect 42116 13815 42156 13821
rect 42150 13812 42156 13815
rect 42208 13812 42214 13864
rect 42308 13855 42366 13861
rect 42308 13821 42320 13855
rect 42354 13821 42366 13855
rect 42444 13852 42472 13892
rect 42518 13880 42524 13932
rect 42576 13920 42582 13932
rect 43073 13923 43131 13929
rect 43073 13920 43085 13923
rect 42576 13892 43085 13920
rect 42576 13880 42582 13892
rect 43073 13889 43085 13892
rect 43119 13920 43131 13923
rect 43119 13892 43852 13920
rect 43119 13889 43131 13892
rect 43073 13883 43131 13889
rect 43530 13852 43536 13864
rect 42444 13824 43536 13852
rect 42308 13815 42366 13821
rect 35250 13744 35256 13796
rect 35308 13784 35314 13796
rect 38838 13784 38844 13796
rect 35308 13756 35353 13784
rect 38799 13756 38844 13784
rect 35308 13744 35314 13756
rect 38838 13744 38844 13756
rect 38896 13744 38902 13796
rect 41414 13744 41420 13796
rect 41472 13784 41478 13796
rect 42323 13784 42351 13815
rect 43530 13812 43536 13824
rect 43588 13812 43594 13864
rect 43622 13812 43628 13864
rect 43680 13861 43686 13864
rect 43680 13855 43738 13861
rect 43680 13821 43692 13855
rect 43726 13821 43738 13855
rect 43824 13852 43852 13892
rect 43898 13880 43904 13932
rect 43956 13920 43962 13932
rect 43956 13892 44001 13920
rect 43956 13880 43962 13892
rect 46584 13861 46612 14028
rect 47486 14016 47492 14028
rect 47544 14016 47550 14068
rect 48314 14056 48320 14068
rect 48275 14028 48320 14056
rect 48314 14016 48320 14028
rect 48372 14016 48378 14068
rect 48958 14016 48964 14068
rect 49016 14056 49022 14068
rect 49053 14059 49111 14065
rect 49053 14056 49065 14059
rect 49016 14028 49065 14056
rect 49016 14016 49022 14028
rect 49053 14025 49065 14028
rect 49099 14025 49111 14059
rect 49053 14019 49111 14025
rect 49142 14016 49148 14068
rect 49200 14056 49206 14068
rect 49881 14059 49939 14065
rect 49881 14056 49893 14059
rect 49200 14028 49893 14056
rect 49200 14016 49206 14028
rect 49881 14025 49893 14028
rect 49927 14056 49939 14059
rect 50065 14059 50123 14065
rect 50065 14056 50077 14059
rect 49927 14028 50077 14056
rect 49927 14025 49939 14028
rect 49881 14019 49939 14025
rect 50065 14025 50077 14028
rect 50111 14056 50123 14059
rect 50893 14059 50951 14065
rect 50111 14028 50292 14056
rect 50111 14025 50123 14028
rect 50065 14019 50123 14025
rect 46842 13948 46848 14000
rect 46900 13988 46906 14000
rect 47765 13991 47823 13997
rect 47765 13988 47777 13991
rect 46900 13960 47777 13988
rect 46900 13948 46906 13960
rect 47765 13957 47777 13960
rect 47811 13988 47823 13991
rect 49789 13991 49847 13997
rect 49789 13988 49801 13991
rect 47811 13960 49801 13988
rect 47811 13957 47823 13960
rect 47765 13951 47823 13957
rect 49789 13957 49801 13960
rect 49835 13957 49847 13991
rect 50264 13988 50292 14028
rect 50893 14025 50905 14059
rect 50939 14056 50951 14059
rect 51077 14059 51135 14065
rect 51077 14056 51089 14059
rect 50939 14028 51089 14056
rect 50939 14025 50951 14028
rect 50893 14019 50951 14025
rect 51077 14025 51089 14028
rect 51123 14025 51135 14059
rect 51077 14019 51135 14025
rect 51442 14016 51448 14068
rect 51500 14056 51506 14068
rect 51905 14059 51963 14065
rect 51905 14056 51917 14059
rect 51500 14028 51917 14056
rect 51500 14016 51506 14028
rect 51905 14025 51917 14028
rect 51951 14025 51963 14059
rect 51905 14019 51963 14025
rect 52270 14016 52276 14068
rect 52328 14056 52334 14068
rect 53009 14059 53067 14065
rect 53009 14056 53021 14059
rect 52328 14028 53021 14056
rect 52328 14016 52334 14028
rect 53009 14025 53021 14028
rect 53055 14025 53067 14059
rect 55674 14056 55680 14068
rect 53009 14019 53067 14025
rect 53300 14028 55680 14056
rect 53300 14000 53328 14028
rect 55674 14016 55680 14028
rect 55732 14016 55738 14068
rect 55766 14016 55772 14068
rect 55824 14056 55830 14068
rect 56137 14059 56195 14065
rect 56137 14056 56149 14059
rect 55824 14028 56149 14056
rect 55824 14016 55830 14028
rect 56137 14025 56149 14028
rect 56183 14025 56195 14059
rect 56137 14019 56195 14025
rect 56410 14016 56416 14068
rect 56468 14056 56474 14068
rect 57057 14059 57115 14065
rect 57057 14056 57069 14059
rect 56468 14028 57069 14056
rect 56468 14016 56474 14028
rect 57057 14025 57069 14028
rect 57103 14025 57115 14059
rect 57057 14019 57115 14025
rect 58713 14059 58771 14065
rect 58713 14025 58725 14059
rect 58759 14056 58771 14059
rect 58894 14056 58900 14068
rect 58759 14028 58900 14056
rect 58759 14025 58771 14028
rect 58713 14019 58771 14025
rect 53282 13988 53288 14000
rect 50264 13960 53288 13988
rect 49789 13951 49847 13957
rect 53282 13948 53288 13960
rect 53340 13948 53346 14000
rect 53742 13948 53748 14000
rect 53800 13988 53806 14000
rect 54297 13991 54355 13997
rect 54297 13988 54309 13991
rect 53800 13960 54309 13988
rect 53800 13948 53806 13960
rect 54297 13957 54309 13960
rect 54343 13957 54355 13991
rect 55122 13988 55128 14000
rect 55083 13960 55128 13988
rect 54297 13951 54355 13957
rect 48222 13929 48228 13932
rect 48188 13923 48228 13929
rect 48188 13889 48200 13923
rect 48188 13883 48228 13889
rect 48222 13880 48228 13883
rect 48280 13880 48286 13932
rect 48406 13920 48412 13932
rect 48367 13892 48412 13920
rect 48406 13880 48412 13892
rect 48464 13880 48470 13932
rect 48501 13923 48559 13929
rect 48501 13889 48513 13923
rect 48547 13889 48559 13923
rect 48501 13883 48559 13889
rect 49605 13923 49663 13929
rect 49605 13889 49617 13923
rect 49651 13920 49663 13923
rect 52454 13920 52460 13932
rect 49651 13892 52460 13920
rect 49651 13889 49663 13892
rect 49605 13883 49663 13889
rect 46569 13855 46627 13861
rect 43824 13824 46244 13852
rect 43680 13815 43738 13821
rect 43680 13812 43686 13815
rect 43257 13787 43315 13793
rect 43257 13784 43269 13787
rect 41472 13756 43269 13784
rect 41472 13744 41478 13756
rect 43257 13753 43269 13756
rect 43303 13784 43315 13787
rect 43898 13784 43904 13796
rect 43303 13756 43904 13784
rect 43303 13753 43315 13756
rect 43257 13747 43315 13753
rect 43898 13744 43904 13756
rect 43956 13784 43962 13796
rect 44545 13787 44603 13793
rect 44545 13784 44557 13787
rect 43956 13756 44557 13784
rect 43956 13744 43962 13756
rect 44545 13753 44557 13756
rect 44591 13753 44603 13787
rect 44545 13747 44603 13753
rect 45646 13744 45652 13796
rect 45704 13784 45710 13796
rect 46106 13784 46112 13796
rect 45704 13756 46112 13784
rect 45704 13744 45710 13756
rect 46106 13744 46112 13756
rect 46164 13744 46170 13796
rect 46216 13784 46244 13824
rect 46569 13821 46581 13855
rect 46615 13821 46627 13855
rect 46750 13852 46756 13864
rect 46711 13824 46756 13852
rect 46569 13815 46627 13821
rect 46750 13812 46756 13824
rect 46808 13812 46814 13864
rect 46842 13812 46848 13864
rect 46900 13852 46906 13864
rect 46937 13855 46995 13861
rect 46937 13852 46949 13855
rect 46900 13824 46949 13852
rect 46900 13812 46906 13824
rect 46937 13821 46949 13824
rect 46983 13821 46995 13855
rect 48516 13852 48544 13883
rect 50246 13852 50252 13864
rect 46937 13815 46995 13821
rect 47044 13824 48544 13852
rect 50207 13824 50252 13852
rect 47044 13784 47072 13824
rect 50246 13812 50252 13824
rect 50304 13812 50310 13864
rect 50356 13861 50384 13892
rect 52454 13880 52460 13892
rect 52512 13880 52518 13932
rect 54312 13920 54340 13951
rect 55122 13948 55128 13960
rect 55180 13948 55186 14000
rect 55582 13988 55588 14000
rect 55232 13960 55588 13988
rect 55232 13920 55260 13960
rect 55582 13948 55588 13960
rect 55640 13948 55646 14000
rect 55784 13920 55812 14016
rect 57609 13991 57667 13997
rect 57609 13957 57621 13991
rect 57655 13988 57667 13991
rect 58434 13988 58440 14000
rect 57655 13960 58440 13988
rect 57655 13957 57667 13960
rect 57609 13951 57667 13957
rect 58434 13948 58440 13960
rect 58492 13948 58498 14000
rect 58728 13920 58756 14019
rect 58894 14016 58900 14028
rect 58952 14016 58958 14068
rect 54312 13892 55260 13920
rect 55324 13892 55812 13920
rect 57808 13892 58756 13920
rect 50341 13855 50399 13861
rect 50341 13821 50353 13855
rect 50387 13821 50399 13855
rect 50341 13815 50399 13821
rect 50522 13812 50528 13864
rect 50580 13852 50586 13864
rect 50801 13855 50859 13861
rect 50801 13852 50813 13855
rect 50580 13824 50813 13852
rect 50580 13812 50586 13824
rect 50801 13821 50813 13824
rect 50847 13852 50859 13855
rect 50893 13855 50951 13861
rect 50893 13852 50905 13855
rect 50847 13824 50905 13852
rect 50847 13821 50859 13824
rect 50801 13815 50859 13821
rect 50893 13821 50905 13824
rect 50939 13821 50951 13855
rect 50893 13815 50951 13821
rect 51721 13855 51779 13861
rect 51721 13821 51733 13855
rect 51767 13852 51779 13855
rect 52086 13852 52092 13864
rect 51767 13824 52092 13852
rect 51767 13821 51779 13824
rect 51721 13815 51779 13821
rect 52086 13812 52092 13824
rect 52144 13812 52150 13864
rect 52178 13812 52184 13864
rect 52236 13852 52242 13864
rect 52638 13852 52644 13864
rect 52236 13824 52644 13852
rect 52236 13812 52242 13824
rect 52638 13812 52644 13824
rect 52696 13812 52702 13864
rect 52730 13812 52736 13864
rect 52788 13852 52794 13864
rect 52825 13855 52883 13861
rect 52825 13852 52837 13855
rect 52788 13824 52837 13852
rect 52788 13812 52794 13824
rect 52825 13821 52837 13824
rect 52871 13852 52883 13855
rect 53377 13855 53435 13861
rect 53377 13852 53389 13855
rect 52871 13824 53389 13852
rect 52871 13821 52883 13824
rect 52825 13815 52883 13821
rect 53377 13821 53389 13824
rect 53423 13821 53435 13855
rect 53377 13815 53435 13821
rect 54757 13855 54815 13861
rect 54757 13821 54769 13855
rect 54803 13852 54815 13855
rect 55214 13852 55220 13864
rect 54803 13824 55220 13852
rect 54803 13821 54815 13824
rect 54757 13815 54815 13821
rect 55214 13812 55220 13824
rect 55272 13812 55278 13864
rect 55324 13861 55352 13892
rect 55309 13855 55367 13861
rect 55309 13821 55321 13855
rect 55355 13821 55367 13855
rect 55490 13852 55496 13864
rect 55451 13824 55496 13852
rect 55309 13815 55367 13821
rect 55490 13812 55496 13824
rect 55548 13812 55554 13864
rect 55677 13855 55735 13861
rect 55677 13821 55689 13855
rect 55723 13852 55735 13855
rect 55858 13852 55864 13864
rect 55723 13824 55864 13852
rect 55723 13821 55735 13824
rect 55677 13815 55735 13821
rect 55858 13812 55864 13824
rect 55916 13852 55922 13864
rect 56505 13855 56563 13861
rect 56505 13852 56517 13855
rect 55916 13824 56517 13852
rect 55916 13812 55922 13824
rect 56505 13821 56517 13824
rect 56551 13821 56563 13855
rect 56505 13815 56563 13821
rect 56962 13812 56968 13864
rect 57020 13852 57026 13864
rect 57808 13861 57836 13892
rect 57793 13855 57851 13861
rect 57020 13824 57744 13852
rect 57020 13812 57026 13824
rect 46216 13756 47072 13784
rect 47302 13744 47308 13796
rect 47360 13784 47366 13796
rect 48041 13787 48099 13793
rect 48041 13784 48053 13787
rect 47360 13756 48053 13784
rect 47360 13744 47366 13756
rect 48041 13753 48053 13756
rect 48087 13753 48099 13787
rect 52362 13784 52368 13796
rect 48041 13747 48099 13753
rect 48148 13756 52368 13784
rect 35069 13719 35127 13725
rect 35069 13716 35081 13719
rect 34624 13688 35081 13716
rect 35069 13685 35081 13688
rect 35115 13685 35127 13719
rect 35069 13679 35127 13685
rect 35161 13719 35219 13725
rect 35161 13685 35173 13719
rect 35207 13716 35219 13719
rect 35342 13716 35348 13728
rect 35207 13688 35348 13716
rect 35207 13685 35219 13688
rect 35161 13679 35219 13685
rect 35342 13676 35348 13688
rect 35400 13676 35406 13728
rect 35526 13676 35532 13728
rect 35584 13716 35590 13728
rect 39206 13716 39212 13728
rect 35584 13688 39212 13716
rect 35584 13676 35590 13688
rect 39206 13676 39212 13688
rect 39264 13676 39270 13728
rect 39298 13676 39304 13728
rect 39356 13716 39362 13728
rect 43349 13719 43407 13725
rect 43349 13716 43361 13719
rect 39356 13688 43361 13716
rect 39356 13676 39362 13688
rect 43349 13685 43361 13688
rect 43395 13716 43407 13719
rect 43438 13716 43444 13728
rect 43395 13688 43444 13716
rect 43395 13685 43407 13688
rect 43349 13679 43407 13685
rect 43438 13676 43444 13688
rect 43496 13716 43502 13728
rect 45094 13716 45100 13728
rect 43496 13688 45100 13716
rect 43496 13676 43502 13688
rect 45094 13676 45100 13688
rect 45152 13676 45158 13728
rect 45554 13716 45560 13728
rect 45515 13688 45560 13716
rect 45554 13676 45560 13688
rect 45612 13676 45618 13728
rect 46198 13676 46204 13728
rect 46256 13716 46262 13728
rect 48148 13716 48176 13756
rect 52362 13744 52368 13756
rect 52420 13744 52426 13796
rect 57716 13784 57744 13824
rect 57793 13821 57805 13855
rect 57839 13821 57851 13855
rect 57977 13855 58035 13861
rect 57977 13852 57989 13855
rect 57793 13815 57851 13821
rect 57900 13824 57989 13852
rect 57900 13796 57928 13824
rect 57977 13821 57989 13824
rect 58023 13821 58035 13855
rect 58158 13852 58164 13864
rect 58119 13824 58164 13852
rect 57977 13815 58035 13821
rect 58158 13812 58164 13824
rect 58216 13852 58222 13864
rect 58989 13855 59047 13861
rect 58989 13852 59001 13855
rect 58216 13824 59001 13852
rect 58216 13812 58222 13824
rect 58989 13821 59001 13824
rect 59035 13821 59047 13855
rect 58989 13815 59047 13821
rect 57882 13784 57888 13796
rect 57716 13756 57888 13784
rect 57882 13744 57888 13756
rect 57940 13744 57946 13796
rect 46256 13688 48176 13716
rect 49789 13719 49847 13725
rect 46256 13676 46262 13688
rect 49789 13685 49801 13719
rect 49835 13716 49847 13719
rect 50982 13716 50988 13728
rect 49835 13688 50988 13716
rect 49835 13685 49847 13688
rect 49789 13679 49847 13685
rect 50982 13676 50988 13688
rect 51040 13676 51046 13728
rect 51074 13676 51080 13728
rect 51132 13716 51138 13728
rect 51445 13719 51503 13725
rect 51445 13716 51457 13719
rect 51132 13688 51457 13716
rect 51132 13676 51138 13688
rect 51445 13685 51457 13688
rect 51491 13685 51503 13719
rect 51445 13679 51503 13685
rect 52086 13676 52092 13728
rect 52144 13716 52150 13728
rect 52273 13719 52331 13725
rect 52273 13716 52285 13719
rect 52144 13688 52285 13716
rect 52144 13676 52150 13688
rect 52273 13685 52285 13688
rect 52319 13685 52331 13719
rect 52273 13679 52331 13685
rect 1104 13626 63480 13648
rect 1104 13574 21774 13626
rect 21826 13574 21838 13626
rect 21890 13574 21902 13626
rect 21954 13574 21966 13626
rect 22018 13574 42566 13626
rect 42618 13574 42630 13626
rect 42682 13574 42694 13626
rect 42746 13574 42758 13626
rect 42810 13574 63480 13626
rect 1104 13552 63480 13574
rect 4522 13472 4528 13524
rect 4580 13512 4586 13524
rect 5442 13512 5448 13524
rect 4580 13484 5448 13512
rect 4580 13472 4586 13484
rect 5442 13472 5448 13484
rect 5500 13512 5506 13524
rect 6089 13515 6147 13521
rect 6089 13512 6101 13515
rect 5500 13484 6101 13512
rect 5500 13472 5506 13484
rect 6089 13481 6101 13484
rect 6135 13481 6147 13515
rect 7561 13515 7619 13521
rect 7561 13512 7573 13515
rect 6089 13475 6147 13481
rect 6840 13484 7573 13512
rect 5534 13404 5540 13456
rect 5592 13444 5598 13456
rect 6273 13447 6331 13453
rect 6273 13444 6285 13447
rect 5592 13416 6285 13444
rect 5592 13404 5598 13416
rect 6273 13413 6285 13416
rect 6319 13413 6331 13447
rect 6273 13407 6331 13413
rect 4982 13376 4988 13388
rect 4943 13348 4988 13376
rect 4982 13336 4988 13348
rect 5040 13376 5046 13388
rect 6840 13376 6868 13484
rect 7561 13481 7573 13484
rect 7607 13481 7619 13515
rect 7742 13512 7748 13524
rect 7703 13484 7748 13512
rect 7561 13475 7619 13481
rect 7742 13472 7748 13484
rect 7800 13472 7806 13524
rect 8110 13472 8116 13524
rect 8168 13512 8174 13524
rect 8941 13515 8999 13521
rect 8941 13512 8953 13515
rect 8168 13484 8953 13512
rect 8168 13472 8174 13484
rect 8941 13481 8953 13484
rect 8987 13512 8999 13515
rect 13722 13512 13728 13524
rect 8987 13484 13728 13512
rect 8987 13481 8999 13484
rect 8941 13475 8999 13481
rect 13722 13472 13728 13484
rect 13780 13472 13786 13524
rect 14734 13512 14740 13524
rect 13832 13484 14740 13512
rect 10594 13444 10600 13456
rect 7300 13416 9904 13444
rect 10555 13416 10600 13444
rect 7300 13388 7328 13416
rect 5040 13348 6868 13376
rect 6917 13379 6975 13385
rect 5040 13336 5046 13348
rect 6917 13345 6929 13379
rect 6963 13376 6975 13379
rect 7006 13376 7012 13388
rect 6963 13348 7012 13376
rect 6963 13345 6975 13348
rect 6917 13339 6975 13345
rect 7006 13336 7012 13348
rect 7064 13376 7070 13388
rect 7064 13348 7236 13376
rect 7064 13336 7070 13348
rect 4893 13311 4951 13317
rect 4893 13308 4905 13311
rect 4724 13280 4905 13308
rect 4724 13184 4752 13280
rect 4893 13277 4905 13280
rect 4939 13277 4951 13311
rect 4893 13271 4951 13277
rect 5445 13311 5503 13317
rect 5445 13277 5457 13311
rect 5491 13308 5503 13311
rect 6546 13308 6552 13320
rect 5491 13280 6552 13308
rect 5491 13277 5503 13280
rect 5445 13271 5503 13277
rect 6546 13268 6552 13280
rect 6604 13268 6610 13320
rect 6825 13311 6883 13317
rect 6825 13277 6837 13311
rect 6871 13308 6883 13311
rect 6871 13280 6960 13308
rect 6871 13277 6883 13280
rect 6825 13271 6883 13277
rect 6932 13252 6960 13280
rect 6914 13200 6920 13252
rect 6972 13200 6978 13252
rect 7208 13240 7236 13348
rect 7282 13336 7288 13388
rect 7340 13376 7346 13388
rect 7561 13379 7619 13385
rect 7340 13348 7433 13376
rect 7340 13336 7346 13348
rect 7561 13345 7573 13379
rect 7607 13376 7619 13379
rect 9766 13376 9772 13388
rect 7607 13348 9772 13376
rect 7607 13345 7619 13348
rect 7561 13339 7619 13345
rect 9766 13336 9772 13348
rect 9824 13336 9830 13388
rect 9876 13376 9904 13416
rect 10594 13404 10600 13416
rect 10652 13404 10658 13456
rect 11698 13444 11704 13456
rect 11659 13416 11704 13444
rect 11698 13404 11704 13416
rect 11756 13404 11762 13456
rect 13832 13444 13860 13484
rect 14734 13472 14740 13484
rect 14792 13472 14798 13524
rect 14918 13472 14924 13524
rect 14976 13512 14982 13524
rect 15657 13515 15715 13521
rect 15657 13512 15669 13515
rect 14976 13484 15669 13512
rect 14976 13472 14982 13484
rect 15657 13481 15669 13484
rect 15703 13481 15715 13515
rect 15657 13475 15715 13481
rect 16393 13515 16451 13521
rect 16393 13481 16405 13515
rect 16439 13512 16451 13515
rect 16850 13512 16856 13524
rect 16439 13484 16856 13512
rect 16439 13481 16451 13484
rect 16393 13475 16451 13481
rect 16850 13472 16856 13484
rect 16908 13472 16914 13524
rect 18230 13472 18236 13524
rect 18288 13512 18294 13524
rect 20990 13512 20996 13524
rect 18288 13484 20996 13512
rect 18288 13472 18294 13484
rect 20990 13472 20996 13484
rect 21048 13472 21054 13524
rect 25038 13472 25044 13524
rect 25096 13512 25102 13524
rect 25133 13515 25191 13521
rect 25133 13512 25145 13515
rect 25096 13484 25145 13512
rect 25096 13472 25102 13484
rect 25133 13481 25145 13484
rect 25179 13481 25191 13515
rect 25133 13475 25191 13481
rect 25501 13515 25559 13521
rect 25501 13481 25513 13515
rect 25547 13512 25559 13515
rect 25547 13484 26188 13512
rect 25547 13481 25559 13484
rect 25501 13475 25559 13481
rect 11808 13416 13860 13444
rect 11808 13376 11836 13416
rect 13906 13404 13912 13456
rect 13964 13444 13970 13456
rect 16761 13447 16819 13453
rect 16761 13444 16773 13447
rect 13964 13416 16773 13444
rect 13964 13404 13970 13416
rect 16761 13413 16773 13416
rect 16807 13413 16819 13447
rect 17586 13444 17592 13456
rect 16761 13407 16819 13413
rect 17236 13416 17592 13444
rect 9876 13348 11836 13376
rect 11974 13336 11980 13388
rect 12032 13376 12038 13388
rect 12161 13379 12219 13385
rect 12161 13376 12173 13379
rect 12032 13348 12173 13376
rect 12032 13336 12038 13348
rect 12161 13345 12173 13348
rect 12207 13345 12219 13379
rect 12161 13339 12219 13345
rect 12529 13379 12587 13385
rect 12529 13345 12541 13379
rect 12575 13345 12587 13379
rect 12529 13339 12587 13345
rect 7374 13308 7380 13320
rect 7335 13280 7380 13308
rect 7374 13268 7380 13280
rect 7432 13268 7438 13320
rect 7653 13311 7711 13317
rect 7653 13277 7665 13311
rect 7699 13308 7711 13311
rect 9582 13308 9588 13320
rect 7699 13280 9588 13308
rect 7699 13277 7711 13280
rect 7653 13271 7711 13277
rect 9582 13268 9588 13280
rect 9640 13268 9646 13320
rect 9674 13268 9680 13320
rect 9732 13317 9738 13320
rect 9732 13311 9745 13317
rect 9733 13308 9745 13311
rect 10229 13311 10287 13317
rect 9733 13280 10180 13308
rect 9733 13277 9745 13280
rect 9732 13271 9745 13277
rect 9732 13268 9738 13271
rect 10152 13240 10180 13280
rect 10229 13277 10241 13311
rect 10275 13308 10287 13311
rect 10686 13308 10692 13320
rect 10275 13280 10692 13308
rect 10275 13277 10287 13280
rect 10229 13271 10287 13277
rect 10686 13268 10692 13280
rect 10744 13268 10750 13320
rect 12544 13308 12572 13339
rect 12618 13336 12624 13388
rect 12676 13376 12682 13388
rect 13078 13376 13084 13388
rect 12676 13348 12721 13376
rect 13039 13348 13084 13376
rect 12676 13336 12682 13348
rect 13078 13336 13084 13348
rect 13136 13336 13142 13388
rect 13817 13379 13875 13385
rect 13817 13345 13829 13379
rect 13863 13345 13875 13379
rect 13817 13339 13875 13345
rect 14001 13379 14059 13385
rect 14001 13345 14013 13379
rect 14047 13376 14059 13379
rect 14090 13376 14096 13388
rect 14047 13348 14096 13376
rect 14047 13345 14059 13348
rect 14001 13339 14059 13345
rect 13096 13308 13124 13336
rect 12544 13280 13124 13308
rect 13832 13308 13860 13339
rect 14090 13336 14096 13348
rect 14148 13376 14154 13388
rect 14642 13376 14648 13388
rect 14148 13348 14648 13376
rect 14148 13336 14154 13348
rect 14642 13336 14648 13348
rect 14700 13336 14706 13388
rect 14737 13379 14795 13385
rect 14737 13345 14749 13379
rect 14783 13376 14795 13379
rect 14918 13376 14924 13388
rect 14783 13348 14924 13376
rect 14783 13345 14795 13348
rect 14737 13339 14795 13345
rect 14918 13336 14924 13348
rect 14976 13336 14982 13388
rect 15289 13379 15347 13385
rect 15289 13345 15301 13379
rect 15335 13376 15347 13379
rect 16022 13376 16028 13388
rect 15335 13348 16028 13376
rect 15335 13345 15347 13348
rect 15289 13339 15347 13345
rect 16022 13336 16028 13348
rect 16080 13336 16086 13388
rect 16574 13376 16580 13388
rect 16487 13348 16580 13376
rect 16574 13336 16580 13348
rect 16632 13376 16638 13388
rect 17236 13376 17264 13416
rect 17586 13404 17592 13416
rect 17644 13404 17650 13456
rect 17862 13404 17868 13456
rect 17920 13404 17926 13456
rect 19610 13404 19616 13456
rect 19668 13444 19674 13456
rect 20806 13444 20812 13456
rect 19668 13416 20812 13444
rect 19668 13404 19674 13416
rect 20806 13404 20812 13416
rect 20864 13404 20870 13456
rect 22094 13444 22100 13456
rect 21100 13416 22100 13444
rect 17402 13376 17408 13388
rect 16632 13348 17264 13376
rect 17363 13348 17408 13376
rect 16632 13336 16638 13348
rect 17402 13336 17408 13348
rect 17460 13336 17466 13388
rect 17678 13336 17684 13388
rect 17736 13376 17742 13388
rect 17773 13379 17831 13385
rect 17773 13376 17785 13379
rect 17736 13348 17785 13376
rect 17736 13336 17742 13348
rect 17773 13345 17785 13348
rect 17819 13345 17831 13379
rect 17880 13376 17908 13404
rect 21100 13385 21128 13416
rect 22094 13404 22100 13416
rect 22152 13404 22158 13456
rect 17957 13379 18015 13385
rect 17957 13376 17969 13379
rect 17880 13348 17969 13376
rect 17773 13339 17831 13345
rect 17957 13345 17969 13348
rect 18003 13376 18015 13379
rect 18969 13379 19027 13385
rect 18969 13376 18981 13379
rect 18003 13348 18981 13376
rect 18003 13345 18015 13348
rect 17957 13339 18015 13345
rect 18969 13345 18981 13348
rect 19015 13345 19027 13379
rect 18969 13339 19027 13345
rect 19797 13379 19855 13385
rect 19797 13345 19809 13379
rect 19843 13376 19855 13379
rect 21085 13379 21143 13385
rect 21085 13376 21097 13379
rect 19843 13348 21097 13376
rect 19843 13345 19855 13348
rect 19797 13339 19855 13345
rect 21085 13345 21097 13348
rect 21131 13345 21143 13379
rect 21085 13339 21143 13345
rect 21542 13336 21548 13388
rect 21600 13376 21606 13388
rect 21818 13376 21824 13388
rect 21600 13348 21824 13376
rect 21600 13336 21606 13348
rect 21818 13336 21824 13348
rect 21876 13336 21882 13388
rect 21910 13336 21916 13388
rect 21968 13376 21974 13388
rect 22005 13379 22063 13385
rect 22005 13376 22017 13379
rect 21968 13348 22017 13376
rect 21968 13336 21974 13348
rect 22005 13345 22017 13348
rect 22051 13345 22063 13379
rect 22005 13339 22063 13345
rect 22189 13379 22247 13385
rect 22189 13345 22201 13379
rect 22235 13376 22247 13379
rect 23109 13379 23167 13385
rect 23109 13376 23121 13379
rect 22235 13348 23121 13376
rect 22235 13345 22247 13348
rect 22189 13339 22247 13345
rect 23109 13345 23121 13348
rect 23155 13376 23167 13379
rect 23382 13376 23388 13388
rect 23155 13348 23388 13376
rect 23155 13345 23167 13348
rect 23109 13339 23167 13345
rect 23382 13336 23388 13348
rect 23440 13376 23446 13388
rect 24029 13379 24087 13385
rect 24029 13376 24041 13379
rect 23440 13348 24041 13376
rect 23440 13336 23446 13348
rect 24029 13345 24041 13348
rect 24075 13376 24087 13379
rect 25056 13376 25084 13472
rect 25516 13444 25544 13475
rect 24075 13348 25084 13376
rect 25240 13416 25544 13444
rect 24075 13345 24087 13348
rect 24029 13339 24087 13345
rect 14182 13308 14188 13320
rect 13832 13280 14188 13308
rect 12636 13252 12664 13280
rect 14182 13268 14188 13280
rect 14240 13268 14246 13320
rect 14369 13311 14427 13317
rect 14369 13277 14381 13311
rect 14415 13308 14427 13311
rect 14826 13308 14832 13320
rect 14415 13280 14832 13308
rect 14415 13277 14427 13280
rect 14369 13271 14427 13277
rect 14826 13268 14832 13280
rect 14884 13308 14890 13320
rect 15013 13311 15071 13317
rect 15013 13308 15025 13311
rect 14884 13280 15025 13308
rect 14884 13268 14890 13280
rect 15013 13277 15025 13280
rect 15059 13277 15071 13311
rect 15013 13271 15071 13277
rect 15562 13268 15568 13320
rect 15620 13308 15626 13320
rect 15933 13311 15991 13317
rect 15933 13308 15945 13311
rect 15620 13280 15945 13308
rect 15620 13268 15626 13280
rect 15933 13277 15945 13280
rect 15979 13308 15991 13311
rect 17310 13308 17316 13320
rect 15979 13280 17172 13308
rect 17271 13280 17316 13308
rect 15979 13277 15991 13280
rect 15933 13271 15991 13277
rect 10502 13240 10508 13252
rect 7208 13212 7788 13240
rect 2406 13172 2412 13184
rect 2367 13144 2412 13172
rect 2406 13132 2412 13144
rect 2464 13132 2470 13184
rect 3878 13172 3884 13184
rect 3839 13144 3884 13172
rect 3878 13132 3884 13144
rect 3936 13132 3942 13184
rect 4706 13172 4712 13184
rect 4667 13144 4712 13172
rect 4706 13132 4712 13144
rect 4764 13132 4770 13184
rect 5166 13132 5172 13184
rect 5224 13172 5230 13184
rect 5813 13175 5871 13181
rect 5813 13172 5825 13175
rect 5224 13144 5825 13172
rect 5224 13132 5230 13144
rect 5813 13141 5825 13144
rect 5859 13172 5871 13175
rect 7653 13175 7711 13181
rect 7653 13172 7665 13175
rect 5859 13144 7665 13172
rect 5859 13141 5871 13144
rect 5813 13135 5871 13141
rect 7653 13141 7665 13144
rect 7699 13141 7711 13175
rect 7760 13172 7788 13212
rect 7944 13212 9536 13240
rect 10152 13212 10508 13240
rect 7944 13172 7972 13212
rect 7760 13144 7972 13172
rect 7653 13135 7711 13141
rect 8018 13132 8024 13184
rect 8076 13172 8082 13184
rect 8113 13175 8171 13181
rect 8113 13172 8125 13175
rect 8076 13144 8125 13172
rect 8076 13132 8082 13144
rect 8113 13141 8125 13144
rect 8159 13141 8171 13175
rect 8478 13172 8484 13184
rect 8439 13144 8484 13172
rect 8113 13135 8171 13141
rect 8478 13132 8484 13144
rect 8536 13132 8542 13184
rect 9398 13172 9404 13184
rect 9359 13144 9404 13172
rect 9398 13132 9404 13144
rect 9456 13132 9462 13184
rect 9508 13172 9536 13212
rect 10502 13200 10508 13212
rect 10560 13240 10566 13252
rect 11425 13243 11483 13249
rect 11425 13240 11437 13243
rect 10560 13212 11437 13240
rect 10560 13200 10566 13212
rect 11425 13209 11437 13212
rect 11471 13209 11483 13243
rect 11425 13203 11483 13209
rect 10226 13172 10232 13184
rect 9508 13144 10232 13172
rect 10226 13132 10232 13144
rect 10284 13132 10290 13184
rect 11146 13172 11152 13184
rect 11107 13144 11152 13172
rect 11146 13132 11152 13144
rect 11204 13132 11210 13184
rect 11440 13172 11468 13203
rect 12618 13200 12624 13252
rect 12676 13200 12682 13252
rect 12710 13200 12716 13252
rect 12768 13240 12774 13252
rect 13449 13243 13507 13249
rect 13449 13240 13461 13243
rect 12768 13212 13461 13240
rect 12768 13200 12774 13212
rect 13449 13209 13461 13212
rect 13495 13240 13507 13243
rect 15473 13243 15531 13249
rect 15473 13240 15485 13243
rect 13495 13212 15485 13240
rect 13495 13209 13507 13212
rect 13449 13203 13507 13209
rect 15473 13209 15485 13212
rect 15519 13209 15531 13243
rect 17144 13240 17172 13280
rect 17310 13268 17316 13280
rect 17368 13268 17374 13320
rect 19518 13308 19524 13320
rect 19479 13280 19524 13308
rect 19518 13268 19524 13280
rect 19576 13268 19582 13320
rect 19981 13311 20039 13317
rect 19981 13277 19993 13311
rect 20027 13308 20039 13311
rect 20625 13311 20683 13317
rect 20625 13308 20637 13311
rect 20027 13280 20637 13308
rect 20027 13277 20039 13280
rect 19981 13271 20039 13277
rect 20625 13277 20637 13280
rect 20671 13308 20683 13311
rect 21269 13311 21327 13317
rect 21269 13308 21281 13311
rect 20671 13280 21281 13308
rect 20671 13277 20683 13280
rect 20625 13271 20683 13277
rect 21269 13277 21281 13280
rect 21315 13277 21327 13311
rect 23201 13311 23259 13317
rect 23201 13308 23213 13311
rect 21269 13271 21327 13277
rect 21376 13280 23213 13308
rect 20349 13243 20407 13249
rect 17144 13212 18736 13240
rect 15473 13203 15531 13209
rect 12066 13172 12072 13184
rect 11440 13144 12072 13172
rect 12066 13132 12072 13144
rect 12124 13132 12130 13184
rect 15657 13175 15715 13181
rect 15657 13141 15669 13175
rect 15703 13172 15715 13175
rect 16301 13175 16359 13181
rect 16301 13172 16313 13175
rect 15703 13144 16313 13172
rect 15703 13141 15715 13144
rect 15657 13135 15715 13141
rect 16301 13141 16313 13144
rect 16347 13172 16359 13175
rect 17034 13172 17040 13184
rect 16347 13144 17040 13172
rect 16347 13141 16359 13144
rect 16301 13135 16359 13141
rect 17034 13132 17040 13144
rect 17092 13132 17098 13184
rect 18598 13172 18604 13184
rect 18559 13144 18604 13172
rect 18598 13132 18604 13144
rect 18656 13132 18662 13184
rect 18708 13172 18736 13212
rect 20349 13209 20361 13243
rect 20395 13240 20407 13243
rect 20898 13240 20904 13252
rect 20395 13212 20904 13240
rect 20395 13209 20407 13212
rect 20349 13203 20407 13209
rect 20898 13200 20904 13212
rect 20956 13200 20962 13252
rect 21376 13240 21404 13280
rect 23201 13277 23213 13280
rect 23247 13277 23259 13311
rect 23201 13271 23259 13277
rect 23290 13268 23296 13320
rect 23348 13308 23354 13320
rect 23753 13311 23811 13317
rect 23753 13308 23765 13311
rect 23348 13280 23765 13308
rect 23348 13268 23354 13280
rect 23753 13277 23765 13280
rect 23799 13277 23811 13311
rect 24210 13308 24216 13320
rect 24123 13280 24216 13308
rect 23753 13271 23811 13277
rect 24210 13268 24216 13280
rect 24268 13308 24274 13320
rect 25240 13308 25268 13416
rect 25317 13379 25375 13385
rect 25317 13345 25329 13379
rect 25363 13376 25375 13379
rect 26050 13376 26056 13388
rect 25363 13348 26056 13376
rect 25363 13345 25375 13348
rect 25317 13339 25375 13345
rect 26050 13336 26056 13348
rect 26108 13336 26114 13388
rect 26160 13376 26188 13484
rect 26234 13472 26240 13524
rect 26292 13512 26298 13524
rect 26292 13484 27200 13512
rect 26292 13472 26298 13484
rect 27172 13453 27200 13484
rect 27706 13472 27712 13524
rect 27764 13512 27770 13524
rect 27801 13515 27859 13521
rect 27801 13512 27813 13515
rect 27764 13484 27813 13512
rect 27764 13472 27770 13484
rect 27801 13481 27813 13484
rect 27847 13481 27859 13515
rect 28166 13512 28172 13524
rect 28127 13484 28172 13512
rect 27801 13475 27859 13481
rect 28166 13472 28172 13484
rect 28224 13472 28230 13524
rect 28534 13512 28540 13524
rect 28495 13484 28540 13512
rect 28534 13472 28540 13484
rect 28592 13472 28598 13524
rect 28810 13472 28816 13524
rect 28868 13512 28874 13524
rect 28905 13515 28963 13521
rect 28905 13512 28917 13515
rect 28868 13484 28917 13512
rect 28868 13472 28874 13484
rect 28905 13481 28917 13484
rect 28951 13481 28963 13515
rect 29270 13512 29276 13524
rect 29231 13484 29276 13512
rect 28905 13475 28963 13481
rect 27157 13447 27215 13453
rect 27157 13413 27169 13447
rect 27203 13413 27215 13447
rect 28920 13444 28948 13475
rect 29270 13472 29276 13484
rect 29328 13472 29334 13524
rect 29730 13512 29736 13524
rect 29691 13484 29736 13512
rect 29730 13472 29736 13484
rect 29788 13472 29794 13524
rect 30466 13512 30472 13524
rect 30427 13484 30472 13512
rect 30466 13472 30472 13484
rect 30524 13472 30530 13524
rect 31113 13515 31171 13521
rect 31113 13481 31125 13515
rect 31159 13512 31171 13515
rect 31202 13512 31208 13524
rect 31159 13484 31208 13512
rect 31159 13481 31171 13484
rect 31113 13475 31171 13481
rect 31202 13472 31208 13484
rect 31260 13472 31266 13524
rect 35526 13512 35532 13524
rect 31312 13484 35532 13512
rect 30484 13444 30512 13472
rect 31312 13444 31340 13484
rect 35526 13472 35532 13484
rect 35584 13472 35590 13524
rect 36633 13515 36691 13521
rect 36633 13481 36645 13515
rect 36679 13512 36691 13515
rect 41046 13512 41052 13524
rect 36679 13484 41052 13512
rect 36679 13481 36691 13484
rect 36633 13475 36691 13481
rect 41046 13472 41052 13484
rect 41104 13472 41110 13524
rect 41138 13472 41144 13524
rect 41196 13512 41202 13524
rect 41601 13515 41659 13521
rect 41601 13512 41613 13515
rect 41196 13484 41613 13512
rect 41196 13472 41202 13484
rect 41601 13481 41613 13484
rect 41647 13481 41659 13515
rect 41601 13475 41659 13481
rect 41690 13472 41696 13524
rect 41748 13512 41754 13524
rect 42337 13515 42395 13521
rect 42337 13512 42349 13515
rect 41748 13484 42349 13512
rect 41748 13472 41754 13484
rect 42337 13481 42349 13484
rect 42383 13481 42395 13515
rect 42337 13475 42395 13481
rect 42797 13515 42855 13521
rect 42797 13481 42809 13515
rect 42843 13512 42855 13515
rect 42978 13512 42984 13524
rect 42843 13484 42984 13512
rect 42843 13481 42855 13484
rect 42797 13475 42855 13481
rect 42978 13472 42984 13484
rect 43036 13472 43042 13524
rect 43530 13472 43536 13524
rect 43588 13512 43594 13524
rect 44177 13515 44235 13521
rect 44177 13512 44189 13515
rect 43588 13484 44189 13512
rect 43588 13472 43594 13484
rect 44177 13481 44189 13484
rect 44223 13481 44235 13515
rect 44177 13475 44235 13481
rect 46661 13515 46719 13521
rect 46661 13481 46673 13515
rect 46707 13512 46719 13515
rect 47857 13515 47915 13521
rect 46707 13484 47624 13512
rect 46707 13481 46719 13484
rect 46661 13475 46719 13481
rect 27157 13407 27215 13413
rect 27264 13416 28856 13444
rect 28920 13416 30512 13444
rect 30852 13416 31340 13444
rect 31573 13447 31631 13453
rect 27264 13376 27292 13416
rect 28718 13376 28724 13388
rect 26160 13348 27292 13376
rect 28679 13348 28724 13376
rect 28718 13336 28724 13348
rect 28776 13336 28782 13388
rect 28828 13376 28856 13416
rect 29822 13376 29828 13388
rect 28828 13348 29684 13376
rect 29783 13348 29828 13376
rect 24268 13280 25268 13308
rect 27525 13311 27583 13317
rect 24268 13268 24274 13280
rect 27525 13277 27537 13311
rect 27571 13308 27583 13311
rect 28166 13308 28172 13320
rect 27571 13280 28172 13308
rect 27571 13277 27583 13280
rect 27525 13271 27583 13277
rect 28166 13268 28172 13280
rect 28224 13268 28230 13320
rect 28736 13308 28764 13336
rect 29086 13308 29092 13320
rect 28736 13280 29092 13308
rect 29086 13268 29092 13280
rect 29144 13268 29150 13320
rect 29656 13308 29684 13348
rect 29822 13336 29828 13348
rect 29880 13336 29886 13388
rect 30852 13308 30880 13416
rect 31573 13413 31585 13447
rect 31619 13444 31631 13447
rect 31619 13416 32444 13444
rect 31619 13413 31631 13416
rect 31573 13407 31631 13413
rect 30926 13336 30932 13388
rect 30984 13376 30990 13388
rect 32416 13385 32444 13416
rect 33042 13404 33048 13456
rect 33100 13444 33106 13456
rect 33689 13447 33747 13453
rect 33689 13444 33701 13447
rect 33100 13416 33701 13444
rect 33100 13404 33106 13416
rect 33689 13413 33701 13416
rect 33735 13413 33747 13447
rect 35434 13444 35440 13456
rect 33689 13407 33747 13413
rect 34440 13416 35440 13444
rect 31941 13379 31999 13385
rect 30984 13348 31029 13376
rect 30984 13336 30990 13348
rect 31941 13345 31953 13379
rect 31987 13376 31999 13379
rect 32309 13379 32367 13385
rect 32309 13376 32321 13379
rect 31987 13348 32321 13376
rect 31987 13345 31999 13348
rect 31941 13339 31999 13345
rect 32309 13345 32321 13348
rect 32355 13345 32367 13379
rect 32309 13339 32367 13345
rect 32401 13379 32459 13385
rect 32401 13345 32413 13379
rect 32447 13376 32459 13379
rect 32490 13376 32496 13388
rect 32447 13348 32496 13376
rect 32447 13345 32459 13348
rect 32401 13339 32459 13345
rect 29656 13280 30880 13308
rect 31662 13268 31668 13320
rect 31720 13308 31726 13320
rect 32324 13308 32352 13339
rect 32490 13336 32496 13348
rect 32548 13336 32554 13388
rect 33502 13376 33508 13388
rect 33463 13348 33508 13376
rect 33502 13336 33508 13348
rect 33560 13336 33566 13388
rect 34238 13376 34244 13388
rect 33612 13348 34244 13376
rect 32674 13308 32680 13320
rect 31720 13280 32260 13308
rect 32324 13280 32680 13308
rect 31720 13268 31726 13280
rect 21008 13212 21404 13240
rect 21637 13243 21695 13249
rect 21008 13172 21036 13212
rect 21637 13209 21649 13243
rect 21683 13240 21695 13243
rect 22554 13240 22560 13252
rect 21683 13212 22560 13240
rect 21683 13209 21695 13212
rect 21637 13203 21695 13209
rect 22554 13200 22560 13212
rect 22612 13200 22618 13252
rect 22741 13243 22799 13249
rect 22741 13209 22753 13243
rect 22787 13240 22799 13243
rect 22830 13240 22836 13252
rect 22787 13212 22836 13240
rect 22787 13209 22799 13212
rect 22741 13203 22799 13209
rect 22830 13200 22836 13212
rect 22888 13200 22894 13252
rect 23658 13200 23664 13252
rect 23716 13240 23722 13252
rect 25869 13243 25927 13249
rect 25869 13240 25881 13243
rect 23716 13212 25881 13240
rect 23716 13200 23722 13212
rect 25869 13209 25881 13212
rect 25915 13240 25927 13243
rect 27154 13240 27160 13252
rect 25915 13212 27160 13240
rect 25915 13209 25927 13212
rect 25869 13203 25927 13209
rect 27154 13200 27160 13212
rect 27212 13200 27218 13252
rect 27322 13243 27380 13249
rect 27322 13209 27334 13243
rect 27368 13240 27380 13243
rect 29178 13240 29184 13252
rect 27368 13212 29184 13240
rect 27368 13209 27380 13212
rect 27322 13203 27380 13209
rect 29178 13200 29184 13212
rect 29236 13200 29242 13252
rect 32232 13240 32260 13280
rect 32674 13268 32680 13280
rect 32732 13268 32738 13320
rect 33226 13268 33232 13320
rect 33284 13308 33290 13320
rect 33612 13308 33640 13348
rect 34238 13336 34244 13348
rect 34296 13336 34302 13388
rect 34440 13385 34468 13416
rect 35434 13404 35440 13416
rect 35492 13404 35498 13456
rect 37553 13447 37611 13453
rect 37553 13413 37565 13447
rect 37599 13444 37611 13447
rect 38194 13444 38200 13456
rect 37599 13416 38200 13444
rect 37599 13413 37611 13416
rect 37553 13407 37611 13413
rect 38194 13404 38200 13416
rect 38252 13404 38258 13456
rect 39025 13447 39083 13453
rect 39025 13413 39037 13447
rect 39071 13444 39083 13447
rect 39298 13444 39304 13456
rect 39071 13416 39304 13444
rect 39071 13413 39083 13416
rect 39025 13407 39083 13413
rect 39298 13404 39304 13416
rect 39356 13404 39362 13456
rect 39482 13404 39488 13456
rect 39540 13444 39546 13456
rect 39577 13447 39635 13453
rect 39577 13444 39589 13447
rect 39540 13416 39589 13444
rect 39540 13404 39546 13416
rect 39577 13413 39589 13416
rect 39623 13413 39635 13447
rect 40126 13444 40132 13456
rect 40087 13416 40132 13444
rect 39577 13407 39635 13413
rect 40126 13404 40132 13416
rect 40184 13404 40190 13456
rect 42245 13447 42303 13453
rect 42245 13444 42257 13447
rect 40236 13416 42257 13444
rect 34425 13379 34483 13385
rect 34425 13345 34437 13379
rect 34471 13345 34483 13379
rect 34606 13376 34612 13388
rect 34567 13348 34612 13376
rect 34425 13339 34483 13345
rect 34606 13336 34612 13348
rect 34664 13336 34670 13388
rect 35894 13336 35900 13388
rect 35952 13376 35958 13388
rect 35989 13379 36047 13385
rect 35989 13376 36001 13379
rect 35952 13348 36001 13376
rect 35952 13336 35958 13348
rect 35989 13345 36001 13348
rect 36035 13345 36047 13379
rect 38102 13376 38108 13388
rect 38063 13348 38108 13376
rect 35989 13339 36047 13345
rect 38102 13336 38108 13348
rect 38160 13336 38166 13388
rect 38286 13336 38292 13388
rect 38344 13376 38350 13388
rect 39390 13376 39396 13388
rect 38344 13348 39396 13376
rect 38344 13336 38350 13348
rect 39390 13336 39396 13348
rect 39448 13336 39454 13388
rect 39666 13336 39672 13388
rect 39724 13376 39730 13388
rect 39724 13348 39769 13376
rect 39724 13336 39730 13348
rect 33284 13280 33640 13308
rect 33284 13268 33290 13280
rect 34146 13268 34152 13320
rect 34204 13308 34210 13320
rect 34793 13311 34851 13317
rect 34793 13308 34805 13311
rect 34204 13280 34805 13308
rect 34204 13268 34210 13280
rect 34793 13277 34805 13280
rect 34839 13277 34851 13311
rect 34793 13271 34851 13277
rect 35069 13311 35127 13317
rect 35069 13277 35081 13311
rect 35115 13277 35127 13311
rect 36354 13308 36360 13320
rect 36315 13280 36360 13308
rect 35069 13271 35127 13277
rect 33042 13240 33048 13252
rect 32232 13212 33048 13240
rect 33042 13200 33048 13212
rect 33100 13200 33106 13252
rect 34330 13200 34336 13252
rect 34388 13240 34394 13252
rect 35084 13240 35112 13271
rect 36354 13268 36360 13280
rect 36412 13308 36418 13320
rect 36814 13308 36820 13320
rect 36412 13280 36820 13308
rect 36412 13268 36418 13280
rect 36814 13268 36820 13280
rect 36872 13308 36878 13320
rect 37001 13311 37059 13317
rect 37001 13308 37013 13311
rect 36872 13280 37013 13308
rect 36872 13268 36878 13280
rect 37001 13277 37013 13280
rect 37047 13277 37059 13311
rect 37001 13271 37059 13277
rect 37918 13268 37924 13320
rect 37976 13308 37982 13320
rect 38013 13311 38071 13317
rect 38013 13308 38025 13311
rect 37976 13280 38025 13308
rect 37976 13268 37982 13280
rect 38013 13277 38025 13280
rect 38059 13277 38071 13311
rect 38013 13271 38071 13277
rect 38565 13311 38623 13317
rect 38565 13277 38577 13311
rect 38611 13308 38623 13311
rect 39942 13308 39948 13320
rect 38611 13280 39948 13308
rect 38611 13277 38623 13280
rect 38565 13271 38623 13277
rect 39942 13268 39948 13280
rect 40000 13268 40006 13320
rect 35437 13243 35495 13249
rect 35437 13240 35449 13243
rect 34388 13212 35449 13240
rect 34388 13200 34394 13212
rect 35437 13209 35449 13212
rect 35483 13209 35495 13243
rect 35437 13203 35495 13209
rect 36630 13200 36636 13252
rect 36688 13240 36694 13252
rect 40236 13240 40264 13416
rect 42245 13413 42257 13416
rect 42291 13413 42303 13447
rect 45005 13447 45063 13453
rect 45005 13444 45017 13447
rect 42245 13407 42303 13413
rect 42904 13416 45017 13444
rect 40402 13376 40408 13388
rect 40363 13348 40408 13376
rect 40402 13336 40408 13348
rect 40460 13336 40466 13388
rect 40678 13336 40684 13388
rect 40736 13376 40742 13388
rect 40957 13379 41015 13385
rect 40957 13376 40969 13379
rect 40736 13348 40969 13376
rect 40736 13336 40742 13348
rect 40957 13345 40969 13348
rect 41003 13345 41015 13379
rect 40957 13339 41015 13345
rect 41046 13336 41052 13388
rect 41104 13376 41110 13388
rect 42904 13376 42932 13416
rect 45005 13413 45017 13416
rect 45051 13413 45063 13447
rect 45005 13407 45063 13413
rect 45373 13447 45431 13453
rect 45373 13413 45385 13447
rect 45419 13444 45431 13447
rect 45646 13444 45652 13456
rect 45419 13416 45652 13444
rect 45419 13413 45431 13416
rect 45373 13407 45431 13413
rect 41104 13348 42932 13376
rect 42981 13379 43039 13385
rect 41104 13336 41110 13348
rect 42981 13345 42993 13379
rect 43027 13376 43039 13379
rect 43073 13379 43131 13385
rect 43073 13376 43085 13379
rect 43027 13348 43085 13376
rect 43027 13345 43039 13348
rect 42981 13339 43039 13345
rect 43073 13345 43085 13348
rect 43119 13345 43131 13379
rect 43346 13376 43352 13388
rect 43307 13348 43352 13376
rect 43073 13339 43131 13345
rect 43346 13336 43352 13348
rect 43404 13336 43410 13388
rect 43441 13379 43499 13385
rect 43441 13345 43453 13379
rect 43487 13376 43499 13379
rect 43530 13376 43536 13388
rect 43487 13348 43536 13376
rect 43487 13345 43499 13348
rect 43441 13339 43499 13345
rect 43530 13336 43536 13348
rect 43588 13336 43594 13388
rect 43901 13379 43959 13385
rect 43901 13345 43913 13379
rect 43947 13376 43959 13379
rect 43993 13379 44051 13385
rect 43993 13376 44005 13379
rect 43947 13348 44005 13376
rect 43947 13345 43959 13348
rect 43901 13339 43959 13345
rect 43993 13345 44005 13348
rect 44039 13345 44051 13379
rect 44542 13376 44548 13388
rect 44503 13348 44548 13376
rect 43993 13339 44051 13345
rect 44542 13336 44548 13348
rect 44600 13336 44606 13388
rect 45020 13376 45048 13407
rect 45646 13404 45652 13416
rect 45704 13404 45710 13456
rect 45830 13404 45836 13456
rect 45888 13444 45894 13456
rect 45925 13447 45983 13453
rect 45925 13444 45937 13447
rect 45888 13416 45937 13444
rect 45888 13404 45894 13416
rect 45925 13413 45937 13416
rect 45971 13413 45983 13447
rect 45925 13407 45983 13413
rect 46293 13447 46351 13453
rect 46293 13413 46305 13447
rect 46339 13444 46351 13447
rect 47302 13444 47308 13456
rect 46339 13416 47308 13444
rect 46339 13413 46351 13416
rect 46293 13407 46351 13413
rect 47302 13404 47308 13416
rect 47360 13404 47366 13456
rect 47596 13444 47624 13484
rect 47857 13481 47869 13515
rect 47903 13512 47915 13515
rect 48314 13512 48320 13524
rect 47903 13484 48320 13512
rect 47903 13481 47915 13484
rect 47857 13475 47915 13481
rect 48314 13472 48320 13484
rect 48372 13472 48378 13524
rect 48501 13515 48559 13521
rect 48501 13481 48513 13515
rect 48547 13512 48559 13515
rect 49605 13515 49663 13521
rect 48547 13484 49188 13512
rect 48547 13481 48559 13484
rect 48501 13475 48559 13481
rect 48222 13444 48228 13456
rect 47596 13416 48228 13444
rect 48222 13404 48228 13416
rect 48280 13404 48286 13456
rect 49160 13444 49188 13484
rect 49605 13481 49617 13515
rect 49651 13512 49663 13515
rect 49786 13512 49792 13524
rect 49651 13484 49792 13512
rect 49651 13481 49663 13484
rect 49605 13475 49663 13481
rect 49786 13472 49792 13484
rect 49844 13472 49850 13524
rect 50246 13512 50252 13524
rect 50207 13484 50252 13512
rect 50246 13472 50252 13484
rect 50304 13472 50310 13524
rect 50982 13472 50988 13524
rect 51040 13512 51046 13524
rect 54757 13515 54815 13521
rect 54757 13512 54769 13515
rect 51040 13484 54769 13512
rect 51040 13472 51046 13484
rect 54757 13481 54769 13484
rect 54803 13481 54815 13515
rect 54757 13475 54815 13481
rect 55122 13472 55128 13524
rect 55180 13512 55186 13524
rect 55493 13515 55551 13521
rect 55493 13512 55505 13515
rect 55180 13484 55505 13512
rect 55180 13472 55186 13484
rect 55493 13481 55505 13484
rect 55539 13481 55551 13515
rect 57146 13512 57152 13524
rect 57107 13484 57152 13512
rect 55493 13475 55551 13481
rect 57146 13472 57152 13484
rect 57204 13472 57210 13524
rect 53745 13447 53803 13453
rect 53745 13444 53757 13447
rect 49160 13416 53757 13444
rect 53745 13413 53757 13416
rect 53791 13413 53803 13447
rect 53745 13407 53803 13413
rect 56778 13404 56784 13456
rect 56836 13444 56842 13456
rect 57701 13447 57759 13453
rect 57701 13444 57713 13447
rect 56836 13416 57713 13444
rect 56836 13404 56842 13416
rect 57701 13413 57713 13416
rect 57747 13444 57759 13447
rect 57790 13444 57796 13456
rect 57747 13416 57796 13444
rect 57747 13413 57759 13416
rect 57701 13407 57759 13413
rect 57790 13404 57796 13416
rect 57848 13444 57854 13456
rect 58069 13447 58127 13453
rect 58069 13444 58081 13447
rect 57848 13416 58081 13444
rect 57848 13404 57854 13416
rect 58069 13413 58081 13416
rect 58115 13413 58127 13447
rect 58434 13444 58440 13456
rect 58395 13416 58440 13444
rect 58069 13407 58127 13413
rect 58434 13404 58440 13416
rect 58492 13404 58498 13456
rect 45465 13379 45523 13385
rect 45465 13376 45477 13379
rect 45020 13348 45477 13376
rect 45465 13345 45477 13348
rect 45511 13345 45523 13379
rect 46842 13376 46848 13388
rect 46803 13348 46848 13376
rect 45465 13339 45523 13345
rect 46842 13336 46848 13348
rect 46900 13336 46906 13388
rect 46934 13336 46940 13388
rect 46992 13376 46998 13388
rect 48317 13379 48375 13385
rect 48317 13376 48329 13379
rect 46992 13348 48329 13376
rect 46992 13336 46998 13348
rect 48317 13345 48329 13348
rect 48363 13376 48375 13379
rect 48501 13379 48559 13385
rect 48501 13376 48513 13379
rect 48363 13348 48513 13376
rect 48363 13345 48375 13348
rect 48317 13339 48375 13345
rect 48501 13345 48513 13348
rect 48547 13345 48559 13379
rect 48958 13376 48964 13388
rect 48919 13348 48964 13376
rect 48501 13339 48559 13345
rect 48958 13336 48964 13348
rect 49016 13336 49022 13388
rect 51074 13336 51080 13388
rect 51132 13376 51138 13388
rect 51353 13379 51411 13385
rect 51132 13348 51177 13376
rect 51132 13336 51138 13348
rect 51353 13345 51365 13379
rect 51399 13376 51411 13379
rect 52362 13376 52368 13388
rect 51399 13348 52040 13376
rect 52323 13348 52368 13376
rect 51399 13345 51411 13348
rect 51353 13339 51411 13345
rect 40865 13311 40923 13317
rect 40865 13277 40877 13311
rect 40911 13308 40923 13311
rect 41325 13311 41383 13317
rect 40911 13280 41276 13308
rect 40911 13277 40923 13280
rect 40865 13271 40923 13277
rect 41138 13249 41144 13252
rect 36688 13212 40264 13240
rect 41122 13243 41144 13249
rect 36688 13200 36694 13212
rect 41122 13209 41134 13243
rect 41122 13203 41144 13209
rect 41138 13200 41144 13203
rect 41196 13200 41202 13252
rect 41248 13240 41276 13280
rect 41325 13277 41337 13311
rect 41371 13308 41383 13311
rect 41414 13308 41420 13320
rect 41371 13280 41420 13308
rect 41371 13277 41383 13280
rect 41325 13271 41383 13277
rect 41414 13268 41420 13280
rect 41472 13268 41478 13320
rect 41966 13268 41972 13320
rect 42024 13268 42030 13320
rect 42245 13311 42303 13317
rect 42245 13277 42257 13311
rect 42291 13308 42303 13311
rect 46198 13308 46204 13320
rect 42291 13280 46204 13308
rect 42291 13277 42303 13280
rect 42245 13271 42303 13277
rect 46198 13268 46204 13280
rect 46256 13268 46262 13320
rect 46566 13268 46572 13320
rect 46624 13308 46630 13320
rect 46753 13311 46811 13317
rect 46753 13308 46765 13311
rect 46624 13280 46765 13308
rect 46624 13268 46630 13280
rect 46753 13277 46765 13280
rect 46799 13277 46811 13311
rect 46753 13271 46811 13277
rect 47026 13268 47032 13320
rect 47084 13308 47090 13320
rect 47084 13280 48360 13308
rect 47084 13268 47090 13280
rect 41984 13240 42012 13268
rect 43993 13243 44051 13249
rect 43993 13240 44005 13243
rect 41248 13212 44005 13240
rect 43993 13209 44005 13212
rect 44039 13209 44051 13243
rect 48332 13240 48360 13280
rect 48406 13268 48412 13320
rect 48464 13308 48470 13320
rect 48682 13308 48688 13320
rect 48464 13280 48688 13308
rect 48464 13268 48470 13280
rect 48682 13268 48688 13280
rect 48740 13308 48746 13320
rect 49329 13311 49387 13317
rect 49329 13308 49341 13311
rect 48740 13280 49341 13308
rect 48740 13268 48746 13280
rect 49329 13277 49341 13280
rect 49375 13277 49387 13311
rect 49329 13271 49387 13277
rect 49418 13268 49424 13320
rect 49476 13308 49482 13320
rect 50525 13311 50583 13317
rect 50525 13308 50537 13311
rect 49476 13280 50537 13308
rect 49476 13268 49482 13280
rect 50525 13277 50537 13280
rect 50571 13277 50583 13311
rect 50525 13271 50583 13277
rect 51537 13311 51595 13317
rect 51537 13277 51549 13311
rect 51583 13308 51595 13311
rect 51583 13280 51764 13308
rect 51583 13277 51595 13280
rect 51537 13271 51595 13277
rect 51736 13240 51764 13280
rect 48332 13212 51764 13240
rect 52012 13240 52040 13348
rect 52362 13336 52368 13348
rect 52420 13336 52426 13388
rect 54573 13379 54631 13385
rect 54573 13345 54585 13379
rect 54619 13345 54631 13379
rect 54573 13339 54631 13345
rect 52086 13268 52092 13320
rect 52144 13308 52150 13320
rect 54588 13308 54616 13339
rect 55674 13336 55680 13388
rect 55732 13376 55738 13388
rect 58250 13376 58256 13388
rect 55732 13348 58256 13376
rect 55732 13336 55738 13348
rect 58250 13336 58256 13348
rect 58308 13336 58314 13388
rect 58529 13379 58587 13385
rect 58529 13345 58541 13379
rect 58575 13376 58587 13379
rect 59170 13376 59176 13388
rect 58575 13348 59176 13376
rect 58575 13345 58587 13348
rect 58529 13339 58587 13345
rect 59170 13336 59176 13348
rect 59228 13336 59234 13388
rect 55125 13311 55183 13317
rect 55125 13308 55137 13311
rect 52144 13280 55137 13308
rect 52144 13268 52150 13280
rect 55125 13277 55137 13280
rect 55171 13277 55183 13311
rect 55125 13271 55183 13277
rect 55582 13268 55588 13320
rect 55640 13308 55646 13320
rect 55769 13311 55827 13317
rect 55769 13308 55781 13311
rect 55640 13280 55781 13308
rect 55640 13268 55646 13280
rect 55769 13277 55781 13280
rect 55815 13277 55827 13311
rect 56042 13308 56048 13320
rect 56003 13280 56048 13308
rect 55769 13271 55827 13277
rect 56042 13268 56048 13280
rect 56100 13268 56106 13320
rect 53466 13240 53472 13252
rect 52012 13212 53052 13240
rect 53379 13212 53472 13240
rect 43993 13203 44051 13209
rect 51736 13184 51764 13212
rect 18708 13144 21036 13172
rect 21269 13175 21327 13181
rect 21269 13141 21281 13175
rect 21315 13172 21327 13175
rect 24210 13172 24216 13184
rect 21315 13144 24216 13172
rect 21315 13141 21327 13144
rect 21269 13135 21327 13141
rect 24210 13132 24216 13144
rect 24268 13132 24274 13184
rect 24854 13172 24860 13184
rect 24815 13144 24860 13172
rect 24854 13132 24860 13144
rect 24912 13132 24918 13184
rect 26326 13132 26332 13184
rect 26384 13172 26390 13184
rect 26697 13175 26755 13181
rect 26697 13172 26709 13175
rect 26384 13144 26709 13172
rect 26384 13132 26390 13144
rect 26697 13141 26709 13144
rect 26743 13141 26755 13175
rect 27430 13172 27436 13184
rect 27391 13144 27436 13172
rect 26697 13135 26755 13141
rect 27430 13132 27436 13144
rect 27488 13132 27494 13184
rect 28258 13132 28264 13184
rect 28316 13172 28322 13184
rect 29730 13172 29736 13184
rect 28316 13144 29736 13172
rect 28316 13132 28322 13144
rect 29730 13132 29736 13144
rect 29788 13132 29794 13184
rect 30006 13172 30012 13184
rect 29967 13144 30012 13172
rect 30006 13132 30012 13144
rect 30064 13132 30070 13184
rect 32030 13132 32036 13184
rect 32088 13172 32094 13184
rect 32125 13175 32183 13181
rect 32125 13172 32137 13175
rect 32088 13144 32137 13172
rect 32088 13132 32094 13144
rect 32125 13141 32137 13144
rect 32171 13141 32183 13175
rect 32582 13172 32588 13184
rect 32543 13144 32588 13172
rect 32125 13135 32183 13141
rect 32582 13132 32588 13144
rect 32640 13132 32646 13184
rect 33229 13175 33287 13181
rect 33229 13141 33241 13175
rect 33275 13172 33287 13175
rect 33410 13172 33416 13184
rect 33275 13144 33416 13172
rect 33275 13141 33287 13144
rect 33229 13135 33287 13141
rect 33410 13132 33416 13144
rect 33468 13132 33474 13184
rect 34054 13132 34060 13184
rect 34112 13172 34118 13184
rect 34882 13172 34888 13184
rect 34112 13144 34888 13172
rect 34112 13132 34118 13144
rect 34882 13132 34888 13144
rect 34940 13132 34946 13184
rect 34974 13132 34980 13184
rect 35032 13172 35038 13184
rect 35250 13172 35256 13184
rect 35032 13144 35256 13172
rect 35032 13132 35038 13144
rect 35250 13132 35256 13144
rect 35308 13172 35314 13184
rect 36170 13181 36176 13184
rect 35805 13175 35863 13181
rect 35805 13172 35817 13175
rect 35308 13144 35817 13172
rect 35308 13132 35314 13144
rect 35805 13141 35817 13144
rect 35851 13141 35863 13175
rect 35805 13135 35863 13141
rect 36154 13175 36176 13181
rect 36154 13141 36166 13175
rect 36154 13135 36176 13141
rect 36170 13132 36176 13135
rect 36228 13132 36234 13184
rect 36265 13175 36323 13181
rect 36265 13141 36277 13175
rect 36311 13172 36323 13175
rect 36446 13172 36452 13184
rect 36311 13144 36452 13172
rect 36311 13141 36323 13144
rect 36265 13135 36323 13141
rect 36446 13132 36452 13144
rect 36504 13132 36510 13184
rect 36814 13132 36820 13184
rect 36872 13172 36878 13184
rect 39025 13175 39083 13181
rect 39025 13172 39037 13175
rect 36872 13144 39037 13172
rect 36872 13132 36878 13144
rect 39025 13141 39037 13144
rect 39071 13141 39083 13175
rect 39206 13172 39212 13184
rect 39119 13144 39212 13172
rect 39025 13135 39083 13141
rect 39206 13132 39212 13144
rect 39264 13172 39270 13184
rect 40586 13172 40592 13184
rect 39264 13144 40592 13172
rect 39264 13132 39270 13144
rect 40586 13132 40592 13144
rect 40644 13132 40650 13184
rect 41230 13172 41236 13184
rect 41191 13144 41236 13172
rect 41230 13132 41236 13144
rect 41288 13172 41294 13184
rect 41782 13172 41788 13184
rect 41288 13144 41788 13172
rect 41288 13132 41294 13144
rect 41782 13132 41788 13144
rect 41840 13132 41846 13184
rect 41966 13172 41972 13184
rect 41927 13144 41972 13172
rect 41966 13132 41972 13144
rect 42024 13132 42030 13184
rect 43070 13172 43076 13184
rect 42983 13144 43076 13172
rect 43070 13132 43076 13144
rect 43128 13172 43134 13184
rect 43714 13172 43720 13184
rect 43128 13144 43720 13172
rect 43128 13132 43134 13144
rect 43714 13132 43720 13144
rect 43772 13132 43778 13184
rect 45186 13172 45192 13184
rect 45147 13144 45192 13172
rect 45186 13132 45192 13144
rect 45244 13132 45250 13184
rect 47210 13132 47216 13184
rect 47268 13172 47274 13184
rect 47581 13175 47639 13181
rect 47581 13172 47593 13175
rect 47268 13144 47593 13172
rect 47268 13132 47274 13144
rect 47581 13141 47593 13144
rect 47627 13172 47639 13175
rect 47857 13175 47915 13181
rect 47857 13172 47869 13175
rect 47627 13144 47869 13172
rect 47627 13141 47639 13144
rect 47581 13135 47639 13141
rect 47857 13141 47869 13144
rect 47903 13141 47915 13175
rect 48038 13172 48044 13184
rect 47999 13144 48044 13172
rect 47857 13135 47915 13141
rect 48038 13132 48044 13144
rect 48096 13132 48102 13184
rect 48130 13132 48136 13184
rect 48188 13172 48194 13184
rect 48682 13172 48688 13184
rect 48188 13144 48233 13172
rect 48643 13144 48688 13172
rect 48188 13132 48194 13144
rect 48682 13132 48688 13144
rect 48740 13132 48746 13184
rect 48774 13132 48780 13184
rect 48832 13172 48838 13184
rect 49099 13175 49157 13181
rect 49099 13172 49111 13175
rect 48832 13144 49111 13172
rect 48832 13132 48838 13144
rect 49099 13141 49111 13144
rect 49145 13141 49157 13175
rect 49234 13172 49240 13184
rect 49195 13144 49240 13172
rect 49099 13135 49157 13141
rect 49234 13132 49240 13144
rect 49292 13132 49298 13184
rect 51718 13132 51724 13184
rect 51776 13172 51782 13184
rect 51813 13175 51871 13181
rect 51813 13172 51825 13175
rect 51776 13144 51825 13172
rect 51776 13132 51782 13144
rect 51813 13141 51825 13144
rect 51859 13141 51871 13175
rect 51813 13135 51871 13141
rect 51902 13132 51908 13184
rect 51960 13172 51966 13184
rect 52181 13175 52239 13181
rect 52181 13172 52193 13175
rect 51960 13144 52193 13172
rect 51960 13132 51966 13144
rect 52181 13141 52193 13144
rect 52227 13141 52239 13175
rect 52546 13172 52552 13184
rect 52507 13144 52552 13172
rect 52181 13135 52239 13141
rect 52546 13132 52552 13144
rect 52604 13132 52610 13184
rect 53024 13181 53052 13212
rect 53466 13200 53472 13212
rect 53524 13240 53530 13252
rect 54202 13240 54208 13252
rect 53524 13212 54208 13240
rect 53524 13200 53530 13212
rect 54202 13200 54208 13212
rect 54260 13200 54266 13252
rect 57330 13240 57336 13252
rect 56704 13212 57336 13240
rect 53009 13175 53067 13181
rect 53009 13141 53021 13175
rect 53055 13172 53067 13175
rect 56704 13172 56732 13212
rect 57330 13200 57336 13212
rect 57388 13200 57394 13252
rect 58710 13172 58716 13184
rect 53055 13144 56732 13172
rect 58671 13144 58716 13172
rect 53055 13141 53067 13144
rect 53009 13135 53067 13141
rect 58710 13132 58716 13144
rect 58768 13132 58774 13184
rect 59262 13172 59268 13184
rect 59223 13144 59268 13172
rect 59262 13132 59268 13144
rect 59320 13132 59326 13184
rect 1104 13082 63480 13104
rect 1104 13030 11378 13082
rect 11430 13030 11442 13082
rect 11494 13030 11506 13082
rect 11558 13030 11570 13082
rect 11622 13030 32170 13082
rect 32222 13030 32234 13082
rect 32286 13030 32298 13082
rect 32350 13030 32362 13082
rect 32414 13030 52962 13082
rect 53014 13030 53026 13082
rect 53078 13030 53090 13082
rect 53142 13030 53154 13082
rect 53206 13030 63480 13082
rect 1104 13008 63480 13030
rect 3145 12971 3203 12977
rect 3145 12968 3157 12971
rect 2608 12940 3157 12968
rect 2406 12764 2412 12776
rect 2367 12736 2412 12764
rect 2406 12724 2412 12736
rect 2464 12724 2470 12776
rect 2608 12773 2636 12940
rect 3145 12937 3157 12940
rect 3191 12937 3203 12971
rect 3145 12931 3203 12937
rect 4065 12971 4123 12977
rect 4065 12937 4077 12971
rect 4111 12968 4123 12971
rect 8478 12968 8484 12980
rect 4111 12940 8484 12968
rect 4111 12937 4123 12940
rect 4065 12931 4123 12937
rect 2976 12872 7972 12900
rect 2976 12841 3004 12872
rect 2961 12835 3019 12841
rect 2961 12801 2973 12835
rect 3007 12801 3019 12835
rect 3878 12832 3884 12844
rect 3791 12804 3884 12832
rect 2961 12795 3019 12801
rect 3804 12773 3832 12804
rect 3878 12792 3884 12804
rect 3936 12832 3942 12844
rect 5718 12832 5724 12844
rect 3936 12804 5724 12832
rect 3936 12792 3942 12804
rect 5718 12792 5724 12804
rect 5776 12792 5782 12844
rect 6641 12835 6699 12841
rect 6641 12801 6653 12835
rect 6687 12832 6699 12835
rect 7374 12832 7380 12844
rect 6687 12804 7380 12832
rect 6687 12801 6699 12804
rect 6641 12795 6699 12801
rect 7374 12792 7380 12804
rect 7432 12832 7438 12844
rect 7653 12835 7711 12841
rect 7653 12832 7665 12835
rect 7432 12804 7665 12832
rect 7432 12792 7438 12804
rect 7653 12801 7665 12804
rect 7699 12801 7711 12835
rect 7653 12795 7711 12801
rect 2593 12767 2651 12773
rect 2593 12733 2605 12767
rect 2639 12733 2651 12767
rect 2593 12727 2651 12733
rect 3789 12767 3847 12773
rect 3789 12733 3801 12767
rect 3835 12733 3847 12767
rect 3789 12727 3847 12733
rect 3973 12767 4031 12773
rect 3973 12733 3985 12767
rect 4019 12764 4031 12767
rect 4433 12767 4491 12773
rect 4433 12764 4445 12767
rect 4019 12736 4445 12764
rect 4019 12733 4031 12736
rect 3973 12727 4031 12733
rect 4433 12733 4445 12736
rect 4479 12733 4491 12767
rect 4982 12764 4988 12776
rect 4943 12736 4988 12764
rect 4433 12727 4491 12733
rect 4982 12724 4988 12736
rect 5040 12724 5046 12776
rect 5166 12764 5172 12776
rect 5127 12736 5172 12764
rect 5166 12724 5172 12736
rect 5224 12724 5230 12776
rect 5442 12764 5448 12776
rect 5403 12736 5448 12764
rect 5442 12724 5448 12736
rect 5500 12724 5506 12776
rect 5905 12767 5963 12773
rect 5905 12733 5917 12767
rect 5951 12764 5963 12767
rect 6914 12764 6920 12776
rect 5951 12736 6920 12764
rect 5951 12733 5963 12736
rect 5905 12727 5963 12733
rect 6914 12724 6920 12736
rect 6972 12724 6978 12776
rect 7193 12767 7251 12773
rect 7193 12733 7205 12767
rect 7239 12764 7251 12767
rect 7282 12764 7288 12776
rect 7239 12736 7288 12764
rect 7239 12733 7251 12736
rect 7193 12727 7251 12733
rect 7282 12724 7288 12736
rect 7340 12724 7346 12776
rect 2424 12628 2452 12724
rect 5258 12696 5264 12708
rect 3068 12668 5264 12696
rect 3068 12628 3096 12668
rect 5258 12656 5264 12668
rect 5316 12656 5322 12708
rect 5350 12656 5356 12708
rect 5408 12696 5414 12708
rect 6181 12699 6239 12705
rect 6181 12696 6193 12699
rect 5408 12668 6193 12696
rect 5408 12656 5414 12668
rect 6181 12665 6193 12668
rect 6227 12665 6239 12699
rect 7944 12696 7972 12872
rect 8110 12764 8116 12776
rect 8071 12736 8116 12764
rect 8110 12724 8116 12736
rect 8168 12724 8174 12776
rect 8220 12764 8248 12940
rect 8478 12928 8484 12940
rect 8536 12928 8542 12980
rect 9766 12968 9772 12980
rect 9727 12940 9772 12968
rect 9766 12928 9772 12940
rect 9824 12928 9830 12980
rect 11057 12971 11115 12977
rect 11057 12968 11069 12971
rect 10152 12940 11069 12968
rect 8496 12872 10088 12900
rect 8297 12767 8355 12773
rect 8297 12764 8309 12767
rect 8220 12736 8309 12764
rect 8297 12733 8309 12736
rect 8343 12733 8355 12767
rect 8297 12727 8355 12733
rect 8496 12696 8524 12872
rect 8754 12832 8760 12844
rect 8715 12804 8760 12832
rect 8754 12792 8760 12804
rect 8812 12792 8818 12844
rect 9950 12832 9956 12844
rect 9911 12804 9956 12832
rect 9950 12792 9956 12804
rect 10008 12792 10014 12844
rect 8573 12767 8631 12773
rect 8573 12733 8585 12767
rect 8619 12733 8631 12767
rect 9122 12764 9128 12776
rect 9083 12736 9128 12764
rect 8573 12727 8631 12733
rect 7944 12668 8524 12696
rect 8588 12696 8616 12727
rect 9122 12724 9128 12736
rect 9180 12724 9186 12776
rect 8588 12668 9536 12696
rect 6181 12659 6239 12665
rect 9508 12640 9536 12668
rect 2424 12600 3096 12628
rect 3145 12631 3203 12637
rect 3145 12597 3157 12631
rect 3191 12628 3203 12631
rect 3329 12631 3387 12637
rect 3329 12628 3341 12631
rect 3191 12600 3341 12628
rect 3191 12597 3203 12600
rect 3145 12591 3203 12597
rect 3329 12597 3341 12600
rect 3375 12628 3387 12631
rect 4154 12628 4160 12640
rect 3375 12600 4160 12628
rect 3375 12597 3387 12600
rect 3329 12591 3387 12597
rect 4154 12588 4160 12600
rect 4212 12588 4218 12640
rect 4433 12631 4491 12637
rect 4433 12597 4445 12631
rect 4479 12628 4491 12631
rect 4709 12631 4767 12637
rect 4709 12628 4721 12631
rect 4479 12600 4721 12628
rect 4479 12597 4491 12600
rect 4433 12591 4491 12597
rect 4709 12597 4721 12600
rect 4755 12628 4767 12631
rect 5810 12628 5816 12640
rect 4755 12600 5816 12628
rect 4755 12597 4767 12600
rect 4709 12591 4767 12597
rect 5810 12588 5816 12600
rect 5868 12588 5874 12640
rect 7561 12631 7619 12637
rect 7561 12597 7573 12631
rect 7607 12628 7619 12631
rect 8662 12628 8668 12640
rect 7607 12600 8668 12628
rect 7607 12597 7619 12600
rect 7561 12591 7619 12597
rect 8662 12588 8668 12600
rect 8720 12588 8726 12640
rect 9490 12628 9496 12640
rect 9451 12600 9496 12628
rect 9490 12588 9496 12600
rect 9548 12588 9554 12640
rect 10060 12628 10088 12872
rect 10152 12773 10180 12940
rect 11057 12937 11069 12940
rect 11103 12968 11115 12971
rect 11103 12940 13584 12968
rect 11103 12937 11115 12940
rect 11057 12931 11115 12937
rect 12526 12900 12532 12912
rect 11808 12872 12532 12900
rect 10226 12792 10232 12844
rect 10284 12832 10290 12844
rect 10689 12835 10747 12841
rect 10689 12832 10701 12835
rect 10284 12804 10701 12832
rect 10284 12792 10290 12804
rect 10689 12801 10701 12804
rect 10735 12801 10747 12835
rect 10689 12795 10747 12801
rect 10137 12767 10195 12773
rect 10137 12733 10149 12767
rect 10183 12733 10195 12767
rect 10137 12727 10195 12733
rect 10318 12696 10324 12708
rect 10279 12668 10324 12696
rect 10318 12656 10324 12668
rect 10376 12656 10382 12708
rect 11238 12656 11244 12708
rect 11296 12696 11302 12708
rect 11808 12705 11836 12872
rect 12526 12860 12532 12872
rect 12584 12860 12590 12912
rect 12710 12900 12716 12912
rect 12671 12872 12716 12900
rect 12710 12860 12716 12872
rect 12768 12860 12774 12912
rect 11974 12792 11980 12844
rect 12032 12832 12038 12844
rect 12161 12835 12219 12841
rect 12161 12832 12173 12835
rect 12032 12804 12173 12832
rect 12032 12792 12038 12804
rect 12161 12801 12173 12804
rect 12207 12801 12219 12835
rect 12802 12832 12808 12844
rect 12715 12804 12808 12832
rect 12161 12795 12219 12801
rect 12802 12792 12808 12804
rect 12860 12832 12866 12844
rect 13449 12835 13507 12841
rect 13449 12832 13461 12835
rect 12860 12804 13461 12832
rect 12860 12792 12866 12804
rect 13449 12801 13461 12804
rect 13495 12801 13507 12835
rect 13556 12832 13584 12940
rect 13630 12928 13636 12980
rect 13688 12968 13694 12980
rect 13688 12940 14228 12968
rect 13688 12928 13694 12940
rect 14090 12900 14096 12912
rect 14051 12872 14096 12900
rect 14090 12860 14096 12872
rect 14148 12860 14154 12912
rect 14200 12900 14228 12940
rect 14458 12928 14464 12980
rect 14516 12968 14522 12980
rect 14553 12971 14611 12977
rect 14553 12968 14565 12971
rect 14516 12940 14565 12968
rect 14516 12928 14522 12940
rect 14553 12937 14565 12940
rect 14599 12968 14611 12971
rect 14918 12968 14924 12980
rect 14599 12940 14924 12968
rect 14599 12937 14611 12940
rect 14553 12931 14611 12937
rect 14918 12928 14924 12940
rect 14976 12928 14982 12980
rect 17402 12968 17408 12980
rect 17363 12940 17408 12968
rect 17402 12928 17408 12940
rect 17460 12928 17466 12980
rect 18509 12971 18567 12977
rect 18509 12937 18521 12971
rect 18555 12968 18567 12971
rect 19426 12968 19432 12980
rect 18555 12940 19432 12968
rect 18555 12937 18567 12940
rect 18509 12931 18567 12937
rect 19426 12928 19432 12940
rect 19484 12928 19490 12980
rect 19518 12928 19524 12980
rect 19576 12968 19582 12980
rect 22373 12971 22431 12977
rect 22373 12968 22385 12971
rect 19576 12940 22385 12968
rect 19576 12928 19582 12940
rect 22373 12937 22385 12940
rect 22419 12937 22431 12971
rect 22922 12968 22928 12980
rect 22883 12940 22928 12968
rect 22373 12931 22431 12937
rect 22922 12928 22928 12940
rect 22980 12928 22986 12980
rect 23382 12968 23388 12980
rect 23343 12940 23388 12968
rect 23382 12928 23388 12940
rect 23440 12928 23446 12980
rect 24210 12968 24216 12980
rect 24171 12940 24216 12968
rect 24210 12928 24216 12940
rect 24268 12928 24274 12980
rect 25593 12971 25651 12977
rect 25593 12968 25605 12971
rect 24688 12940 25605 12968
rect 16393 12903 16451 12909
rect 16393 12900 16405 12903
rect 14200 12872 16405 12900
rect 16393 12869 16405 12872
rect 16439 12869 16451 12903
rect 17420 12900 17448 12928
rect 17420 12872 19564 12900
rect 16393 12863 16451 12869
rect 19536 12844 19564 12872
rect 20806 12860 20812 12912
rect 20864 12900 20870 12912
rect 22462 12900 22468 12912
rect 20864 12872 22468 12900
rect 20864 12860 20870 12872
rect 22462 12860 22468 12872
rect 22520 12860 22526 12912
rect 22646 12860 22652 12912
rect 22704 12900 22710 12912
rect 23290 12900 23296 12912
rect 22704 12872 23296 12900
rect 22704 12860 22710 12872
rect 23290 12860 23296 12872
rect 23348 12900 23354 12912
rect 24489 12903 24547 12909
rect 24489 12900 24501 12903
rect 23348 12872 24501 12900
rect 23348 12860 23354 12872
rect 24489 12869 24501 12872
rect 24535 12869 24547 12903
rect 24489 12863 24547 12869
rect 13556 12804 18552 12832
rect 13449 12795 13507 12801
rect 12584 12767 12642 12773
rect 12584 12733 12596 12767
rect 12630 12764 12642 12767
rect 13078 12764 13084 12776
rect 12630 12736 13084 12764
rect 12630 12733 12642 12736
rect 12584 12727 12642 12733
rect 13078 12724 13084 12736
rect 13136 12724 13142 12776
rect 14734 12764 14740 12776
rect 14695 12736 14740 12764
rect 14734 12724 14740 12736
rect 14792 12724 14798 12776
rect 14829 12767 14887 12773
rect 14829 12733 14841 12767
rect 14875 12733 14887 12767
rect 15286 12764 15292 12776
rect 15247 12736 15292 12764
rect 14829 12727 14887 12733
rect 11793 12699 11851 12705
rect 11793 12696 11805 12699
rect 11296 12668 11805 12696
rect 11296 12656 11302 12668
rect 11793 12665 11805 12668
rect 11839 12665 11851 12699
rect 11793 12659 11851 12665
rect 11882 12656 11888 12708
rect 11940 12696 11946 12708
rect 12437 12699 12495 12705
rect 12437 12696 12449 12699
rect 11940 12668 12449 12696
rect 11940 12656 11946 12668
rect 12437 12665 12449 12668
rect 12483 12665 12495 12699
rect 12437 12659 12495 12665
rect 14461 12699 14519 12705
rect 14461 12665 14473 12699
rect 14507 12696 14519 12699
rect 14844 12696 14872 12727
rect 15286 12724 15292 12736
rect 15344 12724 15350 12776
rect 16025 12767 16083 12773
rect 16025 12733 16037 12767
rect 16071 12764 16083 12767
rect 16577 12767 16635 12773
rect 16577 12764 16589 12767
rect 16071 12736 16589 12764
rect 16071 12733 16083 12736
rect 16025 12727 16083 12733
rect 16577 12733 16589 12736
rect 16623 12733 16635 12767
rect 16942 12764 16948 12776
rect 16903 12736 16948 12764
rect 16577 12727 16635 12733
rect 15194 12696 15200 12708
rect 14507 12668 15200 12696
rect 14507 12665 14519 12668
rect 14461 12659 14519 12665
rect 15194 12656 15200 12668
rect 15252 12656 15258 12708
rect 10229 12631 10287 12637
rect 10229 12628 10241 12631
rect 10060 12600 10241 12628
rect 10229 12597 10241 12600
rect 10275 12628 10287 12631
rect 11333 12631 11391 12637
rect 11333 12628 11345 12631
rect 10275 12600 11345 12628
rect 10275 12597 10287 12600
rect 10229 12591 10287 12597
rect 11333 12597 11345 12600
rect 11379 12597 11391 12631
rect 11333 12591 11391 12597
rect 12250 12588 12256 12640
rect 12308 12628 12314 12640
rect 13081 12631 13139 12637
rect 13081 12628 13093 12631
rect 12308 12600 13093 12628
rect 12308 12588 12314 12600
rect 13081 12597 13093 12600
rect 13127 12597 13139 12631
rect 13081 12591 13139 12597
rect 13722 12588 13728 12640
rect 13780 12628 13786 12640
rect 15470 12628 15476 12640
rect 13780 12600 15476 12628
rect 13780 12588 13786 12600
rect 15470 12588 15476 12600
rect 15528 12588 15534 12640
rect 15657 12631 15715 12637
rect 15657 12597 15669 12631
rect 15703 12628 15715 12631
rect 16022 12628 16028 12640
rect 15703 12600 16028 12628
rect 15703 12597 15715 12600
rect 15657 12591 15715 12597
rect 16022 12588 16028 12600
rect 16080 12588 16086 12640
rect 16592 12628 16620 12727
rect 16942 12724 16948 12736
rect 17000 12724 17006 12776
rect 17037 12767 17095 12773
rect 17037 12733 17049 12767
rect 17083 12764 17095 12767
rect 17494 12764 17500 12776
rect 17083 12736 17500 12764
rect 17083 12733 17095 12736
rect 17037 12727 17095 12733
rect 17494 12724 17500 12736
rect 17552 12724 17558 12776
rect 18230 12764 18236 12776
rect 18191 12736 18236 12764
rect 18230 12724 18236 12736
rect 18288 12724 18294 12776
rect 18322 12724 18328 12776
rect 18380 12764 18386 12776
rect 18417 12767 18475 12773
rect 18417 12764 18429 12767
rect 18380 12736 18429 12764
rect 18380 12724 18386 12736
rect 18417 12733 18429 12736
rect 18463 12733 18475 12767
rect 18524 12764 18552 12804
rect 19518 12792 19524 12844
rect 19576 12792 19582 12844
rect 24688 12841 24716 12940
rect 25593 12937 25605 12940
rect 25639 12968 25651 12971
rect 27706 12968 27712 12980
rect 25639 12940 27712 12968
rect 25639 12937 25651 12940
rect 25593 12931 25651 12937
rect 27706 12928 27712 12940
rect 27764 12928 27770 12980
rect 28077 12971 28135 12977
rect 28077 12937 28089 12971
rect 28123 12968 28135 12971
rect 28166 12968 28172 12980
rect 28123 12940 28172 12968
rect 28123 12937 28135 12940
rect 28077 12931 28135 12937
rect 28166 12928 28172 12940
rect 28224 12928 28230 12980
rect 28445 12971 28503 12977
rect 28445 12937 28457 12971
rect 28491 12968 28503 12971
rect 28810 12968 28816 12980
rect 28491 12940 28816 12968
rect 28491 12937 28503 12940
rect 28445 12931 28503 12937
rect 28810 12928 28816 12940
rect 28868 12928 28874 12980
rect 30926 12968 30932 12980
rect 30887 12940 30932 12968
rect 30926 12928 30932 12940
rect 30984 12928 30990 12980
rect 32582 12968 32588 12980
rect 31128 12940 32588 12968
rect 25961 12903 26019 12909
rect 25961 12869 25973 12903
rect 26007 12900 26019 12903
rect 26050 12900 26056 12912
rect 26007 12872 26056 12900
rect 26007 12869 26019 12872
rect 25961 12863 26019 12869
rect 26050 12860 26056 12872
rect 26108 12860 26114 12912
rect 27154 12860 27160 12912
rect 27212 12900 27218 12912
rect 27433 12903 27491 12909
rect 27433 12900 27445 12903
rect 27212 12872 27445 12900
rect 27212 12860 27218 12872
rect 27433 12869 27445 12872
rect 27479 12900 27491 12903
rect 27801 12903 27859 12909
rect 27801 12900 27813 12903
rect 27479 12872 27813 12900
rect 27479 12869 27491 12872
rect 27433 12863 27491 12869
rect 27801 12869 27813 12872
rect 27847 12869 27859 12903
rect 27801 12863 27859 12869
rect 28350 12860 28356 12912
rect 28408 12900 28414 12912
rect 29457 12903 29515 12909
rect 29457 12900 29469 12903
rect 28408 12872 29469 12900
rect 28408 12860 28414 12872
rect 29457 12869 29469 12872
rect 29503 12900 29515 12903
rect 29733 12903 29791 12909
rect 29733 12900 29745 12903
rect 29503 12872 29745 12900
rect 29503 12869 29515 12872
rect 29457 12863 29515 12869
rect 29733 12869 29745 12872
rect 29779 12869 29791 12903
rect 29733 12863 29791 12869
rect 29822 12860 29828 12912
rect 29880 12900 29886 12912
rect 29917 12903 29975 12909
rect 29917 12900 29929 12903
rect 29880 12872 29929 12900
rect 29880 12860 29886 12872
rect 29917 12869 29929 12872
rect 29963 12900 29975 12903
rect 31128 12900 31156 12940
rect 32582 12928 32588 12940
rect 32640 12928 32646 12980
rect 32674 12928 32680 12980
rect 32732 12968 32738 12980
rect 32732 12940 32777 12968
rect 32732 12928 32738 12940
rect 33502 12928 33508 12980
rect 33560 12968 33566 12980
rect 35161 12971 35219 12977
rect 35161 12968 35173 12971
rect 33560 12940 35173 12968
rect 33560 12928 33566 12940
rect 35161 12937 35173 12940
rect 35207 12937 35219 12971
rect 35161 12931 35219 12937
rect 36170 12928 36176 12980
rect 36228 12968 36234 12980
rect 36354 12968 36360 12980
rect 36228 12940 36360 12968
rect 36228 12928 36234 12940
rect 36354 12928 36360 12940
rect 36412 12928 36418 12980
rect 38102 12968 38108 12980
rect 38063 12940 38108 12968
rect 38102 12928 38108 12940
rect 38160 12928 38166 12980
rect 38565 12971 38623 12977
rect 38565 12937 38577 12971
rect 38611 12968 38623 12971
rect 38838 12968 38844 12980
rect 38611 12940 38844 12968
rect 38611 12937 38623 12940
rect 38565 12931 38623 12937
rect 38838 12928 38844 12940
rect 38896 12968 38902 12980
rect 39301 12971 39359 12977
rect 39301 12968 39313 12971
rect 38896 12940 39313 12968
rect 38896 12928 38902 12940
rect 39301 12937 39313 12940
rect 39347 12937 39359 12971
rect 39301 12931 39359 12937
rect 39390 12928 39396 12980
rect 39448 12968 39454 12980
rect 39853 12971 39911 12977
rect 39853 12968 39865 12971
rect 39448 12940 39865 12968
rect 39448 12928 39454 12940
rect 39853 12937 39865 12940
rect 39899 12937 39911 12971
rect 39853 12931 39911 12937
rect 40402 12928 40408 12980
rect 40460 12968 40466 12980
rect 40681 12971 40739 12977
rect 40681 12968 40693 12971
rect 40460 12940 40693 12968
rect 40460 12928 40466 12940
rect 40681 12937 40693 12940
rect 40727 12937 40739 12971
rect 40681 12931 40739 12937
rect 40862 12928 40868 12980
rect 40920 12968 40926 12980
rect 41049 12971 41107 12977
rect 41049 12968 41061 12971
rect 40920 12940 41061 12968
rect 40920 12928 40926 12940
rect 41049 12937 41061 12940
rect 41095 12937 41107 12971
rect 41506 12968 41512 12980
rect 41467 12940 41512 12968
rect 41049 12931 41107 12937
rect 41506 12928 41512 12940
rect 41564 12928 41570 12980
rect 44545 12971 44603 12977
rect 44545 12968 44557 12971
rect 41616 12940 44557 12968
rect 34974 12900 34980 12912
rect 29963 12872 31156 12900
rect 32968 12872 34980 12900
rect 29963 12869 29975 12872
rect 29917 12863 29975 12869
rect 24673 12835 24731 12841
rect 24673 12801 24685 12835
rect 24719 12801 24731 12835
rect 24673 12795 24731 12801
rect 25225 12835 25283 12841
rect 25225 12801 25237 12835
rect 25271 12832 25283 12835
rect 26326 12832 26332 12844
rect 25271 12804 26332 12832
rect 25271 12801 25283 12804
rect 25225 12795 25283 12801
rect 26326 12792 26332 12804
rect 26384 12792 26390 12844
rect 31662 12832 31668 12844
rect 26436 12804 31668 12832
rect 19617 12773 19623 12776
rect 19613 12764 19623 12773
rect 18524 12736 19472 12764
rect 19578 12736 19623 12764
rect 18417 12727 18475 12733
rect 17512 12696 17540 12724
rect 18690 12696 18696 12708
rect 17512 12668 18696 12696
rect 18690 12656 18696 12668
rect 18748 12656 18754 12708
rect 16942 12628 16948 12640
rect 16592 12600 16948 12628
rect 16942 12588 16948 12600
rect 17000 12588 17006 12640
rect 17678 12588 17684 12640
rect 17736 12628 17742 12640
rect 17865 12631 17923 12637
rect 17865 12628 17877 12631
rect 17736 12600 17877 12628
rect 17736 12588 17742 12600
rect 17865 12597 17877 12600
rect 17911 12628 17923 12631
rect 18874 12628 18880 12640
rect 17911 12600 18880 12628
rect 17911 12597 17923 12600
rect 17865 12591 17923 12597
rect 18874 12588 18880 12600
rect 18932 12588 18938 12640
rect 18966 12588 18972 12640
rect 19024 12628 19030 12640
rect 19061 12631 19119 12637
rect 19061 12628 19073 12631
rect 19024 12600 19073 12628
rect 19024 12588 19030 12600
rect 19061 12597 19073 12600
rect 19107 12597 19119 12631
rect 19444 12628 19472 12736
rect 19613 12727 19623 12736
rect 19617 12724 19623 12727
rect 19675 12724 19681 12776
rect 19889 12767 19947 12773
rect 19889 12733 19901 12767
rect 19935 12764 19947 12767
rect 20898 12764 20904 12776
rect 19935 12736 20904 12764
rect 19935 12733 19947 12736
rect 19889 12727 19947 12733
rect 20898 12724 20904 12736
rect 20956 12724 20962 12776
rect 22281 12767 22339 12773
rect 22281 12733 22293 12767
rect 22327 12764 22339 12767
rect 22830 12764 22836 12776
rect 22327 12736 22836 12764
rect 22327 12733 22339 12736
rect 22281 12727 22339 12733
rect 22830 12724 22836 12736
rect 22888 12724 22894 12776
rect 23658 12764 23664 12776
rect 23619 12736 23664 12764
rect 23658 12724 23664 12736
rect 23716 12724 23722 12776
rect 24765 12767 24823 12773
rect 24765 12733 24777 12767
rect 24811 12764 24823 12767
rect 24854 12764 24860 12776
rect 24811 12736 24860 12764
rect 24811 12733 24823 12736
rect 24765 12727 24823 12733
rect 24854 12724 24860 12736
rect 24912 12724 24918 12776
rect 25958 12724 25964 12776
rect 26016 12764 26022 12776
rect 26053 12767 26111 12773
rect 26053 12764 26065 12767
rect 26016 12736 26065 12764
rect 26016 12724 26022 12736
rect 26053 12733 26065 12736
rect 26099 12733 26111 12767
rect 26436 12764 26464 12804
rect 31662 12792 31668 12804
rect 31720 12792 31726 12844
rect 31757 12835 31815 12841
rect 31757 12801 31769 12835
rect 31803 12832 31815 12835
rect 32968 12832 32996 12872
rect 34974 12860 34980 12872
rect 35032 12860 35038 12912
rect 35250 12860 35256 12912
rect 35308 12900 35314 12912
rect 41322 12900 41328 12912
rect 35308 12872 41328 12900
rect 35308 12860 35314 12872
rect 41322 12860 41328 12872
rect 41380 12860 41386 12912
rect 41616 12900 41644 12940
rect 44545 12937 44557 12940
rect 44591 12937 44603 12971
rect 45186 12968 45192 12980
rect 45147 12940 45192 12968
rect 44545 12931 44603 12937
rect 45186 12928 45192 12940
rect 45244 12928 45250 12980
rect 45649 12971 45707 12977
rect 45649 12937 45661 12971
rect 45695 12968 45707 12971
rect 46934 12968 46940 12980
rect 45695 12940 46940 12968
rect 45695 12937 45707 12940
rect 45649 12931 45707 12937
rect 43530 12900 43536 12912
rect 41432 12872 41644 12900
rect 43491 12872 43536 12900
rect 33134 12832 33140 12844
rect 31803 12804 32996 12832
rect 33095 12804 33140 12832
rect 31803 12801 31815 12804
rect 31757 12795 31815 12801
rect 33134 12792 33140 12804
rect 33192 12792 33198 12844
rect 33410 12792 33416 12844
rect 33468 12832 33474 12844
rect 33689 12835 33747 12841
rect 33689 12832 33701 12835
rect 33468 12804 33701 12832
rect 33468 12792 33474 12804
rect 33689 12801 33701 12804
rect 33735 12832 33747 12835
rect 33778 12832 33784 12844
rect 33735 12804 33784 12832
rect 33735 12801 33747 12804
rect 33689 12795 33747 12801
rect 33778 12792 33784 12804
rect 33836 12792 33842 12844
rect 34238 12792 34244 12844
rect 34296 12832 34302 12844
rect 36265 12835 36323 12841
rect 36265 12832 36277 12835
rect 34296 12804 36277 12832
rect 34296 12792 34302 12804
rect 36265 12801 36277 12804
rect 36311 12801 36323 12835
rect 36265 12795 36323 12801
rect 37553 12835 37611 12841
rect 37553 12801 37565 12835
rect 37599 12832 37611 12835
rect 38746 12832 38752 12844
rect 37599 12804 38752 12832
rect 37599 12801 37611 12804
rect 37553 12795 37611 12801
rect 38746 12792 38752 12804
rect 38804 12792 38810 12844
rect 41432 12832 41460 12872
rect 43530 12860 43536 12872
rect 43588 12860 43594 12912
rect 43714 12860 43720 12912
rect 43772 12900 43778 12912
rect 45664 12900 45692 12931
rect 46934 12928 46940 12940
rect 46992 12928 46998 12980
rect 47210 12968 47216 12980
rect 47171 12940 47216 12968
rect 47210 12928 47216 12940
rect 47268 12928 47274 12980
rect 47578 12968 47584 12980
rect 47539 12940 47584 12968
rect 47578 12928 47584 12940
rect 47636 12928 47642 12980
rect 48038 12928 48044 12980
rect 48096 12968 48102 12980
rect 48639 12971 48697 12977
rect 48639 12968 48651 12971
rect 48096 12940 48651 12968
rect 48096 12928 48102 12940
rect 48639 12937 48651 12940
rect 48685 12937 48697 12971
rect 48639 12931 48697 12937
rect 49145 12971 49203 12977
rect 49145 12937 49157 12971
rect 49191 12968 49203 12971
rect 49602 12968 49608 12980
rect 49191 12940 49608 12968
rect 49191 12937 49203 12940
rect 49145 12931 49203 12937
rect 49602 12928 49608 12940
rect 49660 12928 49666 12980
rect 50706 12968 50712 12980
rect 50667 12940 50712 12968
rect 50706 12928 50712 12940
rect 50764 12928 50770 12980
rect 52546 12928 52552 12980
rect 52604 12968 52610 12980
rect 58250 12968 58256 12980
rect 52604 12940 57376 12968
rect 58211 12940 58256 12968
rect 52604 12928 52610 12940
rect 47118 12909 47124 12912
rect 43772 12872 45692 12900
rect 46477 12903 46535 12909
rect 43772 12860 43778 12872
rect 46477 12869 46489 12903
rect 46523 12900 46535 12903
rect 47075 12903 47124 12909
rect 47075 12900 47087 12903
rect 46523 12872 47087 12900
rect 46523 12869 46535 12872
rect 46477 12863 46535 12869
rect 47075 12869 47087 12872
rect 47121 12869 47124 12903
rect 47075 12863 47124 12869
rect 47118 12860 47124 12863
rect 47176 12860 47182 12912
rect 47228 12900 47256 12928
rect 48777 12903 48835 12909
rect 48777 12900 48789 12903
rect 47228 12872 48789 12900
rect 48777 12869 48789 12872
rect 48823 12900 48835 12903
rect 49234 12900 49240 12912
rect 48823 12872 49240 12900
rect 48823 12869 48835 12872
rect 48777 12863 48835 12869
rect 49234 12860 49240 12872
rect 49292 12900 49298 12912
rect 49881 12903 49939 12909
rect 49881 12900 49893 12903
rect 49292 12872 49893 12900
rect 49292 12860 49298 12872
rect 49881 12869 49893 12872
rect 49927 12900 49939 12903
rect 50246 12900 50252 12912
rect 49927 12872 50252 12900
rect 49927 12869 49939 12872
rect 49881 12863 49939 12869
rect 50246 12860 50252 12872
rect 50304 12900 50310 12912
rect 50341 12903 50399 12909
rect 50341 12900 50353 12903
rect 50304 12872 50353 12900
rect 50304 12860 50310 12872
rect 50341 12869 50353 12872
rect 50387 12869 50399 12903
rect 51077 12903 51135 12909
rect 51077 12900 51089 12903
rect 50341 12863 50399 12869
rect 50448 12872 51089 12900
rect 42978 12832 42984 12844
rect 40236 12804 41460 12832
rect 41623 12804 42984 12832
rect 26053 12727 26111 12733
rect 26160 12736 26464 12764
rect 27801 12767 27859 12773
rect 19518 12656 19524 12708
rect 19576 12696 19582 12708
rect 19576 12668 19621 12696
rect 20548 12668 21404 12696
rect 19576 12656 19582 12668
rect 20548 12628 20576 12668
rect 19444 12600 20576 12628
rect 19061 12591 19119 12597
rect 21174 12588 21180 12640
rect 21232 12628 21238 12640
rect 21376 12628 21404 12668
rect 21818 12656 21824 12708
rect 21876 12696 21882 12708
rect 22097 12699 22155 12705
rect 21876 12668 21921 12696
rect 21876 12656 21882 12668
rect 22097 12665 22109 12699
rect 22143 12696 22155 12699
rect 22186 12696 22192 12708
rect 22143 12668 22192 12696
rect 22143 12665 22155 12668
rect 22097 12659 22155 12665
rect 22186 12656 22192 12668
rect 22244 12656 22250 12708
rect 22462 12656 22468 12708
rect 22520 12696 22526 12708
rect 23753 12699 23811 12705
rect 23753 12696 23765 12699
rect 22520 12668 23765 12696
rect 22520 12656 22526 12668
rect 23753 12665 23765 12668
rect 23799 12696 23811 12699
rect 26160 12696 26188 12736
rect 27801 12733 27813 12767
rect 27847 12764 27859 12767
rect 28534 12764 28540 12776
rect 27847 12736 28540 12764
rect 27847 12733 27859 12736
rect 27801 12727 27859 12733
rect 28534 12724 28540 12736
rect 28592 12764 28598 12776
rect 29273 12767 29331 12773
rect 29273 12764 29285 12767
rect 28592 12736 29285 12764
rect 28592 12724 28598 12736
rect 29273 12733 29285 12736
rect 29319 12764 29331 12767
rect 30190 12764 30196 12776
rect 29319 12736 30196 12764
rect 29319 12733 29331 12736
rect 29273 12727 29331 12733
rect 30190 12724 30196 12736
rect 30248 12724 30254 12776
rect 31386 12724 31392 12776
rect 31444 12764 31450 12776
rect 31444 12736 31489 12764
rect 31444 12724 31450 12736
rect 31570 12724 31576 12776
rect 31628 12764 31634 12776
rect 31628 12736 32536 12764
rect 31628 12724 31634 12736
rect 30006 12696 30012 12708
rect 23799 12668 26188 12696
rect 28552 12668 30012 12696
rect 23799 12665 23811 12668
rect 23753 12659 23811 12665
rect 22554 12628 22560 12640
rect 21232 12600 21277 12628
rect 21376 12600 22560 12628
rect 21232 12588 21238 12600
rect 22554 12588 22560 12600
rect 22612 12588 22618 12640
rect 24762 12588 24768 12640
rect 24820 12628 24826 12640
rect 28552 12628 28580 12668
rect 30006 12656 30012 12668
rect 30064 12656 30070 12708
rect 30653 12699 30711 12705
rect 30653 12665 30665 12699
rect 30699 12696 30711 12699
rect 31202 12696 31208 12708
rect 30699 12668 31208 12696
rect 30699 12665 30711 12668
rect 30653 12659 30711 12665
rect 31202 12656 31208 12668
rect 31260 12656 31266 12708
rect 32122 12696 32128 12708
rect 32083 12668 32128 12696
rect 32122 12656 32128 12668
rect 32180 12656 32186 12708
rect 28718 12628 28724 12640
rect 24820 12600 28580 12628
rect 28679 12600 28724 12628
rect 24820 12588 24826 12600
rect 28718 12588 28724 12600
rect 28776 12588 28782 12640
rect 29733 12631 29791 12637
rect 29733 12597 29745 12631
rect 29779 12628 29791 12631
rect 31386 12628 31392 12640
rect 29779 12600 31392 12628
rect 29779 12597 29791 12600
rect 29733 12591 29791 12597
rect 31386 12588 31392 12600
rect 31444 12588 31450 12640
rect 32030 12588 32036 12640
rect 32088 12628 32094 12640
rect 32401 12631 32459 12637
rect 32401 12628 32413 12631
rect 32088 12600 32413 12628
rect 32088 12588 32094 12600
rect 32401 12597 32413 12600
rect 32447 12597 32459 12631
rect 32508 12628 32536 12736
rect 33042 12724 33048 12776
rect 33100 12764 33106 12776
rect 33229 12767 33287 12773
rect 33229 12764 33241 12767
rect 33100 12736 33241 12764
rect 33100 12724 33106 12736
rect 33229 12733 33241 12736
rect 33275 12733 33287 12767
rect 33229 12727 33287 12733
rect 33598 12767 33656 12773
rect 33598 12733 33610 12767
rect 33644 12764 33656 12767
rect 33962 12764 33968 12776
rect 33644 12736 33968 12764
rect 33644 12733 33656 12736
rect 33598 12727 33656 12733
rect 33244 12696 33272 12727
rect 33962 12724 33968 12736
rect 34020 12764 34026 12776
rect 34514 12764 34520 12776
rect 34020 12736 34520 12764
rect 34020 12724 34026 12736
rect 34514 12724 34520 12736
rect 34572 12724 34578 12776
rect 35069 12767 35127 12773
rect 35069 12764 35081 12767
rect 34624 12736 35081 12764
rect 34054 12696 34060 12708
rect 33244 12668 34060 12696
rect 34054 12656 34060 12668
rect 34112 12656 34118 12708
rect 34624 12696 34652 12736
rect 35069 12733 35081 12736
rect 35115 12733 35127 12767
rect 35069 12727 35127 12733
rect 34164 12668 34652 12696
rect 34164 12628 34192 12668
rect 34790 12656 34796 12708
rect 34848 12696 34854 12708
rect 34885 12699 34943 12705
rect 34885 12696 34897 12699
rect 34848 12668 34897 12696
rect 34848 12656 34854 12668
rect 34885 12665 34897 12668
rect 34931 12665 34943 12699
rect 34885 12659 34943 12665
rect 34606 12628 34612 12640
rect 32508 12600 34192 12628
rect 34567 12600 34612 12628
rect 32401 12591 32459 12597
rect 34606 12588 34612 12600
rect 34664 12588 34670 12640
rect 35084 12628 35112 12727
rect 36170 12724 36176 12776
rect 36228 12764 36234 12776
rect 36722 12764 36728 12776
rect 36228 12736 36728 12764
rect 36228 12724 36234 12736
rect 36722 12724 36728 12736
rect 36780 12724 36786 12776
rect 36998 12764 37004 12776
rect 36959 12736 37004 12764
rect 36998 12724 37004 12736
rect 37056 12724 37062 12776
rect 37182 12764 37188 12776
rect 37143 12736 37188 12764
rect 37182 12724 37188 12736
rect 37240 12724 37246 12776
rect 37734 12764 37740 12776
rect 37695 12736 37740 12764
rect 37734 12724 37740 12736
rect 37792 12724 37798 12776
rect 38654 12724 38660 12776
rect 38712 12764 38718 12776
rect 39206 12773 39212 12776
rect 39025 12767 39083 12773
rect 39025 12764 39037 12767
rect 38712 12736 39037 12764
rect 38712 12724 38718 12736
rect 39025 12733 39037 12736
rect 39071 12733 39083 12767
rect 39025 12727 39083 12733
rect 39158 12767 39212 12773
rect 39158 12733 39170 12767
rect 39204 12733 39212 12767
rect 39158 12727 39212 12733
rect 39206 12724 39212 12727
rect 39264 12724 39270 12776
rect 35342 12656 35348 12708
rect 35400 12696 35406 12708
rect 40236 12696 40264 12804
rect 40497 12767 40555 12773
rect 40497 12733 40509 12767
rect 40543 12764 40555 12767
rect 40862 12764 40868 12776
rect 40543 12736 40868 12764
rect 40543 12733 40555 12736
rect 40497 12727 40555 12733
rect 40862 12724 40868 12736
rect 40920 12724 40926 12776
rect 41414 12724 41420 12776
rect 41472 12724 41478 12776
rect 41623 12773 41651 12804
rect 42978 12792 42984 12804
rect 43036 12792 43042 12844
rect 43257 12835 43315 12841
rect 43257 12801 43269 12835
rect 43303 12832 43315 12835
rect 43346 12832 43352 12844
rect 43303 12804 43352 12832
rect 43303 12801 43315 12804
rect 43257 12795 43315 12801
rect 43346 12792 43352 12804
rect 43404 12792 43410 12844
rect 43548 12832 43576 12860
rect 46753 12835 46811 12841
rect 46753 12832 46765 12835
rect 43548 12804 46765 12832
rect 46753 12801 46765 12804
rect 46799 12832 46811 12835
rect 46842 12832 46848 12844
rect 46799 12804 46848 12832
rect 46799 12801 46811 12804
rect 46753 12795 46811 12801
rect 46842 12792 46848 12804
rect 46900 12792 46906 12844
rect 47302 12832 47308 12844
rect 47263 12804 47308 12832
rect 47302 12792 47308 12804
rect 47360 12832 47366 12844
rect 47949 12835 48007 12841
rect 47949 12832 47961 12835
rect 47360 12804 47961 12832
rect 47360 12792 47366 12804
rect 47949 12801 47961 12804
rect 47995 12832 48007 12835
rect 48317 12835 48375 12841
rect 48317 12832 48329 12835
rect 47995 12804 48329 12832
rect 47995 12801 48007 12804
rect 47949 12795 48007 12801
rect 48317 12801 48329 12804
rect 48363 12832 48375 12835
rect 48682 12832 48688 12844
rect 48363 12804 48688 12832
rect 48363 12801 48375 12804
rect 48317 12795 48375 12801
rect 48682 12792 48688 12804
rect 48740 12832 48746 12844
rect 50448 12841 50476 12872
rect 51077 12869 51089 12872
rect 51123 12869 51135 12903
rect 51077 12863 51135 12869
rect 52362 12860 52368 12912
rect 52420 12900 52426 12912
rect 52641 12903 52699 12909
rect 52641 12900 52653 12903
rect 52420 12872 52653 12900
rect 52420 12860 52426 12872
rect 52641 12869 52653 12872
rect 52687 12900 52699 12903
rect 53650 12900 53656 12912
rect 52687 12872 53656 12900
rect 52687 12869 52699 12872
rect 52641 12863 52699 12869
rect 53650 12860 53656 12872
rect 53708 12860 53714 12912
rect 56042 12900 56048 12912
rect 53852 12872 56048 12900
rect 48869 12835 48927 12841
rect 48869 12832 48881 12835
rect 48740 12804 48881 12832
rect 48740 12792 48746 12804
rect 48869 12801 48881 12804
rect 48915 12832 48927 12835
rect 49513 12835 49571 12841
rect 49513 12832 49525 12835
rect 48915 12804 49525 12832
rect 48915 12801 48927 12804
rect 48869 12795 48927 12801
rect 49513 12801 49525 12804
rect 49559 12832 49571 12835
rect 50433 12835 50491 12841
rect 50433 12832 50445 12835
rect 49559 12804 50445 12832
rect 49559 12801 49571 12804
rect 49513 12795 49571 12801
rect 50433 12801 50445 12804
rect 50479 12801 50491 12835
rect 50433 12795 50491 12801
rect 50522 12792 50528 12844
rect 50580 12832 50586 12844
rect 53852 12841 53880 12872
rect 56042 12860 56048 12872
rect 56100 12860 56106 12912
rect 56778 12900 56784 12912
rect 56739 12872 56784 12900
rect 56778 12860 56784 12872
rect 56836 12860 56842 12912
rect 50893 12835 50951 12841
rect 50580 12804 50752 12832
rect 50580 12792 50586 12804
rect 41601 12767 41659 12773
rect 41601 12733 41613 12767
rect 41647 12733 41659 12767
rect 41877 12767 41935 12773
rect 41877 12764 41889 12767
rect 41601 12727 41659 12733
rect 41708 12736 41889 12764
rect 35400 12668 40264 12696
rect 40313 12699 40371 12705
rect 35400 12656 35406 12668
rect 40313 12665 40325 12699
rect 40359 12696 40371 12699
rect 41432 12696 41460 12724
rect 40359 12668 41460 12696
rect 40359 12665 40371 12668
rect 40313 12659 40371 12665
rect 35802 12628 35808 12640
rect 35084 12600 35808 12628
rect 35802 12588 35808 12600
rect 35860 12588 35866 12640
rect 36173 12631 36231 12637
rect 36173 12597 36185 12631
rect 36219 12628 36231 12631
rect 36446 12628 36452 12640
rect 36219 12600 36452 12628
rect 36219 12597 36231 12600
rect 36173 12591 36231 12597
rect 36446 12588 36452 12600
rect 36504 12588 36510 12640
rect 38102 12588 38108 12640
rect 38160 12628 38166 12640
rect 38838 12628 38844 12640
rect 38160 12600 38844 12628
rect 38160 12588 38166 12600
rect 38838 12588 38844 12600
rect 38896 12588 38902 12640
rect 38933 12631 38991 12637
rect 38933 12597 38945 12631
rect 38979 12628 38991 12631
rect 39022 12628 39028 12640
rect 38979 12600 39028 12628
rect 38979 12597 38991 12600
rect 38933 12591 38991 12597
rect 39022 12588 39028 12600
rect 39080 12628 39086 12640
rect 39482 12628 39488 12640
rect 39080 12600 39488 12628
rect 39080 12588 39086 12600
rect 39482 12588 39488 12600
rect 39540 12588 39546 12640
rect 41708 12628 41736 12736
rect 41877 12733 41889 12736
rect 41923 12733 41935 12767
rect 41877 12727 41935 12733
rect 44453 12767 44511 12773
rect 44453 12733 44465 12767
rect 44499 12764 44511 12767
rect 44542 12764 44548 12776
rect 44499 12736 44548 12764
rect 44499 12733 44511 12736
rect 44453 12727 44511 12733
rect 44542 12724 44548 12736
rect 44600 12724 44606 12776
rect 45554 12724 45560 12776
rect 45612 12764 45618 12776
rect 45830 12764 45836 12776
rect 45612 12736 45836 12764
rect 45612 12724 45618 12736
rect 45830 12724 45836 12736
rect 45888 12724 45894 12776
rect 45922 12724 45928 12776
rect 45980 12764 45986 12776
rect 49418 12764 49424 12776
rect 45980 12736 49424 12764
rect 45980 12724 45986 12736
rect 49418 12724 49424 12736
rect 49476 12724 49482 12776
rect 50212 12767 50270 12773
rect 50212 12733 50224 12767
rect 50258 12764 50270 12767
rect 50724 12764 50752 12804
rect 50893 12801 50905 12835
rect 50939 12832 50951 12835
rect 53837 12835 53895 12841
rect 50939 12804 53788 12832
rect 50939 12801 50951 12804
rect 50893 12795 50951 12801
rect 51902 12764 51908 12776
rect 50258 12736 50660 12764
rect 50724 12736 51908 12764
rect 50258 12733 50270 12736
rect 50212 12727 50270 12733
rect 43346 12656 43352 12708
rect 43404 12696 43410 12708
rect 43901 12699 43959 12705
rect 43901 12696 43913 12699
rect 43404 12668 43913 12696
rect 43404 12656 43410 12668
rect 43901 12665 43913 12668
rect 43947 12665 43959 12699
rect 44266 12696 44272 12708
rect 44227 12668 44272 12696
rect 43901 12659 43959 12665
rect 44266 12656 44272 12668
rect 44324 12656 44330 12708
rect 46934 12696 46940 12708
rect 46895 12668 46940 12696
rect 46934 12656 46940 12668
rect 46992 12656 46998 12708
rect 48498 12696 48504 12708
rect 48459 12668 48504 12696
rect 48498 12656 48504 12668
rect 48556 12656 48562 12708
rect 50062 12696 50068 12708
rect 50023 12668 50068 12696
rect 50062 12656 50068 12668
rect 50120 12656 50126 12708
rect 50632 12696 50660 12736
rect 51902 12724 51908 12736
rect 51960 12724 51966 12776
rect 53282 12764 53288 12776
rect 53243 12736 53288 12764
rect 53282 12724 53288 12736
rect 53340 12724 53346 12776
rect 53377 12767 53435 12773
rect 53377 12733 53389 12767
rect 53423 12764 53435 12767
rect 53466 12764 53472 12776
rect 53423 12736 53472 12764
rect 53423 12733 53435 12736
rect 53377 12727 53435 12733
rect 53466 12724 53472 12736
rect 53524 12724 53530 12776
rect 51445 12699 51503 12705
rect 51445 12696 51457 12699
rect 50632 12668 51457 12696
rect 51445 12665 51457 12668
rect 51491 12696 51503 12699
rect 51534 12696 51540 12708
rect 51491 12668 51540 12696
rect 51491 12665 51503 12668
rect 51445 12659 51503 12665
rect 51534 12656 51540 12668
rect 51592 12656 51598 12708
rect 51721 12699 51779 12705
rect 51721 12665 51733 12699
rect 51767 12696 51779 12699
rect 52917 12699 52975 12705
rect 52917 12696 52929 12699
rect 51767 12668 52929 12696
rect 51767 12665 51779 12668
rect 51721 12659 51779 12665
rect 52917 12665 52929 12668
rect 52963 12696 52975 12699
rect 53760 12696 53788 12804
rect 53837 12801 53849 12835
rect 53883 12801 53895 12835
rect 53837 12795 53895 12801
rect 55214 12792 55220 12844
rect 55272 12832 55278 12844
rect 55401 12835 55459 12841
rect 55401 12832 55413 12835
rect 55272 12804 55413 12832
rect 55272 12792 55278 12804
rect 55401 12801 55413 12804
rect 55447 12801 55459 12835
rect 55401 12795 55459 12801
rect 57348 12773 57376 12940
rect 58250 12928 58256 12940
rect 58308 12928 58314 12980
rect 57790 12792 57796 12844
rect 57848 12832 57854 12844
rect 58621 12835 58679 12841
rect 58621 12832 58633 12835
rect 57848 12804 58633 12832
rect 57848 12792 57854 12804
rect 58621 12801 58633 12804
rect 58667 12801 58679 12835
rect 58894 12832 58900 12844
rect 58807 12804 58900 12832
rect 58621 12795 58679 12801
rect 58894 12792 58900 12804
rect 58952 12832 58958 12844
rect 59262 12832 59268 12844
rect 58952 12804 59268 12832
rect 58952 12792 58958 12804
rect 59262 12792 59268 12804
rect 59320 12792 59326 12844
rect 54389 12767 54447 12773
rect 54389 12733 54401 12767
rect 54435 12764 54447 12767
rect 54665 12767 54723 12773
rect 54665 12764 54677 12767
rect 54435 12736 54677 12764
rect 54435 12733 54447 12736
rect 54389 12727 54447 12733
rect 54665 12733 54677 12736
rect 54711 12733 54723 12767
rect 54665 12727 54723 12733
rect 54941 12767 54999 12773
rect 54941 12733 54953 12767
rect 54987 12764 54999 12767
rect 57333 12767 57391 12773
rect 54987 12736 55904 12764
rect 54987 12733 54999 12736
rect 54941 12727 54999 12733
rect 55876 12708 55904 12736
rect 57333 12733 57345 12767
rect 57379 12764 57391 12767
rect 57885 12767 57943 12773
rect 57885 12764 57897 12767
rect 57379 12736 57897 12764
rect 57379 12733 57391 12736
rect 57333 12727 57391 12733
rect 57885 12733 57897 12736
rect 57931 12733 57943 12767
rect 57885 12727 57943 12733
rect 54849 12699 54907 12705
rect 52963 12668 53328 12696
rect 53760 12668 54616 12696
rect 52963 12665 52975 12668
rect 52917 12659 52975 12665
rect 53300 12640 53328 12668
rect 41966 12628 41972 12640
rect 41708 12600 41972 12628
rect 41966 12588 41972 12600
rect 42024 12588 42030 12640
rect 50246 12588 50252 12640
rect 50304 12628 50310 12640
rect 50893 12631 50951 12637
rect 50893 12628 50905 12631
rect 50304 12600 50905 12628
rect 50304 12588 50310 12600
rect 50893 12597 50905 12600
rect 50939 12597 50951 12631
rect 50893 12591 50951 12597
rect 51626 12588 51632 12640
rect 51684 12628 51690 12640
rect 51997 12631 52055 12637
rect 51997 12628 52009 12631
rect 51684 12600 52009 12628
rect 51684 12588 51690 12600
rect 51997 12597 52009 12600
rect 52043 12597 52055 12631
rect 51997 12591 52055 12597
rect 53282 12588 53288 12640
rect 53340 12588 53346 12640
rect 53374 12588 53380 12640
rect 53432 12628 53438 12640
rect 54113 12631 54171 12637
rect 54113 12628 54125 12631
rect 53432 12600 54125 12628
rect 53432 12588 53438 12600
rect 54113 12597 54125 12600
rect 54159 12628 54171 12631
rect 54389 12631 54447 12637
rect 54389 12628 54401 12631
rect 54159 12600 54401 12628
rect 54159 12597 54171 12600
rect 54113 12591 54171 12597
rect 54389 12597 54401 12600
rect 54435 12628 54447 12631
rect 54481 12631 54539 12637
rect 54481 12628 54493 12631
rect 54435 12600 54493 12628
rect 54435 12597 54447 12600
rect 54389 12591 54447 12597
rect 54481 12597 54493 12600
rect 54527 12597 54539 12631
rect 54588 12628 54616 12668
rect 54849 12665 54861 12699
rect 54895 12696 54907 12699
rect 55122 12696 55128 12708
rect 54895 12668 55128 12696
rect 54895 12665 54907 12668
rect 54849 12659 54907 12665
rect 55122 12656 55128 12668
rect 55180 12656 55186 12708
rect 55232 12668 55812 12696
rect 55232 12628 55260 12668
rect 55674 12628 55680 12640
rect 54588 12600 55260 12628
rect 55635 12600 55680 12628
rect 54481 12591 54539 12597
rect 55674 12588 55680 12600
rect 55732 12588 55738 12640
rect 55784 12628 55812 12668
rect 55858 12656 55864 12708
rect 55916 12696 55922 12708
rect 56413 12699 56471 12705
rect 56413 12696 56425 12699
rect 55916 12668 56425 12696
rect 55916 12656 55922 12668
rect 56413 12665 56425 12668
rect 56459 12665 56471 12699
rect 56413 12659 56471 12665
rect 57517 12631 57575 12637
rect 57517 12628 57529 12631
rect 55784 12600 57529 12628
rect 57517 12597 57529 12600
rect 57563 12597 57575 12631
rect 59998 12628 60004 12640
rect 59959 12600 60004 12628
rect 57517 12591 57575 12597
rect 59998 12588 60004 12600
rect 60056 12588 60062 12640
rect 1104 12538 63480 12560
rect 1104 12486 21774 12538
rect 21826 12486 21838 12538
rect 21890 12486 21902 12538
rect 21954 12486 21966 12538
rect 22018 12486 42566 12538
rect 42618 12486 42630 12538
rect 42682 12486 42694 12538
rect 42746 12486 42758 12538
rect 42810 12486 63480 12538
rect 1104 12464 63480 12486
rect 4062 12384 4068 12436
rect 4120 12424 4126 12436
rect 5902 12424 5908 12436
rect 4120 12396 5908 12424
rect 4120 12384 4126 12396
rect 5902 12384 5908 12396
rect 5960 12384 5966 12436
rect 6549 12427 6607 12433
rect 6549 12393 6561 12427
rect 6595 12424 6607 12427
rect 7006 12424 7012 12436
rect 6595 12396 7012 12424
rect 6595 12393 6607 12396
rect 6549 12387 6607 12393
rect 7006 12384 7012 12396
rect 7064 12384 7070 12436
rect 7285 12427 7343 12433
rect 7285 12393 7297 12427
rect 7331 12424 7343 12427
rect 7558 12424 7564 12436
rect 7331 12396 7564 12424
rect 7331 12393 7343 12396
rect 7285 12387 7343 12393
rect 7558 12384 7564 12396
rect 7616 12424 7622 12436
rect 7616 12396 8432 12424
rect 7616 12384 7622 12396
rect 3145 12359 3203 12365
rect 3145 12325 3157 12359
rect 3191 12356 3203 12359
rect 5350 12356 5356 12368
rect 3191 12328 5356 12356
rect 3191 12325 3203 12328
rect 3145 12319 3203 12325
rect 5350 12316 5356 12328
rect 5408 12316 5414 12368
rect 8113 12359 8171 12365
rect 8113 12325 8125 12359
rect 8159 12356 8171 12359
rect 8294 12356 8300 12368
rect 8159 12328 8300 12356
rect 8159 12325 8171 12328
rect 8113 12319 8171 12325
rect 8294 12316 8300 12328
rect 8352 12316 8358 12368
rect 8404 12356 8432 12396
rect 8754 12384 8760 12436
rect 8812 12424 8818 12436
rect 8849 12427 8907 12433
rect 8849 12424 8861 12427
rect 8812 12396 8861 12424
rect 8812 12384 8818 12396
rect 8849 12393 8861 12396
rect 8895 12393 8907 12427
rect 9858 12424 9864 12436
rect 8849 12387 8907 12393
rect 8956 12396 9864 12424
rect 8956 12356 8984 12396
rect 9858 12384 9864 12396
rect 9916 12384 9922 12436
rect 10229 12427 10287 12433
rect 10229 12393 10241 12427
rect 10275 12424 10287 12427
rect 10318 12424 10324 12436
rect 10275 12396 10324 12424
rect 10275 12393 10287 12396
rect 10229 12387 10287 12393
rect 10318 12384 10324 12396
rect 10376 12384 10382 12436
rect 11146 12384 11152 12436
rect 11204 12424 11210 12436
rect 11333 12427 11391 12433
rect 11333 12424 11345 12427
rect 11204 12396 11345 12424
rect 11204 12384 11210 12396
rect 11333 12393 11345 12396
rect 11379 12393 11391 12427
rect 12066 12424 12072 12436
rect 12027 12396 12072 12424
rect 11333 12387 11391 12393
rect 12066 12384 12072 12396
rect 12124 12384 12130 12436
rect 12158 12384 12164 12436
rect 12216 12424 12222 12436
rect 12437 12427 12495 12433
rect 12437 12424 12449 12427
rect 12216 12396 12449 12424
rect 12216 12384 12222 12396
rect 12437 12393 12449 12396
rect 12483 12424 12495 12427
rect 12802 12424 12808 12436
rect 12483 12396 12808 12424
rect 12483 12393 12495 12396
rect 12437 12387 12495 12393
rect 12802 12384 12808 12396
rect 12860 12384 12866 12436
rect 15470 12384 15476 12436
rect 15528 12424 15534 12436
rect 15565 12427 15623 12433
rect 15565 12424 15577 12427
rect 15528 12396 15577 12424
rect 15528 12384 15534 12396
rect 15565 12393 15577 12396
rect 15611 12393 15623 12427
rect 15565 12387 15623 12393
rect 16298 12384 16304 12436
rect 16356 12424 16362 12436
rect 17681 12427 17739 12433
rect 17681 12424 17693 12427
rect 16356 12396 17693 12424
rect 16356 12384 16362 12396
rect 17681 12393 17693 12396
rect 17727 12393 17739 12427
rect 17681 12387 17739 12393
rect 17770 12384 17776 12436
rect 17828 12424 17834 12436
rect 18049 12427 18107 12433
rect 18049 12424 18061 12427
rect 17828 12396 18061 12424
rect 17828 12384 17834 12396
rect 18049 12393 18061 12396
rect 18095 12393 18107 12427
rect 18049 12387 18107 12393
rect 19334 12384 19340 12436
rect 19392 12424 19398 12436
rect 19521 12427 19579 12433
rect 19521 12424 19533 12427
rect 19392 12396 19533 12424
rect 19392 12384 19398 12396
rect 19521 12393 19533 12396
rect 19567 12393 19579 12427
rect 19521 12387 19579 12393
rect 20254 12384 20260 12436
rect 20312 12424 20318 12436
rect 20312 12396 21036 12424
rect 20312 12384 20318 12396
rect 8404 12328 8984 12356
rect 9122 12316 9128 12368
rect 9180 12356 9186 12368
rect 9309 12359 9367 12365
rect 9309 12356 9321 12359
rect 9180 12328 9321 12356
rect 9180 12316 9186 12328
rect 9309 12325 9321 12328
rect 9355 12356 9367 12359
rect 13357 12359 13415 12365
rect 13357 12356 13369 12359
rect 9355 12328 13369 12356
rect 9355 12325 9367 12328
rect 9309 12319 9367 12325
rect 13357 12325 13369 12328
rect 13403 12325 13415 12359
rect 13357 12319 13415 12325
rect 15194 12316 15200 12368
rect 15252 12356 15258 12368
rect 17221 12359 17279 12365
rect 17221 12356 17233 12359
rect 15252 12328 17233 12356
rect 15252 12316 15258 12328
rect 17221 12325 17233 12328
rect 17267 12325 17279 12359
rect 17221 12319 17279 12325
rect 17310 12316 17316 12368
rect 17368 12356 17374 12368
rect 20898 12356 20904 12368
rect 17368 12328 20760 12356
rect 20859 12328 20904 12356
rect 17368 12316 17374 12328
rect 2593 12291 2651 12297
rect 2593 12257 2605 12291
rect 2639 12288 2651 12291
rect 2682 12288 2688 12300
rect 2639 12260 2688 12288
rect 2639 12257 2651 12260
rect 2593 12251 2651 12257
rect 2682 12248 2688 12260
rect 2740 12248 2746 12300
rect 2777 12291 2835 12297
rect 2777 12257 2789 12291
rect 2823 12257 2835 12291
rect 5074 12288 5080 12300
rect 5035 12260 5080 12288
rect 2777 12251 2835 12257
rect 2792 12152 2820 12251
rect 5074 12248 5080 12260
rect 5132 12248 5138 12300
rect 5442 12288 5448 12300
rect 5403 12260 5448 12288
rect 5442 12248 5448 12260
rect 5500 12248 5506 12300
rect 6546 12248 6552 12300
rect 6604 12288 6610 12300
rect 7377 12291 7435 12297
rect 7377 12288 7389 12291
rect 6604 12260 7389 12288
rect 6604 12248 6610 12260
rect 7377 12257 7389 12260
rect 7423 12257 7435 12291
rect 10686 12288 10692 12300
rect 10647 12260 10692 12288
rect 7377 12251 7435 12257
rect 10686 12248 10692 12260
rect 10744 12248 10750 12300
rect 11793 12291 11851 12297
rect 11793 12288 11805 12291
rect 11072 12260 11805 12288
rect 3326 12180 3332 12232
rect 3384 12220 3390 12232
rect 3513 12223 3571 12229
rect 3513 12220 3525 12223
rect 3384 12192 3525 12220
rect 3384 12180 3390 12192
rect 3513 12189 3525 12192
rect 3559 12220 3571 12223
rect 4617 12223 4675 12229
rect 4617 12220 4629 12223
rect 3559 12192 4629 12220
rect 3559 12189 3571 12192
rect 3513 12183 3571 12189
rect 4617 12189 4629 12192
rect 4663 12189 4675 12223
rect 5534 12220 5540 12232
rect 5495 12192 5540 12220
rect 4617 12183 4675 12189
rect 5534 12180 5540 12192
rect 5592 12180 5598 12232
rect 7558 12229 7564 12232
rect 7524 12223 7564 12229
rect 7524 12189 7536 12223
rect 7524 12183 7564 12189
rect 7558 12180 7564 12183
rect 7616 12180 7622 12232
rect 7745 12223 7803 12229
rect 7745 12189 7757 12223
rect 7791 12220 7803 12223
rect 8202 12220 8208 12232
rect 7791 12192 8208 12220
rect 7791 12189 7803 12192
rect 7745 12183 7803 12189
rect 8202 12180 8208 12192
rect 8260 12220 8266 12232
rect 11072 12229 11100 12260
rect 11793 12257 11805 12260
rect 11839 12288 11851 12291
rect 12158 12288 12164 12300
rect 11839 12260 12164 12288
rect 11839 12257 11851 12260
rect 11793 12251 11851 12257
rect 12158 12248 12164 12260
rect 12216 12248 12222 12300
rect 12253 12291 12311 12297
rect 12253 12257 12265 12291
rect 12299 12288 12311 12291
rect 12526 12288 12532 12300
rect 12299 12260 12532 12288
rect 12299 12257 12311 12260
rect 12253 12251 12311 12257
rect 12526 12248 12532 12260
rect 12584 12248 12590 12300
rect 14185 12291 14243 12297
rect 14185 12257 14197 12291
rect 14231 12288 14243 12291
rect 14274 12288 14280 12300
rect 14231 12260 14280 12288
rect 14231 12257 14243 12260
rect 14185 12251 14243 12257
rect 14274 12248 14280 12260
rect 14332 12288 14338 12300
rect 15013 12291 15071 12297
rect 15013 12288 15025 12291
rect 14332 12260 15025 12288
rect 14332 12248 14338 12260
rect 15013 12257 15025 12260
rect 15059 12257 15071 12291
rect 15013 12251 15071 12257
rect 15289 12291 15347 12297
rect 15289 12257 15301 12291
rect 15335 12257 15347 12291
rect 15289 12251 15347 12257
rect 15473 12291 15531 12297
rect 15473 12257 15485 12291
rect 15519 12288 15531 12291
rect 15654 12288 15660 12300
rect 15519 12260 15660 12288
rect 15519 12257 15531 12260
rect 15473 12251 15531 12257
rect 8481 12223 8539 12229
rect 8481 12220 8493 12223
rect 8260 12192 8493 12220
rect 8260 12180 8266 12192
rect 8481 12189 8493 12192
rect 8527 12220 8539 12223
rect 11057 12223 11115 12229
rect 11057 12220 11069 12223
rect 8527 12192 11069 12220
rect 8527 12189 8539 12192
rect 8481 12183 8539 12189
rect 11057 12189 11069 12192
rect 11103 12189 11115 12223
rect 11057 12183 11115 12189
rect 11882 12180 11888 12232
rect 11940 12220 11946 12232
rect 13173 12223 13231 12229
rect 13173 12220 13185 12223
rect 11940 12192 13185 12220
rect 11940 12180 11946 12192
rect 13173 12189 13185 12192
rect 13219 12189 13231 12223
rect 13173 12183 13231 12189
rect 13909 12223 13967 12229
rect 13909 12189 13921 12223
rect 13955 12220 13967 12223
rect 13955 12192 14044 12220
rect 13955 12189 13967 12192
rect 13909 12183 13967 12189
rect 2866 12152 2872 12164
rect 2779 12124 2872 12152
rect 2866 12112 2872 12124
rect 2924 12152 2930 12164
rect 9398 12152 9404 12164
rect 2924 12124 9404 12152
rect 2924 12112 2930 12124
rect 9398 12112 9404 12124
rect 9456 12112 9462 12164
rect 10854 12155 10912 12161
rect 10854 12121 10866 12155
rect 10900 12152 10912 12155
rect 12158 12152 12164 12164
rect 10900 12124 12164 12152
rect 10900 12121 10912 12124
rect 10854 12115 10912 12121
rect 12158 12112 12164 12124
rect 12216 12112 12222 12164
rect 6914 12084 6920 12096
rect 6875 12056 6920 12084
rect 6914 12044 6920 12056
rect 6972 12044 6978 12096
rect 7558 12044 7564 12096
rect 7616 12084 7622 12096
rect 7653 12087 7711 12093
rect 7653 12084 7665 12087
rect 7616 12056 7665 12084
rect 7616 12044 7622 12056
rect 7653 12053 7665 12056
rect 7699 12053 7711 12087
rect 10594 12084 10600 12096
rect 10555 12056 10600 12084
rect 7653 12047 7711 12053
rect 10594 12044 10600 12056
rect 10652 12044 10658 12096
rect 10962 12084 10968 12096
rect 10875 12056 10968 12084
rect 10962 12044 10968 12056
rect 11020 12084 11026 12096
rect 12710 12084 12716 12096
rect 11020 12056 12716 12084
rect 11020 12044 11026 12056
rect 12710 12044 12716 12056
rect 12768 12044 12774 12096
rect 12897 12087 12955 12093
rect 12897 12053 12909 12087
rect 12943 12084 12955 12087
rect 13078 12084 13084 12096
rect 12943 12056 13084 12084
rect 12943 12053 12955 12056
rect 12897 12047 12955 12053
rect 13078 12044 13084 12056
rect 13136 12044 13142 12096
rect 14016 12084 14044 12192
rect 14090 12180 14096 12232
rect 14148 12220 14154 12232
rect 14369 12223 14427 12229
rect 14369 12220 14381 12223
rect 14148 12192 14381 12220
rect 14148 12180 14154 12192
rect 14369 12189 14381 12192
rect 14415 12189 14427 12223
rect 14369 12183 14427 12189
rect 14384 12152 14412 12183
rect 14918 12180 14924 12232
rect 14976 12220 14982 12232
rect 15304 12220 15332 12251
rect 15654 12248 15660 12260
rect 15712 12288 15718 12300
rect 16206 12288 16212 12300
rect 15712 12260 16212 12288
rect 15712 12248 15718 12260
rect 16206 12248 16212 12260
rect 16264 12248 16270 12300
rect 16666 12288 16672 12300
rect 16627 12260 16672 12288
rect 16666 12248 16672 12260
rect 16724 12248 16730 12300
rect 16850 12288 16856 12300
rect 16811 12260 16856 12288
rect 16850 12248 16856 12260
rect 16908 12248 16914 12300
rect 16117 12223 16175 12229
rect 16117 12220 16129 12223
rect 14976 12192 16129 12220
rect 14976 12180 14982 12192
rect 16117 12189 16129 12192
rect 16163 12189 16175 12223
rect 16117 12183 16175 12189
rect 16577 12223 16635 12229
rect 16577 12189 16589 12223
rect 16623 12220 16635 12223
rect 17328 12220 17356 12316
rect 17681 12291 17739 12297
rect 17681 12257 17693 12291
rect 17727 12288 17739 12291
rect 18233 12291 18291 12297
rect 18233 12288 18245 12291
rect 17727 12260 18245 12288
rect 17727 12257 17739 12260
rect 17681 12251 17739 12257
rect 18233 12257 18245 12260
rect 18279 12257 18291 12291
rect 18233 12251 18291 12257
rect 18690 12248 18696 12300
rect 18748 12288 18754 12300
rect 18877 12291 18935 12297
rect 18877 12288 18889 12291
rect 18748 12260 18889 12288
rect 18748 12248 18754 12260
rect 18877 12257 18889 12260
rect 18923 12288 18935 12291
rect 19518 12288 19524 12300
rect 18923 12260 19524 12288
rect 18923 12257 18935 12260
rect 18877 12251 18935 12257
rect 19518 12248 19524 12260
rect 19576 12248 19582 12300
rect 20622 12288 20628 12300
rect 20583 12260 20628 12288
rect 20622 12248 20628 12260
rect 20680 12248 20686 12300
rect 16623 12192 17356 12220
rect 16623 12189 16635 12192
rect 16577 12183 16635 12189
rect 19150 12180 19156 12232
rect 19208 12220 19214 12232
rect 19245 12223 19303 12229
rect 19245 12220 19257 12223
rect 19208 12192 19257 12220
rect 19208 12180 19214 12192
rect 19245 12189 19257 12192
rect 19291 12189 19303 12223
rect 19245 12183 19303 12189
rect 14737 12155 14795 12161
rect 14737 12152 14749 12155
rect 14384 12124 14749 12152
rect 14737 12121 14749 12124
rect 14783 12152 14795 12155
rect 17957 12155 18015 12161
rect 17957 12152 17969 12155
rect 14783 12124 17969 12152
rect 14783 12121 14795 12124
rect 14737 12115 14795 12121
rect 17957 12121 17969 12124
rect 18003 12152 18015 12155
rect 18322 12152 18328 12164
rect 18003 12124 18328 12152
rect 18003 12121 18015 12124
rect 17957 12115 18015 12121
rect 18322 12112 18328 12124
rect 18380 12112 18386 12164
rect 18414 12112 18420 12164
rect 18472 12152 18478 12164
rect 18966 12152 18972 12164
rect 18472 12124 18972 12152
rect 18472 12112 18478 12124
rect 18966 12112 18972 12124
rect 19024 12161 19030 12164
rect 19024 12155 19073 12161
rect 19024 12121 19027 12155
rect 19061 12121 19073 12155
rect 19024 12115 19073 12121
rect 19024 12112 19030 12115
rect 19610 12112 19616 12164
rect 19668 12152 19674 12164
rect 20441 12155 20499 12161
rect 20441 12152 20453 12155
rect 19668 12124 20453 12152
rect 19668 12112 19674 12124
rect 20441 12121 20453 12124
rect 20487 12152 20499 12155
rect 20530 12152 20536 12164
rect 20487 12124 20536 12152
rect 20487 12121 20499 12124
rect 20441 12115 20499 12121
rect 20530 12112 20536 12124
rect 20588 12112 20594 12164
rect 20732 12152 20760 12328
rect 20898 12316 20904 12328
rect 20956 12316 20962 12368
rect 21008 12220 21036 12396
rect 21082 12384 21088 12436
rect 21140 12424 21146 12436
rect 24486 12424 24492 12436
rect 21140 12396 23060 12424
rect 24447 12396 24492 12424
rect 21140 12384 21146 12396
rect 22005 12359 22063 12365
rect 22005 12325 22017 12359
rect 22051 12356 22063 12359
rect 22189 12359 22247 12365
rect 22189 12356 22201 12359
rect 22051 12328 22201 12356
rect 22051 12325 22063 12328
rect 22005 12319 22063 12325
rect 22189 12325 22201 12328
rect 22235 12325 22247 12359
rect 22189 12319 22247 12325
rect 21361 12291 21419 12297
rect 21361 12257 21373 12291
rect 21407 12288 21419 12291
rect 21450 12288 21456 12300
rect 21407 12260 21456 12288
rect 21407 12257 21419 12260
rect 21361 12251 21419 12257
rect 21450 12248 21456 12260
rect 21508 12248 21514 12300
rect 21726 12288 21732 12300
rect 21687 12260 21732 12288
rect 21726 12248 21732 12260
rect 21784 12248 21790 12300
rect 21821 12291 21879 12297
rect 21821 12257 21833 12291
rect 21867 12288 21879 12291
rect 22094 12288 22100 12300
rect 21867 12260 22100 12288
rect 21867 12257 21879 12260
rect 21821 12251 21879 12257
rect 22094 12248 22100 12260
rect 22152 12248 22158 12300
rect 22922 12288 22928 12300
rect 22204 12260 22928 12288
rect 22204 12220 22232 12260
rect 22922 12248 22928 12260
rect 22980 12248 22986 12300
rect 23032 12297 23060 12396
rect 24486 12384 24492 12396
rect 24544 12384 24550 12436
rect 24854 12384 24860 12436
rect 24912 12424 24918 12436
rect 24949 12427 25007 12433
rect 24949 12424 24961 12427
rect 24912 12396 24961 12424
rect 24912 12384 24918 12396
rect 24949 12393 24961 12396
rect 24995 12393 25007 12427
rect 24949 12387 25007 12393
rect 25774 12384 25780 12436
rect 25832 12424 25838 12436
rect 26050 12424 26056 12436
rect 25832 12396 26056 12424
rect 25832 12384 25838 12396
rect 26050 12384 26056 12396
rect 26108 12384 26114 12436
rect 26234 12424 26240 12436
rect 26195 12396 26240 12424
rect 26234 12384 26240 12396
rect 26292 12384 26298 12436
rect 27706 12424 27712 12436
rect 27667 12396 27712 12424
rect 27706 12384 27712 12396
rect 27764 12384 27770 12436
rect 27985 12427 28043 12433
rect 27985 12393 27997 12427
rect 28031 12424 28043 12427
rect 33134 12424 33140 12436
rect 28031 12396 33140 12424
rect 28031 12393 28043 12396
rect 27985 12387 28043 12393
rect 33134 12384 33140 12396
rect 33192 12384 33198 12436
rect 33229 12427 33287 12433
rect 33229 12393 33241 12427
rect 33275 12424 33287 12427
rect 33318 12424 33324 12436
rect 33275 12396 33324 12424
rect 33275 12393 33287 12396
rect 33229 12387 33287 12393
rect 33318 12384 33324 12396
rect 33376 12384 33382 12436
rect 33502 12424 33508 12436
rect 33463 12396 33508 12424
rect 33502 12384 33508 12396
rect 33560 12384 33566 12436
rect 35250 12424 35256 12436
rect 35211 12396 35256 12424
rect 35250 12384 35256 12396
rect 35308 12384 35314 12436
rect 36262 12384 36268 12436
rect 36320 12424 36326 12436
rect 36357 12427 36415 12433
rect 36357 12424 36369 12427
rect 36320 12396 36369 12424
rect 36320 12384 36326 12396
rect 36357 12393 36369 12396
rect 36403 12393 36415 12427
rect 37182 12424 37188 12436
rect 37143 12396 37188 12424
rect 36357 12387 36415 12393
rect 37182 12384 37188 12396
rect 37240 12384 37246 12436
rect 39574 12384 39580 12436
rect 39632 12424 39638 12436
rect 40221 12427 40279 12433
rect 40221 12424 40233 12427
rect 39632 12396 40233 12424
rect 39632 12384 39638 12396
rect 40221 12393 40233 12396
rect 40267 12393 40279 12427
rect 40678 12424 40684 12436
rect 40639 12396 40684 12424
rect 40221 12387 40279 12393
rect 40678 12384 40684 12396
rect 40736 12384 40742 12436
rect 41601 12427 41659 12433
rect 41601 12393 41613 12427
rect 41647 12424 41659 12427
rect 41782 12424 41788 12436
rect 41647 12396 41788 12424
rect 41647 12393 41659 12396
rect 41601 12387 41659 12393
rect 41782 12384 41788 12396
rect 41840 12384 41846 12436
rect 43070 12424 43076 12436
rect 43031 12396 43076 12424
rect 43070 12384 43076 12396
rect 43128 12384 43134 12436
rect 52546 12424 52552 12436
rect 48700 12396 52552 12424
rect 23106 12316 23112 12368
rect 23164 12356 23170 12368
rect 23477 12359 23535 12365
rect 23477 12356 23489 12359
rect 23164 12328 23489 12356
rect 23164 12316 23170 12328
rect 23477 12325 23489 12328
rect 23523 12325 23535 12359
rect 23477 12319 23535 12325
rect 23934 12316 23940 12368
rect 23992 12356 23998 12368
rect 31481 12359 31539 12365
rect 31481 12356 31493 12359
rect 23992 12328 31493 12356
rect 23992 12316 23998 12328
rect 31481 12325 31493 12328
rect 31527 12356 31539 12359
rect 31665 12359 31723 12365
rect 31665 12356 31677 12359
rect 31527 12328 31677 12356
rect 31527 12325 31539 12328
rect 31481 12319 31539 12325
rect 31665 12325 31677 12328
rect 31711 12325 31723 12359
rect 31665 12319 31723 12325
rect 32490 12316 32496 12368
rect 32548 12356 32554 12368
rect 33689 12359 33747 12365
rect 33689 12356 33701 12359
rect 32548 12328 33701 12356
rect 32548 12316 32554 12328
rect 33689 12325 33701 12328
rect 33735 12325 33747 12359
rect 34146 12356 34152 12368
rect 33689 12319 33747 12325
rect 33796 12328 34152 12356
rect 23017 12291 23075 12297
rect 23017 12257 23029 12291
rect 23063 12288 23075 12291
rect 23842 12288 23848 12300
rect 23063 12260 23848 12288
rect 23063 12257 23075 12260
rect 23017 12251 23075 12257
rect 23842 12248 23848 12260
rect 23900 12248 23906 12300
rect 24946 12288 24952 12300
rect 24907 12260 24952 12288
rect 24946 12248 24952 12260
rect 25004 12248 25010 12300
rect 25314 12288 25320 12300
rect 25275 12260 25320 12288
rect 25314 12248 25320 12260
rect 25372 12248 25378 12300
rect 26234 12248 26240 12300
rect 26292 12288 26298 12300
rect 26682 12291 26740 12297
rect 26682 12288 26694 12291
rect 26292 12260 26694 12288
rect 26292 12248 26298 12260
rect 26682 12257 26694 12260
rect 26728 12257 26740 12291
rect 26682 12251 26740 12257
rect 26786 12248 26792 12300
rect 26844 12288 26850 12300
rect 27246 12288 27252 12300
rect 26844 12260 26889 12288
rect 27207 12260 27252 12288
rect 26844 12248 26850 12260
rect 27246 12248 27252 12260
rect 27304 12248 27310 12300
rect 27338 12248 27344 12300
rect 27396 12288 27402 12300
rect 27433 12291 27491 12297
rect 27433 12288 27445 12291
rect 27396 12260 27445 12288
rect 27396 12248 27402 12260
rect 27433 12257 27445 12260
rect 27479 12257 27491 12291
rect 27433 12251 27491 12257
rect 28534 12248 28540 12300
rect 28592 12288 28598 12300
rect 28721 12291 28779 12297
rect 28721 12288 28733 12291
rect 28592 12260 28733 12288
rect 28592 12248 28598 12260
rect 28721 12257 28733 12260
rect 28767 12257 28779 12291
rect 28721 12251 28779 12257
rect 28813 12291 28871 12297
rect 28813 12257 28825 12291
rect 28859 12288 28871 12291
rect 29549 12291 29607 12297
rect 29549 12288 29561 12291
rect 28859 12260 29561 12288
rect 28859 12257 28871 12260
rect 28813 12251 28871 12257
rect 29549 12257 29561 12260
rect 29595 12257 29607 12291
rect 30098 12288 30104 12300
rect 30059 12260 30104 12288
rect 29549 12251 29607 12257
rect 21008 12192 22232 12220
rect 22554 12180 22560 12232
rect 22612 12220 22618 12232
rect 22741 12223 22799 12229
rect 22741 12220 22753 12223
rect 22612 12192 22753 12220
rect 22612 12180 22618 12192
rect 22741 12189 22753 12192
rect 22787 12220 22799 12223
rect 23290 12220 23296 12232
rect 22787 12192 23296 12220
rect 22787 12189 22799 12192
rect 22741 12183 22799 12189
rect 23290 12180 23296 12192
rect 23348 12180 23354 12232
rect 28828 12220 28856 12251
rect 30098 12248 30104 12260
rect 30156 12288 30162 12300
rect 30282 12288 30288 12300
rect 30156 12260 30288 12288
rect 30156 12248 30162 12260
rect 30282 12248 30288 12260
rect 30340 12288 30346 12300
rect 30653 12291 30711 12297
rect 30653 12288 30665 12291
rect 30340 12260 30665 12288
rect 30340 12248 30346 12260
rect 30653 12257 30665 12260
rect 30699 12257 30711 12291
rect 30653 12251 30711 12257
rect 31757 12291 31815 12297
rect 31757 12257 31769 12291
rect 31803 12288 31815 12291
rect 32309 12291 32367 12297
rect 32309 12288 32321 12291
rect 31803 12260 32321 12288
rect 31803 12257 31815 12260
rect 31757 12251 31815 12257
rect 32309 12257 32321 12260
rect 32355 12257 32367 12291
rect 32309 12251 32367 12257
rect 32401 12291 32459 12297
rect 32401 12257 32413 12291
rect 32447 12288 32459 12291
rect 32582 12288 32588 12300
rect 32447 12260 32588 12288
rect 32447 12257 32459 12260
rect 32401 12251 32459 12257
rect 32582 12248 32588 12260
rect 32640 12248 32646 12300
rect 33796 12288 33824 12328
rect 34146 12316 34152 12328
rect 34204 12316 34210 12368
rect 32784 12260 33824 12288
rect 27632 12192 28856 12220
rect 23106 12152 23112 12164
rect 20732 12124 23112 12152
rect 23106 12112 23112 12124
rect 23164 12112 23170 12164
rect 24210 12112 24216 12164
rect 24268 12152 24274 12164
rect 24268 12124 26004 12152
rect 24268 12112 24274 12124
rect 14458 12084 14464 12096
rect 14016 12056 14464 12084
rect 14458 12044 14464 12056
rect 14516 12084 14522 12096
rect 17310 12084 17316 12096
rect 14516 12056 17316 12084
rect 14516 12044 14522 12056
rect 17310 12044 17316 12056
rect 17368 12044 17374 12096
rect 17494 12084 17500 12096
rect 17455 12056 17500 12084
rect 17494 12044 17500 12056
rect 17552 12044 17558 12096
rect 17678 12044 17684 12096
rect 17736 12084 17742 12096
rect 18785 12087 18843 12093
rect 18785 12084 18797 12087
rect 17736 12056 18797 12084
rect 17736 12044 17742 12056
rect 18785 12053 18797 12056
rect 18831 12084 18843 12087
rect 19153 12087 19211 12093
rect 19153 12084 19165 12087
rect 18831 12056 19165 12084
rect 18831 12053 18843 12056
rect 18785 12047 18843 12053
rect 19153 12053 19165 12056
rect 19199 12084 19211 12087
rect 19518 12084 19524 12096
rect 19199 12056 19524 12084
rect 19199 12053 19211 12056
rect 19153 12047 19211 12053
rect 19518 12044 19524 12056
rect 19576 12044 19582 12096
rect 19794 12044 19800 12096
rect 19852 12084 19858 12096
rect 19981 12087 20039 12093
rect 19981 12084 19993 12087
rect 19852 12056 19993 12084
rect 19852 12044 19858 12056
rect 19981 12053 19993 12056
rect 20027 12053 20039 12087
rect 19981 12047 20039 12053
rect 21450 12044 21456 12096
rect 21508 12084 21514 12096
rect 22005 12087 22063 12093
rect 22005 12084 22017 12087
rect 21508 12056 22017 12084
rect 21508 12044 21514 12056
rect 22005 12053 22017 12056
rect 22051 12053 22063 12087
rect 22005 12047 22063 12053
rect 22186 12044 22192 12096
rect 22244 12084 22250 12096
rect 22557 12087 22615 12093
rect 22557 12084 22569 12087
rect 22244 12056 22569 12084
rect 22244 12044 22250 12056
rect 22557 12053 22569 12056
rect 22603 12084 22615 12087
rect 23753 12087 23811 12093
rect 23753 12084 23765 12087
rect 22603 12056 23765 12084
rect 22603 12053 22615 12056
rect 22557 12047 22615 12053
rect 23753 12053 23765 12056
rect 23799 12053 23811 12087
rect 24118 12084 24124 12096
rect 24079 12056 24124 12084
rect 23753 12047 23811 12053
rect 24118 12044 24124 12056
rect 24176 12044 24182 12096
rect 25774 12044 25780 12096
rect 25832 12084 25838 12096
rect 25869 12087 25927 12093
rect 25869 12084 25881 12087
rect 25832 12056 25881 12084
rect 25832 12044 25838 12056
rect 25869 12053 25881 12056
rect 25915 12053 25927 12087
rect 25976 12084 26004 12124
rect 27154 12112 27160 12164
rect 27212 12152 27218 12164
rect 27632 12152 27660 12192
rect 28902 12180 28908 12232
rect 28960 12220 28966 12232
rect 31205 12223 31263 12229
rect 28960 12192 30328 12220
rect 28960 12180 28966 12192
rect 27212 12124 27660 12152
rect 27212 12112 27218 12124
rect 27706 12112 27712 12164
rect 27764 12152 27770 12164
rect 28261 12155 28319 12161
rect 27764 12124 28212 12152
rect 27764 12112 27770 12124
rect 27985 12087 28043 12093
rect 27985 12084 27997 12087
rect 25976 12056 27997 12084
rect 25869 12047 25927 12053
rect 27985 12053 27997 12056
rect 28031 12053 28043 12087
rect 28184 12084 28212 12124
rect 28261 12121 28273 12155
rect 28307 12152 28319 12155
rect 29178 12152 29184 12164
rect 28307 12124 29184 12152
rect 28307 12121 28319 12124
rect 28261 12115 28319 12121
rect 29178 12112 29184 12124
rect 29236 12112 29242 12164
rect 29454 12112 29460 12164
rect 29512 12152 29518 12164
rect 30300 12161 30328 12192
rect 31205 12189 31217 12223
rect 31251 12220 31263 12223
rect 31941 12223 31999 12229
rect 31251 12192 31892 12220
rect 31251 12189 31263 12192
rect 31205 12183 31263 12189
rect 29917 12155 29975 12161
rect 29917 12152 29929 12155
rect 29512 12124 29929 12152
rect 29512 12112 29518 12124
rect 29917 12121 29929 12124
rect 29963 12121 29975 12155
rect 29917 12115 29975 12121
rect 30285 12155 30343 12161
rect 30285 12121 30297 12155
rect 30331 12152 30343 12155
rect 31570 12152 31576 12164
rect 30331 12124 31576 12152
rect 30331 12121 30343 12124
rect 30285 12115 30343 12121
rect 31570 12112 31576 12124
rect 31628 12112 31634 12164
rect 28537 12087 28595 12093
rect 28537 12084 28549 12087
rect 28184 12056 28549 12084
rect 27985 12047 28043 12053
rect 28537 12053 28549 12056
rect 28583 12053 28595 12087
rect 28994 12084 29000 12096
rect 28955 12056 29000 12084
rect 28537 12047 28595 12053
rect 28994 12044 29000 12056
rect 29052 12044 29058 12096
rect 31864 12084 31892 12192
rect 31941 12189 31953 12223
rect 31987 12220 31999 12223
rect 32784 12220 32812 12260
rect 33962 12248 33968 12300
rect 34020 12288 34026 12300
rect 34330 12288 34336 12300
rect 34020 12260 34336 12288
rect 34020 12248 34026 12260
rect 34330 12248 34336 12260
rect 34388 12248 34394 12300
rect 34514 12248 34520 12300
rect 34572 12288 34578 12300
rect 34701 12291 34759 12297
rect 34701 12288 34713 12291
rect 34572 12260 34713 12288
rect 34572 12248 34578 12260
rect 34701 12257 34713 12260
rect 34747 12257 34759 12291
rect 34701 12251 34759 12257
rect 34885 12291 34943 12297
rect 34885 12257 34897 12291
rect 34931 12288 34943 12291
rect 35268 12288 35296 12384
rect 37734 12356 37740 12368
rect 37695 12328 37740 12356
rect 37734 12316 37740 12328
rect 37792 12316 37798 12368
rect 37826 12316 37832 12368
rect 37884 12356 37890 12368
rect 39758 12356 39764 12368
rect 37884 12328 38792 12356
rect 39671 12328 39764 12356
rect 37884 12316 37890 12328
rect 35710 12288 35716 12300
rect 34931 12260 35296 12288
rect 35671 12260 35716 12288
rect 34931 12257 34943 12260
rect 34885 12251 34943 12257
rect 35710 12248 35716 12260
rect 35768 12248 35774 12300
rect 38764 12297 38792 12328
rect 39684 12297 39712 12328
rect 39758 12316 39764 12328
rect 39816 12356 39822 12368
rect 46106 12356 46112 12368
rect 39816 12328 42012 12356
rect 46067 12328 46112 12356
rect 39816 12316 39822 12328
rect 38565 12291 38623 12297
rect 38565 12257 38577 12291
rect 38611 12257 38623 12291
rect 38565 12251 38623 12257
rect 38749 12291 38807 12297
rect 38749 12257 38761 12291
rect 38795 12288 38807 12291
rect 39025 12291 39083 12297
rect 39025 12288 39037 12291
rect 38795 12260 39037 12288
rect 38795 12257 38807 12260
rect 38749 12251 38807 12257
rect 39025 12257 39037 12260
rect 39071 12257 39083 12291
rect 39025 12251 39083 12257
rect 39669 12291 39727 12297
rect 39669 12257 39681 12291
rect 39715 12257 39727 12291
rect 39669 12251 39727 12257
rect 31987 12192 32812 12220
rect 32861 12223 32919 12229
rect 31987 12189 31999 12192
rect 31941 12183 31999 12189
rect 32861 12189 32873 12223
rect 32907 12189 32919 12223
rect 32861 12183 32919 12189
rect 32876 12152 32904 12183
rect 33686 12180 33692 12232
rect 33744 12220 33750 12232
rect 34241 12223 34299 12229
rect 34241 12220 34253 12223
rect 33744 12192 34253 12220
rect 33744 12180 33750 12192
rect 34241 12189 34253 12192
rect 34287 12189 34299 12223
rect 34241 12183 34299 12189
rect 34790 12180 34796 12232
rect 34848 12220 34854 12232
rect 34848 12192 36032 12220
rect 34848 12180 34854 12192
rect 35526 12152 35532 12164
rect 32876 12124 35532 12152
rect 35526 12112 35532 12124
rect 35584 12152 35590 12164
rect 35851 12155 35909 12161
rect 35851 12152 35863 12155
rect 35584 12124 35863 12152
rect 35584 12112 35590 12124
rect 35851 12121 35863 12124
rect 35897 12121 35909 12155
rect 36004 12152 36032 12192
rect 36078 12180 36084 12232
rect 36136 12220 36142 12232
rect 36814 12220 36820 12232
rect 36136 12192 36820 12220
rect 36136 12180 36142 12192
rect 36814 12180 36820 12192
rect 36872 12180 36878 12232
rect 38286 12220 38292 12232
rect 38247 12192 38292 12220
rect 38286 12180 38292 12192
rect 38344 12180 38350 12232
rect 38580 12220 38608 12251
rect 39942 12248 39948 12300
rect 40000 12288 40006 12300
rect 40773 12291 40831 12297
rect 40773 12288 40785 12291
rect 40000 12260 40785 12288
rect 40000 12248 40006 12260
rect 40773 12257 40785 12260
rect 40819 12257 40831 12291
rect 40773 12251 40831 12257
rect 40920 12291 40978 12297
rect 40920 12257 40932 12291
rect 40966 12288 40978 12291
rect 41874 12288 41880 12300
rect 40966 12260 41880 12288
rect 40966 12257 40978 12260
rect 40920 12251 40978 12257
rect 41874 12248 41880 12260
rect 41932 12248 41938 12300
rect 39850 12220 39856 12232
rect 38580 12192 39856 12220
rect 39850 12180 39856 12192
rect 39908 12180 39914 12232
rect 41141 12223 41199 12229
rect 41141 12189 41153 12223
rect 41187 12220 41199 12223
rect 41506 12220 41512 12232
rect 41187 12192 41512 12220
rect 41187 12189 41199 12192
rect 41141 12183 41199 12189
rect 41506 12180 41512 12192
rect 41564 12180 41570 12232
rect 37826 12152 37832 12164
rect 36004 12124 37832 12152
rect 35851 12115 35909 12121
rect 37826 12112 37832 12124
rect 37884 12112 37890 12164
rect 39577 12155 39635 12161
rect 39577 12121 39589 12155
rect 39623 12152 39635 12155
rect 39666 12152 39672 12164
rect 39623 12124 39672 12152
rect 39623 12121 39635 12124
rect 39577 12115 39635 12121
rect 39666 12112 39672 12124
rect 39724 12152 39730 12164
rect 41233 12155 41291 12161
rect 41233 12152 41245 12155
rect 39724 12124 41245 12152
rect 39724 12112 39730 12124
rect 41233 12121 41245 12124
rect 41279 12121 41291 12155
rect 41984 12152 42012 12328
rect 46106 12316 46112 12328
rect 46164 12316 46170 12368
rect 46293 12359 46351 12365
rect 46293 12325 46305 12359
rect 46339 12356 46351 12359
rect 48700 12356 48728 12396
rect 52546 12384 52552 12396
rect 52604 12384 52610 12436
rect 57072 12396 58388 12424
rect 46339 12328 48728 12356
rect 48777 12359 48835 12365
rect 46339 12325 46351 12328
rect 46293 12319 46351 12325
rect 48777 12325 48789 12359
rect 48823 12356 48835 12359
rect 49234 12356 49240 12368
rect 48823 12328 49240 12356
rect 48823 12325 48835 12328
rect 48777 12319 48835 12325
rect 49234 12316 49240 12328
rect 49292 12316 49298 12368
rect 50246 12316 50252 12368
rect 50304 12356 50310 12368
rect 50341 12359 50399 12365
rect 50341 12356 50353 12359
rect 50304 12328 50353 12356
rect 50304 12316 50310 12328
rect 50341 12325 50353 12328
rect 50387 12325 50399 12359
rect 50341 12319 50399 12325
rect 54849 12359 54907 12365
rect 54849 12325 54861 12359
rect 54895 12356 54907 12359
rect 55398 12356 55404 12368
rect 54895 12328 55404 12356
rect 54895 12325 54907 12328
rect 54849 12319 54907 12325
rect 55398 12316 55404 12328
rect 55456 12316 55462 12368
rect 55858 12356 55864 12368
rect 55819 12328 55864 12356
rect 55858 12316 55864 12328
rect 55916 12316 55922 12368
rect 42978 12248 42984 12300
rect 43036 12288 43042 12300
rect 43533 12291 43591 12297
rect 43533 12288 43545 12291
rect 43036 12260 43545 12288
rect 43036 12248 43042 12260
rect 43533 12257 43545 12260
rect 43579 12257 43591 12291
rect 43533 12251 43591 12257
rect 44085 12291 44143 12297
rect 44085 12257 44097 12291
rect 44131 12288 44143 12291
rect 44266 12288 44272 12300
rect 44131 12260 44272 12288
rect 44131 12257 44143 12260
rect 44085 12251 44143 12257
rect 42150 12180 42156 12232
rect 42208 12220 42214 12232
rect 42245 12223 42303 12229
rect 42245 12220 42257 12223
rect 42208 12192 42257 12220
rect 42208 12180 42214 12192
rect 42245 12189 42257 12192
rect 42291 12220 42303 12223
rect 43438 12220 43444 12232
rect 42291 12192 43444 12220
rect 42291 12189 42303 12192
rect 42245 12183 42303 12189
rect 43438 12180 43444 12192
rect 43496 12180 43502 12232
rect 43548 12220 43576 12251
rect 44266 12248 44272 12260
rect 44324 12288 44330 12300
rect 44910 12288 44916 12300
rect 44324 12260 44916 12288
rect 44324 12248 44330 12260
rect 44910 12248 44916 12260
rect 44968 12288 44974 12300
rect 46753 12291 46811 12297
rect 44968 12260 45600 12288
rect 44968 12248 44974 12260
rect 44174 12220 44180 12232
rect 43548 12192 44180 12220
rect 44174 12180 44180 12192
rect 44232 12180 44238 12232
rect 44450 12220 44456 12232
rect 44411 12192 44456 12220
rect 44450 12180 44456 12192
rect 44508 12180 44514 12232
rect 45572 12229 45600 12260
rect 46753 12257 46765 12291
rect 46799 12288 46811 12291
rect 46842 12288 46848 12300
rect 46799 12260 46848 12288
rect 46799 12257 46811 12260
rect 46753 12251 46811 12257
rect 46842 12248 46848 12260
rect 46900 12288 46906 12300
rect 47026 12288 47032 12300
rect 46900 12260 47032 12288
rect 46900 12248 46906 12260
rect 47026 12248 47032 12260
rect 47084 12248 47090 12300
rect 48041 12291 48099 12297
rect 48041 12257 48053 12291
rect 48087 12288 48099 12291
rect 48314 12288 48320 12300
rect 48087 12260 48320 12288
rect 48087 12257 48099 12260
rect 48041 12251 48099 12257
rect 48314 12248 48320 12260
rect 48372 12288 48378 12300
rect 48866 12288 48872 12300
rect 48372 12260 48872 12288
rect 48372 12248 48378 12260
rect 48866 12248 48872 12260
rect 48924 12248 48930 12300
rect 49050 12288 49056 12300
rect 49011 12260 49056 12288
rect 49050 12248 49056 12260
rect 49108 12248 49114 12300
rect 50706 12288 50712 12300
rect 50667 12260 50712 12288
rect 50706 12248 50712 12260
rect 50764 12248 50770 12300
rect 51442 12248 51448 12300
rect 51500 12288 51506 12300
rect 51537 12291 51595 12297
rect 51537 12288 51549 12291
rect 51500 12260 51549 12288
rect 51500 12248 51506 12260
rect 51537 12257 51549 12260
rect 51583 12257 51595 12291
rect 51537 12251 51595 12257
rect 52822 12248 52828 12300
rect 52880 12288 52886 12300
rect 53193 12291 53251 12297
rect 53193 12288 53205 12291
rect 52880 12260 53205 12288
rect 52880 12248 52886 12260
rect 53193 12257 53205 12260
rect 53239 12288 53251 12291
rect 53466 12288 53472 12300
rect 53239 12260 53472 12288
rect 53239 12257 53251 12260
rect 53193 12251 53251 12257
rect 53466 12248 53472 12260
rect 53524 12248 53530 12300
rect 54389 12291 54447 12297
rect 54389 12257 54401 12291
rect 54435 12288 54447 12291
rect 55122 12288 55128 12300
rect 54435 12260 55128 12288
rect 54435 12257 54447 12260
rect 54389 12251 54447 12257
rect 55122 12248 55128 12260
rect 55180 12248 55186 12300
rect 56870 12248 56876 12300
rect 56928 12288 56934 12300
rect 57072 12297 57100 12396
rect 58066 12356 58072 12368
rect 57808 12328 58072 12356
rect 57808 12297 57836 12328
rect 58066 12316 58072 12328
rect 58124 12316 58130 12368
rect 58360 12356 58388 12396
rect 58434 12384 58440 12436
rect 58492 12424 58498 12436
rect 58805 12427 58863 12433
rect 58805 12424 58817 12427
rect 58492 12396 58817 12424
rect 58492 12384 58498 12396
rect 58805 12393 58817 12396
rect 58851 12393 58863 12427
rect 58805 12387 58863 12393
rect 59998 12356 60004 12368
rect 58360 12328 60004 12356
rect 59998 12316 60004 12328
rect 60056 12356 60062 12368
rect 61013 12359 61071 12365
rect 61013 12356 61025 12359
rect 60056 12328 61025 12356
rect 60056 12316 60062 12328
rect 60200 12297 60228 12328
rect 61013 12325 61025 12328
rect 61059 12325 61071 12359
rect 61013 12319 61071 12325
rect 57057 12291 57115 12297
rect 57057 12288 57069 12291
rect 56928 12260 57069 12288
rect 56928 12248 56934 12260
rect 57057 12257 57069 12260
rect 57103 12257 57115 12291
rect 57057 12251 57115 12257
rect 57793 12291 57851 12297
rect 57793 12257 57805 12291
rect 57839 12257 57851 12291
rect 57793 12251 57851 12257
rect 60185 12291 60243 12297
rect 60185 12257 60197 12291
rect 60231 12257 60243 12291
rect 60185 12251 60243 12257
rect 60277 12291 60335 12297
rect 60277 12257 60289 12291
rect 60323 12288 60335 12291
rect 60550 12288 60556 12300
rect 60323 12260 60556 12288
rect 60323 12257 60335 12260
rect 60277 12251 60335 12257
rect 60550 12248 60556 12260
rect 60608 12248 60614 12300
rect 45557 12223 45615 12229
rect 45557 12189 45569 12223
rect 45603 12220 45615 12223
rect 46477 12223 46535 12229
rect 46477 12220 46489 12223
rect 45603 12192 46489 12220
rect 45603 12189 45615 12192
rect 45557 12183 45615 12189
rect 46477 12189 46489 12192
rect 46523 12220 46535 12223
rect 46566 12220 46572 12232
rect 46523 12192 46572 12220
rect 46523 12189 46535 12192
rect 46477 12183 46535 12189
rect 46566 12180 46572 12192
rect 46624 12180 46630 12232
rect 46658 12180 46664 12232
rect 46716 12220 46722 12232
rect 46716 12192 46761 12220
rect 46716 12180 46722 12192
rect 46934 12180 46940 12232
rect 46992 12220 46998 12232
rect 47213 12223 47271 12229
rect 47213 12220 47225 12223
rect 46992 12192 47225 12220
rect 46992 12180 46998 12192
rect 47213 12189 47225 12192
rect 47259 12220 47271 12223
rect 47489 12223 47547 12229
rect 47489 12220 47501 12223
rect 47259 12192 47501 12220
rect 47259 12189 47271 12192
rect 47213 12183 47271 12189
rect 47489 12189 47501 12192
rect 47535 12189 47547 12223
rect 48958 12220 48964 12232
rect 48919 12192 48964 12220
rect 47489 12183 47547 12189
rect 48958 12180 48964 12192
rect 49016 12180 49022 12232
rect 51258 12220 51264 12232
rect 51219 12192 51264 12220
rect 51258 12180 51264 12192
rect 51316 12180 51322 12232
rect 51718 12220 51724 12232
rect 51679 12192 51724 12220
rect 51718 12180 51724 12192
rect 51776 12180 51782 12232
rect 53101 12223 53159 12229
rect 53101 12189 53113 12223
rect 53147 12220 53159 12223
rect 53282 12220 53288 12232
rect 53147 12192 53288 12220
rect 53147 12189 53159 12192
rect 53101 12183 53159 12189
rect 53282 12180 53288 12192
rect 53340 12180 53346 12232
rect 53653 12223 53711 12229
rect 53653 12189 53665 12223
rect 53699 12220 53711 12223
rect 54110 12220 54116 12232
rect 53699 12192 54116 12220
rect 53699 12189 53711 12192
rect 53653 12183 53711 12189
rect 54110 12180 54116 12192
rect 54168 12180 54174 12232
rect 55490 12220 55496 12232
rect 55451 12192 55496 12220
rect 55490 12180 55496 12192
rect 55548 12180 55554 12232
rect 57882 12180 57888 12232
rect 57940 12220 57946 12232
rect 58069 12223 58127 12229
rect 58069 12220 58081 12223
rect 57940 12192 58081 12220
rect 57940 12180 57946 12192
rect 58069 12189 58081 12192
rect 58115 12220 58127 12223
rect 58437 12223 58495 12229
rect 58437 12220 58449 12223
rect 58115 12192 58449 12220
rect 58115 12189 58127 12192
rect 58069 12183 58127 12189
rect 58437 12189 58449 12192
rect 58483 12189 58495 12223
rect 58437 12183 58495 12189
rect 41984 12124 42656 12152
rect 41233 12115 41291 12121
rect 34790 12084 34796 12096
rect 31864 12056 34796 12084
rect 34790 12044 34796 12056
rect 34848 12044 34854 12096
rect 35618 12084 35624 12096
rect 35579 12056 35624 12084
rect 35618 12044 35624 12056
rect 35676 12044 35682 12096
rect 35989 12087 36047 12093
rect 35989 12053 36001 12087
rect 36035 12084 36047 12087
rect 36446 12084 36452 12096
rect 36035 12056 36452 12084
rect 36035 12053 36047 12056
rect 35989 12047 36047 12053
rect 36446 12044 36452 12056
rect 36504 12044 36510 12096
rect 36814 12084 36820 12096
rect 36775 12056 36820 12084
rect 36814 12044 36820 12056
rect 36872 12044 36878 12096
rect 39853 12087 39911 12093
rect 39853 12053 39865 12087
rect 39899 12084 39911 12087
rect 40862 12084 40868 12096
rect 39899 12056 40868 12084
rect 39899 12053 39911 12056
rect 39853 12047 39911 12053
rect 40862 12044 40868 12056
rect 40920 12084 40926 12096
rect 41049 12087 41107 12093
rect 41049 12084 41061 12087
rect 40920 12056 41061 12084
rect 40920 12044 40926 12056
rect 41049 12053 41061 12056
rect 41095 12084 41107 12087
rect 41601 12087 41659 12093
rect 41601 12084 41613 12087
rect 41095 12056 41613 12084
rect 41095 12053 41107 12056
rect 41049 12047 41107 12053
rect 41601 12053 41613 12056
rect 41647 12053 41659 12087
rect 41601 12047 41659 12053
rect 41782 12044 41788 12096
rect 41840 12084 41846 12096
rect 42521 12087 42579 12093
rect 42521 12084 42533 12087
rect 41840 12056 42533 12084
rect 41840 12044 41846 12056
rect 42521 12053 42533 12056
rect 42567 12053 42579 12087
rect 42628 12084 42656 12124
rect 47026 12112 47032 12164
rect 47084 12152 47090 12164
rect 49050 12152 49056 12164
rect 47084 12124 49056 12152
rect 47084 12112 47090 12124
rect 49050 12112 49056 12124
rect 49108 12112 49114 12164
rect 50246 12112 50252 12164
rect 50304 12152 50310 12164
rect 51276 12152 51304 12180
rect 51626 12152 51632 12164
rect 50304 12124 51212 12152
rect 51276 12124 51632 12152
rect 50304 12112 50310 12124
rect 46293 12087 46351 12093
rect 46293 12084 46305 12087
rect 42628 12056 46305 12084
rect 42521 12047 42579 12053
rect 46293 12053 46305 12056
rect 46339 12053 46351 12087
rect 46293 12047 46351 12053
rect 48409 12087 48467 12093
rect 48409 12053 48421 12087
rect 48455 12084 48467 12087
rect 48498 12084 48504 12096
rect 48455 12056 48504 12084
rect 48455 12053 48467 12056
rect 48409 12047 48467 12053
rect 48498 12044 48504 12056
rect 48556 12084 48562 12096
rect 49237 12087 49295 12093
rect 49237 12084 49249 12087
rect 48556 12056 49249 12084
rect 48556 12044 48562 12056
rect 49237 12053 49249 12056
rect 49283 12053 49295 12087
rect 50062 12084 50068 12096
rect 49975 12056 50068 12084
rect 49237 12047 49295 12053
rect 50062 12044 50068 12056
rect 50120 12084 50126 12096
rect 50522 12084 50528 12096
rect 50120 12056 50528 12084
rect 50120 12044 50126 12056
rect 50522 12044 50528 12056
rect 50580 12044 50586 12096
rect 50614 12044 50620 12096
rect 50672 12084 50678 12096
rect 51074 12084 51080 12096
rect 50672 12056 51080 12084
rect 50672 12044 50678 12056
rect 51074 12044 51080 12056
rect 51132 12044 51138 12096
rect 51184 12084 51212 12124
rect 51626 12112 51632 12124
rect 51684 12112 51690 12164
rect 51902 12112 51908 12164
rect 51960 12152 51966 12164
rect 52270 12152 52276 12164
rect 51960 12124 52276 12152
rect 51960 12112 51966 12124
rect 52270 12112 52276 12124
rect 52328 12152 52334 12164
rect 52733 12155 52791 12161
rect 52733 12152 52745 12155
rect 52328 12124 52745 12152
rect 52328 12112 52334 12124
rect 52733 12121 52745 12124
rect 52779 12121 52791 12155
rect 52733 12115 52791 12121
rect 54202 12112 54208 12164
rect 54260 12152 54266 12164
rect 57333 12155 57391 12161
rect 54260 12124 57284 12152
rect 54260 12112 54266 12124
rect 51997 12087 52055 12093
rect 51997 12084 52009 12087
rect 51184 12056 52009 12084
rect 51997 12053 52009 12056
rect 52043 12053 52055 12087
rect 52362 12084 52368 12096
rect 52323 12056 52368 12084
rect 51997 12047 52055 12053
rect 52362 12044 52368 12056
rect 52420 12044 52426 12096
rect 53926 12084 53932 12096
rect 53887 12056 53932 12084
rect 53926 12044 53932 12056
rect 53984 12044 53990 12096
rect 55214 12044 55220 12096
rect 55272 12093 55278 12096
rect 55272 12087 55321 12093
rect 55272 12053 55275 12087
rect 55309 12053 55321 12087
rect 55272 12047 55321 12053
rect 55272 12044 55278 12047
rect 55398 12044 55404 12096
rect 55456 12084 55462 12096
rect 55950 12084 55956 12096
rect 55456 12056 55956 12084
rect 55456 12044 55462 12056
rect 55950 12044 55956 12056
rect 56008 12084 56014 12096
rect 56229 12087 56287 12093
rect 56229 12084 56241 12087
rect 56008 12056 56241 12084
rect 56008 12044 56014 12056
rect 56229 12053 56241 12056
rect 56275 12084 56287 12087
rect 56597 12087 56655 12093
rect 56597 12084 56609 12087
rect 56275 12056 56609 12084
rect 56275 12053 56287 12056
rect 56229 12047 56287 12053
rect 56597 12053 56609 12056
rect 56643 12084 56655 12087
rect 56686 12084 56692 12096
rect 56643 12056 56692 12084
rect 56643 12053 56655 12056
rect 56597 12047 56655 12053
rect 56686 12044 56692 12056
rect 56744 12044 56750 12096
rect 56870 12084 56876 12096
rect 56831 12056 56876 12084
rect 56870 12044 56876 12056
rect 56928 12044 56934 12096
rect 57256 12084 57284 12124
rect 57333 12121 57345 12155
rect 57379 12152 57391 12155
rect 57790 12152 57796 12164
rect 57379 12124 57796 12152
rect 57379 12121 57391 12124
rect 57333 12115 57391 12121
rect 57790 12112 57796 12124
rect 57848 12112 57854 12164
rect 58176 12124 60504 12152
rect 58176 12096 58204 12124
rect 58158 12084 58164 12096
rect 57256 12056 58164 12084
rect 58158 12044 58164 12056
rect 58216 12044 58222 12096
rect 59170 12084 59176 12096
rect 59131 12056 59176 12084
rect 59170 12044 59176 12056
rect 59228 12044 59234 12096
rect 59722 12084 59728 12096
rect 59683 12056 59728 12084
rect 59722 12044 59728 12056
rect 59780 12044 59786 12096
rect 60476 12093 60504 12124
rect 60461 12087 60519 12093
rect 60461 12053 60473 12087
rect 60507 12053 60519 12087
rect 60461 12047 60519 12053
rect 1104 11994 63480 12016
rect 1104 11942 11378 11994
rect 11430 11942 11442 11994
rect 11494 11942 11506 11994
rect 11558 11942 11570 11994
rect 11622 11942 32170 11994
rect 32222 11942 32234 11994
rect 32286 11942 32298 11994
rect 32350 11942 32362 11994
rect 32414 11942 52962 11994
rect 53014 11942 53026 11994
rect 53078 11942 53090 11994
rect 53142 11942 53154 11994
rect 53206 11942 63480 11994
rect 1104 11920 63480 11942
rect 2866 11880 2872 11892
rect 2827 11852 2872 11880
rect 2866 11840 2872 11852
rect 2924 11840 2930 11892
rect 4617 11883 4675 11889
rect 4617 11849 4629 11883
rect 4663 11880 4675 11883
rect 4706 11880 4712 11892
rect 4663 11852 4712 11880
rect 4663 11849 4675 11852
rect 4617 11843 4675 11849
rect 4706 11840 4712 11852
rect 4764 11880 4770 11892
rect 5442 11880 5448 11892
rect 4764 11852 5448 11880
rect 4764 11840 4770 11852
rect 5442 11840 5448 11852
rect 5500 11880 5506 11892
rect 5813 11883 5871 11889
rect 5813 11880 5825 11883
rect 5500 11852 5825 11880
rect 5500 11840 5506 11852
rect 5813 11849 5825 11852
rect 5859 11849 5871 11883
rect 6546 11880 6552 11892
rect 6507 11852 6552 11880
rect 5813 11843 5871 11849
rect 6546 11840 6552 11852
rect 6604 11840 6610 11892
rect 7929 11883 7987 11889
rect 7929 11849 7941 11883
rect 7975 11880 7987 11883
rect 8018 11880 8024 11892
rect 7975 11852 8024 11880
rect 7975 11849 7987 11852
rect 7929 11843 7987 11849
rect 8018 11840 8024 11852
rect 8076 11840 8082 11892
rect 8386 11840 8392 11892
rect 8444 11880 8450 11892
rect 8757 11883 8815 11889
rect 8757 11880 8769 11883
rect 8444 11852 8769 11880
rect 8444 11840 8450 11852
rect 8757 11849 8769 11852
rect 8803 11880 8815 11883
rect 10321 11883 10379 11889
rect 10321 11880 10333 11883
rect 8803 11852 10333 11880
rect 8803 11849 8815 11852
rect 8757 11843 8815 11849
rect 10321 11849 10333 11852
rect 10367 11880 10379 11883
rect 10962 11880 10968 11892
rect 10367 11852 10968 11880
rect 10367 11849 10379 11852
rect 10321 11843 10379 11849
rect 10962 11840 10968 11852
rect 11020 11840 11026 11892
rect 12158 11880 12164 11892
rect 12119 11852 12164 11880
rect 12158 11840 12164 11852
rect 12216 11840 12222 11892
rect 12526 11840 12532 11892
rect 12584 11880 12590 11892
rect 14277 11883 14335 11889
rect 12584 11852 12756 11880
rect 12584 11840 12590 11852
rect 7193 11815 7251 11821
rect 7193 11781 7205 11815
rect 7239 11812 7251 11815
rect 7558 11812 7564 11824
rect 7239 11784 7564 11812
rect 7239 11781 7251 11784
rect 7193 11775 7251 11781
rect 7558 11772 7564 11784
rect 7616 11812 7622 11824
rect 8404 11812 8432 11840
rect 7616 11784 8432 11812
rect 11885 11815 11943 11821
rect 7616 11772 7622 11784
rect 11885 11781 11897 11815
rect 11931 11812 11943 11815
rect 12618 11812 12624 11824
rect 11931 11784 12624 11812
rect 11931 11781 11943 11784
rect 11885 11775 11943 11781
rect 3326 11744 3332 11756
rect 3287 11716 3332 11744
rect 3326 11704 3332 11716
rect 3384 11704 3390 11756
rect 7650 11744 7656 11756
rect 7563 11716 7656 11744
rect 7650 11704 7656 11716
rect 7708 11744 7714 11756
rect 8202 11744 8208 11756
rect 7708 11716 8208 11744
rect 7708 11704 7714 11716
rect 8202 11704 8208 11716
rect 8260 11744 8266 11756
rect 8297 11747 8355 11753
rect 8297 11744 8309 11747
rect 8260 11716 8309 11744
rect 8260 11704 8266 11716
rect 8297 11713 8309 11716
rect 8343 11713 8355 11747
rect 8297 11707 8355 11713
rect 8478 11704 8484 11756
rect 8536 11744 8542 11756
rect 10689 11747 10747 11753
rect 10689 11744 10701 11747
rect 8536 11716 10701 11744
rect 8536 11704 8542 11716
rect 10689 11713 10701 11716
rect 10735 11744 10747 11747
rect 10781 11747 10839 11753
rect 10781 11744 10793 11747
rect 10735 11716 10793 11744
rect 10735 11713 10747 11716
rect 10689 11707 10747 11713
rect 10781 11713 10793 11716
rect 10827 11713 10839 11747
rect 11900 11744 11928 11775
rect 12618 11772 12624 11784
rect 12676 11772 12682 11824
rect 12728 11821 12756 11852
rect 14277 11849 14289 11883
rect 14323 11880 14335 11883
rect 14458 11880 14464 11892
rect 14323 11852 14464 11880
rect 14323 11849 14335 11852
rect 14277 11843 14335 11849
rect 14458 11840 14464 11852
rect 14516 11840 14522 11892
rect 15654 11880 15660 11892
rect 15615 11852 15660 11880
rect 15654 11840 15660 11852
rect 15712 11840 15718 11892
rect 16761 11883 16819 11889
rect 16761 11849 16773 11883
rect 16807 11880 16819 11883
rect 16850 11880 16856 11892
rect 16807 11852 16856 11880
rect 16807 11849 16819 11852
rect 16761 11843 16819 11849
rect 16850 11840 16856 11852
rect 16908 11840 16914 11892
rect 17037 11883 17095 11889
rect 17037 11849 17049 11883
rect 17083 11880 17095 11883
rect 17494 11880 17500 11892
rect 17083 11852 17500 11880
rect 17083 11849 17095 11852
rect 17037 11843 17095 11849
rect 17494 11840 17500 11852
rect 17552 11840 17558 11892
rect 17586 11840 17592 11892
rect 17644 11880 17650 11892
rect 21821 11883 21879 11889
rect 17644 11852 21220 11880
rect 17644 11840 17650 11852
rect 12713 11815 12771 11821
rect 12713 11781 12725 11815
rect 12759 11812 12771 11815
rect 15381 11815 15439 11821
rect 15381 11812 15393 11815
rect 12759 11784 15393 11812
rect 12759 11781 12771 11784
rect 12713 11775 12771 11781
rect 15381 11781 15393 11784
rect 15427 11781 15439 11815
rect 15381 11775 15439 11781
rect 15838 11772 15844 11824
rect 15896 11812 15902 11824
rect 15933 11815 15991 11821
rect 15933 11812 15945 11815
rect 15896 11784 15945 11812
rect 15896 11772 15902 11784
rect 15933 11781 15945 11784
rect 15979 11812 15991 11815
rect 19150 11812 19156 11824
rect 15979 11784 19156 11812
rect 15979 11781 15991 11784
rect 15933 11775 15991 11781
rect 19150 11772 19156 11784
rect 19208 11772 19214 11824
rect 21082 11812 21088 11824
rect 21043 11784 21088 11812
rect 21082 11772 21088 11784
rect 21140 11772 21146 11824
rect 21192 11812 21220 11852
rect 21821 11849 21833 11883
rect 21867 11880 21879 11883
rect 22094 11880 22100 11892
rect 21867 11852 22100 11880
rect 21867 11849 21879 11852
rect 21821 11843 21879 11849
rect 22094 11840 22100 11852
rect 22152 11840 22158 11892
rect 23842 11880 23848 11892
rect 23803 11852 23848 11880
rect 23842 11840 23848 11852
rect 23900 11840 23906 11892
rect 23952 11852 26464 11880
rect 23952 11812 23980 11852
rect 21192 11784 23980 11812
rect 26436 11812 26464 11852
rect 27246 11840 27252 11892
rect 27304 11880 27310 11892
rect 27433 11883 27491 11889
rect 27433 11880 27445 11883
rect 27304 11852 27445 11880
rect 27304 11840 27310 11852
rect 27433 11849 27445 11852
rect 27479 11880 27491 11883
rect 28994 11880 29000 11892
rect 27479 11852 29000 11880
rect 27479 11849 27491 11852
rect 27433 11843 27491 11849
rect 28994 11840 29000 11852
rect 29052 11840 29058 11892
rect 30190 11840 30196 11892
rect 30248 11880 30254 11892
rect 30469 11883 30527 11889
rect 30469 11880 30481 11883
rect 30248 11852 30481 11880
rect 30248 11840 30254 11852
rect 30469 11849 30481 11852
rect 30515 11849 30527 11883
rect 30469 11843 30527 11849
rect 33137 11883 33195 11889
rect 33137 11849 33149 11883
rect 33183 11880 33195 11883
rect 33318 11880 33324 11892
rect 33183 11852 33324 11880
rect 33183 11849 33195 11852
rect 33137 11843 33195 11849
rect 33318 11840 33324 11852
rect 33376 11840 33382 11892
rect 34146 11880 34152 11892
rect 33428 11852 34152 11880
rect 30742 11812 30748 11824
rect 26436 11784 30748 11812
rect 30742 11772 30748 11784
rect 30800 11772 30806 11824
rect 30837 11815 30895 11821
rect 30837 11781 30849 11815
rect 30883 11812 30895 11815
rect 33428 11812 33456 11852
rect 34146 11840 34152 11852
rect 34204 11840 34210 11892
rect 34330 11880 34336 11892
rect 34291 11852 34336 11880
rect 34330 11840 34336 11852
rect 34388 11840 34394 11892
rect 34514 11840 34520 11892
rect 34572 11880 34578 11892
rect 35069 11883 35127 11889
rect 35069 11880 35081 11883
rect 34572 11852 35081 11880
rect 34572 11840 34578 11852
rect 35069 11849 35081 11852
rect 35115 11849 35127 11883
rect 35526 11880 35532 11892
rect 35487 11852 35532 11880
rect 35069 11843 35127 11849
rect 35526 11840 35532 11852
rect 35584 11840 35590 11892
rect 36173 11883 36231 11889
rect 36173 11849 36185 11883
rect 36219 11849 36231 11883
rect 36173 11843 36231 11849
rect 30883 11784 33456 11812
rect 30883 11781 30895 11784
rect 30837 11775 30895 11781
rect 33686 11772 33692 11824
rect 33744 11812 33750 11824
rect 36188 11812 36216 11843
rect 36998 11840 37004 11892
rect 37056 11880 37062 11892
rect 38933 11883 38991 11889
rect 38933 11880 38945 11883
rect 37056 11852 38945 11880
rect 37056 11840 37062 11852
rect 38933 11849 38945 11852
rect 38979 11849 38991 11883
rect 39758 11880 39764 11892
rect 39719 11852 39764 11880
rect 38933 11843 38991 11849
rect 39758 11840 39764 11852
rect 39816 11840 39822 11892
rect 39942 11840 39948 11892
rect 40000 11880 40006 11892
rect 40221 11883 40279 11889
rect 40221 11880 40233 11883
rect 40000 11852 40233 11880
rect 40000 11840 40006 11852
rect 40221 11849 40233 11852
rect 40267 11849 40279 11883
rect 40862 11880 40868 11892
rect 40823 11852 40868 11880
rect 40221 11843 40279 11849
rect 40862 11840 40868 11852
rect 40920 11840 40926 11892
rect 41233 11883 41291 11889
rect 41233 11849 41245 11883
rect 41279 11880 41291 11883
rect 41506 11880 41512 11892
rect 41279 11852 41512 11880
rect 41279 11849 41291 11852
rect 41233 11843 41291 11849
rect 41506 11840 41512 11852
rect 41564 11840 41570 11892
rect 42429 11883 42487 11889
rect 42429 11849 42441 11883
rect 42475 11880 42487 11883
rect 43073 11883 43131 11889
rect 43073 11880 43085 11883
rect 42475 11852 43085 11880
rect 42475 11849 42487 11852
rect 42429 11843 42487 11849
rect 43073 11849 43085 11852
rect 43119 11880 43131 11883
rect 43346 11880 43352 11892
rect 43119 11852 43352 11880
rect 43119 11849 43131 11852
rect 43073 11843 43131 11849
rect 43346 11840 43352 11852
rect 43404 11840 43410 11892
rect 43438 11840 43444 11892
rect 43496 11880 43502 11892
rect 48406 11880 48412 11892
rect 43496 11852 44588 11880
rect 48367 11852 48412 11880
rect 43496 11840 43502 11852
rect 33744 11784 36216 11812
rect 33744 11772 33750 11784
rect 36446 11772 36452 11824
rect 36504 11812 36510 11824
rect 36725 11815 36783 11821
rect 36725 11812 36737 11815
rect 36504 11784 36737 11812
rect 36504 11772 36510 11784
rect 36725 11781 36737 11784
rect 36771 11812 36783 11815
rect 39776 11812 39804 11840
rect 36771 11784 39804 11812
rect 41601 11815 41659 11821
rect 36771 11781 36783 11784
rect 36725 11775 36783 11781
rect 41601 11781 41613 11815
rect 41647 11812 41659 11815
rect 41966 11812 41972 11824
rect 41647 11784 41972 11812
rect 41647 11781 41659 11784
rect 41601 11775 41659 11781
rect 41966 11772 41972 11784
rect 42024 11772 42030 11824
rect 44085 11815 44143 11821
rect 44085 11781 44097 11815
rect 44131 11812 44143 11815
rect 44450 11812 44456 11824
rect 44131 11784 44456 11812
rect 44131 11781 44143 11784
rect 44085 11775 44143 11781
rect 44450 11772 44456 11784
rect 44508 11772 44514 11824
rect 44560 11812 44588 11852
rect 48406 11840 48412 11852
rect 48464 11840 48470 11892
rect 48774 11880 48780 11892
rect 48735 11852 48780 11880
rect 48774 11840 48780 11852
rect 48832 11840 48838 11892
rect 49050 11840 49056 11892
rect 49108 11880 49114 11892
rect 49697 11883 49755 11889
rect 49697 11880 49709 11883
rect 49108 11852 49709 11880
rect 49108 11840 49114 11852
rect 49697 11849 49709 11852
rect 49743 11849 49755 11883
rect 50522 11880 50528 11892
rect 50483 11852 50528 11880
rect 49697 11843 49755 11849
rect 50522 11840 50528 11852
rect 50580 11840 50586 11892
rect 51537 11883 51595 11889
rect 51537 11849 51549 11883
rect 51583 11880 51595 11883
rect 51718 11880 51724 11892
rect 51583 11852 51724 11880
rect 51583 11849 51595 11852
rect 51537 11843 51595 11849
rect 51718 11840 51724 11852
rect 51776 11840 51782 11892
rect 51902 11840 51908 11892
rect 51960 11880 51966 11892
rect 52227 11883 52285 11889
rect 52227 11880 52239 11883
rect 51960 11852 52239 11880
rect 51960 11840 51966 11852
rect 52227 11849 52239 11852
rect 52273 11849 52285 11883
rect 52362 11880 52368 11892
rect 52323 11852 52368 11880
rect 52227 11843 52285 11849
rect 52362 11840 52368 11852
rect 52420 11840 52426 11892
rect 52454 11840 52460 11892
rect 52512 11880 52518 11892
rect 52549 11883 52607 11889
rect 52549 11880 52561 11883
rect 52512 11852 52561 11880
rect 52512 11840 52518 11852
rect 52549 11849 52561 11852
rect 52595 11849 52607 11883
rect 53466 11880 53472 11892
rect 53427 11852 53472 11880
rect 52549 11843 52607 11849
rect 53466 11840 53472 11852
rect 53524 11840 53530 11892
rect 54570 11880 54576 11892
rect 54531 11852 54576 11880
rect 54570 11840 54576 11852
rect 54628 11840 54634 11892
rect 55490 11840 55496 11892
rect 55548 11880 55554 11892
rect 55548 11852 56088 11880
rect 55548 11840 55554 11852
rect 50890 11812 50896 11824
rect 44560 11784 50896 11812
rect 50890 11772 50896 11784
rect 50948 11772 50954 11824
rect 51994 11812 52000 11824
rect 51907 11784 52000 11812
rect 51994 11772 52000 11784
rect 52052 11812 52058 11824
rect 53558 11812 53564 11824
rect 52052 11784 53564 11812
rect 52052 11772 52058 11784
rect 53558 11772 53564 11784
rect 53616 11812 53622 11824
rect 54389 11815 54447 11821
rect 54389 11812 54401 11815
rect 53616 11784 54401 11812
rect 53616 11772 53622 11784
rect 54389 11781 54401 11784
rect 54435 11812 54447 11815
rect 55398 11812 55404 11824
rect 54435 11784 55404 11812
rect 54435 11781 54447 11784
rect 54389 11775 54447 11781
rect 55398 11772 55404 11784
rect 55456 11772 55462 11824
rect 55766 11812 55772 11824
rect 55692 11784 55772 11812
rect 10781 11707 10839 11713
rect 10980 11716 11928 11744
rect 11977 11747 12035 11753
rect 3053 11679 3111 11685
rect 3053 11645 3065 11679
rect 3099 11676 3111 11679
rect 4246 11676 4252 11688
rect 3099 11648 4252 11676
rect 3099 11645 3111 11648
rect 3053 11639 3111 11645
rect 4246 11636 4252 11648
rect 4304 11636 4310 11688
rect 7432 11679 7490 11685
rect 7432 11645 7444 11679
rect 7478 11676 7490 11679
rect 8662 11676 8668 11688
rect 7478 11648 8668 11676
rect 7478 11645 7490 11648
rect 7432 11639 7490 11645
rect 8662 11636 8668 11648
rect 8720 11636 8726 11688
rect 8846 11676 8852 11688
rect 8807 11648 8852 11676
rect 8846 11636 8852 11648
rect 8904 11636 8910 11688
rect 8941 11679 8999 11685
rect 8941 11645 8953 11679
rect 8987 11676 8999 11679
rect 9766 11676 9772 11688
rect 8987 11648 9772 11676
rect 8987 11645 8999 11648
rect 8941 11639 8999 11645
rect 9766 11636 9772 11648
rect 9824 11636 9830 11688
rect 10594 11636 10600 11688
rect 10652 11676 10658 11688
rect 10980 11685 11008 11716
rect 11977 11713 11989 11747
rect 12023 11744 12035 11747
rect 23934 11744 23940 11756
rect 12023 11716 23940 11744
rect 12023 11713 12035 11716
rect 11977 11707 12035 11713
rect 23934 11704 23940 11716
rect 23992 11704 23998 11756
rect 25774 11744 25780 11756
rect 25735 11716 25780 11744
rect 25774 11704 25780 11716
rect 25832 11704 25838 11756
rect 27154 11744 27160 11756
rect 27115 11716 27160 11744
rect 27154 11704 27160 11716
rect 27212 11704 27218 11756
rect 27430 11704 27436 11756
rect 27488 11744 27494 11756
rect 31573 11747 31631 11753
rect 31573 11744 31585 11747
rect 27488 11716 31585 11744
rect 27488 11704 27494 11716
rect 31573 11713 31585 11716
rect 31619 11744 31631 11747
rect 31662 11744 31668 11756
rect 31619 11716 31668 11744
rect 31619 11713 31631 11716
rect 31573 11707 31631 11713
rect 31662 11704 31668 11716
rect 31720 11704 31726 11756
rect 31754 11704 31760 11756
rect 31812 11744 31818 11756
rect 31812 11716 32076 11744
rect 31812 11704 31818 11716
rect 10965 11679 11023 11685
rect 10652 11648 10916 11676
rect 10652 11636 10658 11648
rect 3988 11580 5580 11608
rect 2501 11543 2559 11549
rect 2501 11509 2513 11543
rect 2547 11540 2559 11543
rect 2866 11540 2872 11552
rect 2547 11512 2872 11540
rect 2547 11509 2559 11512
rect 2501 11503 2559 11509
rect 2866 11500 2872 11512
rect 2924 11500 2930 11552
rect 2958 11500 2964 11552
rect 3016 11540 3022 11552
rect 3988 11540 4016 11580
rect 5552 11552 5580 11580
rect 6914 11568 6920 11620
rect 6972 11608 6978 11620
rect 7285 11611 7343 11617
rect 7285 11608 7297 11611
rect 6972 11580 7297 11608
rect 6972 11568 6978 11580
rect 7285 11577 7297 11580
rect 7331 11608 7343 11611
rect 9401 11611 9459 11617
rect 9401 11608 9413 11611
rect 7331 11580 9413 11608
rect 7331 11577 7343 11580
rect 7285 11571 7343 11577
rect 9401 11577 9413 11580
rect 9447 11577 9459 11611
rect 10888 11608 10916 11648
rect 10965 11645 10977 11679
rect 11011 11645 11023 11679
rect 10965 11639 11023 11645
rect 11057 11679 11115 11685
rect 11057 11645 11069 11679
rect 11103 11676 11115 11679
rect 11238 11676 11244 11688
rect 11103 11648 11244 11676
rect 11103 11645 11115 11648
rect 11057 11639 11115 11645
rect 11238 11636 11244 11648
rect 11296 11636 11302 11688
rect 13081 11679 13139 11685
rect 11348 11648 12664 11676
rect 11149 11611 11207 11617
rect 11149 11608 11161 11611
rect 9401 11571 9459 11577
rect 9508 11580 10732 11608
rect 10888 11580 11161 11608
rect 3016 11512 4016 11540
rect 3016 11500 3022 11512
rect 4614 11500 4620 11552
rect 4672 11540 4678 11552
rect 5074 11540 5080 11552
rect 4672 11512 5080 11540
rect 4672 11500 4678 11512
rect 5074 11500 5080 11512
rect 5132 11500 5138 11552
rect 5534 11540 5540 11552
rect 5447 11512 5540 11540
rect 5534 11500 5540 11512
rect 5592 11540 5598 11552
rect 7006 11540 7012 11552
rect 5592 11512 7012 11540
rect 5592 11500 5598 11512
rect 7006 11500 7012 11512
rect 7064 11500 7070 11552
rect 7190 11500 7196 11552
rect 7248 11540 7254 11552
rect 9508 11540 9536 11580
rect 9766 11540 9772 11552
rect 7248 11512 9536 11540
rect 9679 11512 9772 11540
rect 7248 11500 7254 11512
rect 9766 11500 9772 11512
rect 9824 11540 9830 11552
rect 9950 11540 9956 11552
rect 9824 11512 9956 11540
rect 9824 11500 9830 11512
rect 9950 11500 9956 11512
rect 10008 11500 10014 11552
rect 10704 11540 10732 11580
rect 11149 11577 11161 11580
rect 11195 11608 11207 11611
rect 11348 11608 11376 11648
rect 11195 11580 11376 11608
rect 11517 11611 11575 11617
rect 11195 11577 11207 11580
rect 11149 11571 11207 11577
rect 11517 11577 11529 11611
rect 11563 11608 11575 11611
rect 12342 11608 12348 11620
rect 11563 11580 12348 11608
rect 11563 11577 11575 11580
rect 11517 11571 11575 11577
rect 12342 11568 12348 11580
rect 12400 11568 12406 11620
rect 12636 11608 12664 11648
rect 13081 11645 13093 11679
rect 13127 11645 13139 11679
rect 13081 11639 13139 11645
rect 13357 11679 13415 11685
rect 13357 11645 13369 11679
rect 13403 11676 13415 11679
rect 13403 11648 13952 11676
rect 13403 11645 13415 11648
rect 13357 11639 13415 11645
rect 13096 11608 13124 11639
rect 13722 11608 13728 11620
rect 12636 11580 12940 11608
rect 13096 11580 13728 11608
rect 12912 11549 12940 11580
rect 13722 11568 13728 11580
rect 13780 11568 13786 11620
rect 13924 11617 13952 11648
rect 14274 11636 14280 11688
rect 14332 11676 14338 11688
rect 14369 11679 14427 11685
rect 14369 11676 14381 11679
rect 14332 11648 14381 11676
rect 14332 11636 14338 11648
rect 14369 11645 14381 11648
rect 14415 11645 14427 11679
rect 14369 11639 14427 11645
rect 14458 11636 14464 11688
rect 14516 11676 14522 11688
rect 15194 11676 15200 11688
rect 14516 11648 14561 11676
rect 14844 11648 15200 11676
rect 14516 11636 14522 11648
rect 13909 11611 13967 11617
rect 13909 11577 13921 11611
rect 13955 11608 13967 11611
rect 14844 11608 14872 11648
rect 15194 11636 15200 11648
rect 15252 11636 15258 11688
rect 15381 11679 15439 11685
rect 15381 11645 15393 11679
rect 15427 11676 15439 11679
rect 15749 11679 15807 11685
rect 15749 11676 15761 11679
rect 15427 11648 15761 11676
rect 15427 11645 15439 11648
rect 15381 11639 15439 11645
rect 15749 11645 15761 11648
rect 15795 11676 15807 11679
rect 16390 11676 16396 11688
rect 15795 11648 16396 11676
rect 15795 11645 15807 11648
rect 15749 11639 15807 11645
rect 16390 11636 16396 11648
rect 16448 11636 16454 11688
rect 16853 11679 16911 11685
rect 16853 11645 16865 11679
rect 16899 11676 16911 11679
rect 17405 11679 17463 11685
rect 17405 11676 17417 11679
rect 16899 11648 17417 11676
rect 16899 11645 16911 11648
rect 16853 11639 16911 11645
rect 17405 11645 17417 11648
rect 17451 11676 17463 11679
rect 17954 11676 17960 11688
rect 17451 11648 17960 11676
rect 17451 11645 17463 11648
rect 17405 11639 17463 11645
rect 17954 11636 17960 11648
rect 18012 11636 18018 11688
rect 18322 11676 18328 11688
rect 18283 11648 18328 11676
rect 18322 11636 18328 11648
rect 18380 11636 18386 11688
rect 18417 11679 18475 11685
rect 18417 11645 18429 11679
rect 18463 11645 18475 11679
rect 18417 11639 18475 11645
rect 13955 11580 14872 11608
rect 14921 11611 14979 11617
rect 13955 11577 13967 11580
rect 13909 11571 13967 11577
rect 14921 11577 14933 11611
rect 14967 11608 14979 11611
rect 15286 11608 15292 11620
rect 14967 11580 15292 11608
rect 14967 11577 14979 11580
rect 14921 11571 14979 11577
rect 15286 11568 15292 11580
rect 15344 11568 15350 11620
rect 18046 11608 18052 11620
rect 15396 11580 18052 11608
rect 11977 11543 12035 11549
rect 11977 11540 11989 11543
rect 10704 11512 11989 11540
rect 11977 11509 11989 11512
rect 12023 11509 12035 11543
rect 11977 11503 12035 11509
rect 12897 11543 12955 11549
rect 12897 11509 12909 11543
rect 12943 11509 12955 11543
rect 12897 11503 12955 11509
rect 14458 11500 14464 11552
rect 14516 11540 14522 11552
rect 15102 11540 15108 11552
rect 14516 11512 15108 11540
rect 14516 11500 14522 11512
rect 15102 11500 15108 11512
rect 15160 11540 15166 11552
rect 15197 11543 15255 11549
rect 15197 11540 15209 11543
rect 15160 11512 15209 11540
rect 15160 11500 15166 11512
rect 15197 11509 15209 11512
rect 15243 11540 15255 11543
rect 15396 11540 15424 11580
rect 17788 11552 17816 11580
rect 18046 11568 18052 11580
rect 18104 11568 18110 11620
rect 18230 11568 18236 11620
rect 18288 11608 18294 11620
rect 18432 11608 18460 11639
rect 19610 11636 19616 11688
rect 19668 11676 19674 11688
rect 19705 11679 19763 11685
rect 19705 11676 19717 11679
rect 19668 11648 19717 11676
rect 19668 11636 19674 11648
rect 19705 11645 19717 11648
rect 19751 11645 19763 11679
rect 19705 11639 19763 11645
rect 19794 11636 19800 11688
rect 19852 11676 19858 11688
rect 19981 11679 20039 11685
rect 19981 11676 19993 11679
rect 19852 11648 19993 11676
rect 19852 11636 19858 11648
rect 19981 11645 19993 11648
rect 20027 11645 20039 11679
rect 19981 11639 20039 11645
rect 21082 11636 21088 11688
rect 21140 11676 21146 11688
rect 22186 11676 22192 11688
rect 21140 11648 22192 11676
rect 21140 11636 21146 11648
rect 22186 11636 22192 11648
rect 22244 11636 22250 11688
rect 22281 11679 22339 11685
rect 22281 11645 22293 11679
rect 22327 11676 22339 11679
rect 23014 11676 23020 11688
rect 22327 11648 23020 11676
rect 22327 11645 22339 11648
rect 22281 11639 22339 11645
rect 23014 11636 23020 11648
rect 23072 11636 23078 11688
rect 23290 11636 23296 11688
rect 23348 11676 23354 11688
rect 23477 11679 23535 11685
rect 23477 11676 23489 11679
rect 23348 11648 23489 11676
rect 23348 11636 23354 11648
rect 23477 11645 23489 11648
rect 23523 11676 23535 11679
rect 24305 11679 24363 11685
rect 24305 11676 24317 11679
rect 23523 11648 24317 11676
rect 23523 11645 23535 11648
rect 23477 11639 23535 11645
rect 24305 11645 24317 11648
rect 24351 11676 24363 11679
rect 24486 11676 24492 11688
rect 24351 11648 24492 11676
rect 24351 11645 24363 11648
rect 24305 11639 24363 11645
rect 24486 11636 24492 11648
rect 24544 11636 24550 11688
rect 25501 11679 25559 11685
rect 25501 11645 25513 11679
rect 25547 11645 25559 11679
rect 25501 11639 25559 11645
rect 18874 11608 18880 11620
rect 18288 11580 18460 11608
rect 18835 11580 18880 11608
rect 18288 11568 18294 11580
rect 18874 11568 18880 11580
rect 18932 11568 18938 11620
rect 20898 11568 20904 11620
rect 20956 11608 20962 11620
rect 22741 11611 22799 11617
rect 22741 11608 22753 11611
rect 20956 11580 22753 11608
rect 20956 11568 20962 11580
rect 22741 11577 22753 11580
rect 22787 11577 22799 11611
rect 22741 11571 22799 11577
rect 24118 11568 24124 11620
rect 24176 11608 24182 11620
rect 24673 11611 24731 11617
rect 24176 11580 24221 11608
rect 24176 11568 24182 11580
rect 24673 11577 24685 11611
rect 24719 11608 24731 11611
rect 25130 11608 25136 11620
rect 24719 11580 25136 11608
rect 24719 11577 24731 11580
rect 24673 11571 24731 11577
rect 25130 11568 25136 11580
rect 25188 11568 25194 11620
rect 16390 11540 16396 11552
rect 15243 11512 15424 11540
rect 16351 11512 16396 11540
rect 15243 11509 15255 11512
rect 15197 11503 15255 11509
rect 16390 11500 16396 11512
rect 16448 11500 16454 11552
rect 17770 11540 17776 11552
rect 17731 11512 17776 11540
rect 17770 11500 17776 11512
rect 17828 11500 17834 11552
rect 19150 11500 19156 11552
rect 19208 11540 19214 11552
rect 19245 11543 19303 11549
rect 19245 11540 19257 11543
rect 19208 11512 19257 11540
rect 19208 11500 19214 11512
rect 19245 11509 19257 11512
rect 19291 11509 19303 11543
rect 23014 11540 23020 11552
rect 22975 11512 23020 11540
rect 19245 11503 19303 11509
rect 23014 11500 23020 11512
rect 23072 11500 23078 11552
rect 24946 11500 24952 11552
rect 25004 11540 25010 11552
rect 25041 11543 25099 11549
rect 25041 11540 25053 11543
rect 25004 11512 25053 11540
rect 25004 11500 25010 11512
rect 25041 11509 25053 11512
rect 25087 11540 25099 11543
rect 25406 11540 25412 11552
rect 25087 11512 25412 11540
rect 25087 11509 25099 11512
rect 25041 11503 25099 11509
rect 25406 11500 25412 11512
rect 25464 11500 25470 11552
rect 25516 11540 25544 11639
rect 27798 11636 27804 11688
rect 27856 11676 27862 11688
rect 27985 11679 28043 11685
rect 27985 11676 27997 11679
rect 27856 11648 27997 11676
rect 27856 11636 27862 11648
rect 27985 11645 27997 11648
rect 28031 11676 28043 11679
rect 28537 11679 28595 11685
rect 28537 11676 28549 11679
rect 28031 11648 28549 11676
rect 28031 11645 28043 11648
rect 27985 11639 28043 11645
rect 28537 11645 28549 11648
rect 28583 11676 28595 11679
rect 28902 11676 28908 11688
rect 28583 11648 28908 11676
rect 28583 11645 28595 11648
rect 28537 11639 28595 11645
rect 28902 11636 28908 11648
rect 28960 11636 28966 11688
rect 28994 11636 29000 11688
rect 29052 11676 29058 11688
rect 29273 11679 29331 11685
rect 29273 11676 29285 11679
rect 29052 11648 29285 11676
rect 29052 11636 29058 11648
rect 29273 11645 29285 11648
rect 29319 11645 29331 11679
rect 29273 11639 29331 11645
rect 29457 11679 29515 11685
rect 29457 11645 29469 11679
rect 29503 11676 29515 11679
rect 30653 11679 30711 11685
rect 29503 11648 30236 11676
rect 29503 11645 29515 11648
rect 29457 11639 29515 11645
rect 29086 11608 29092 11620
rect 28184 11580 29092 11608
rect 25866 11540 25872 11552
rect 25516 11512 25872 11540
rect 25866 11500 25872 11512
rect 25924 11500 25930 11552
rect 26786 11500 26792 11552
rect 26844 11540 26850 11552
rect 27522 11540 27528 11552
rect 26844 11512 27528 11540
rect 26844 11500 26850 11512
rect 27522 11500 27528 11512
rect 27580 11540 27586 11552
rect 28184 11549 28212 11580
rect 29086 11568 29092 11580
rect 29144 11608 29150 11620
rect 29472 11608 29500 11639
rect 29144 11580 29500 11608
rect 29144 11568 29150 11580
rect 30208 11552 30236 11648
rect 30653 11645 30665 11679
rect 30699 11645 30711 11679
rect 30653 11639 30711 11645
rect 31941 11679 31999 11685
rect 31941 11645 31953 11679
rect 31987 11676 31999 11679
rect 32048 11676 32076 11716
rect 32398 11704 32404 11756
rect 32456 11744 32462 11756
rect 33870 11744 33876 11756
rect 32456 11716 33732 11744
rect 33831 11716 33876 11744
rect 32456 11704 32462 11716
rect 32858 11676 32864 11688
rect 31987 11648 32864 11676
rect 31987 11645 31999 11648
rect 31941 11639 31999 11645
rect 30668 11608 30696 11639
rect 32858 11636 32864 11648
rect 32916 11636 32922 11688
rect 33045 11679 33103 11685
rect 33045 11645 33057 11679
rect 33091 11676 33103 11679
rect 33410 11676 33416 11688
rect 33091 11648 33416 11676
rect 33091 11645 33103 11648
rect 33045 11639 33103 11645
rect 33410 11636 33416 11648
rect 33468 11636 33474 11688
rect 33704 11676 33732 11716
rect 33870 11704 33876 11716
rect 33928 11704 33934 11756
rect 36814 11744 36820 11756
rect 35912 11716 36820 11744
rect 35912 11685 35940 11716
rect 36814 11704 36820 11716
rect 36872 11704 36878 11756
rect 37737 11747 37795 11753
rect 37737 11744 37749 11747
rect 36924 11716 37749 11744
rect 35713 11679 35771 11685
rect 35713 11676 35725 11679
rect 33704 11648 35725 11676
rect 31297 11611 31355 11617
rect 31297 11608 31309 11611
rect 30668 11580 31309 11608
rect 31297 11577 31309 11580
rect 31343 11608 31355 11611
rect 31343 11580 31708 11608
rect 31343 11577 31355 11580
rect 31297 11571 31355 11577
rect 27801 11543 27859 11549
rect 27801 11540 27813 11543
rect 27580 11512 27813 11540
rect 27580 11500 27586 11512
rect 27801 11509 27813 11512
rect 27847 11509 27859 11543
rect 27801 11503 27859 11509
rect 28169 11543 28227 11549
rect 28169 11509 28181 11543
rect 28215 11509 28227 11543
rect 28169 11503 28227 11509
rect 28258 11500 28264 11552
rect 28316 11540 28322 11552
rect 29549 11543 29607 11549
rect 29549 11540 29561 11543
rect 28316 11512 29561 11540
rect 28316 11500 28322 11512
rect 29549 11509 29561 11512
rect 29595 11509 29607 11543
rect 30190 11540 30196 11552
rect 30103 11512 30196 11540
rect 29549 11503 29607 11509
rect 30190 11500 30196 11512
rect 30248 11540 30254 11552
rect 31478 11540 31484 11552
rect 30248 11512 31484 11540
rect 30248 11500 30254 11512
rect 31478 11500 31484 11512
rect 31536 11500 31542 11552
rect 31680 11540 31708 11580
rect 31754 11568 31760 11620
rect 31812 11608 31818 11620
rect 32309 11611 32367 11617
rect 31812 11580 31857 11608
rect 31812 11568 31818 11580
rect 32309 11577 32321 11611
rect 32355 11608 32367 11611
rect 33321 11611 33379 11617
rect 33321 11608 33333 11611
rect 32355 11580 33333 11608
rect 32355 11577 32367 11580
rect 32309 11571 32367 11577
rect 33321 11577 33333 11580
rect 33367 11608 33379 11611
rect 33502 11608 33508 11620
rect 33367 11580 33508 11608
rect 33367 11577 33379 11580
rect 33321 11571 33379 11577
rect 33502 11568 33508 11580
rect 33560 11568 33566 11620
rect 33594 11568 33600 11620
rect 33652 11608 33658 11620
rect 35158 11608 35164 11620
rect 33652 11580 35164 11608
rect 33652 11568 33658 11580
rect 35158 11568 35164 11580
rect 35216 11568 35222 11620
rect 32490 11540 32496 11552
rect 31680 11512 32496 11540
rect 32490 11500 32496 11512
rect 32548 11500 32554 11552
rect 32582 11500 32588 11552
rect 32640 11540 32646 11552
rect 32677 11543 32735 11549
rect 32677 11540 32689 11543
rect 32640 11512 32689 11540
rect 32640 11500 32646 11512
rect 32677 11509 32689 11512
rect 32723 11540 32735 11543
rect 33042 11540 33048 11552
rect 32723 11512 33048 11540
rect 32723 11509 32735 11512
rect 32677 11503 32735 11509
rect 33042 11500 33048 11512
rect 33100 11500 33106 11552
rect 33134 11500 33140 11552
rect 33192 11540 33198 11552
rect 35342 11540 35348 11552
rect 33192 11512 35348 11540
rect 33192 11500 33198 11512
rect 35342 11500 35348 11512
rect 35400 11500 35406 11552
rect 35544 11540 35572 11648
rect 35713 11645 35725 11648
rect 35759 11645 35771 11679
rect 35713 11639 35771 11645
rect 35897 11679 35955 11685
rect 35897 11645 35909 11679
rect 35943 11645 35955 11679
rect 35897 11639 35955 11645
rect 35989 11679 36047 11685
rect 35989 11645 36001 11679
rect 36035 11676 36047 11679
rect 36924 11676 36952 11716
rect 37737 11713 37749 11716
rect 37783 11713 37795 11747
rect 37737 11707 37795 11713
rect 37826 11704 37832 11756
rect 37884 11744 37890 11756
rect 37884 11716 41651 11744
rect 37884 11704 37890 11716
rect 37458 11676 37464 11688
rect 36035 11648 36952 11676
rect 37419 11648 37464 11676
rect 36035 11645 36047 11648
rect 35989 11639 36047 11645
rect 35618 11568 35624 11620
rect 35676 11608 35682 11620
rect 36004 11608 36032 11639
rect 37458 11636 37464 11648
rect 37516 11676 37522 11688
rect 38841 11679 38899 11685
rect 38841 11676 38853 11679
rect 37516 11648 38853 11676
rect 37516 11636 37522 11648
rect 38841 11645 38853 11648
rect 38887 11645 38899 11679
rect 38841 11639 38899 11645
rect 37093 11611 37151 11617
rect 37093 11608 37105 11611
rect 35676 11580 36032 11608
rect 36188 11580 37105 11608
rect 35676 11568 35682 11580
rect 36188 11540 36216 11580
rect 37093 11577 37105 11580
rect 37139 11577 37151 11611
rect 37274 11608 37280 11620
rect 37235 11580 37280 11608
rect 37093 11571 37151 11577
rect 35544 11512 36216 11540
rect 37108 11540 37136 11571
rect 37274 11568 37280 11580
rect 37332 11568 37338 11620
rect 38654 11568 38660 11620
rect 38712 11608 38718 11620
rect 40402 11608 40408 11620
rect 38712 11580 40408 11608
rect 38712 11568 38718 11580
rect 40402 11568 40408 11580
rect 40460 11568 40466 11620
rect 41623 11608 41651 11716
rect 41690 11704 41696 11756
rect 41748 11744 41754 11756
rect 42245 11747 42303 11753
rect 42245 11744 42257 11747
rect 41748 11716 42257 11744
rect 41748 11704 41754 11716
rect 42245 11713 42257 11716
rect 42291 11744 42303 11747
rect 42613 11747 42671 11753
rect 42613 11744 42625 11747
rect 42291 11716 42625 11744
rect 42291 11713 42303 11716
rect 42245 11707 42303 11713
rect 42613 11713 42625 11716
rect 42659 11744 42671 11747
rect 45278 11744 45284 11756
rect 42659 11716 45284 11744
rect 42659 11713 42671 11716
rect 42613 11707 42671 11713
rect 41782 11676 41788 11688
rect 41743 11648 41788 11676
rect 41782 11636 41788 11648
rect 41840 11676 41846 11688
rect 41966 11676 41972 11688
rect 41840 11648 41972 11676
rect 41840 11636 41846 11648
rect 41966 11636 41972 11648
rect 42024 11636 42030 11688
rect 44836 11685 44864 11716
rect 45278 11704 45284 11716
rect 45336 11744 45342 11756
rect 45465 11747 45523 11753
rect 45465 11744 45477 11747
rect 45336 11716 45477 11744
rect 45336 11704 45342 11716
rect 45465 11713 45477 11716
rect 45511 11713 45523 11747
rect 45465 11707 45523 11713
rect 47397 11747 47455 11753
rect 47397 11713 47409 11747
rect 47443 11744 47455 11747
rect 48314 11744 48320 11756
rect 47443 11716 48320 11744
rect 47443 11713 47455 11716
rect 47397 11707 47455 11713
rect 48314 11704 48320 11716
rect 48372 11704 48378 11756
rect 49421 11747 49479 11753
rect 49421 11713 49433 11747
rect 49467 11744 49479 11747
rect 50614 11744 50620 11756
rect 49467 11716 50620 11744
rect 49467 11713 49479 11716
rect 49421 11707 49479 11713
rect 50614 11704 50620 11716
rect 50672 11704 50678 11756
rect 52454 11744 52460 11756
rect 52415 11716 52460 11744
rect 52454 11704 52460 11716
rect 52512 11744 52518 11756
rect 53101 11747 53159 11753
rect 53101 11744 53113 11747
rect 52512 11716 53113 11744
rect 52512 11704 52518 11716
rect 53101 11713 53113 11716
rect 53147 11713 53159 11747
rect 54481 11747 54539 11753
rect 54481 11744 54493 11747
rect 53101 11707 53159 11713
rect 53944 11716 54493 11744
rect 42153 11679 42211 11685
rect 42153 11645 42165 11679
rect 42199 11676 42211 11679
rect 42429 11679 42487 11685
rect 42429 11676 42441 11679
rect 42199 11648 42441 11676
rect 42199 11645 42211 11648
rect 42153 11639 42211 11645
rect 42429 11645 42441 11648
rect 42475 11645 42487 11679
rect 42429 11639 42487 11645
rect 44637 11679 44695 11685
rect 44637 11645 44649 11679
rect 44683 11645 44695 11679
rect 44637 11639 44695 11645
rect 44821 11679 44879 11685
rect 44821 11645 44833 11679
rect 44867 11645 44879 11679
rect 44821 11639 44879 11645
rect 43438 11608 43444 11620
rect 41623 11580 43444 11608
rect 43438 11568 43444 11580
rect 43496 11568 43502 11620
rect 44542 11568 44548 11620
rect 44600 11608 44606 11620
rect 44652 11608 44680 11639
rect 44910 11636 44916 11688
rect 44968 11676 44974 11688
rect 45005 11679 45063 11685
rect 45005 11676 45017 11679
rect 44968 11648 45017 11676
rect 44968 11636 44974 11648
rect 45005 11645 45017 11648
rect 45051 11676 45063 11679
rect 46293 11679 46351 11685
rect 46293 11676 46305 11679
rect 45051 11648 46305 11676
rect 45051 11645 45063 11648
rect 45005 11639 45063 11645
rect 46293 11645 46305 11648
rect 46339 11645 46351 11679
rect 46842 11676 46848 11688
rect 46803 11648 46848 11676
rect 46293 11639 46351 11645
rect 46842 11636 46848 11648
rect 46900 11636 46906 11688
rect 46937 11679 46995 11685
rect 46937 11645 46949 11679
rect 46983 11676 46995 11679
rect 47026 11676 47032 11688
rect 46983 11648 47032 11676
rect 46983 11645 46995 11648
rect 46937 11639 46995 11645
rect 45833 11611 45891 11617
rect 45833 11608 45845 11611
rect 44600 11580 45845 11608
rect 44600 11568 44606 11580
rect 45833 11577 45845 11580
rect 45879 11577 45891 11611
rect 45833 11571 45891 11577
rect 46753 11611 46811 11617
rect 46753 11577 46765 11611
rect 46799 11608 46811 11611
rect 46952 11608 46980 11639
rect 47026 11636 47032 11648
rect 47084 11676 47090 11688
rect 47673 11679 47731 11685
rect 47673 11676 47685 11679
rect 47084 11648 47685 11676
rect 47084 11636 47090 11648
rect 47673 11645 47685 11648
rect 47719 11645 47731 11679
rect 47673 11639 47731 11645
rect 48406 11636 48412 11688
rect 48464 11676 48470 11688
rect 49053 11679 49111 11685
rect 49053 11676 49065 11679
rect 48464 11648 49065 11676
rect 48464 11636 48470 11648
rect 49053 11645 49065 11648
rect 49099 11645 49111 11679
rect 50246 11676 50252 11688
rect 50207 11648 50252 11676
rect 49053 11639 49111 11645
rect 50246 11636 50252 11648
rect 50304 11636 50310 11688
rect 50341 11679 50399 11685
rect 50341 11645 50353 11679
rect 50387 11676 50399 11679
rect 50387 11648 51212 11676
rect 50387 11645 50399 11648
rect 50341 11639 50399 11645
rect 46799 11580 46980 11608
rect 46799 11577 46811 11580
rect 46753 11571 46811 11577
rect 47486 11568 47492 11620
rect 47544 11608 47550 11620
rect 48869 11611 48927 11617
rect 47544 11580 48820 11608
rect 47544 11568 47550 11580
rect 38286 11540 38292 11552
rect 37108 11512 38292 11540
rect 38286 11500 38292 11512
rect 38344 11500 38350 11552
rect 43717 11543 43775 11549
rect 43717 11509 43729 11543
rect 43763 11540 43775 11543
rect 43898 11540 43904 11552
rect 43763 11512 43904 11540
rect 43763 11509 43775 11512
rect 43717 11503 43775 11509
rect 43898 11500 43904 11512
rect 43956 11500 43962 11552
rect 48792 11540 48820 11580
rect 48869 11577 48881 11611
rect 48915 11608 48927 11611
rect 48958 11608 48964 11620
rect 48915 11580 48964 11608
rect 48915 11577 48927 11580
rect 48869 11571 48927 11577
rect 48958 11568 48964 11580
rect 49016 11608 49022 11620
rect 49418 11608 49424 11620
rect 49016 11580 49424 11608
rect 49016 11568 49022 11580
rect 49418 11568 49424 11580
rect 49476 11608 49482 11620
rect 50065 11611 50123 11617
rect 50065 11608 50077 11611
rect 49476 11580 50077 11608
rect 49476 11568 49482 11580
rect 50065 11577 50077 11580
rect 50111 11577 50123 11611
rect 50065 11571 50123 11577
rect 50264 11540 50292 11636
rect 51184 11617 51212 11648
rect 51994 11636 52000 11688
rect 52052 11676 52058 11688
rect 52089 11679 52147 11685
rect 52089 11676 52101 11679
rect 52052 11648 52101 11676
rect 52052 11636 52058 11648
rect 52089 11645 52101 11648
rect 52135 11645 52147 11679
rect 52089 11639 52147 11645
rect 52270 11636 52276 11688
rect 52328 11676 52334 11688
rect 53944 11676 53972 11716
rect 54481 11713 54493 11716
rect 54527 11744 54539 11747
rect 55125 11747 55183 11753
rect 55125 11744 55137 11747
rect 54527 11716 55137 11744
rect 54527 11713 54539 11716
rect 54481 11707 54539 11713
rect 55125 11713 55137 11716
rect 55171 11744 55183 11747
rect 55490 11744 55496 11756
rect 55171 11716 55496 11744
rect 55171 11713 55183 11716
rect 55125 11707 55183 11713
rect 55490 11704 55496 11716
rect 55548 11704 55554 11756
rect 54110 11676 54116 11688
rect 52328 11648 53972 11676
rect 54071 11648 54116 11676
rect 52328 11636 52334 11648
rect 54110 11636 54116 11648
rect 54168 11636 54174 11688
rect 54260 11679 54318 11685
rect 54260 11645 54272 11679
rect 54306 11676 54318 11679
rect 54306 11645 54340 11676
rect 54260 11639 54340 11645
rect 51169 11611 51227 11617
rect 51169 11577 51181 11611
rect 51215 11608 51227 11611
rect 52822 11608 52828 11620
rect 51215 11580 52828 11608
rect 51215 11577 51227 11580
rect 51169 11571 51227 11577
rect 52822 11568 52828 11580
rect 52880 11568 52886 11620
rect 48792 11512 50292 11540
rect 54021 11543 54079 11549
rect 54021 11509 54033 11543
rect 54067 11540 54079 11543
rect 54312 11540 54340 11639
rect 55692 11617 55720 11784
rect 55766 11772 55772 11784
rect 55824 11772 55830 11824
rect 55950 11812 55956 11824
rect 55911 11784 55956 11812
rect 55950 11772 55956 11784
rect 56008 11772 56014 11824
rect 56060 11753 56088 11852
rect 56226 11840 56232 11892
rect 56284 11880 56290 11892
rect 56321 11883 56379 11889
rect 56321 11880 56333 11883
rect 56284 11852 56333 11880
rect 56284 11840 56290 11852
rect 56321 11849 56333 11852
rect 56367 11849 56379 11883
rect 56321 11843 56379 11849
rect 58437 11883 58495 11889
rect 58437 11849 58449 11883
rect 58483 11880 58495 11883
rect 58894 11880 58900 11892
rect 58483 11852 58900 11880
rect 58483 11849 58495 11852
rect 58437 11843 58495 11849
rect 58894 11840 58900 11852
rect 58952 11840 58958 11892
rect 59538 11812 59544 11824
rect 59499 11784 59544 11812
rect 59538 11772 59544 11784
rect 59596 11772 59602 11824
rect 56045 11747 56103 11753
rect 56045 11713 56057 11747
rect 56091 11744 56103 11747
rect 56689 11747 56747 11753
rect 56689 11744 56701 11747
rect 56091 11716 56701 11744
rect 56091 11713 56103 11716
rect 56045 11707 56103 11713
rect 56689 11713 56701 11716
rect 56735 11744 56747 11747
rect 56778 11744 56784 11756
rect 56735 11716 56784 11744
rect 56735 11713 56747 11716
rect 56689 11707 56747 11713
rect 56778 11704 56784 11716
rect 56836 11704 56842 11756
rect 58713 11747 58771 11753
rect 58713 11744 58725 11747
rect 57808 11716 58725 11744
rect 57808 11688 57836 11716
rect 58713 11713 58725 11716
rect 58759 11713 58771 11747
rect 61102 11744 61108 11756
rect 58713 11707 58771 11713
rect 59924 11716 61108 11744
rect 55824 11679 55882 11685
rect 55824 11645 55836 11679
rect 55870 11676 55882 11679
rect 56134 11676 56140 11688
rect 55870 11648 56140 11676
rect 55870 11645 55882 11648
rect 55824 11639 55882 11645
rect 56134 11636 56140 11648
rect 56192 11676 56198 11688
rect 57057 11679 57115 11685
rect 57057 11676 57069 11679
rect 56192 11648 57069 11676
rect 56192 11636 56198 11648
rect 57057 11645 57069 11648
rect 57103 11645 57115 11679
rect 57422 11676 57428 11688
rect 57383 11648 57428 11676
rect 57057 11639 57115 11645
rect 57422 11636 57428 11648
rect 57480 11636 57486 11688
rect 57790 11676 57796 11688
rect 57751 11648 57796 11676
rect 57790 11636 57796 11648
rect 57848 11636 57854 11688
rect 58158 11676 58164 11688
rect 58119 11648 58164 11676
rect 58158 11636 58164 11648
rect 58216 11676 58222 11688
rect 59081 11679 59139 11685
rect 59081 11676 59093 11679
rect 58216 11648 59093 11676
rect 58216 11636 58222 11648
rect 59081 11645 59093 11648
rect 59127 11645 59139 11679
rect 59722 11676 59728 11688
rect 59683 11648 59728 11676
rect 59081 11639 59139 11645
rect 59722 11636 59728 11648
rect 59780 11636 59786 11688
rect 59924 11685 59952 11716
rect 61102 11704 61108 11716
rect 61160 11704 61166 11756
rect 59909 11679 59967 11685
rect 59909 11645 59921 11679
rect 59955 11645 59967 11679
rect 59909 11639 59967 11645
rect 60093 11679 60151 11685
rect 60093 11645 60105 11679
rect 60139 11645 60151 11679
rect 60093 11639 60151 11645
rect 55677 11611 55735 11617
rect 55677 11577 55689 11611
rect 55723 11608 55735 11611
rect 57606 11608 57612 11620
rect 55723 11580 57612 11608
rect 55723 11577 55735 11580
rect 55677 11571 55735 11577
rect 57606 11568 57612 11580
rect 57664 11568 57670 11620
rect 59262 11568 59268 11620
rect 59320 11608 59326 11620
rect 59924 11608 59952 11639
rect 59320 11580 59952 11608
rect 60108 11608 60136 11639
rect 60826 11608 60832 11620
rect 60108 11580 60832 11608
rect 59320 11568 59326 11580
rect 54846 11540 54852 11552
rect 54067 11512 54852 11540
rect 54067 11509 54079 11512
rect 54021 11503 54079 11509
rect 54846 11500 54852 11512
rect 54904 11500 54910 11552
rect 55030 11500 55036 11552
rect 55088 11540 55094 11552
rect 60108 11540 60136 11580
rect 60826 11568 60832 11580
rect 60884 11608 60890 11620
rect 61289 11611 61347 11617
rect 61289 11608 61301 11611
rect 60884 11580 61301 11608
rect 60884 11568 60890 11580
rect 61289 11577 61301 11580
rect 61335 11577 61347 11611
rect 61289 11571 61347 11577
rect 60550 11540 60556 11552
rect 55088 11512 60136 11540
rect 60511 11512 60556 11540
rect 55088 11500 55094 11512
rect 60550 11500 60556 11512
rect 60608 11500 60614 11552
rect 61013 11543 61071 11549
rect 61013 11509 61025 11543
rect 61059 11540 61071 11543
rect 61102 11540 61108 11552
rect 61059 11512 61108 11540
rect 61059 11509 61071 11512
rect 61013 11503 61071 11509
rect 61102 11500 61108 11512
rect 61160 11500 61166 11552
rect 1104 11450 63480 11472
rect 1104 11398 21774 11450
rect 21826 11398 21838 11450
rect 21890 11398 21902 11450
rect 21954 11398 21966 11450
rect 22018 11398 42566 11450
rect 42618 11398 42630 11450
rect 42682 11398 42694 11450
rect 42746 11398 42758 11450
rect 42810 11398 63480 11450
rect 1104 11376 63480 11398
rect 5626 11296 5632 11348
rect 5684 11336 5690 11348
rect 5997 11339 6055 11345
rect 5997 11336 6009 11339
rect 5684 11308 6009 11336
rect 5684 11296 5690 11308
rect 5997 11305 6009 11308
rect 6043 11305 6055 11339
rect 5997 11299 6055 11305
rect 6012 11268 6040 11299
rect 7098 11296 7104 11348
rect 7156 11336 7162 11348
rect 7929 11339 7987 11345
rect 7929 11336 7941 11339
rect 7156 11308 7941 11336
rect 7156 11296 7162 11308
rect 7929 11305 7941 11308
rect 7975 11305 7987 11339
rect 8386 11336 8392 11348
rect 8347 11308 8392 11336
rect 7929 11299 7987 11305
rect 8386 11296 8392 11308
rect 8444 11296 8450 11348
rect 9766 11296 9772 11348
rect 9824 11296 9830 11348
rect 10686 11336 10692 11348
rect 10647 11308 10692 11336
rect 10686 11296 10692 11308
rect 10744 11296 10750 11348
rect 11149 11339 11207 11345
rect 11149 11305 11161 11339
rect 11195 11336 11207 11339
rect 11238 11336 11244 11348
rect 11195 11308 11244 11336
rect 11195 11305 11207 11308
rect 11149 11299 11207 11305
rect 11238 11296 11244 11308
rect 11296 11296 11302 11348
rect 13998 11296 14004 11348
rect 14056 11336 14062 11348
rect 14277 11339 14335 11345
rect 14277 11336 14289 11339
rect 14056 11308 14289 11336
rect 14056 11296 14062 11308
rect 14277 11305 14289 11308
rect 14323 11305 14335 11339
rect 15102 11336 15108 11348
rect 15063 11308 15108 11336
rect 14277 11299 14335 11305
rect 15102 11296 15108 11308
rect 15160 11296 15166 11348
rect 17034 11336 17040 11348
rect 16995 11308 17040 11336
rect 17034 11296 17040 11308
rect 17092 11296 17098 11348
rect 18785 11339 18843 11345
rect 18785 11305 18797 11339
rect 18831 11336 18843 11339
rect 18874 11336 18880 11348
rect 18831 11308 18880 11336
rect 18831 11305 18843 11308
rect 18785 11299 18843 11305
rect 18874 11296 18880 11308
rect 18932 11296 18938 11348
rect 21174 11336 21180 11348
rect 19168 11308 21180 11336
rect 8846 11268 8852 11280
rect 6012 11240 8852 11268
rect 8846 11228 8852 11240
rect 8904 11228 8910 11280
rect 9784 11268 9812 11296
rect 13173 11271 13231 11277
rect 13173 11268 13185 11271
rect 9692 11240 9812 11268
rect 11992 11240 13185 11268
rect 2866 11160 2872 11212
rect 2924 11200 2930 11212
rect 9692 11209 9720 11240
rect 11992 11212 12020 11240
rect 13173 11237 13185 11240
rect 13219 11237 13231 11271
rect 14918 11268 14924 11280
rect 13173 11231 13231 11237
rect 13556 11240 14924 11268
rect 7285 11203 7343 11209
rect 2924 11172 5396 11200
rect 2924 11160 2930 11172
rect 5368 11144 5396 11172
rect 7285 11169 7297 11203
rect 7331 11169 7343 11203
rect 7285 11163 7343 11169
rect 9677 11203 9735 11209
rect 9677 11169 9689 11203
rect 9723 11169 9735 11203
rect 9677 11163 9735 11169
rect 9769 11203 9827 11209
rect 9769 11169 9781 11203
rect 9815 11169 9827 11203
rect 11974 11200 11980 11212
rect 11935 11172 11980 11200
rect 9769 11163 9827 11169
rect 4617 11135 4675 11141
rect 4617 11132 4629 11135
rect 4264 11104 4629 11132
rect 3145 11067 3203 11073
rect 3145 11033 3157 11067
rect 3191 11064 3203 11067
rect 4264 11064 4292 11104
rect 4617 11101 4629 11104
rect 4663 11101 4675 11135
rect 4617 11095 4675 11101
rect 4893 11135 4951 11141
rect 4893 11101 4905 11135
rect 4939 11132 4951 11135
rect 4982 11132 4988 11144
rect 4939 11104 4988 11132
rect 4939 11101 4951 11104
rect 4893 11095 4951 11101
rect 4982 11092 4988 11104
rect 5040 11092 5046 11144
rect 5350 11092 5356 11144
rect 5408 11132 5414 11144
rect 7190 11132 7196 11144
rect 5408 11104 7196 11132
rect 5408 11092 5414 11104
rect 7190 11092 7196 11104
rect 7248 11092 7254 11144
rect 3191 11036 4292 11064
rect 3191 11033 3203 11036
rect 3145 11027 3203 11033
rect 4264 11008 4292 11036
rect 6825 11067 6883 11073
rect 6825 11033 6837 11067
rect 6871 11064 6883 11067
rect 7299 11064 7327 11163
rect 7466 11141 7472 11144
rect 7432 11135 7472 11141
rect 7432 11101 7444 11135
rect 7432 11095 7472 11101
rect 7466 11092 7472 11095
rect 7524 11092 7530 11144
rect 7650 11132 7656 11144
rect 7611 11104 7656 11132
rect 7650 11092 7656 11104
rect 7708 11092 7714 11144
rect 9784 11132 9812 11163
rect 11974 11160 11980 11172
rect 12032 11160 12038 11212
rect 12066 11160 12072 11212
rect 12124 11200 12130 11212
rect 12161 11203 12219 11209
rect 12161 11200 12173 11203
rect 12124 11172 12173 11200
rect 12124 11160 12130 11172
rect 12161 11169 12173 11172
rect 12207 11169 12219 11203
rect 12161 11163 12219 11169
rect 12250 11160 12256 11212
rect 12308 11200 12314 11212
rect 12345 11203 12403 11209
rect 12345 11200 12357 11203
rect 12308 11172 12357 11200
rect 12308 11160 12314 11172
rect 12345 11169 12357 11172
rect 12391 11200 12403 11203
rect 13556 11200 13584 11240
rect 14918 11228 14924 11240
rect 14976 11228 14982 11280
rect 15286 11268 15292 11280
rect 15247 11240 15292 11268
rect 15286 11228 15292 11240
rect 15344 11228 15350 11280
rect 16025 11271 16083 11277
rect 16025 11237 16037 11271
rect 16071 11268 16083 11271
rect 16114 11268 16120 11280
rect 16071 11240 16120 11268
rect 16071 11237 16083 11240
rect 16025 11231 16083 11237
rect 16114 11228 16120 11240
rect 16172 11228 16178 11280
rect 16850 11228 16856 11280
rect 16908 11268 16914 11280
rect 19168 11268 19196 11308
rect 21174 11296 21180 11308
rect 21232 11296 21238 11348
rect 21821 11339 21879 11345
rect 21821 11305 21833 11339
rect 21867 11336 21879 11339
rect 22005 11339 22063 11345
rect 22005 11336 22017 11339
rect 21867 11308 22017 11336
rect 21867 11305 21879 11308
rect 21821 11299 21879 11305
rect 22005 11305 22017 11308
rect 22051 11336 22063 11339
rect 22097 11339 22155 11345
rect 22097 11336 22109 11339
rect 22051 11308 22109 11336
rect 22051 11305 22063 11308
rect 22005 11299 22063 11305
rect 22097 11305 22109 11308
rect 22143 11305 22155 11339
rect 22097 11299 22155 11305
rect 22557 11339 22615 11345
rect 22557 11305 22569 11339
rect 22603 11336 22615 11339
rect 22738 11336 22744 11348
rect 22603 11308 22744 11336
rect 22603 11305 22615 11308
rect 22557 11299 22615 11305
rect 22738 11296 22744 11308
rect 22796 11296 22802 11348
rect 22922 11336 22928 11348
rect 22883 11308 22928 11336
rect 22922 11296 22928 11308
rect 22980 11296 22986 11348
rect 23198 11296 23204 11348
rect 23256 11336 23262 11348
rect 23293 11339 23351 11345
rect 23293 11336 23305 11339
rect 23256 11308 23305 11336
rect 23256 11296 23262 11308
rect 23293 11305 23305 11308
rect 23339 11305 23351 11339
rect 23293 11299 23351 11305
rect 23474 11296 23480 11348
rect 23532 11336 23538 11348
rect 26697 11339 26755 11345
rect 26697 11336 26709 11339
rect 23532 11308 26709 11336
rect 23532 11296 23538 11308
rect 26697 11305 26709 11308
rect 26743 11336 26755 11339
rect 26743 11308 28580 11336
rect 26743 11305 26755 11308
rect 26697 11299 26755 11305
rect 19978 11268 19984 11280
rect 16908 11240 19196 11268
rect 19939 11240 19984 11268
rect 16908 11228 16914 11240
rect 19978 11228 19984 11240
rect 20036 11228 20042 11280
rect 20717 11271 20775 11277
rect 20717 11237 20729 11271
rect 20763 11268 20775 11271
rect 20898 11268 20904 11280
rect 20763 11240 20904 11268
rect 20763 11237 20775 11240
rect 20717 11231 20775 11237
rect 20898 11228 20904 11240
rect 20956 11228 20962 11280
rect 21637 11271 21695 11277
rect 21637 11237 21649 11271
rect 21683 11268 21695 11271
rect 23566 11268 23572 11280
rect 21683 11240 23572 11268
rect 21683 11237 21695 11240
rect 21637 11231 21695 11237
rect 23566 11228 23572 11240
rect 23624 11228 23630 11280
rect 24305 11271 24363 11277
rect 24305 11268 24317 11271
rect 23676 11240 24317 11268
rect 23676 11212 23704 11240
rect 24305 11237 24317 11240
rect 24351 11268 24363 11271
rect 24762 11268 24768 11280
rect 24351 11240 24768 11268
rect 24351 11237 24363 11240
rect 24305 11231 24363 11237
rect 24762 11228 24768 11240
rect 24820 11228 24826 11280
rect 25593 11271 25651 11277
rect 25593 11237 25605 11271
rect 25639 11268 25651 11271
rect 25774 11268 25780 11280
rect 25639 11240 25780 11268
rect 25639 11237 25651 11240
rect 25593 11231 25651 11237
rect 25774 11228 25780 11240
rect 25832 11228 25838 11280
rect 28552 11268 28580 11308
rect 28994 11296 29000 11348
rect 29052 11336 29058 11348
rect 29362 11336 29368 11348
rect 29052 11308 29368 11336
rect 29052 11296 29058 11308
rect 29362 11296 29368 11308
rect 29420 11336 29426 11348
rect 29549 11339 29607 11345
rect 29549 11336 29561 11339
rect 29420 11308 29561 11336
rect 29420 11296 29426 11308
rect 29549 11305 29561 11308
rect 29595 11305 29607 11339
rect 29549 11299 29607 11305
rect 30742 11296 30748 11348
rect 30800 11336 30806 11348
rect 31113 11339 31171 11345
rect 31113 11336 31125 11339
rect 30800 11308 31125 11336
rect 30800 11296 30806 11308
rect 31113 11305 31125 11308
rect 31159 11336 31171 11339
rect 33226 11336 33232 11348
rect 31159 11308 32536 11336
rect 33187 11308 33232 11336
rect 31159 11305 31171 11308
rect 31113 11299 31171 11305
rect 32398 11268 32404 11280
rect 28552 11240 32404 11268
rect 32398 11228 32404 11240
rect 32456 11228 32462 11280
rect 12391 11172 13584 11200
rect 13633 11203 13691 11209
rect 12391 11169 12403 11172
rect 12345 11163 12403 11169
rect 13633 11169 13645 11203
rect 13679 11200 13691 11203
rect 14182 11200 14188 11212
rect 13679 11172 14188 11200
rect 13679 11169 13691 11172
rect 13633 11163 13691 11169
rect 14182 11160 14188 11172
rect 14240 11160 14246 11212
rect 14274 11160 14280 11212
rect 14332 11200 14338 11212
rect 14645 11203 14703 11209
rect 14645 11200 14657 11203
rect 14332 11172 14657 11200
rect 14332 11160 14338 11172
rect 14645 11169 14657 11172
rect 14691 11169 14703 11203
rect 14645 11163 14703 11169
rect 16206 11160 16212 11212
rect 16264 11200 16270 11212
rect 17678 11200 17684 11212
rect 16264 11172 17684 11200
rect 16264 11160 16270 11172
rect 17678 11160 17684 11172
rect 17736 11160 17742 11212
rect 17770 11160 17776 11212
rect 17828 11200 17834 11212
rect 17957 11203 18015 11209
rect 17957 11200 17969 11203
rect 17828 11172 17969 11200
rect 17828 11160 17834 11172
rect 17957 11169 17969 11172
rect 18003 11169 18015 11203
rect 17957 11163 18015 11169
rect 18417 11203 18475 11209
rect 18417 11169 18429 11203
rect 18463 11200 18475 11203
rect 18690 11200 18696 11212
rect 18463 11172 18696 11200
rect 18463 11169 18475 11172
rect 18417 11163 18475 11169
rect 18690 11160 18696 11172
rect 18748 11160 18754 11212
rect 19245 11203 19303 11209
rect 19245 11169 19257 11203
rect 19291 11169 19303 11203
rect 19245 11163 19303 11169
rect 9950 11132 9956 11144
rect 9784 11104 9956 11132
rect 9950 11092 9956 11104
rect 10008 11132 10014 11144
rect 14001 11135 14059 11141
rect 10008 11104 11928 11132
rect 10008 11092 10014 11104
rect 8294 11064 8300 11076
rect 6871 11036 7236 11064
rect 7299 11036 8300 11064
rect 6871 11033 6883 11036
rect 6825 11027 6883 11033
rect 4246 10996 4252 11008
rect 4207 10968 4252 10996
rect 4246 10956 4252 10968
rect 4304 10956 4310 11008
rect 7098 10996 7104 11008
rect 7059 10968 7104 10996
rect 7098 10956 7104 10968
rect 7156 10956 7162 11008
rect 7208 10996 7236 11036
rect 8294 11024 8300 11036
rect 8352 11064 8358 11076
rect 11790 11064 11796 11076
rect 8352 11036 9996 11064
rect 11751 11036 11796 11064
rect 8352 11024 8358 11036
rect 7374 10996 7380 11008
rect 7208 10968 7380 10996
rect 7374 10956 7380 10968
rect 7432 10956 7438 11008
rect 7561 10999 7619 11005
rect 7561 10965 7573 10999
rect 7607 10996 7619 10999
rect 8386 10996 8392 11008
rect 7607 10968 8392 10996
rect 7607 10965 7619 10968
rect 7561 10959 7619 10965
rect 8386 10956 8392 10968
rect 8444 10956 8450 11008
rect 8754 10956 8760 11008
rect 8812 10996 8818 11008
rect 9968 11005 9996 11036
rect 11790 11024 11796 11036
rect 11848 11024 11854 11076
rect 11900 11064 11928 11104
rect 14001 11101 14013 11135
rect 14047 11132 14059 11135
rect 15657 11135 15715 11141
rect 15657 11132 15669 11135
rect 14047 11104 15669 11132
rect 14047 11101 14059 11104
rect 14001 11095 14059 11101
rect 15657 11101 15669 11104
rect 15703 11132 15715 11135
rect 15838 11132 15844 11144
rect 15703 11104 15844 11132
rect 15703 11101 15715 11104
rect 15657 11095 15715 11101
rect 15838 11092 15844 11104
rect 15896 11092 15902 11144
rect 16666 11092 16672 11144
rect 16724 11132 16730 11144
rect 16761 11135 16819 11141
rect 16761 11132 16773 11135
rect 16724 11104 16773 11132
rect 16724 11092 16730 11104
rect 16761 11101 16773 11104
rect 16807 11132 16819 11135
rect 17862 11132 17868 11144
rect 16807 11104 17724 11132
rect 17823 11104 17868 11132
rect 16807 11101 16819 11104
rect 16761 11095 16819 11101
rect 17586 11064 17592 11076
rect 11900 11036 17592 11064
rect 17586 11024 17592 11036
rect 17644 11024 17650 11076
rect 17696 11064 17724 11104
rect 17862 11092 17868 11104
rect 17920 11092 17926 11144
rect 18874 11092 18880 11144
rect 18932 11132 18938 11144
rect 19260 11132 19288 11163
rect 22462 11160 22468 11212
rect 22520 11200 22526 11212
rect 23474 11200 23480 11212
rect 22520 11172 22565 11200
rect 23435 11172 23480 11200
rect 22520 11160 22526 11172
rect 23474 11160 23480 11172
rect 23532 11160 23538 11212
rect 23658 11200 23664 11212
rect 23619 11172 23664 11200
rect 23658 11160 23664 11172
rect 23716 11160 23722 11212
rect 24029 11203 24087 11209
rect 24029 11169 24041 11203
rect 24075 11200 24087 11203
rect 24854 11200 24860 11212
rect 24075 11172 24860 11200
rect 24075 11169 24087 11172
rect 24029 11163 24087 11169
rect 24854 11160 24860 11172
rect 24912 11200 24918 11212
rect 25041 11203 25099 11209
rect 25041 11200 25053 11203
rect 24912 11172 25053 11200
rect 24912 11160 24918 11172
rect 25041 11169 25053 11172
rect 25087 11169 25099 11203
rect 25041 11163 25099 11169
rect 25130 11160 25136 11212
rect 25188 11200 25194 11212
rect 26237 11203 26295 11209
rect 26237 11200 26249 11203
rect 25188 11172 26249 11200
rect 25188 11160 25194 11172
rect 26237 11169 26249 11172
rect 26283 11169 26295 11203
rect 26237 11163 26295 11169
rect 26326 11160 26332 11212
rect 26384 11200 26390 11212
rect 26513 11203 26571 11209
rect 26513 11200 26525 11203
rect 26384 11172 26525 11200
rect 26384 11160 26390 11172
rect 26513 11169 26525 11172
rect 26559 11200 26571 11203
rect 27154 11200 27160 11212
rect 26559 11172 27160 11200
rect 26559 11169 26571 11172
rect 26513 11163 26571 11169
rect 27154 11160 27160 11172
rect 27212 11160 27218 11212
rect 29454 11200 29460 11212
rect 27632 11172 29460 11200
rect 18932 11104 19288 11132
rect 19613 11135 19671 11141
rect 18932 11092 18938 11104
rect 19613 11101 19625 11135
rect 19659 11132 19671 11135
rect 21266 11132 21272 11144
rect 19659 11104 21272 11132
rect 19659 11101 19671 11104
rect 19613 11095 19671 11101
rect 21266 11092 21272 11104
rect 21324 11092 21330 11144
rect 22097 11135 22155 11141
rect 22097 11101 22109 11135
rect 22143 11132 22155 11135
rect 25314 11132 25320 11144
rect 22143 11104 25320 11132
rect 22143 11101 22155 11104
rect 22097 11095 22155 11101
rect 25314 11092 25320 11104
rect 25372 11092 25378 11144
rect 25866 11092 25872 11144
rect 25924 11132 25930 11144
rect 27632 11141 27660 11172
rect 29454 11160 29460 11172
rect 29512 11200 29518 11212
rect 29917 11203 29975 11209
rect 29917 11200 29929 11203
rect 29512 11172 29929 11200
rect 29512 11160 29518 11172
rect 29917 11169 29929 11172
rect 29963 11169 29975 11203
rect 29917 11163 29975 11169
rect 30929 11203 30987 11209
rect 30929 11169 30941 11203
rect 30975 11200 30987 11203
rect 31570 11200 31576 11212
rect 30975 11172 31576 11200
rect 30975 11169 30987 11172
rect 30929 11163 30987 11169
rect 31570 11160 31576 11172
rect 31628 11160 31634 11212
rect 32508 11209 32536 11308
rect 33226 11296 33232 11308
rect 33284 11296 33290 11348
rect 33686 11336 33692 11348
rect 33647 11308 33692 11336
rect 33686 11296 33692 11308
rect 33744 11296 33750 11348
rect 35894 11336 35900 11348
rect 33888 11308 35900 11336
rect 32953 11271 33011 11277
rect 32953 11237 32965 11271
rect 32999 11268 33011 11271
rect 33888 11268 33916 11308
rect 35894 11296 35900 11308
rect 35952 11296 35958 11348
rect 36078 11336 36084 11348
rect 36039 11308 36084 11336
rect 36078 11296 36084 11308
rect 36136 11296 36142 11348
rect 37458 11336 37464 11348
rect 36188 11308 37464 11336
rect 35434 11268 35440 11280
rect 32999 11240 33916 11268
rect 35395 11240 35440 11268
rect 32999 11237 33011 11240
rect 32953 11231 33011 11237
rect 35434 11228 35440 11240
rect 35492 11228 35498 11280
rect 32493 11203 32551 11209
rect 32493 11169 32505 11203
rect 32539 11200 32551 11203
rect 32582 11200 32588 11212
rect 32539 11172 32588 11200
rect 32539 11169 32551 11172
rect 32493 11163 32551 11169
rect 32582 11160 32588 11172
rect 32640 11160 32646 11212
rect 32858 11160 32864 11212
rect 32916 11200 32922 11212
rect 34057 11203 34115 11209
rect 32916 11172 34008 11200
rect 32916 11160 32922 11172
rect 27617 11135 27675 11141
rect 27617 11132 27629 11135
rect 25924 11104 27629 11132
rect 25924 11092 25930 11104
rect 27617 11101 27629 11104
rect 27663 11101 27675 11135
rect 27617 11095 27675 11101
rect 27798 11092 27804 11144
rect 27856 11132 27862 11144
rect 27893 11135 27951 11141
rect 27893 11132 27905 11135
rect 27856 11104 27905 11132
rect 27856 11092 27862 11104
rect 27893 11101 27905 11104
rect 27939 11101 27951 11135
rect 27893 11095 27951 11101
rect 32401 11135 32459 11141
rect 32401 11101 32413 11135
rect 32447 11101 32459 11135
rect 32401 11095 32459 11101
rect 17773 11067 17831 11073
rect 17773 11064 17785 11067
rect 17696 11036 17785 11064
rect 17773 11033 17785 11036
rect 17819 11064 17831 11067
rect 18322 11064 18328 11076
rect 17819 11036 18328 11064
rect 17819 11033 17831 11036
rect 17773 11027 17831 11033
rect 18322 11024 18328 11036
rect 18380 11064 18386 11076
rect 19058 11064 19064 11076
rect 18380 11036 18920 11064
rect 19019 11036 19064 11064
rect 18380 11024 18386 11036
rect 9217 10999 9275 11005
rect 9217 10996 9229 10999
rect 8812 10968 9229 10996
rect 8812 10956 8818 10968
rect 9217 10965 9229 10968
rect 9263 10965 9275 10999
rect 9217 10959 9275 10965
rect 9953 10999 10011 11005
rect 9953 10965 9965 10999
rect 9999 10965 10011 10999
rect 12802 10996 12808 11008
rect 12763 10968 12808 10996
rect 9953 10959 10011 10965
rect 12802 10956 12808 10968
rect 12860 10956 12866 11008
rect 13814 11005 13820 11008
rect 13798 10999 13820 11005
rect 13798 10965 13810 10999
rect 13798 10959 13820 10965
rect 13814 10956 13820 10959
rect 13872 10956 13878 11008
rect 13909 10999 13967 11005
rect 13909 10965 13921 10999
rect 13955 10996 13967 10999
rect 15194 10996 15200 11008
rect 13955 10968 15200 10996
rect 13955 10965 13967 10968
rect 13909 10959 13967 10965
rect 15194 10956 15200 10968
rect 15252 10956 15258 11008
rect 15470 11005 15476 11008
rect 15454 10999 15476 11005
rect 15454 10965 15466 10999
rect 15454 10959 15476 10965
rect 15470 10956 15476 10959
rect 15528 10956 15534 11008
rect 15562 10956 15568 11008
rect 15620 10996 15626 11008
rect 16206 10996 16212 11008
rect 15620 10968 16212 10996
rect 15620 10956 15626 10968
rect 16206 10956 16212 10968
rect 16264 10956 16270 11008
rect 16298 10956 16304 11008
rect 16356 10996 16362 11008
rect 16356 10968 16401 10996
rect 16356 10956 16362 10968
rect 17954 10956 17960 11008
rect 18012 10996 18018 11008
rect 18690 10996 18696 11008
rect 18012 10968 18696 10996
rect 18012 10956 18018 10968
rect 18690 10956 18696 10968
rect 18748 10956 18754 11008
rect 18892 10996 18920 11036
rect 19058 11024 19064 11036
rect 19116 11064 19122 11076
rect 19383 11067 19441 11073
rect 19383 11064 19395 11067
rect 19116 11036 19395 11064
rect 19116 11024 19122 11036
rect 19383 11033 19395 11036
rect 19429 11033 19441 11067
rect 21066 11067 21124 11073
rect 19383 11027 19441 11033
rect 19812 11036 20484 11064
rect 19242 10996 19248 11008
rect 18892 10968 19248 10996
rect 19242 10956 19248 10968
rect 19300 10956 19306 11008
rect 19518 10996 19524 11008
rect 19431 10968 19524 10996
rect 19518 10956 19524 10968
rect 19576 10996 19582 11008
rect 19812 10996 19840 11036
rect 20456 11008 20484 11036
rect 21066 11033 21078 11067
rect 21112 11064 21124 11067
rect 21821 11067 21879 11073
rect 21821 11064 21833 11067
rect 21112 11036 21833 11064
rect 21112 11033 21124 11036
rect 21066 11027 21124 11033
rect 21821 11033 21833 11036
rect 21867 11033 21879 11067
rect 21821 11027 21879 11033
rect 24765 11067 24823 11073
rect 24765 11033 24777 11067
rect 24811 11064 24823 11067
rect 24946 11064 24952 11076
rect 24811 11036 24952 11064
rect 24811 11033 24823 11036
rect 24765 11027 24823 11033
rect 24946 11024 24952 11036
rect 25004 11024 25010 11076
rect 28997 11067 29055 11073
rect 27080 11036 27384 11064
rect 20346 10996 20352 11008
rect 19576 10968 19840 10996
rect 20307 10968 20352 10996
rect 19576 10956 19582 10968
rect 20346 10956 20352 10968
rect 20404 10956 20410 11008
rect 20438 10956 20444 11008
rect 20496 10996 20502 11008
rect 21177 10999 21235 11005
rect 21177 10996 21189 10999
rect 20496 10968 21189 10996
rect 20496 10956 20502 10968
rect 21177 10965 21189 10968
rect 21223 10996 21235 10999
rect 21726 10996 21732 11008
rect 21223 10968 21732 10996
rect 21223 10965 21235 10968
rect 21177 10959 21235 10965
rect 21726 10956 21732 10968
rect 21784 10956 21790 11008
rect 22094 10956 22100 11008
rect 22152 10996 22158 11008
rect 22281 10999 22339 11005
rect 22281 10996 22293 10999
rect 22152 10968 22293 10996
rect 22152 10956 22158 10968
rect 22281 10965 22293 10968
rect 22327 10965 22339 10999
rect 22281 10959 22339 10965
rect 24670 10956 24676 11008
rect 24728 10996 24734 11008
rect 24857 10999 24915 11005
rect 24857 10996 24869 10999
rect 24728 10968 24869 10996
rect 24728 10956 24734 10968
rect 24857 10965 24869 10968
rect 24903 10965 24915 10999
rect 24964 10996 24992 11024
rect 25774 10996 25780 11008
rect 24964 10968 25780 10996
rect 24857 10959 24915 10965
rect 25774 10956 25780 10968
rect 25832 10956 25838 11008
rect 25958 10996 25964 11008
rect 25919 10968 25964 10996
rect 25958 10956 25964 10968
rect 26016 10956 26022 11008
rect 26050 10956 26056 11008
rect 26108 10996 26114 11008
rect 27080 10996 27108 11036
rect 26108 10968 27108 10996
rect 26108 10956 26114 10968
rect 27154 10956 27160 11008
rect 27212 10996 27218 11008
rect 27356 10996 27384 11036
rect 28997 11033 29009 11067
rect 29043 11064 29055 11067
rect 30098 11064 30104 11076
rect 29043 11036 30104 11064
rect 29043 11033 29055 11036
rect 28997 11027 29055 11033
rect 29012 10996 29040 11027
rect 30098 11024 30104 11036
rect 30156 11024 30162 11076
rect 31573 11067 31631 11073
rect 31573 11033 31585 11067
rect 31619 11064 31631 11067
rect 31754 11064 31760 11076
rect 31619 11036 31760 11064
rect 31619 11033 31631 11036
rect 31573 11027 31631 11033
rect 31754 11024 31760 11036
rect 31812 11064 31818 11076
rect 31938 11064 31944 11076
rect 31812 11036 31944 11064
rect 31812 11024 31818 11036
rect 31938 11024 31944 11036
rect 31996 11064 32002 11076
rect 32416 11064 32444 11095
rect 32766 11092 32772 11144
rect 32824 11132 32830 11144
rect 33134 11132 33140 11144
rect 32824 11104 33140 11132
rect 32824 11092 32830 11104
rect 33134 11092 33140 11104
rect 33192 11132 33198 11144
rect 33778 11132 33784 11144
rect 33192 11104 33784 11132
rect 33192 11092 33198 11104
rect 33778 11092 33784 11104
rect 33836 11092 33842 11144
rect 33980 11132 34008 11172
rect 34057 11169 34069 11203
rect 34103 11200 34115 11203
rect 34330 11200 34336 11212
rect 34103 11172 34336 11200
rect 34103 11169 34115 11172
rect 34057 11163 34115 11169
rect 34330 11160 34336 11172
rect 34388 11160 34394 11212
rect 35342 11160 35348 11212
rect 35400 11200 35406 11212
rect 36188 11200 36216 11308
rect 37458 11296 37464 11308
rect 37516 11336 37522 11348
rect 38289 11339 38347 11345
rect 38289 11336 38301 11339
rect 37516 11308 38301 11336
rect 37516 11296 37522 11308
rect 38289 11305 38301 11308
rect 38335 11305 38347 11339
rect 38289 11299 38347 11305
rect 38470 11296 38476 11348
rect 38528 11336 38534 11348
rect 39758 11336 39764 11348
rect 38528 11308 39764 11336
rect 38528 11296 38534 11308
rect 39758 11296 39764 11308
rect 39816 11296 39822 11348
rect 39850 11296 39856 11348
rect 39908 11336 39914 11348
rect 39908 11308 42012 11336
rect 39908 11296 39914 11308
rect 36265 11271 36323 11277
rect 36265 11237 36277 11271
rect 36311 11268 36323 11271
rect 36814 11268 36820 11280
rect 36311 11240 36676 11268
rect 36775 11240 36820 11268
rect 36311 11237 36323 11240
rect 36265 11231 36323 11237
rect 35400 11172 36216 11200
rect 36449 11203 36507 11209
rect 35400 11160 35406 11172
rect 36449 11169 36461 11203
rect 36495 11169 36507 11203
rect 36449 11163 36507 11169
rect 36354 11132 36360 11144
rect 33980 11104 36360 11132
rect 36354 11092 36360 11104
rect 36412 11132 36418 11144
rect 36464 11132 36492 11163
rect 36412 11104 36492 11132
rect 36648 11132 36676 11240
rect 36814 11228 36820 11240
rect 36872 11228 36878 11280
rect 37366 11228 37372 11280
rect 37424 11268 37430 11280
rect 38488 11268 38516 11296
rect 37424 11240 38516 11268
rect 40129 11271 40187 11277
rect 37424 11228 37430 11240
rect 40129 11237 40141 11271
rect 40175 11268 40187 11271
rect 40494 11268 40500 11280
rect 40175 11240 40500 11268
rect 40175 11237 40187 11240
rect 40129 11231 40187 11237
rect 40494 11228 40500 11240
rect 40552 11228 40558 11280
rect 40586 11228 40592 11280
rect 40644 11268 40650 11280
rect 41984 11268 42012 11308
rect 43438 11296 43444 11348
rect 43496 11336 43502 11348
rect 51258 11336 51264 11348
rect 43496 11308 51120 11336
rect 51219 11308 51264 11336
rect 43496 11296 43502 11308
rect 40644 11240 41914 11268
rect 40644 11228 40650 11240
rect 38013 11203 38071 11209
rect 38013 11169 38025 11203
rect 38059 11200 38071 11203
rect 38838 11200 38844 11212
rect 38059 11172 38844 11200
rect 38059 11169 38071 11172
rect 38013 11163 38071 11169
rect 38838 11160 38844 11172
rect 38896 11200 38902 11212
rect 39390 11200 39396 11212
rect 38896 11172 39396 11200
rect 38896 11160 38902 11172
rect 39390 11160 39396 11172
rect 39448 11160 39454 11212
rect 40402 11200 40408 11212
rect 40363 11172 40408 11200
rect 40402 11160 40408 11172
rect 40460 11160 40466 11212
rect 41506 11160 41512 11212
rect 41564 11200 41570 11212
rect 41601 11203 41659 11209
rect 41601 11200 41613 11203
rect 41564 11172 41613 11200
rect 41564 11160 41570 11172
rect 41601 11169 41613 11172
rect 41647 11169 41659 11203
rect 41601 11163 41659 11169
rect 41690 11160 41696 11212
rect 41748 11200 41754 11212
rect 41785 11203 41843 11209
rect 41785 11200 41797 11203
rect 41748 11172 41797 11200
rect 41748 11160 41754 11172
rect 41785 11169 41797 11172
rect 41831 11169 41843 11203
rect 41785 11163 41843 11169
rect 38286 11132 38292 11144
rect 36648 11104 38292 11132
rect 36412 11092 36418 11104
rect 38286 11092 38292 11104
rect 38344 11092 38350 11144
rect 38473 11135 38531 11141
rect 38473 11101 38485 11135
rect 38519 11101 38531 11135
rect 38746 11132 38752 11144
rect 38707 11104 38752 11132
rect 38473 11095 38531 11101
rect 31996 11036 32444 11064
rect 31996 11024 32002 11036
rect 32490 11024 32496 11076
rect 32548 11064 32554 11076
rect 33594 11064 33600 11076
rect 32548 11036 33600 11064
rect 32548 11024 32554 11036
rect 33594 11024 33600 11036
rect 33652 11024 33658 11076
rect 35710 11064 35716 11076
rect 34716 11036 35716 11064
rect 27212 10968 27257 10996
rect 27356 10968 29040 10996
rect 30377 10999 30435 11005
rect 27212 10956 27218 10968
rect 30377 10965 30389 10999
rect 30423 10996 30435 10999
rect 30466 10996 30472 11008
rect 30423 10968 30472 10996
rect 30423 10965 30435 10968
rect 30377 10959 30435 10965
rect 30466 10956 30472 10968
rect 30524 10956 30530 11008
rect 30745 10999 30803 11005
rect 30745 10965 30757 10999
rect 30791 10996 30803 10999
rect 30926 10996 30932 11008
rect 30791 10968 30932 10996
rect 30791 10965 30803 10968
rect 30745 10959 30803 10965
rect 30926 10956 30932 10968
rect 30984 10956 30990 11008
rect 34422 10956 34428 11008
rect 34480 10996 34486 11008
rect 34716 10996 34744 11036
rect 35710 11024 35716 11036
rect 35768 11024 35774 11076
rect 36446 11024 36452 11076
rect 36504 11064 36510 11076
rect 38010 11064 38016 11076
rect 36504 11036 38016 11064
rect 36504 11024 36510 11036
rect 38010 11024 38016 11036
rect 38068 11064 38074 11076
rect 38488 11064 38516 11095
rect 38746 11092 38752 11104
rect 38804 11092 38810 11144
rect 41049 11135 41107 11141
rect 41049 11101 41061 11135
rect 41095 11132 41107 11135
rect 41886 11132 41914 11240
rect 41984 11240 42932 11268
rect 41984 11209 42012 11240
rect 41969 11203 42027 11209
rect 41969 11169 41981 11203
rect 42015 11169 42027 11203
rect 41969 11163 42027 11169
rect 42904 11141 42932 11240
rect 46658 11228 46664 11280
rect 46716 11268 46722 11280
rect 47213 11271 47271 11277
rect 47213 11268 47225 11271
rect 46716 11240 47225 11268
rect 46716 11228 46722 11240
rect 47213 11237 47225 11240
rect 47259 11237 47271 11271
rect 48038 11268 48044 11280
rect 47999 11240 48044 11268
rect 47213 11231 47271 11237
rect 48038 11228 48044 11240
rect 48096 11228 48102 11280
rect 48774 11228 48780 11280
rect 48832 11268 48838 11280
rect 49513 11271 49571 11277
rect 49513 11268 49525 11271
rect 48832 11240 49525 11268
rect 48832 11228 48838 11240
rect 49513 11237 49525 11240
rect 49559 11237 49571 11271
rect 50890 11268 50896 11280
rect 50851 11240 50896 11268
rect 49513 11231 49571 11237
rect 50890 11228 50896 11240
rect 50948 11228 50954 11280
rect 51092 11268 51120 11308
rect 51258 11296 51264 11308
rect 51316 11296 51322 11348
rect 52546 11296 52552 11348
rect 52604 11336 52610 11348
rect 53009 11339 53067 11345
rect 53009 11336 53021 11339
rect 52604 11308 53021 11336
rect 52604 11296 52610 11308
rect 53009 11305 53021 11308
rect 53055 11305 53067 11339
rect 53009 11299 53067 11305
rect 53469 11339 53527 11345
rect 53469 11305 53481 11339
rect 53515 11336 53527 11339
rect 53558 11336 53564 11348
rect 53515 11308 53564 11336
rect 53515 11305 53527 11308
rect 53469 11299 53527 11305
rect 53558 11296 53564 11308
rect 53616 11296 53622 11348
rect 54110 11296 54116 11348
rect 54168 11336 54174 11348
rect 54205 11339 54263 11345
rect 54205 11336 54217 11339
rect 54168 11308 54217 11336
rect 54168 11296 54174 11308
rect 54205 11305 54217 11308
rect 54251 11305 54263 11339
rect 54205 11299 54263 11305
rect 54941 11339 54999 11345
rect 54941 11305 54953 11339
rect 54987 11336 54999 11339
rect 55214 11336 55220 11348
rect 54987 11308 55220 11336
rect 54987 11305 54999 11308
rect 54941 11299 54999 11305
rect 55214 11296 55220 11308
rect 55272 11296 55278 11348
rect 57793 11339 57851 11345
rect 57793 11305 57805 11339
rect 57839 11336 57851 11339
rect 58066 11336 58072 11348
rect 57839 11308 58072 11336
rect 57839 11305 57851 11308
rect 57793 11299 57851 11305
rect 58066 11296 58072 11308
rect 58124 11296 58130 11348
rect 59538 11336 59544 11348
rect 59499 11308 59544 11336
rect 59538 11296 59544 11308
rect 59596 11296 59602 11348
rect 61565 11339 61623 11345
rect 61565 11336 61577 11339
rect 59924 11308 61577 11336
rect 51626 11268 51632 11280
rect 51092 11240 51632 11268
rect 51626 11228 51632 11240
rect 51684 11228 51690 11280
rect 52362 11228 52368 11280
rect 52420 11268 52426 11280
rect 52457 11271 52515 11277
rect 52457 11268 52469 11271
rect 52420 11240 52469 11268
rect 52420 11228 52426 11240
rect 52457 11237 52469 11240
rect 52503 11237 52515 11271
rect 52457 11231 52515 11237
rect 52825 11271 52883 11277
rect 52825 11237 52837 11271
rect 52871 11268 52883 11271
rect 55030 11268 55036 11280
rect 52871 11240 55036 11268
rect 52871 11237 52883 11240
rect 52825 11231 52883 11237
rect 43346 11200 43352 11212
rect 43307 11172 43352 11200
rect 43346 11160 43352 11172
rect 43404 11160 43410 11212
rect 44174 11160 44180 11212
rect 44232 11200 44238 11212
rect 44637 11203 44695 11209
rect 44637 11200 44649 11203
rect 44232 11172 44649 11200
rect 44232 11160 44238 11172
rect 44637 11169 44649 11172
rect 44683 11169 44695 11203
rect 46676 11200 46704 11228
rect 47578 11200 47584 11212
rect 44637 11163 44695 11169
rect 44744 11172 46704 11200
rect 47539 11172 47584 11200
rect 42889 11135 42947 11141
rect 41095 11104 41828 11132
rect 41886 11104 42012 11132
rect 41095 11101 41107 11104
rect 41049 11095 41107 11101
rect 38068 11036 38516 11064
rect 41417 11067 41475 11073
rect 38068 11024 38074 11036
rect 41417 11033 41429 11067
rect 41463 11033 41475 11067
rect 41800 11064 41828 11104
rect 41874 11064 41880 11076
rect 41800 11036 41880 11064
rect 41417 11027 41475 11033
rect 37090 10996 37096 11008
rect 34480 10968 34744 10996
rect 37051 10968 37096 10996
rect 34480 10956 34486 10968
rect 37090 10956 37096 10968
rect 37148 10956 37154 11008
rect 41432 10996 41460 11027
rect 41874 11024 41880 11036
rect 41932 11024 41938 11076
rect 41984 11064 42012 11104
rect 42889 11101 42901 11135
rect 42935 11132 42947 11135
rect 43162 11132 43168 11144
rect 42935 11104 43168 11132
rect 42935 11101 42947 11104
rect 42889 11095 42947 11101
rect 43162 11092 43168 11104
rect 43220 11132 43226 11144
rect 44744 11132 44772 11172
rect 47578 11160 47584 11172
rect 47636 11200 47642 11212
rect 49053 11203 49111 11209
rect 49053 11200 49065 11203
rect 47636 11172 49065 11200
rect 47636 11160 47642 11172
rect 49053 11169 49065 11172
rect 49099 11200 49111 11203
rect 49326 11200 49332 11212
rect 49099 11172 49332 11200
rect 49099 11169 49111 11172
rect 49053 11163 49111 11169
rect 49326 11160 49332 11172
rect 49384 11200 49390 11212
rect 49973 11203 50031 11209
rect 49973 11200 49985 11203
rect 49384 11172 49985 11200
rect 49384 11160 49390 11172
rect 49973 11169 49985 11172
rect 50019 11200 50031 11203
rect 50433 11203 50491 11209
rect 50433 11200 50445 11203
rect 50019 11172 50445 11200
rect 50019 11169 50031 11172
rect 49973 11163 50031 11169
rect 50433 11169 50445 11172
rect 50479 11169 50491 11203
rect 50433 11163 50491 11169
rect 51997 11203 52055 11209
rect 51997 11169 52009 11203
rect 52043 11200 52055 11203
rect 52270 11200 52276 11212
rect 52043 11172 52276 11200
rect 52043 11169 52055 11172
rect 51997 11163 52055 11169
rect 52270 11160 52276 11172
rect 52328 11160 52334 11212
rect 43220 11104 44772 11132
rect 44913 11135 44971 11141
rect 43220 11092 43226 11104
rect 44913 11101 44925 11135
rect 44959 11132 44971 11135
rect 45370 11132 45376 11144
rect 44959 11104 45376 11132
rect 44959 11101 44971 11104
rect 44913 11095 44971 11101
rect 45370 11092 45376 11104
rect 45428 11092 45434 11144
rect 45554 11092 45560 11144
rect 45612 11132 45618 11144
rect 46017 11135 46075 11141
rect 46017 11132 46029 11135
rect 45612 11104 46029 11132
rect 45612 11092 45618 11104
rect 46017 11101 46029 11104
rect 46063 11132 46075 11135
rect 46842 11132 46848 11144
rect 46063 11104 46848 11132
rect 46063 11101 46075 11104
rect 46017 11095 46075 11101
rect 46842 11092 46848 11104
rect 46900 11092 46906 11144
rect 47489 11135 47547 11141
rect 47489 11101 47501 11135
rect 47535 11132 47547 11135
rect 47854 11132 47860 11144
rect 47535 11104 47860 11132
rect 47535 11101 47547 11104
rect 47489 11095 47547 11101
rect 47854 11092 47860 11104
rect 47912 11092 47918 11144
rect 48498 11092 48504 11144
rect 48556 11132 48562 11144
rect 48961 11135 49019 11141
rect 48961 11132 48973 11135
rect 48556 11104 48973 11132
rect 48556 11092 48562 11104
rect 48961 11101 48973 11104
rect 49007 11132 49019 11135
rect 50338 11132 50344 11144
rect 49007 11104 49832 11132
rect 50299 11104 50344 11132
rect 49007 11101 49019 11104
rect 48961 11095 49019 11101
rect 43533 11067 43591 11073
rect 43533 11064 43545 11067
rect 41984 11036 43545 11064
rect 43533 11033 43545 11036
rect 43579 11033 43591 11067
rect 43533 11027 43591 11033
rect 48409 11067 48467 11073
rect 48409 11033 48421 11067
rect 48455 11064 48467 11067
rect 48866 11064 48872 11076
rect 48455 11036 48872 11064
rect 48455 11033 48467 11036
rect 48409 11027 48467 11033
rect 48866 11024 48872 11036
rect 48924 11024 48930 11076
rect 42058 10996 42064 11008
rect 41432 10968 42064 10996
rect 42058 10956 42064 10968
rect 42116 10996 42122 11008
rect 42429 10999 42487 11005
rect 42429 10996 42441 10999
rect 42116 10968 42441 10996
rect 42116 10956 42122 10968
rect 42429 10965 42441 10968
rect 42475 10965 42487 10999
rect 43898 10996 43904 11008
rect 43859 10968 43904 10996
rect 42429 10959 42487 10965
rect 43898 10956 43904 10968
rect 43956 10956 43962 11008
rect 44358 10996 44364 11008
rect 44319 10968 44364 10996
rect 44358 10956 44364 10968
rect 44416 10956 44422 11008
rect 48774 10996 48780 11008
rect 48735 10968 48780 10996
rect 48774 10956 48780 10968
rect 48832 10956 48838 11008
rect 49804 10996 49832 11104
rect 50338 11092 50344 11104
rect 50396 11092 50402 11144
rect 51442 11092 51448 11144
rect 51500 11132 51506 11144
rect 51905 11135 51963 11141
rect 51905 11132 51917 11135
rect 51500 11104 51917 11132
rect 51500 11092 51506 11104
rect 51905 11101 51917 11104
rect 51951 11132 51963 11135
rect 52840 11132 52868 11231
rect 55030 11228 55036 11240
rect 55088 11228 55094 11280
rect 57149 11271 57207 11277
rect 57149 11237 57161 11271
rect 57195 11268 57207 11271
rect 59170 11268 59176 11280
rect 57195 11240 59176 11268
rect 57195 11237 57207 11240
rect 57149 11231 57207 11237
rect 59170 11228 59176 11240
rect 59228 11228 59234 11280
rect 53009 11203 53067 11209
rect 53009 11169 53021 11203
rect 53055 11200 53067 11203
rect 53285 11203 53343 11209
rect 53285 11200 53297 11203
rect 53055 11172 53297 11200
rect 53055 11169 53067 11172
rect 53009 11163 53067 11169
rect 53285 11169 53297 11172
rect 53331 11200 53343 11203
rect 53837 11203 53895 11209
rect 53837 11200 53849 11203
rect 53331 11172 53849 11200
rect 53331 11169 53343 11172
rect 53285 11163 53343 11169
rect 53837 11169 53849 11172
rect 53883 11169 53895 11203
rect 54938 11200 54944 11212
rect 54851 11172 54944 11200
rect 53837 11163 53895 11169
rect 53190 11132 53196 11144
rect 51951 11104 52868 11132
rect 53151 11104 53196 11132
rect 51951 11101 51963 11104
rect 51905 11095 51963 11101
rect 53190 11092 53196 11104
rect 53248 11092 53254 11144
rect 53466 11092 53472 11144
rect 53524 11132 53530 11144
rect 54864 11132 54892 11172
rect 54938 11160 54944 11172
rect 54996 11200 55002 11212
rect 55125 11203 55183 11209
rect 55125 11200 55137 11203
rect 54996 11172 55137 11200
rect 54996 11160 55002 11172
rect 55125 11169 55137 11172
rect 55171 11169 55183 11203
rect 55125 11163 55183 11169
rect 55585 11203 55643 11209
rect 55585 11169 55597 11203
rect 55631 11200 55643 11203
rect 56410 11200 56416 11212
rect 55631 11172 56416 11200
rect 55631 11169 55643 11172
rect 55585 11163 55643 11169
rect 56410 11160 56416 11172
rect 56468 11160 56474 11212
rect 57422 11160 57428 11212
rect 57480 11200 57486 11212
rect 58069 11203 58127 11209
rect 58069 11200 58081 11203
rect 57480 11172 58081 11200
rect 57480 11160 57486 11172
rect 58069 11169 58081 11172
rect 58115 11169 58127 11203
rect 58069 11163 58127 11169
rect 58713 11203 58771 11209
rect 58713 11169 58725 11203
rect 58759 11200 58771 11203
rect 58802 11200 58808 11212
rect 58759 11172 58808 11200
rect 58759 11169 58771 11172
rect 58713 11163 58771 11169
rect 58802 11160 58808 11172
rect 58860 11160 58866 11212
rect 59924 11209 59952 11308
rect 61565 11305 61577 11308
rect 61611 11305 61623 11339
rect 61565 11299 61623 11305
rect 59081 11203 59139 11209
rect 59081 11169 59093 11203
rect 59127 11200 59139 11203
rect 59909 11203 59967 11209
rect 59909 11200 59921 11203
rect 59127 11172 59921 11200
rect 59127 11169 59139 11172
rect 59081 11163 59139 11169
rect 59909 11169 59921 11172
rect 59955 11169 59967 11203
rect 60458 11200 60464 11212
rect 59909 11163 59967 11169
rect 60108 11172 60464 11200
rect 53524 11104 54892 11132
rect 55033 11135 55091 11141
rect 53524 11092 53530 11104
rect 55033 11101 55045 11135
rect 55079 11101 55091 11135
rect 56778 11132 56784 11144
rect 56739 11104 56784 11132
rect 55033 11095 55091 11101
rect 51350 11024 51356 11076
rect 51408 11064 51414 11076
rect 55048 11064 55076 11095
rect 56778 11092 56784 11104
rect 56836 11092 56842 11144
rect 57330 11092 57336 11144
rect 57388 11132 57394 11144
rect 59096 11132 59124 11163
rect 57388 11104 59124 11132
rect 57388 11092 57394 11104
rect 59170 11092 59176 11144
rect 59228 11132 59234 11144
rect 59228 11104 59273 11132
rect 59228 11092 59234 11104
rect 55766 11064 55772 11076
rect 51408 11036 55772 11064
rect 51408 11024 51414 11036
rect 55766 11024 55772 11036
rect 55824 11024 55830 11076
rect 58529 11067 58587 11073
rect 58529 11033 58541 11067
rect 58575 11064 58587 11067
rect 60108 11064 60136 11172
rect 60458 11160 60464 11172
rect 60516 11160 60522 11212
rect 60185 11135 60243 11141
rect 60185 11101 60197 11135
rect 60231 11101 60243 11135
rect 60185 11095 60243 11101
rect 58575 11036 60136 11064
rect 58575 11033 58587 11036
rect 58529 11027 58587 11033
rect 51074 10996 51080 11008
rect 49804 10968 51080 10996
rect 51074 10956 51080 10968
rect 51132 10956 51138 11008
rect 51718 10996 51724 11008
rect 51679 10968 51724 10996
rect 51718 10956 51724 10968
rect 51776 10956 51782 11008
rect 55950 10996 55956 11008
rect 55911 10968 55956 10996
rect 55950 10956 55956 10968
rect 56008 10956 56014 11008
rect 56594 11005 56600 11008
rect 56578 10999 56600 11005
rect 56578 10965 56590 10999
rect 56578 10959 56600 10965
rect 56594 10956 56600 10959
rect 56652 10956 56658 11008
rect 56686 10956 56692 11008
rect 56744 10996 56750 11008
rect 57238 10996 57244 11008
rect 56744 10968 57244 10996
rect 56744 10956 56750 10968
rect 57238 10956 57244 10968
rect 57296 10956 57302 11008
rect 59262 10956 59268 11008
rect 59320 10996 59326 11008
rect 60200 10996 60228 11095
rect 59320 10968 60228 10996
rect 59320 10956 59326 10968
rect 1104 10906 63480 10928
rect 1104 10854 11378 10906
rect 11430 10854 11442 10906
rect 11494 10854 11506 10906
rect 11558 10854 11570 10906
rect 11622 10854 32170 10906
rect 32222 10854 32234 10906
rect 32286 10854 32298 10906
rect 32350 10854 32362 10906
rect 32414 10854 52962 10906
rect 53014 10854 53026 10906
rect 53078 10854 53090 10906
rect 53142 10854 53154 10906
rect 53206 10854 63480 10906
rect 1104 10832 63480 10854
rect 5258 10752 5264 10804
rect 5316 10792 5322 10804
rect 5442 10792 5448 10804
rect 5316 10764 5448 10792
rect 5316 10752 5322 10764
rect 5442 10752 5448 10764
rect 5500 10792 5506 10804
rect 5629 10795 5687 10801
rect 5629 10792 5641 10795
rect 5500 10764 5641 10792
rect 5500 10752 5506 10764
rect 5629 10761 5641 10764
rect 5675 10761 5687 10795
rect 5629 10755 5687 10761
rect 3789 10659 3847 10665
rect 3789 10625 3801 10659
rect 3835 10656 3847 10659
rect 5644 10656 5672 10755
rect 7650 10752 7656 10804
rect 7708 10792 7714 10804
rect 8113 10795 8171 10801
rect 8113 10792 8125 10795
rect 7708 10764 8125 10792
rect 7708 10752 7714 10764
rect 8113 10761 8125 10764
rect 8159 10761 8171 10795
rect 8113 10755 8171 10761
rect 8294 10752 8300 10804
rect 8352 10792 8358 10804
rect 8481 10795 8539 10801
rect 8481 10792 8493 10795
rect 8352 10764 8493 10792
rect 8352 10752 8358 10764
rect 8481 10761 8493 10764
rect 8527 10761 8539 10795
rect 8481 10755 8539 10761
rect 8662 10752 8668 10804
rect 8720 10792 8726 10804
rect 8941 10795 8999 10801
rect 8941 10792 8953 10795
rect 8720 10764 8953 10792
rect 8720 10752 8726 10764
rect 8941 10761 8953 10764
rect 8987 10761 8999 10795
rect 9950 10792 9956 10804
rect 9911 10764 9956 10792
rect 8941 10755 8999 10761
rect 9950 10752 9956 10764
rect 10008 10752 10014 10804
rect 11241 10795 11299 10801
rect 11241 10761 11253 10795
rect 11287 10792 11299 10795
rect 11882 10792 11888 10804
rect 11287 10764 11888 10792
rect 11287 10761 11299 10764
rect 11241 10755 11299 10761
rect 11882 10752 11888 10764
rect 11940 10752 11946 10804
rect 12618 10792 12624 10804
rect 12176 10764 12624 10792
rect 7282 10684 7288 10736
rect 7340 10724 7346 10736
rect 9766 10724 9772 10736
rect 7340 10696 9772 10724
rect 7340 10684 7346 10696
rect 9766 10684 9772 10696
rect 9824 10724 9830 10736
rect 10229 10727 10287 10733
rect 10229 10724 10241 10727
rect 9824 10696 10241 10724
rect 9824 10684 9830 10696
rect 10229 10693 10241 10696
rect 10275 10693 10287 10727
rect 10229 10687 10287 10693
rect 10686 10684 10692 10736
rect 10744 10724 10750 10736
rect 12066 10724 12072 10736
rect 10744 10696 12072 10724
rect 10744 10684 10750 10696
rect 12066 10684 12072 10696
rect 12124 10724 12130 10736
rect 12176 10733 12204 10764
rect 12618 10752 12624 10764
rect 12676 10752 12682 10804
rect 14182 10752 14188 10804
rect 14240 10792 14246 10804
rect 15197 10795 15255 10801
rect 15197 10792 15209 10795
rect 14240 10764 15209 10792
rect 14240 10752 14246 10764
rect 15197 10761 15209 10764
rect 15243 10761 15255 10795
rect 15197 10755 15255 10761
rect 15286 10752 15292 10804
rect 15344 10792 15350 10804
rect 16577 10795 16635 10801
rect 16577 10792 16589 10795
rect 15344 10764 16589 10792
rect 15344 10752 15350 10764
rect 16577 10761 16589 10764
rect 16623 10761 16635 10795
rect 16577 10755 16635 10761
rect 18322 10752 18328 10804
rect 18380 10792 18386 10804
rect 18380 10764 19104 10792
rect 18380 10752 18386 10764
rect 12161 10727 12219 10733
rect 12161 10724 12173 10727
rect 12124 10696 12173 10724
rect 12124 10684 12130 10696
rect 12161 10693 12173 10696
rect 12207 10693 12219 10727
rect 12161 10687 12219 10693
rect 14461 10727 14519 10733
rect 14461 10693 14473 10727
rect 14507 10724 14519 10727
rect 15838 10724 15844 10736
rect 14507 10696 15844 10724
rect 14507 10693 14519 10696
rect 14461 10687 14519 10693
rect 15838 10684 15844 10696
rect 15896 10684 15902 10736
rect 16206 10724 16212 10736
rect 16167 10696 16212 10724
rect 16206 10684 16212 10696
rect 16264 10684 16270 10736
rect 17129 10727 17187 10733
rect 17129 10693 17141 10727
rect 17175 10724 17187 10727
rect 17862 10724 17868 10736
rect 17175 10696 17868 10724
rect 17175 10693 17187 10696
rect 17129 10687 17187 10693
rect 17862 10684 17868 10696
rect 17920 10724 17926 10736
rect 19076 10724 19104 10764
rect 19150 10752 19156 10804
rect 19208 10792 19214 10804
rect 19521 10795 19579 10801
rect 19521 10792 19533 10795
rect 19208 10764 19533 10792
rect 19208 10752 19214 10764
rect 19521 10761 19533 10764
rect 19567 10792 19579 10795
rect 21266 10792 21272 10804
rect 19567 10764 21272 10792
rect 19567 10761 19579 10764
rect 19521 10755 19579 10761
rect 21266 10752 21272 10764
rect 21324 10792 21330 10804
rect 21545 10795 21603 10801
rect 21545 10792 21557 10795
rect 21324 10764 21557 10792
rect 21324 10752 21330 10764
rect 21545 10761 21557 10764
rect 21591 10761 21603 10795
rect 21545 10755 21603 10761
rect 21726 10752 21732 10804
rect 21784 10792 21790 10804
rect 21913 10795 21971 10801
rect 21913 10792 21925 10795
rect 21784 10764 21925 10792
rect 21784 10752 21790 10764
rect 21913 10761 21925 10764
rect 21959 10761 21971 10795
rect 21913 10755 21971 10761
rect 22278 10752 22284 10804
rect 22336 10792 22342 10804
rect 30098 10792 30104 10804
rect 22336 10764 30104 10792
rect 22336 10752 22342 10764
rect 30098 10752 30104 10764
rect 30156 10752 30162 10804
rect 30190 10752 30196 10804
rect 30248 10792 30254 10804
rect 30466 10792 30472 10804
rect 30248 10764 30293 10792
rect 30427 10764 30472 10792
rect 30248 10752 30254 10764
rect 30466 10752 30472 10764
rect 30524 10752 30530 10804
rect 31202 10752 31208 10804
rect 31260 10792 31266 10804
rect 33873 10795 33931 10801
rect 33873 10792 33885 10795
rect 31260 10764 33885 10792
rect 31260 10752 31266 10764
rect 33873 10761 33885 10764
rect 33919 10792 33931 10795
rect 34514 10792 34520 10804
rect 33919 10764 34520 10792
rect 33919 10761 33931 10764
rect 33873 10755 33931 10761
rect 34514 10752 34520 10764
rect 34572 10752 34578 10804
rect 36354 10792 36360 10804
rect 36315 10764 36360 10792
rect 36354 10752 36360 10764
rect 36412 10752 36418 10804
rect 36630 10752 36636 10804
rect 36688 10792 36694 10804
rect 37918 10792 37924 10804
rect 36688 10764 37924 10792
rect 36688 10752 36694 10764
rect 37918 10752 37924 10764
rect 37976 10792 37982 10804
rect 38381 10795 38439 10801
rect 38381 10792 38393 10795
rect 37976 10764 38393 10792
rect 37976 10752 37982 10764
rect 38381 10761 38393 10764
rect 38427 10761 38439 10795
rect 38381 10755 38439 10761
rect 38562 10752 38568 10804
rect 38620 10792 38626 10804
rect 44542 10792 44548 10804
rect 38620 10764 44036 10792
rect 44503 10764 44548 10792
rect 38620 10752 38626 10764
rect 19610 10724 19616 10736
rect 17920 10696 18736 10724
rect 19076 10696 19616 10724
rect 17920 10684 17926 10696
rect 10781 10659 10839 10665
rect 10781 10656 10793 10659
rect 3835 10628 4568 10656
rect 5644 10628 10793 10656
rect 3835 10625 3847 10628
rect 3789 10619 3847 10625
rect 4246 10588 4252 10600
rect 4207 10560 4252 10588
rect 4246 10548 4252 10560
rect 4304 10548 4310 10600
rect 4540 10597 4568 10628
rect 4525 10591 4583 10597
rect 4525 10557 4537 10591
rect 4571 10588 4583 10591
rect 6825 10591 6883 10597
rect 6825 10588 6837 10591
rect 4571 10560 6837 10588
rect 4571 10557 4583 10560
rect 4525 10551 4583 10557
rect 6825 10557 6837 10560
rect 6871 10557 6883 10591
rect 6825 10551 6883 10557
rect 7285 10591 7343 10597
rect 7285 10557 7297 10591
rect 7331 10588 7343 10591
rect 7374 10588 7380 10600
rect 7331 10560 7380 10588
rect 7331 10557 7343 10560
rect 7285 10551 7343 10557
rect 7374 10548 7380 10560
rect 7432 10548 7438 10600
rect 7668 10597 7696 10628
rect 10781 10625 10793 10628
rect 10827 10656 10839 10659
rect 10965 10659 11023 10665
rect 10965 10656 10977 10659
rect 10827 10628 10977 10656
rect 10827 10625 10839 10628
rect 10781 10619 10839 10625
rect 10965 10625 10977 10628
rect 11011 10625 11023 10659
rect 10965 10619 11023 10625
rect 12713 10659 12771 10665
rect 12713 10625 12725 10659
rect 12759 10656 12771 10659
rect 12802 10656 12808 10668
rect 12759 10628 12808 10656
rect 12759 10625 12771 10628
rect 12713 10619 12771 10625
rect 12802 10616 12808 10628
rect 12860 10616 12866 10668
rect 12894 10616 12900 10668
rect 12952 10616 12958 10668
rect 14093 10659 14151 10665
rect 14093 10625 14105 10659
rect 14139 10656 14151 10659
rect 14274 10656 14280 10668
rect 14139 10628 14280 10656
rect 14139 10625 14151 10628
rect 14093 10619 14151 10625
rect 14274 10616 14280 10628
rect 14332 10616 14338 10668
rect 14918 10656 14924 10668
rect 14879 10628 14924 10656
rect 14918 10616 14924 10628
rect 14976 10616 14982 10668
rect 18049 10659 18107 10665
rect 18049 10625 18061 10659
rect 18095 10656 18107 10659
rect 18598 10656 18604 10668
rect 18095 10628 18460 10656
rect 18559 10628 18604 10656
rect 18095 10625 18107 10628
rect 18049 10619 18107 10625
rect 7653 10591 7711 10597
rect 7653 10557 7665 10591
rect 7699 10557 7711 10591
rect 7653 10551 7711 10557
rect 7745 10591 7803 10597
rect 7745 10557 7757 10591
rect 7791 10588 7803 10591
rect 7834 10588 7840 10600
rect 7791 10560 7840 10588
rect 7791 10557 7803 10560
rect 7745 10551 7803 10557
rect 7098 10480 7104 10532
rect 7156 10520 7162 10532
rect 7760 10520 7788 10551
rect 7834 10548 7840 10560
rect 7892 10548 7898 10600
rect 8662 10588 8668 10600
rect 8623 10560 8668 10588
rect 8662 10548 8668 10560
rect 8720 10548 8726 10600
rect 8757 10591 8815 10597
rect 8757 10557 8769 10591
rect 8803 10557 8815 10591
rect 8757 10551 8815 10557
rect 11057 10591 11115 10597
rect 11057 10557 11069 10591
rect 11103 10588 11115 10591
rect 11793 10591 11851 10597
rect 11793 10588 11805 10591
rect 11103 10560 11805 10588
rect 11103 10557 11115 10560
rect 11057 10551 11115 10557
rect 11793 10557 11805 10560
rect 11839 10557 11851 10591
rect 11793 10551 11851 10557
rect 12437 10591 12495 10597
rect 12437 10557 12449 10591
rect 12483 10588 12495 10591
rect 12912 10588 12940 10616
rect 13446 10588 13452 10600
rect 12483 10560 13452 10588
rect 12483 10557 12495 10560
rect 12437 10551 12495 10557
rect 7156 10492 7788 10520
rect 7156 10480 7162 10492
rect 4157 10455 4215 10461
rect 4157 10421 4169 10455
rect 4203 10452 4215 10455
rect 4982 10452 4988 10464
rect 4203 10424 4988 10452
rect 4203 10421 4215 10424
rect 4157 10415 4215 10421
rect 4982 10412 4988 10424
rect 5040 10412 5046 10464
rect 6273 10455 6331 10461
rect 6273 10421 6285 10455
rect 6319 10452 6331 10455
rect 6362 10452 6368 10464
rect 6319 10424 6368 10452
rect 6319 10421 6331 10424
rect 6273 10415 6331 10421
rect 6362 10412 6368 10424
rect 6420 10412 6426 10464
rect 6641 10455 6699 10461
rect 6641 10421 6653 10455
rect 6687 10452 6699 10455
rect 7466 10452 7472 10464
rect 6687 10424 7472 10452
rect 6687 10421 6699 10424
rect 6641 10415 6699 10421
rect 7466 10412 7472 10424
rect 7524 10412 7530 10464
rect 8772 10452 8800 10551
rect 9585 10455 9643 10461
rect 9585 10452 9597 10455
rect 8772 10424 9597 10452
rect 9585 10421 9597 10424
rect 9631 10452 9643 10455
rect 9766 10452 9772 10464
rect 9631 10424 9772 10452
rect 9631 10421 9643 10424
rect 9585 10415 9643 10421
rect 9766 10412 9772 10424
rect 9824 10412 9830 10464
rect 11808 10452 11836 10551
rect 13446 10548 13452 10560
rect 13504 10548 13510 10600
rect 15013 10591 15071 10597
rect 15013 10588 15025 10591
rect 14752 10560 15025 10588
rect 14752 10452 14780 10560
rect 15013 10557 15025 10560
rect 15059 10588 15071 10591
rect 15102 10588 15108 10600
rect 15059 10560 15108 10588
rect 15059 10557 15071 10560
rect 15013 10551 15071 10557
rect 15102 10548 15108 10560
rect 15160 10548 15166 10600
rect 18141 10591 18199 10597
rect 18141 10588 18153 10591
rect 17420 10560 18153 10588
rect 14829 10523 14887 10529
rect 14829 10489 14841 10523
rect 14875 10520 14887 10523
rect 15194 10520 15200 10532
rect 14875 10492 15200 10520
rect 14875 10489 14887 10492
rect 14829 10483 14887 10489
rect 15194 10480 15200 10492
rect 15252 10520 15258 10532
rect 15562 10520 15568 10532
rect 15252 10492 15568 10520
rect 15252 10480 15258 10492
rect 15562 10480 15568 10492
rect 15620 10480 15626 10532
rect 17420 10464 17448 10560
rect 18141 10557 18153 10560
rect 18187 10557 18199 10591
rect 18432 10588 18460 10628
rect 18598 10616 18604 10628
rect 18656 10616 18662 10668
rect 18708 10656 18736 10696
rect 19610 10684 19616 10696
rect 19668 10684 19674 10736
rect 20714 10684 20720 10736
rect 20772 10724 20778 10736
rect 22922 10724 22928 10736
rect 20772 10696 22928 10724
rect 20772 10684 20778 10696
rect 20993 10659 21051 10665
rect 20993 10656 21005 10659
rect 18708 10628 21005 10656
rect 20993 10625 21005 10628
rect 21039 10625 21051 10659
rect 20993 10619 21051 10625
rect 19610 10588 19616 10600
rect 18432 10560 19012 10588
rect 19571 10560 19616 10588
rect 18141 10551 18199 10557
rect 18984 10532 19012 10560
rect 19610 10548 19616 10560
rect 19668 10548 19674 10600
rect 19889 10591 19947 10597
rect 19889 10557 19901 10591
rect 19935 10588 19947 10591
rect 20346 10588 20352 10600
rect 19935 10560 20352 10588
rect 19935 10557 19947 10560
rect 19889 10551 19947 10557
rect 20346 10548 20352 10560
rect 20404 10548 20410 10600
rect 18230 10480 18236 10532
rect 18288 10520 18294 10532
rect 18782 10520 18788 10532
rect 18288 10492 18788 10520
rect 18288 10480 18294 10492
rect 18782 10480 18788 10492
rect 18840 10480 18846 10532
rect 18966 10520 18972 10532
rect 18927 10492 18972 10520
rect 18966 10480 18972 10492
rect 19024 10480 19030 10532
rect 21008 10520 21036 10619
rect 22296 10597 22324 10696
rect 22922 10684 22928 10696
rect 22980 10684 22986 10736
rect 23474 10724 23480 10736
rect 23435 10696 23480 10724
rect 23474 10684 23480 10696
rect 23532 10684 23538 10736
rect 25038 10684 25044 10736
rect 25096 10724 25102 10736
rect 25096 10696 29868 10724
rect 25096 10684 25102 10696
rect 22646 10656 22652 10668
rect 22607 10628 22652 10656
rect 22646 10616 22652 10628
rect 22704 10616 22710 10668
rect 24305 10659 24363 10665
rect 24305 10625 24317 10659
rect 24351 10656 24363 10659
rect 25409 10659 25467 10665
rect 24351 10628 25360 10656
rect 24351 10625 24363 10628
rect 24305 10619 24363 10625
rect 22281 10591 22339 10597
rect 22281 10557 22293 10591
rect 22327 10557 22339 10591
rect 22281 10551 22339 10557
rect 23198 10548 23204 10600
rect 23256 10588 23262 10600
rect 23661 10591 23719 10597
rect 23661 10588 23673 10591
rect 23256 10560 23673 10588
rect 23256 10548 23262 10560
rect 23661 10557 23673 10560
rect 23707 10588 23719 10591
rect 24320 10588 24348 10619
rect 23707 10560 24348 10588
rect 23707 10557 23719 10560
rect 23661 10551 23719 10557
rect 24670 10548 24676 10600
rect 24728 10588 24734 10600
rect 24857 10591 24915 10597
rect 24857 10588 24869 10591
rect 24728 10560 24869 10588
rect 24728 10548 24734 10560
rect 24857 10557 24869 10560
rect 24903 10557 24915 10591
rect 24857 10551 24915 10557
rect 22094 10520 22100 10532
rect 21008 10492 22100 10520
rect 22094 10480 22100 10492
rect 22152 10480 22158 10532
rect 17402 10452 17408 10464
rect 11808 10424 14780 10452
rect 17363 10424 17408 10452
rect 17402 10412 17408 10424
rect 17460 10412 17466 10464
rect 17770 10412 17776 10464
rect 17828 10452 17834 10464
rect 17865 10455 17923 10461
rect 17865 10452 17877 10455
rect 17828 10424 17877 10452
rect 17828 10412 17834 10424
rect 17865 10421 17877 10424
rect 17911 10452 17923 10455
rect 23845 10455 23903 10461
rect 23845 10452 23857 10455
rect 17911 10424 23857 10452
rect 17911 10421 17923 10424
rect 17865 10415 17923 10421
rect 23845 10421 23857 10424
rect 23891 10421 23903 10455
rect 23845 10415 23903 10421
rect 24765 10455 24823 10461
rect 24765 10421 24777 10455
rect 24811 10452 24823 10455
rect 24872 10452 24900 10551
rect 24946 10548 24952 10600
rect 25004 10588 25010 10600
rect 25332 10588 25360 10628
rect 25409 10625 25421 10659
rect 25455 10656 25467 10659
rect 27798 10656 27804 10668
rect 25455 10628 27804 10656
rect 25455 10625 25467 10628
rect 25409 10619 25467 10625
rect 27798 10616 27804 10628
rect 27856 10656 27862 10668
rect 27985 10659 28043 10665
rect 27985 10656 27997 10659
rect 27856 10628 27997 10656
rect 27856 10616 27862 10628
rect 27985 10625 27997 10628
rect 28031 10625 28043 10659
rect 27985 10619 28043 10625
rect 28445 10659 28503 10665
rect 28445 10625 28457 10659
rect 28491 10656 28503 10659
rect 29086 10656 29092 10668
rect 28491 10628 29092 10656
rect 28491 10625 28503 10628
rect 28445 10619 28503 10625
rect 25590 10588 25596 10600
rect 25004 10560 25049 10588
rect 25332 10560 25596 10588
rect 25004 10548 25010 10560
rect 25590 10548 25596 10560
rect 25648 10548 25654 10600
rect 25774 10548 25780 10600
rect 25832 10588 25838 10600
rect 26237 10591 26295 10597
rect 26237 10588 26249 10591
rect 25832 10560 26249 10588
rect 25832 10548 25838 10560
rect 26237 10557 26249 10560
rect 26283 10557 26295 10591
rect 26237 10551 26295 10557
rect 26697 10591 26755 10597
rect 26697 10557 26709 10591
rect 26743 10557 26755 10591
rect 26697 10551 26755 10557
rect 26973 10591 27031 10597
rect 26973 10557 26985 10591
rect 27019 10557 27031 10591
rect 27154 10588 27160 10600
rect 27115 10560 27160 10588
rect 26973 10551 27031 10557
rect 26142 10520 26148 10532
rect 26103 10492 26148 10520
rect 26142 10480 26148 10492
rect 26200 10520 26206 10532
rect 26712 10520 26740 10551
rect 26200 10492 26740 10520
rect 26988 10520 27016 10551
rect 27154 10548 27160 10560
rect 27212 10548 27218 10600
rect 27246 10548 27252 10600
rect 27304 10588 27310 10600
rect 27341 10591 27399 10597
rect 27341 10588 27353 10591
rect 27304 10560 27353 10588
rect 27304 10548 27310 10560
rect 27341 10557 27353 10560
rect 27387 10588 27399 10591
rect 27522 10588 27528 10600
rect 27387 10560 27528 10588
rect 27387 10557 27399 10560
rect 27341 10551 27399 10557
rect 27522 10548 27528 10560
rect 27580 10548 27586 10600
rect 27709 10591 27767 10597
rect 27709 10557 27721 10591
rect 27755 10588 27767 10591
rect 28460 10588 28488 10619
rect 29086 10616 29092 10628
rect 29144 10656 29150 10668
rect 29840 10665 29868 10696
rect 33778 10684 33784 10736
rect 33836 10724 33842 10736
rect 33836 10696 36124 10724
rect 33836 10684 33842 10696
rect 29273 10659 29331 10665
rect 29273 10656 29285 10659
rect 29144 10628 29285 10656
rect 29144 10616 29150 10628
rect 29273 10625 29285 10628
rect 29319 10625 29331 10659
rect 29273 10619 29331 10625
rect 29825 10659 29883 10665
rect 29825 10625 29837 10659
rect 29871 10625 29883 10659
rect 29825 10619 29883 10625
rect 32217 10659 32275 10665
rect 32217 10625 32229 10659
rect 32263 10656 32275 10659
rect 35621 10659 35679 10665
rect 32263 10628 32628 10656
rect 32263 10625 32275 10628
rect 32217 10619 32275 10625
rect 27755 10560 28488 10588
rect 27755 10557 27767 10560
rect 27709 10551 27767 10557
rect 29362 10548 29368 10600
rect 29420 10588 29426 10600
rect 30653 10591 30711 10597
rect 29420 10560 29465 10588
rect 29420 10548 29426 10560
rect 30653 10557 30665 10591
rect 30699 10588 30711 10591
rect 30926 10588 30932 10600
rect 30699 10560 30932 10588
rect 30699 10557 30711 10560
rect 30653 10551 30711 10557
rect 27614 10520 27620 10532
rect 26988 10492 27620 10520
rect 26200 10480 26206 10492
rect 27614 10480 27620 10492
rect 27672 10520 27678 10532
rect 28258 10520 28264 10532
rect 27672 10492 28264 10520
rect 27672 10480 27678 10492
rect 28258 10480 28264 10492
rect 28316 10480 28322 10532
rect 30668 10520 30696 10551
rect 30926 10548 30932 10560
rect 30984 10548 30990 10600
rect 32306 10548 32312 10600
rect 32364 10597 32370 10600
rect 32600 10597 32628 10628
rect 35621 10625 35633 10659
rect 35667 10656 35679 10659
rect 35986 10656 35992 10668
rect 35667 10628 35992 10656
rect 35667 10625 35679 10628
rect 35621 10619 35679 10625
rect 35986 10616 35992 10628
rect 36044 10616 36050 10668
rect 36096 10656 36124 10696
rect 39022 10684 39028 10736
rect 39080 10724 39086 10736
rect 40221 10727 40279 10733
rect 40221 10724 40233 10727
rect 39080 10696 40233 10724
rect 39080 10684 39086 10696
rect 40221 10693 40233 10696
rect 40267 10724 40279 10727
rect 40494 10724 40500 10736
rect 40267 10696 40500 10724
rect 40267 10693 40279 10696
rect 40221 10687 40279 10693
rect 40494 10684 40500 10696
rect 40552 10684 40558 10736
rect 43162 10724 43168 10736
rect 43123 10696 43168 10724
rect 43162 10684 43168 10696
rect 43220 10684 43226 10736
rect 43346 10684 43352 10736
rect 43404 10724 43410 10736
rect 43717 10727 43775 10733
rect 43717 10724 43729 10727
rect 43404 10696 43729 10724
rect 43404 10684 43410 10696
rect 43717 10693 43729 10696
rect 43763 10693 43775 10727
rect 44008 10724 44036 10764
rect 44542 10752 44548 10764
rect 44600 10752 44606 10804
rect 45094 10752 45100 10804
rect 45152 10792 45158 10804
rect 46385 10795 46443 10801
rect 46385 10792 46397 10795
rect 45152 10764 46397 10792
rect 45152 10752 45158 10764
rect 46385 10761 46397 10764
rect 46431 10792 46443 10795
rect 46658 10792 46664 10804
rect 46431 10764 46664 10792
rect 46431 10761 46443 10764
rect 46385 10755 46443 10761
rect 46658 10752 46664 10764
rect 46716 10752 46722 10804
rect 47305 10795 47363 10801
rect 47305 10761 47317 10795
rect 47351 10792 47363 10795
rect 47578 10792 47584 10804
rect 47351 10764 47584 10792
rect 47351 10761 47363 10764
rect 47305 10755 47363 10761
rect 47578 10752 47584 10764
rect 47636 10752 47642 10804
rect 47854 10792 47860 10804
rect 47815 10764 47860 10792
rect 47854 10752 47860 10764
rect 47912 10752 47918 10804
rect 48222 10752 48228 10804
rect 48280 10792 48286 10804
rect 50157 10795 50215 10801
rect 50157 10792 50169 10795
rect 48280 10764 50169 10792
rect 48280 10752 48286 10764
rect 50157 10761 50169 10764
rect 50203 10761 50215 10795
rect 51442 10792 51448 10804
rect 51403 10764 51448 10792
rect 50157 10755 50215 10761
rect 51442 10752 51448 10764
rect 51500 10752 51506 10804
rect 54938 10752 54944 10804
rect 54996 10792 55002 10804
rect 55125 10795 55183 10801
rect 55125 10792 55137 10795
rect 54996 10764 55137 10792
rect 54996 10752 55002 10764
rect 55125 10761 55137 10764
rect 55171 10761 55183 10795
rect 56134 10792 56140 10804
rect 56095 10764 56140 10792
rect 55125 10755 55183 10761
rect 47946 10724 47952 10736
rect 44008 10696 46244 10724
rect 43717 10687 43775 10693
rect 36446 10656 36452 10668
rect 36096 10628 36452 10656
rect 36446 10616 36452 10628
rect 36504 10616 36510 10668
rect 36722 10656 36728 10668
rect 36635 10628 36728 10656
rect 36722 10616 36728 10628
rect 36780 10656 36786 10668
rect 37090 10656 37096 10668
rect 36780 10628 37096 10656
rect 36780 10616 36786 10628
rect 37090 10616 37096 10628
rect 37148 10616 37154 10668
rect 39390 10656 39396 10668
rect 37200 10628 39160 10656
rect 39351 10628 39396 10656
rect 32364 10588 32374 10597
rect 32585 10591 32643 10597
rect 32364 10560 32409 10588
rect 32364 10551 32374 10560
rect 32585 10557 32597 10591
rect 32631 10588 32643 10591
rect 33686 10588 33692 10600
rect 32631 10560 33692 10588
rect 32631 10557 32643 10560
rect 32585 10551 32643 10557
rect 32364 10548 32370 10551
rect 33686 10548 33692 10560
rect 33744 10548 33750 10600
rect 34146 10548 34152 10600
rect 34204 10588 34210 10600
rect 34517 10591 34575 10597
rect 34517 10588 34529 10591
rect 34204 10560 34529 10588
rect 34204 10548 34210 10560
rect 34517 10557 34529 10560
rect 34563 10557 34575 10591
rect 34517 10551 34575 10557
rect 34698 10548 34704 10600
rect 34756 10588 34762 10600
rect 35253 10591 35311 10597
rect 35253 10588 35265 10591
rect 34756 10560 35265 10588
rect 34756 10548 34762 10560
rect 35253 10557 35265 10560
rect 35299 10588 35311 10591
rect 35897 10591 35955 10597
rect 35897 10588 35909 10591
rect 35299 10560 35909 10588
rect 35299 10557 35311 10560
rect 35253 10551 35311 10557
rect 35897 10557 35909 10560
rect 35943 10557 35955 10591
rect 37200 10588 37228 10628
rect 35897 10551 35955 10557
rect 36004 10560 37228 10588
rect 32030 10520 32036 10532
rect 28368 10492 30696 10520
rect 30852 10492 32036 10520
rect 25777 10455 25835 10461
rect 25777 10452 25789 10455
rect 24811 10424 25789 10452
rect 24811 10421 24823 10424
rect 24765 10415 24823 10421
rect 25777 10421 25789 10424
rect 25823 10452 25835 10455
rect 27062 10452 27068 10464
rect 25823 10424 27068 10452
rect 25823 10421 25835 10424
rect 25777 10415 25835 10421
rect 27062 10412 27068 10424
rect 27120 10412 27126 10464
rect 27154 10412 27160 10464
rect 27212 10452 27218 10464
rect 28368 10452 28396 10492
rect 30852 10464 30880 10492
rect 32030 10480 32036 10492
rect 32088 10480 32094 10532
rect 35066 10520 35072 10532
rect 33612 10492 35072 10520
rect 27212 10424 28396 10452
rect 28813 10455 28871 10461
rect 27212 10412 27218 10424
rect 28813 10421 28825 10455
rect 28859 10452 28871 10455
rect 28902 10452 28908 10464
rect 28859 10424 28908 10452
rect 28859 10421 28871 10424
rect 28813 10415 28871 10421
rect 28902 10412 28908 10424
rect 28960 10412 28966 10464
rect 30834 10452 30840 10464
rect 30795 10424 30840 10452
rect 30834 10412 30840 10424
rect 30892 10412 30898 10464
rect 31297 10455 31355 10461
rect 31297 10421 31309 10455
rect 31343 10452 31355 10455
rect 31570 10452 31576 10464
rect 31343 10424 31576 10452
rect 31343 10421 31355 10424
rect 31297 10415 31355 10421
rect 31570 10412 31576 10424
rect 31628 10412 31634 10464
rect 31849 10455 31907 10461
rect 31849 10421 31861 10455
rect 31895 10452 31907 10455
rect 33612 10452 33640 10492
rect 35066 10480 35072 10492
rect 35124 10480 35130 10532
rect 35802 10480 35808 10532
rect 35860 10520 35866 10532
rect 36004 10520 36032 10560
rect 38286 10548 38292 10600
rect 38344 10588 38350 10600
rect 38838 10588 38844 10600
rect 38344 10560 38844 10588
rect 38344 10548 38350 10560
rect 38838 10548 38844 10560
rect 38896 10548 38902 10600
rect 38933 10591 38991 10597
rect 38933 10557 38945 10591
rect 38979 10588 38991 10591
rect 39022 10588 39028 10600
rect 38979 10560 39028 10588
rect 38979 10557 38991 10560
rect 38933 10551 38991 10557
rect 39022 10548 39028 10560
rect 39080 10548 39086 10600
rect 39132 10597 39160 10628
rect 39390 10616 39396 10628
rect 39448 10616 39454 10668
rect 40589 10659 40647 10665
rect 40589 10625 40601 10659
rect 40635 10656 40647 10659
rect 41601 10659 41659 10665
rect 41601 10656 41613 10659
rect 40635 10628 41613 10656
rect 40635 10625 40647 10628
rect 40589 10619 40647 10625
rect 41601 10625 41613 10628
rect 41647 10656 41659 10659
rect 41690 10656 41696 10668
rect 41647 10628 41696 10656
rect 41647 10625 41659 10628
rect 41601 10619 41659 10625
rect 41690 10616 41696 10628
rect 41748 10616 41754 10668
rect 42058 10656 42064 10668
rect 42019 10628 42064 10656
rect 42058 10616 42064 10628
rect 42116 10616 42122 10668
rect 44269 10659 44327 10665
rect 44269 10625 44281 10659
rect 44315 10656 44327 10659
rect 44910 10656 44916 10668
rect 44315 10628 44916 10656
rect 44315 10625 44327 10628
rect 44269 10619 44327 10625
rect 44910 10616 44916 10628
rect 44968 10656 44974 10668
rect 45097 10659 45155 10665
rect 45097 10656 45109 10659
rect 44968 10628 45109 10656
rect 44968 10616 44974 10628
rect 45097 10625 45109 10628
rect 45143 10625 45155 10659
rect 45097 10619 45155 10625
rect 39117 10591 39175 10597
rect 39117 10557 39129 10591
rect 39163 10588 39175 10591
rect 39761 10591 39819 10597
rect 39761 10588 39773 10591
rect 39163 10560 39773 10588
rect 39163 10557 39175 10560
rect 39117 10551 39175 10557
rect 39761 10557 39773 10560
rect 39807 10557 39819 10591
rect 40678 10588 40684 10600
rect 40639 10560 40684 10588
rect 39761 10551 39819 10557
rect 40678 10548 40684 10560
rect 40736 10588 40742 10600
rect 41233 10591 41291 10597
rect 41233 10588 41245 10591
rect 40736 10560 41245 10588
rect 40736 10548 40742 10560
rect 41233 10557 41245 10560
rect 41279 10557 41291 10591
rect 41233 10551 41291 10557
rect 41785 10591 41843 10597
rect 41785 10557 41797 10591
rect 41831 10588 41843 10591
rect 42978 10588 42984 10600
rect 41831 10560 42984 10588
rect 41831 10557 41843 10560
rect 41785 10551 41843 10557
rect 42978 10548 42984 10560
rect 43036 10548 43042 10600
rect 44358 10588 44364 10600
rect 44319 10560 44364 10588
rect 44358 10548 44364 10560
rect 44416 10548 44422 10600
rect 46216 10597 46244 10696
rect 46768 10696 47952 10724
rect 46768 10597 46796 10696
rect 47946 10684 47952 10696
rect 48004 10684 48010 10736
rect 48314 10724 48320 10736
rect 48275 10696 48320 10724
rect 48314 10684 48320 10696
rect 48372 10684 48378 10736
rect 51350 10724 51356 10736
rect 49160 10696 51356 10724
rect 46934 10616 46940 10668
rect 46992 10656 46998 10668
rect 49160 10656 49188 10696
rect 51350 10684 51356 10696
rect 51408 10684 51414 10736
rect 51902 10724 51908 10736
rect 51863 10696 51908 10724
rect 51902 10684 51908 10696
rect 51960 10684 51966 10736
rect 55140 10724 55168 10755
rect 56134 10752 56140 10764
rect 56192 10752 56198 10804
rect 56778 10792 56784 10804
rect 56739 10764 56784 10792
rect 56778 10752 56784 10764
rect 56836 10752 56842 10804
rect 57606 10792 57612 10804
rect 57567 10764 57612 10792
rect 57606 10752 57612 10764
rect 57664 10752 57670 10804
rect 60458 10752 60464 10804
rect 60516 10792 60522 10804
rect 61197 10795 61255 10801
rect 61197 10792 61209 10795
rect 60516 10764 61209 10792
rect 60516 10752 60522 10764
rect 61197 10761 61209 10764
rect 61243 10761 61255 10795
rect 61197 10755 61255 10761
rect 60826 10724 60832 10736
rect 55140 10696 57468 10724
rect 60787 10696 60832 10724
rect 49326 10656 49332 10668
rect 46992 10628 49188 10656
rect 49287 10628 49332 10656
rect 46992 10616 46998 10628
rect 49326 10616 49332 10628
rect 49384 10656 49390 10668
rect 49384 10628 50016 10656
rect 49384 10616 49390 10628
rect 46201 10591 46259 10597
rect 46201 10557 46213 10591
rect 46247 10588 46259 10591
rect 46753 10591 46811 10597
rect 46753 10588 46765 10591
rect 46247 10560 46765 10588
rect 46247 10557 46259 10560
rect 46201 10551 46259 10557
rect 46753 10557 46765 10560
rect 46799 10557 46811 10591
rect 46753 10551 46811 10557
rect 47581 10591 47639 10597
rect 47581 10557 47593 10591
rect 47627 10557 47639 10591
rect 47581 10551 47639 10557
rect 48501 10591 48559 10597
rect 48501 10557 48513 10591
rect 48547 10588 48559 10591
rect 48590 10588 48596 10600
rect 48547 10560 48596 10588
rect 48547 10557 48559 10560
rect 48501 10551 48559 10557
rect 38654 10520 38660 10532
rect 35860 10492 36032 10520
rect 38028 10492 38660 10520
rect 35860 10480 35866 10492
rect 34330 10452 34336 10464
rect 31895 10424 33640 10452
rect 34291 10424 34336 10452
rect 31895 10421 31907 10424
rect 31849 10415 31907 10421
rect 34330 10412 34336 10424
rect 34388 10412 34394 10464
rect 34517 10455 34575 10461
rect 34517 10421 34529 10455
rect 34563 10452 34575 10455
rect 34701 10455 34759 10461
rect 34701 10452 34713 10455
rect 34563 10424 34713 10452
rect 34563 10421 34575 10424
rect 34517 10415 34575 10421
rect 34701 10421 34713 10424
rect 34747 10452 34759 10455
rect 36814 10452 36820 10464
rect 34747 10424 36820 10452
rect 34747 10421 34759 10424
rect 34701 10415 34759 10421
rect 36814 10412 36820 10424
rect 36872 10412 36878 10464
rect 37918 10412 37924 10464
rect 37976 10452 37982 10464
rect 38028 10461 38056 10492
rect 38654 10480 38660 10492
rect 38712 10480 38718 10532
rect 47596 10520 47624 10551
rect 48590 10548 48596 10560
rect 48648 10548 48654 10600
rect 48685 10591 48743 10597
rect 48685 10557 48697 10591
rect 48731 10588 48743 10591
rect 48774 10588 48780 10600
rect 48731 10560 48780 10588
rect 48731 10557 48743 10560
rect 48685 10551 48743 10557
rect 48774 10548 48780 10560
rect 48832 10548 48838 10600
rect 48866 10548 48872 10600
rect 48924 10588 48930 10600
rect 49418 10588 49424 10600
rect 48924 10560 49424 10588
rect 48924 10548 48930 10560
rect 49418 10548 49424 10560
rect 49476 10548 49482 10600
rect 49988 10597 50016 10628
rect 50338 10616 50344 10668
rect 50396 10656 50402 10668
rect 51077 10659 51135 10665
rect 51077 10656 51089 10659
rect 50396 10628 51089 10656
rect 50396 10616 50402 10628
rect 51077 10625 51089 10628
rect 51123 10625 51135 10659
rect 51077 10619 51135 10625
rect 51810 10616 51816 10668
rect 51868 10656 51874 10668
rect 53009 10659 53067 10665
rect 53009 10656 53021 10659
rect 51868 10628 53021 10656
rect 51868 10616 51874 10628
rect 53009 10625 53021 10628
rect 53055 10656 53067 10659
rect 53926 10656 53932 10668
rect 53055 10628 53932 10656
rect 53055 10625 53067 10628
rect 53009 10619 53067 10625
rect 53926 10616 53932 10628
rect 53984 10616 53990 10668
rect 57330 10656 57336 10668
rect 57291 10628 57336 10656
rect 57330 10616 57336 10628
rect 57388 10616 57394 10668
rect 49881 10591 49939 10597
rect 49881 10588 49893 10591
rect 49804 10560 49893 10588
rect 49602 10520 49608 10532
rect 45848 10492 47624 10520
rect 47872 10492 49608 10520
rect 45848 10464 45876 10492
rect 38013 10455 38071 10461
rect 38013 10452 38025 10455
rect 37976 10424 38025 10452
rect 37976 10412 37982 10424
rect 38013 10421 38025 10424
rect 38059 10421 38071 10455
rect 38746 10452 38752 10464
rect 38707 10424 38752 10452
rect 38013 10415 38071 10421
rect 38746 10412 38752 10424
rect 38804 10412 38810 10464
rect 38930 10412 38936 10464
rect 38988 10452 38994 10464
rect 40589 10455 40647 10461
rect 40589 10452 40601 10455
rect 38988 10424 40601 10452
rect 38988 10412 38994 10424
rect 40589 10421 40601 10424
rect 40635 10421 40647 10455
rect 40862 10452 40868 10464
rect 40823 10424 40868 10452
rect 40589 10415 40647 10421
rect 40862 10412 40868 10424
rect 40920 10412 40926 10464
rect 43530 10412 43536 10464
rect 43588 10452 43594 10464
rect 43898 10452 43904 10464
rect 43588 10424 43904 10452
rect 43588 10412 43594 10424
rect 43898 10412 43904 10424
rect 43956 10452 43962 10464
rect 44082 10452 44088 10464
rect 43956 10424 44088 10452
rect 43956 10412 43962 10424
rect 44082 10412 44088 10424
rect 44140 10412 44146 10464
rect 45462 10452 45468 10464
rect 45423 10424 45468 10452
rect 45462 10412 45468 10424
rect 45520 10412 45526 10464
rect 45830 10452 45836 10464
rect 45791 10424 45836 10452
rect 45830 10412 45836 10424
rect 45888 10412 45894 10464
rect 47394 10452 47400 10464
rect 47355 10424 47400 10452
rect 47394 10412 47400 10424
rect 47452 10412 47458 10464
rect 47578 10412 47584 10464
rect 47636 10452 47642 10464
rect 47872 10452 47900 10492
rect 49602 10480 49608 10492
rect 49660 10480 49666 10532
rect 47636 10424 47900 10452
rect 47636 10412 47642 10424
rect 47946 10412 47952 10464
rect 48004 10452 48010 10464
rect 49510 10452 49516 10464
rect 48004 10424 49516 10452
rect 48004 10412 48010 10424
rect 49510 10412 49516 10424
rect 49568 10412 49574 10464
rect 49804 10461 49832 10560
rect 49881 10557 49893 10560
rect 49927 10557 49939 10591
rect 49881 10551 49939 10557
rect 49973 10591 50031 10597
rect 49973 10557 49985 10591
rect 50019 10588 50031 10591
rect 50709 10591 50767 10597
rect 50709 10588 50721 10591
rect 50019 10560 50721 10588
rect 50019 10557 50031 10560
rect 49973 10551 50031 10557
rect 50709 10557 50721 10560
rect 50755 10557 50767 10591
rect 51718 10588 51724 10600
rect 51679 10560 51724 10588
rect 50709 10551 50767 10557
rect 51718 10548 51724 10560
rect 51776 10548 51782 10600
rect 53285 10591 53343 10597
rect 53285 10588 53297 10591
rect 53116 10560 53297 10588
rect 53116 10520 53144 10560
rect 53285 10557 53297 10560
rect 53331 10557 53343 10591
rect 53285 10551 53343 10557
rect 54478 10548 54484 10600
rect 54536 10588 54542 10600
rect 55490 10588 55496 10600
rect 54536 10560 55496 10588
rect 54536 10548 54542 10560
rect 55490 10548 55496 10560
rect 55548 10588 55554 10600
rect 55861 10591 55919 10597
rect 55861 10588 55873 10591
rect 55548 10560 55873 10588
rect 55548 10548 55554 10560
rect 55861 10557 55873 10560
rect 55907 10557 55919 10591
rect 55861 10551 55919 10557
rect 55950 10548 55956 10600
rect 56008 10588 56014 10600
rect 57440 10597 57468 10696
rect 60826 10684 60832 10696
rect 60884 10684 60890 10736
rect 59538 10656 59544 10668
rect 59499 10628 59544 10656
rect 59538 10616 59544 10628
rect 59596 10616 59602 10668
rect 57425 10591 57483 10597
rect 56008 10560 56101 10588
rect 56008 10548 56014 10560
rect 57425 10557 57437 10591
rect 57471 10588 57483 10591
rect 58161 10591 58219 10597
rect 58161 10588 58173 10591
rect 57471 10560 58173 10588
rect 57471 10557 57483 10560
rect 57425 10551 57483 10557
rect 58161 10557 58173 10560
rect 58207 10557 58219 10591
rect 58161 10551 58219 10557
rect 58342 10548 58348 10600
rect 58400 10588 58406 10600
rect 59262 10588 59268 10600
rect 58400 10560 59268 10588
rect 58400 10548 58406 10560
rect 59262 10548 59268 10560
rect 59320 10548 59326 10600
rect 53024 10492 53144 10520
rect 49789 10455 49847 10461
rect 49789 10421 49801 10455
rect 49835 10452 49847 10455
rect 51166 10452 51172 10464
rect 49835 10424 51172 10452
rect 49835 10421 49847 10424
rect 49789 10415 49847 10421
rect 51166 10412 51172 10424
rect 51224 10412 51230 10464
rect 52270 10452 52276 10464
rect 52231 10424 52276 10452
rect 52270 10412 52276 10424
rect 52328 10412 52334 10464
rect 52822 10452 52828 10464
rect 52783 10424 52828 10452
rect 52822 10412 52828 10424
rect 52880 10452 52886 10464
rect 53024 10452 53052 10492
rect 55398 10480 55404 10532
rect 55456 10520 55462 10532
rect 55968 10520 55996 10548
rect 56502 10520 56508 10532
rect 55456 10492 56508 10520
rect 55456 10480 55462 10492
rect 56502 10480 56508 10492
rect 56560 10480 56566 10532
rect 54386 10452 54392 10464
rect 52880 10424 53052 10452
rect 54347 10424 54392 10452
rect 52880 10412 52886 10424
rect 54386 10412 54392 10424
rect 54444 10412 54450 10464
rect 55769 10455 55827 10461
rect 55769 10421 55781 10455
rect 55815 10452 55827 10455
rect 56594 10452 56600 10464
rect 55815 10424 56600 10452
rect 55815 10421 55827 10424
rect 55769 10415 55827 10421
rect 56594 10412 56600 10424
rect 56652 10412 56658 10464
rect 58802 10452 58808 10464
rect 58763 10424 58808 10452
rect 58802 10412 58808 10424
rect 58860 10412 58866 10464
rect 59078 10452 59084 10464
rect 59039 10424 59084 10452
rect 59078 10412 59084 10424
rect 59136 10412 59142 10464
rect 61286 10412 61292 10464
rect 61344 10452 61350 10464
rect 61565 10455 61623 10461
rect 61565 10452 61577 10455
rect 61344 10424 61577 10452
rect 61344 10412 61350 10424
rect 61565 10421 61577 10424
rect 61611 10452 61623 10455
rect 61933 10455 61991 10461
rect 61933 10452 61945 10455
rect 61611 10424 61945 10452
rect 61611 10421 61623 10424
rect 61565 10415 61623 10421
rect 61933 10421 61945 10424
rect 61979 10421 61991 10455
rect 61933 10415 61991 10421
rect 1104 10362 63480 10384
rect 1104 10310 21774 10362
rect 21826 10310 21838 10362
rect 21890 10310 21902 10362
rect 21954 10310 21966 10362
rect 22018 10310 42566 10362
rect 42618 10310 42630 10362
rect 42682 10310 42694 10362
rect 42746 10310 42758 10362
rect 42810 10310 63480 10362
rect 1104 10288 63480 10310
rect 5442 10208 5448 10260
rect 5500 10248 5506 10260
rect 6733 10251 6791 10257
rect 6733 10248 6745 10251
rect 5500 10220 6745 10248
rect 5500 10208 5506 10220
rect 6733 10217 6745 10220
rect 6779 10217 6791 10251
rect 6733 10211 6791 10217
rect 8021 10251 8079 10257
rect 8021 10217 8033 10251
rect 8067 10248 8079 10251
rect 8665 10251 8723 10257
rect 8665 10248 8677 10251
rect 8067 10220 8677 10248
rect 8067 10217 8079 10220
rect 8021 10211 8079 10217
rect 8665 10217 8677 10220
rect 8711 10248 8723 10251
rect 8846 10248 8852 10260
rect 8711 10220 8852 10248
rect 8711 10217 8723 10220
rect 8665 10211 8723 10217
rect 8846 10208 8852 10220
rect 8904 10208 8910 10260
rect 13814 10248 13820 10260
rect 13775 10220 13820 10248
rect 13814 10208 13820 10220
rect 13872 10208 13878 10260
rect 14182 10248 14188 10260
rect 14143 10220 14188 10248
rect 14182 10208 14188 10220
rect 14240 10208 14246 10260
rect 14918 10248 14924 10260
rect 14879 10220 14924 10248
rect 14918 10208 14924 10220
rect 14976 10208 14982 10260
rect 15470 10208 15476 10260
rect 15528 10248 15534 10260
rect 15841 10251 15899 10257
rect 15841 10248 15853 10251
rect 15528 10220 15853 10248
rect 15528 10208 15534 10220
rect 15841 10217 15853 10220
rect 15887 10217 15899 10251
rect 15841 10211 15899 10217
rect 16390 10208 16396 10260
rect 16448 10248 16454 10260
rect 20070 10248 20076 10260
rect 16448 10220 20076 10248
rect 16448 10208 16454 10220
rect 20070 10208 20076 10220
rect 20128 10208 20134 10260
rect 20257 10251 20315 10257
rect 20257 10217 20269 10251
rect 20303 10248 20315 10251
rect 20438 10248 20444 10260
rect 20303 10220 20444 10248
rect 20303 10217 20315 10220
rect 20257 10211 20315 10217
rect 20438 10208 20444 10220
rect 20496 10208 20502 10260
rect 21174 10208 21180 10260
rect 21232 10248 21238 10260
rect 22925 10251 22983 10257
rect 21232 10220 22876 10248
rect 21232 10208 21238 10220
rect 7466 10140 7472 10192
rect 7524 10180 7530 10192
rect 10229 10183 10287 10189
rect 10229 10180 10241 10183
rect 7524 10152 10241 10180
rect 7524 10140 7530 10152
rect 10229 10149 10241 10152
rect 10275 10149 10287 10183
rect 10229 10143 10287 10149
rect 13081 10183 13139 10189
rect 13081 10149 13093 10183
rect 13127 10180 13139 10183
rect 14936 10180 14964 10208
rect 13127 10152 14964 10180
rect 13127 10149 13139 10152
rect 13081 10143 13139 10149
rect 15102 10140 15108 10192
rect 15160 10180 15166 10192
rect 15160 10152 18092 10180
rect 15160 10140 15166 10152
rect 4246 10072 4252 10124
rect 4304 10112 4310 10124
rect 4433 10115 4491 10121
rect 4433 10112 4445 10115
rect 4304 10084 4445 10112
rect 4304 10072 4310 10084
rect 4433 10081 4445 10084
rect 4479 10112 4491 10115
rect 4798 10112 4804 10124
rect 4479 10084 4804 10112
rect 4479 10081 4491 10084
rect 4433 10075 4491 10081
rect 4798 10072 4804 10084
rect 4856 10072 4862 10124
rect 4982 10072 4988 10124
rect 5040 10112 5046 10124
rect 6917 10115 6975 10121
rect 6917 10112 6929 10115
rect 5040 10084 6929 10112
rect 5040 10072 5046 10084
rect 6917 10081 6929 10084
rect 6963 10081 6975 10115
rect 6917 10075 6975 10081
rect 7377 10115 7435 10121
rect 7377 10081 7389 10115
rect 7423 10081 7435 10115
rect 7377 10075 7435 10081
rect 7745 10115 7803 10121
rect 7745 10081 7757 10115
rect 7791 10112 7803 10115
rect 8021 10115 8079 10121
rect 8021 10112 8033 10115
rect 7791 10084 8033 10112
rect 7791 10081 7803 10084
rect 7745 10075 7803 10081
rect 8021 10081 8033 10084
rect 8067 10081 8079 10115
rect 8021 10075 8079 10081
rect 9493 10115 9551 10121
rect 9493 10081 9505 10115
rect 9539 10112 9551 10115
rect 9766 10112 9772 10124
rect 9539 10084 9772 10112
rect 9539 10081 9551 10084
rect 9493 10075 9551 10081
rect 4706 10044 4712 10056
rect 4667 10016 4712 10044
rect 4706 10004 4712 10016
rect 4764 10004 4770 10056
rect 5718 10004 5724 10056
rect 5776 10044 5782 10056
rect 5813 10047 5871 10053
rect 5813 10044 5825 10047
rect 5776 10016 5825 10044
rect 5776 10004 5782 10016
rect 5813 10013 5825 10016
rect 5859 10044 5871 10047
rect 7282 10044 7288 10056
rect 5859 10016 7288 10044
rect 5859 10013 5871 10016
rect 5813 10007 5871 10013
rect 7282 10004 7288 10016
rect 7340 10004 7346 10056
rect 7392 9976 7420 10075
rect 9766 10072 9772 10084
rect 9824 10112 9830 10124
rect 10870 10112 10876 10124
rect 9824 10084 10876 10112
rect 9824 10072 9830 10084
rect 10870 10072 10876 10084
rect 10928 10072 10934 10124
rect 11701 10115 11759 10121
rect 11701 10081 11713 10115
rect 11747 10112 11759 10115
rect 11790 10112 11796 10124
rect 11747 10084 11796 10112
rect 11747 10081 11759 10084
rect 11701 10075 11759 10081
rect 11790 10072 11796 10084
rect 11848 10072 11854 10124
rect 14366 10072 14372 10124
rect 14424 10112 14430 10124
rect 15120 10112 15148 10140
rect 14424 10084 15148 10112
rect 15289 10115 15347 10121
rect 14424 10072 14430 10084
rect 15289 10081 15301 10115
rect 15335 10112 15347 10115
rect 16022 10112 16028 10124
rect 15335 10084 16028 10112
rect 15335 10081 15347 10084
rect 15289 10075 15347 10081
rect 16022 10072 16028 10084
rect 16080 10072 16086 10124
rect 17037 10115 17095 10121
rect 17037 10081 17049 10115
rect 17083 10112 17095 10115
rect 17402 10112 17408 10124
rect 17083 10084 17408 10112
rect 17083 10081 17095 10084
rect 17037 10075 17095 10081
rect 17402 10072 17408 10084
rect 17460 10112 17466 10124
rect 17770 10112 17776 10124
rect 17460 10084 17776 10112
rect 17460 10072 17466 10084
rect 17770 10072 17776 10084
rect 17828 10072 17834 10124
rect 7834 10044 7840 10056
rect 7747 10016 7840 10044
rect 7834 10004 7840 10016
rect 7892 10044 7898 10056
rect 8297 10047 8355 10053
rect 8297 10044 8309 10047
rect 7892 10016 8309 10044
rect 7892 10004 7898 10016
rect 8297 10013 8309 10016
rect 8343 10044 8355 10047
rect 9674 10044 9680 10056
rect 8343 10016 9536 10044
rect 9635 10016 9680 10044
rect 8343 10013 8355 10016
rect 8297 10007 8355 10013
rect 8938 9976 8944 9988
rect 7392 9948 8944 9976
rect 8938 9936 8944 9948
rect 8996 9936 9002 9988
rect 9508 9976 9536 10016
rect 9674 10004 9680 10016
rect 9732 10004 9738 10056
rect 9950 10004 9956 10056
rect 10008 10044 10014 10056
rect 11425 10047 11483 10053
rect 11425 10044 11437 10047
rect 10008 10016 11437 10044
rect 10008 10004 10014 10016
rect 11425 10013 11437 10016
rect 11471 10044 11483 10047
rect 12066 10044 12072 10056
rect 11471 10016 12072 10044
rect 11471 10013 11483 10016
rect 11425 10007 11483 10013
rect 12066 10004 12072 10016
rect 12124 10004 12130 10056
rect 12710 10004 12716 10056
rect 12768 10044 12774 10056
rect 13722 10044 13728 10056
rect 12768 10016 13728 10044
rect 12768 10004 12774 10016
rect 13722 10004 13728 10016
rect 13780 10044 13786 10056
rect 14553 10047 14611 10053
rect 14553 10044 14565 10047
rect 13780 10016 14565 10044
rect 13780 10004 13786 10016
rect 14553 10013 14565 10016
rect 14599 10013 14611 10047
rect 14553 10007 14611 10013
rect 16945 10047 17003 10053
rect 16945 10013 16957 10047
rect 16991 10013 17003 10047
rect 16945 10007 17003 10013
rect 17497 10047 17555 10053
rect 17497 10013 17509 10047
rect 17543 10044 17555 10047
rect 17954 10044 17960 10056
rect 17543 10016 17960 10044
rect 17543 10013 17555 10016
rect 17497 10007 17555 10013
rect 10686 9976 10692 9988
rect 9508 9948 10692 9976
rect 10686 9936 10692 9948
rect 10744 9936 10750 9988
rect 15473 9979 15531 9985
rect 15473 9945 15485 9979
rect 15519 9976 15531 9979
rect 15562 9976 15568 9988
rect 15519 9948 15568 9976
rect 15519 9945 15531 9948
rect 15473 9939 15531 9945
rect 15562 9936 15568 9948
rect 15620 9936 15626 9988
rect 16960 9976 16988 10007
rect 17954 10004 17960 10016
rect 18012 10004 18018 10056
rect 18064 10044 18092 10152
rect 18230 10140 18236 10192
rect 18288 10180 18294 10192
rect 18288 10152 18460 10180
rect 18288 10140 18294 10152
rect 18322 10112 18328 10124
rect 18283 10084 18328 10112
rect 18322 10072 18328 10084
rect 18380 10072 18386 10124
rect 18432 10112 18460 10152
rect 20346 10140 20352 10192
rect 20404 10180 20410 10192
rect 20901 10183 20959 10189
rect 20901 10180 20913 10183
rect 20404 10152 20913 10180
rect 20404 10140 20410 10152
rect 20901 10149 20913 10152
rect 20947 10149 20959 10183
rect 22848 10180 22876 10220
rect 22925 10217 22937 10251
rect 22971 10248 22983 10251
rect 23014 10248 23020 10260
rect 22971 10220 23020 10248
rect 22971 10217 22983 10220
rect 22925 10211 22983 10217
rect 23014 10208 23020 10220
rect 23072 10208 23078 10260
rect 24121 10251 24179 10257
rect 24121 10217 24133 10251
rect 24167 10248 24179 10251
rect 24210 10248 24216 10260
rect 24167 10220 24216 10248
rect 24167 10217 24179 10220
rect 24121 10211 24179 10217
rect 24136 10180 24164 10211
rect 24210 10208 24216 10220
rect 24268 10208 24274 10260
rect 24854 10248 24860 10260
rect 24815 10220 24860 10248
rect 24854 10208 24860 10220
rect 24912 10208 24918 10260
rect 26326 10248 26332 10260
rect 26287 10220 26332 10248
rect 26326 10208 26332 10220
rect 26384 10208 26390 10260
rect 27065 10251 27123 10257
rect 27065 10217 27077 10251
rect 27111 10248 27123 10251
rect 27614 10248 27620 10260
rect 27111 10220 27620 10248
rect 27111 10217 27123 10220
rect 27065 10211 27123 10217
rect 27614 10208 27620 10220
rect 27672 10208 27678 10260
rect 27706 10208 27712 10260
rect 27764 10248 27770 10260
rect 30834 10248 30840 10260
rect 27764 10220 30840 10248
rect 27764 10208 27770 10220
rect 30834 10208 30840 10220
rect 30892 10208 30898 10260
rect 32582 10248 32588 10260
rect 32543 10220 32588 10248
rect 32582 10208 32588 10220
rect 32640 10208 32646 10260
rect 35066 10208 35072 10260
rect 35124 10248 35130 10260
rect 44085 10251 44143 10257
rect 35124 10220 44036 10248
rect 35124 10208 35130 10220
rect 20901 10143 20959 10149
rect 21284 10152 21588 10180
rect 22848 10152 24164 10180
rect 24581 10183 24639 10189
rect 18601 10115 18659 10121
rect 18601 10112 18613 10115
rect 18432 10084 18613 10112
rect 18601 10081 18613 10084
rect 18647 10081 18659 10115
rect 18601 10075 18659 10081
rect 20806 10072 20812 10124
rect 20864 10112 20870 10124
rect 21284 10112 21312 10152
rect 21560 10121 21588 10152
rect 24581 10149 24593 10183
rect 24627 10180 24639 10183
rect 26050 10180 26056 10192
rect 24627 10152 26056 10180
rect 24627 10149 24639 10152
rect 24581 10143 24639 10149
rect 20864 10084 21312 10112
rect 21361 10115 21419 10121
rect 20864 10072 20870 10084
rect 21361 10081 21373 10115
rect 21407 10081 21419 10115
rect 21361 10075 21419 10081
rect 21545 10115 21603 10121
rect 21545 10081 21557 10115
rect 21591 10081 21603 10115
rect 21545 10075 21603 10081
rect 21729 10115 21787 10121
rect 21729 10081 21741 10115
rect 21775 10112 21787 10115
rect 22094 10112 22100 10124
rect 21775 10084 22100 10112
rect 21775 10081 21787 10084
rect 21729 10075 21787 10081
rect 20990 10044 20996 10056
rect 18064 10016 20996 10044
rect 20990 10004 20996 10016
rect 21048 10004 21054 10056
rect 21376 10044 21404 10075
rect 22094 10072 22100 10084
rect 22152 10112 22158 10124
rect 22557 10115 22615 10121
rect 22557 10112 22569 10115
rect 22152 10084 22569 10112
rect 22152 10072 22158 10084
rect 22557 10081 22569 10084
rect 22603 10081 22615 10115
rect 22557 10075 22615 10081
rect 22741 10115 22799 10121
rect 22741 10081 22753 10115
rect 22787 10112 22799 10115
rect 23198 10112 23204 10124
rect 22787 10084 23204 10112
rect 22787 10081 22799 10084
rect 22741 10075 22799 10081
rect 23198 10072 23204 10084
rect 23256 10072 23262 10124
rect 23937 10115 23995 10121
rect 23937 10081 23949 10115
rect 23983 10112 23995 10115
rect 24596 10112 24624 10143
rect 26050 10140 26056 10152
rect 26108 10140 26114 10192
rect 27801 10183 27859 10189
rect 27801 10149 27813 10183
rect 27847 10180 27859 10183
rect 27890 10180 27896 10192
rect 27847 10152 27896 10180
rect 27847 10149 27859 10152
rect 27801 10143 27859 10149
rect 27890 10140 27896 10152
rect 27948 10140 27954 10192
rect 29178 10180 29184 10192
rect 28000 10152 28856 10180
rect 29139 10152 29184 10180
rect 23983 10084 24624 10112
rect 25133 10115 25191 10121
rect 23983 10081 23995 10084
rect 23937 10075 23995 10081
rect 25133 10081 25145 10115
rect 25179 10112 25191 10115
rect 25869 10115 25927 10121
rect 25869 10112 25881 10115
rect 25179 10084 25881 10112
rect 25179 10081 25191 10084
rect 25133 10075 25191 10081
rect 25869 10081 25881 10084
rect 25915 10112 25927 10115
rect 27341 10115 27399 10121
rect 27341 10112 27353 10115
rect 25915 10084 27353 10112
rect 25915 10081 25927 10084
rect 25869 10075 25927 10081
rect 27341 10081 27353 10084
rect 27387 10112 27399 10115
rect 27430 10112 27436 10124
rect 27387 10084 27436 10112
rect 27387 10081 27399 10084
rect 27341 10075 27399 10081
rect 27430 10072 27436 10084
rect 27488 10072 27494 10124
rect 22186 10044 22192 10056
rect 21376 10016 22192 10044
rect 22186 10004 22192 10016
rect 22244 10004 22250 10056
rect 24765 10047 24823 10053
rect 24765 10013 24777 10047
rect 24811 10044 24823 10047
rect 25041 10047 25099 10053
rect 25041 10044 25053 10047
rect 24811 10016 25053 10044
rect 24811 10013 24823 10016
rect 24765 10007 24823 10013
rect 25041 10013 25053 10016
rect 25087 10013 25099 10047
rect 27246 10044 27252 10056
rect 27207 10016 27252 10044
rect 25041 10007 25099 10013
rect 27246 10004 27252 10016
rect 27304 10004 27310 10056
rect 17586 9976 17592 9988
rect 16960 9948 17592 9976
rect 17586 9936 17592 9948
rect 17644 9936 17650 9988
rect 21174 9976 21180 9988
rect 17696 9948 18368 9976
rect 4154 9868 4160 9920
rect 4212 9908 4218 9920
rect 4249 9911 4307 9917
rect 4249 9908 4261 9911
rect 4212 9880 4261 9908
rect 4212 9868 4218 9880
rect 4249 9877 4261 9880
rect 4295 9877 4307 9911
rect 6362 9908 6368 9920
rect 6323 9880 6368 9908
rect 4249 9871 4307 9877
rect 6362 9868 6368 9880
rect 6420 9868 6426 9920
rect 9125 9911 9183 9917
rect 9125 9877 9137 9911
rect 9171 9908 9183 9911
rect 9306 9908 9312 9920
rect 9171 9880 9312 9908
rect 9171 9877 9183 9880
rect 9125 9871 9183 9877
rect 9306 9868 9312 9880
rect 9364 9868 9370 9920
rect 10502 9908 10508 9920
rect 10463 9880 10508 9908
rect 10502 9868 10508 9880
rect 10560 9868 10566 9920
rect 10870 9868 10876 9920
rect 10928 9908 10934 9920
rect 11057 9911 11115 9917
rect 11057 9908 11069 9911
rect 10928 9880 11069 9908
rect 10928 9868 10934 9880
rect 11057 9877 11069 9880
rect 11103 9877 11115 9911
rect 11057 9871 11115 9877
rect 12894 9868 12900 9920
rect 12952 9908 12958 9920
rect 13357 9911 13415 9917
rect 13357 9908 13369 9911
rect 12952 9880 13369 9908
rect 12952 9868 12958 9880
rect 13357 9877 13369 9880
rect 13403 9877 13415 9911
rect 13357 9871 13415 9877
rect 15194 9868 15200 9920
rect 15252 9908 15258 9920
rect 16298 9908 16304 9920
rect 15252 9880 16304 9908
rect 15252 9868 15258 9880
rect 16298 9868 16304 9880
rect 16356 9868 16362 9920
rect 16666 9908 16672 9920
rect 16627 9880 16672 9908
rect 16666 9868 16672 9880
rect 16724 9908 16730 9920
rect 17696 9908 17724 9948
rect 16724 9880 17724 9908
rect 16724 9868 16730 9880
rect 17770 9868 17776 9920
rect 17828 9908 17834 9920
rect 17828 9880 17873 9908
rect 17828 9868 17834 9880
rect 18046 9868 18052 9920
rect 18104 9908 18110 9920
rect 18141 9911 18199 9917
rect 18141 9908 18153 9911
rect 18104 9880 18153 9908
rect 18104 9868 18110 9880
rect 18141 9877 18153 9880
rect 18187 9877 18199 9911
rect 18340 9908 18368 9948
rect 19260 9948 21180 9976
rect 19260 9908 19288 9948
rect 21174 9936 21180 9948
rect 21232 9936 21238 9988
rect 22462 9936 22468 9988
rect 22520 9976 22526 9988
rect 23385 9979 23443 9985
rect 23385 9976 23397 9979
rect 22520 9948 23397 9976
rect 22520 9936 22526 9948
rect 23385 9945 23397 9948
rect 23431 9976 23443 9979
rect 26326 9976 26332 9988
rect 23431 9948 26332 9976
rect 23431 9945 23443 9948
rect 23385 9939 23443 9945
rect 26326 9936 26332 9948
rect 26384 9936 26390 9988
rect 28000 9976 28028 10152
rect 28721 10115 28779 10121
rect 28721 10081 28733 10115
rect 28767 10081 28779 10115
rect 28721 10075 28779 10081
rect 28629 10047 28687 10053
rect 28629 10013 28641 10047
rect 28675 10013 28687 10047
rect 28629 10007 28687 10013
rect 26436 9948 28028 9976
rect 18340 9880 19288 9908
rect 18141 9871 18199 9877
rect 19334 9868 19340 9920
rect 19392 9908 19398 9920
rect 19702 9908 19708 9920
rect 19392 9880 19708 9908
rect 19392 9868 19398 9880
rect 19702 9868 19708 9880
rect 19760 9868 19766 9920
rect 20714 9908 20720 9920
rect 20675 9880 20720 9908
rect 20714 9868 20720 9880
rect 20772 9868 20778 9920
rect 21358 9868 21364 9920
rect 21416 9908 21422 9920
rect 21726 9908 21732 9920
rect 21416 9880 21732 9908
rect 21416 9868 21422 9880
rect 21726 9868 21732 9880
rect 21784 9868 21790 9920
rect 23845 9911 23903 9917
rect 23845 9877 23857 9911
rect 23891 9908 23903 9911
rect 23934 9908 23940 9920
rect 23891 9880 23940 9908
rect 23891 9877 23903 9880
rect 23845 9871 23903 9877
rect 23934 9868 23940 9880
rect 23992 9908 23998 9920
rect 24765 9911 24823 9917
rect 24765 9908 24777 9911
rect 23992 9880 24777 9908
rect 23992 9868 23998 9880
rect 24765 9877 24777 9880
rect 24811 9877 24823 9911
rect 25314 9908 25320 9920
rect 25275 9880 25320 9908
rect 24765 9871 24823 9877
rect 25314 9868 25320 9880
rect 25372 9868 25378 9920
rect 25590 9868 25596 9920
rect 25648 9908 25654 9920
rect 26436 9908 26464 9948
rect 25648 9880 26464 9908
rect 25648 9868 25654 9880
rect 27522 9868 27528 9920
rect 27580 9908 27586 9920
rect 28077 9911 28135 9917
rect 28077 9908 28089 9911
rect 27580 9880 28089 9908
rect 27580 9868 27586 9880
rect 28077 9877 28089 9880
rect 28123 9877 28135 9911
rect 28077 9871 28135 9877
rect 28350 9868 28356 9920
rect 28408 9908 28414 9920
rect 28445 9911 28503 9917
rect 28445 9908 28457 9911
rect 28408 9880 28457 9908
rect 28408 9868 28414 9880
rect 28445 9877 28457 9880
rect 28491 9877 28503 9911
rect 28644 9908 28672 10007
rect 28736 9988 28764 10075
rect 28828 10044 28856 10152
rect 29178 10140 29184 10152
rect 29236 10140 29242 10192
rect 34330 10140 34336 10192
rect 34388 10180 34394 10192
rect 35621 10183 35679 10189
rect 35621 10180 35633 10183
rect 34388 10152 35633 10180
rect 34388 10140 34394 10152
rect 35621 10149 35633 10152
rect 35667 10149 35679 10183
rect 38930 10180 38936 10192
rect 35621 10143 35679 10149
rect 38856 10152 38936 10180
rect 30009 10115 30067 10121
rect 30009 10081 30021 10115
rect 30055 10112 30067 10115
rect 30282 10112 30288 10124
rect 30055 10084 30288 10112
rect 30055 10081 30067 10084
rect 30009 10075 30067 10081
rect 30282 10072 30288 10084
rect 30340 10072 30346 10124
rect 31389 10115 31447 10121
rect 31389 10081 31401 10115
rect 31435 10112 31447 10115
rect 32125 10115 32183 10121
rect 32125 10112 32137 10115
rect 31435 10084 32137 10112
rect 31435 10081 31447 10084
rect 31389 10075 31447 10081
rect 32125 10081 32137 10084
rect 32171 10081 32183 10115
rect 32125 10075 32183 10081
rect 32217 10115 32275 10121
rect 32217 10081 32229 10115
rect 32263 10112 32275 10115
rect 33226 10112 33232 10124
rect 32263 10084 33232 10112
rect 32263 10081 32275 10084
rect 32217 10075 32275 10081
rect 31570 10044 31576 10056
rect 28828 10016 31576 10044
rect 31570 10004 31576 10016
rect 31628 10004 31634 10056
rect 28718 9936 28724 9988
rect 28776 9976 28782 9988
rect 30193 9979 30251 9985
rect 30193 9976 30205 9979
rect 28776 9948 30205 9976
rect 28776 9936 28782 9948
rect 30193 9945 30205 9948
rect 30239 9945 30251 9979
rect 32140 9976 32168 10075
rect 33226 10072 33232 10084
rect 33284 10072 33290 10124
rect 36078 10112 36084 10124
rect 36039 10084 36084 10112
rect 36078 10072 36084 10084
rect 36136 10072 36142 10124
rect 36449 10115 36507 10121
rect 36449 10081 36461 10115
rect 36495 10112 36507 10115
rect 37277 10115 37335 10121
rect 37277 10112 37289 10115
rect 36495 10084 37289 10112
rect 36495 10081 36507 10084
rect 36449 10075 36507 10081
rect 37277 10081 37289 10084
rect 37323 10081 37335 10115
rect 38654 10112 38660 10124
rect 38615 10084 38660 10112
rect 37277 10075 37335 10081
rect 32306 10004 32312 10056
rect 32364 10044 32370 10056
rect 33134 10044 33140 10056
rect 32364 10016 33140 10044
rect 32364 10004 32370 10016
rect 33134 10004 33140 10016
rect 33192 10004 33198 10056
rect 33413 10047 33471 10053
rect 33413 10013 33425 10047
rect 33459 10044 33471 10047
rect 33502 10044 33508 10056
rect 33459 10016 33508 10044
rect 33459 10013 33471 10016
rect 33413 10007 33471 10013
rect 33502 10004 33508 10016
rect 33560 10004 33566 10056
rect 35434 10004 35440 10056
rect 35492 10044 35498 10056
rect 36464 10044 36492 10075
rect 38654 10072 38660 10084
rect 38712 10072 38718 10124
rect 38856 10121 38884 10152
rect 38930 10140 38936 10152
rect 38988 10140 38994 10192
rect 39850 10180 39856 10192
rect 39811 10152 39856 10180
rect 39850 10140 39856 10152
rect 39908 10140 39914 10192
rect 41598 10180 41604 10192
rect 39960 10152 41604 10180
rect 38841 10115 38899 10121
rect 38841 10081 38853 10115
rect 38887 10081 38899 10115
rect 39022 10112 39028 10124
rect 38983 10084 39028 10112
rect 38841 10075 38899 10081
rect 39022 10072 39028 10084
rect 39080 10072 39086 10124
rect 35492 10016 36492 10044
rect 35492 10004 35498 10016
rect 36538 10004 36544 10056
rect 36596 10044 36602 10056
rect 36596 10016 36641 10044
rect 36596 10004 36602 10016
rect 36814 10004 36820 10056
rect 36872 10044 36878 10056
rect 39960 10044 39988 10152
rect 41598 10140 41604 10152
rect 41656 10140 41662 10192
rect 41966 10180 41972 10192
rect 41708 10152 41972 10180
rect 40405 10115 40463 10121
rect 40405 10081 40417 10115
rect 40451 10081 40463 10115
rect 40405 10075 40463 10081
rect 40865 10115 40923 10121
rect 40865 10081 40877 10115
rect 40911 10112 40923 10115
rect 41708 10112 41736 10152
rect 41966 10140 41972 10152
rect 42024 10140 42030 10192
rect 44008 10180 44036 10220
rect 44085 10217 44097 10251
rect 44131 10248 44143 10251
rect 45830 10248 45836 10260
rect 44131 10220 45836 10248
rect 44131 10217 44143 10220
rect 44085 10211 44143 10217
rect 45830 10208 45836 10220
rect 45888 10208 45894 10260
rect 46845 10251 46903 10257
rect 46845 10217 46857 10251
rect 46891 10248 46903 10251
rect 47302 10248 47308 10260
rect 46891 10220 47308 10248
rect 46891 10217 46903 10220
rect 46845 10211 46903 10217
rect 47302 10208 47308 10220
rect 47360 10208 47366 10260
rect 47762 10208 47768 10260
rect 47820 10248 47826 10260
rect 47949 10251 48007 10257
rect 47949 10248 47961 10251
rect 47820 10220 47961 10248
rect 47820 10208 47826 10220
rect 47949 10217 47961 10220
rect 47995 10217 48007 10251
rect 48314 10248 48320 10260
rect 48275 10220 48320 10248
rect 47949 10211 48007 10217
rect 48314 10208 48320 10220
rect 48372 10208 48378 10260
rect 49602 10208 49608 10260
rect 49660 10248 49666 10260
rect 50430 10248 50436 10260
rect 49660 10220 50436 10248
rect 49660 10208 49666 10220
rect 50430 10208 50436 10220
rect 50488 10208 50494 10260
rect 50893 10251 50951 10257
rect 50893 10217 50905 10251
rect 50939 10248 50951 10251
rect 51074 10248 51080 10260
rect 50939 10220 51080 10248
rect 50939 10217 50951 10220
rect 50893 10211 50951 10217
rect 51074 10208 51080 10220
rect 51132 10248 51138 10260
rect 51994 10248 52000 10260
rect 51132 10220 52000 10248
rect 51132 10208 51138 10220
rect 51994 10208 52000 10220
rect 52052 10208 52058 10260
rect 53926 10248 53932 10260
rect 53887 10220 53932 10248
rect 53926 10208 53932 10220
rect 53984 10208 53990 10260
rect 54389 10251 54447 10257
rect 54389 10217 54401 10251
rect 54435 10248 54447 10251
rect 54478 10248 54484 10260
rect 54435 10220 54484 10248
rect 54435 10217 54447 10220
rect 54389 10211 54447 10217
rect 54478 10208 54484 10220
rect 54536 10208 54542 10260
rect 54849 10251 54907 10257
rect 54849 10217 54861 10251
rect 54895 10248 54907 10251
rect 54938 10248 54944 10260
rect 54895 10220 54944 10248
rect 54895 10217 54907 10220
rect 54849 10211 54907 10217
rect 54938 10208 54944 10220
rect 54996 10208 55002 10260
rect 55766 10248 55772 10260
rect 55727 10220 55772 10248
rect 55766 10208 55772 10220
rect 55824 10248 55830 10260
rect 56321 10251 56379 10257
rect 55824 10220 56272 10248
rect 55824 10208 55830 10220
rect 46014 10180 46020 10192
rect 44008 10152 45232 10180
rect 45927 10152 46020 10180
rect 40911 10084 41736 10112
rect 40911 10081 40923 10084
rect 40865 10075 40923 10081
rect 40310 10044 40316 10056
rect 36872 10016 39988 10044
rect 40271 10016 40316 10044
rect 36872 10004 36878 10016
rect 40310 10004 40316 10016
rect 40368 10004 40374 10056
rect 40420 10044 40448 10075
rect 41782 10072 41788 10124
rect 41840 10112 41846 10124
rect 41840 10084 41885 10112
rect 41840 10072 41846 10084
rect 43898 10072 43904 10124
rect 43956 10112 43962 10124
rect 44269 10115 44327 10121
rect 44269 10112 44281 10115
rect 43956 10084 44281 10112
rect 43956 10072 43962 10084
rect 44269 10081 44281 10084
rect 44315 10081 44327 10115
rect 44818 10112 44824 10124
rect 44779 10084 44824 10112
rect 44269 10075 44327 10081
rect 44818 10072 44824 10084
rect 44876 10072 44882 10124
rect 45204 10121 45232 10152
rect 46014 10140 46020 10152
rect 46072 10180 46078 10192
rect 47394 10180 47400 10192
rect 46072 10152 47400 10180
rect 46072 10140 46078 10152
rect 47394 10140 47400 10152
rect 47452 10180 47458 10192
rect 47452 10152 51120 10180
rect 47452 10140 47458 10152
rect 45189 10115 45247 10121
rect 45189 10081 45201 10115
rect 45235 10112 45247 10115
rect 45554 10112 45560 10124
rect 45235 10084 45560 10112
rect 45235 10081 45247 10084
rect 45189 10075 45247 10081
rect 45554 10072 45560 10084
rect 45612 10072 45618 10124
rect 46658 10112 46664 10124
rect 46619 10084 46664 10112
rect 46658 10072 46664 10084
rect 46716 10072 46722 10124
rect 47578 10112 47584 10124
rect 47136 10084 47584 10112
rect 41046 10044 41052 10056
rect 40420 10016 41052 10044
rect 41046 10004 41052 10016
rect 41104 10044 41110 10056
rect 41141 10047 41199 10053
rect 41141 10044 41153 10047
rect 41104 10016 41153 10044
rect 41104 10004 41110 10016
rect 41141 10013 41153 10016
rect 41187 10013 41199 10047
rect 41141 10007 41199 10013
rect 41693 10047 41751 10053
rect 41693 10013 41705 10047
rect 41739 10044 41751 10047
rect 42521 10047 42579 10053
rect 42521 10044 42533 10047
rect 41739 10016 42533 10044
rect 41739 10013 41751 10016
rect 41693 10007 41751 10013
rect 42521 10013 42533 10016
rect 42567 10013 42579 10047
rect 45278 10044 45284 10056
rect 45239 10016 45284 10044
rect 42521 10007 42579 10013
rect 32950 9976 32956 9988
rect 32140 9948 32956 9976
rect 30193 9939 30251 9945
rect 32950 9936 32956 9948
rect 33008 9936 33014 9988
rect 38473 9979 38531 9985
rect 38473 9945 38485 9979
rect 38519 9976 38531 9979
rect 38746 9976 38752 9988
rect 38519 9948 38752 9976
rect 38519 9945 38531 9948
rect 38473 9939 38531 9945
rect 38746 9936 38752 9948
rect 38804 9936 38810 9988
rect 41414 9936 41420 9988
rect 41472 9976 41478 9988
rect 42536 9976 42564 10007
rect 45278 10004 45284 10016
rect 45336 10004 45342 10056
rect 47136 10044 47164 10084
rect 47578 10072 47584 10084
rect 47636 10072 47642 10124
rect 47762 10112 47768 10124
rect 47723 10084 47768 10112
rect 47762 10072 47768 10084
rect 47820 10072 47826 10124
rect 47854 10072 47860 10124
rect 47912 10112 47918 10124
rect 48682 10112 48688 10124
rect 47912 10084 48688 10112
rect 47912 10072 47918 10084
rect 48682 10072 48688 10084
rect 48740 10072 48746 10124
rect 49053 10115 49111 10121
rect 49053 10081 49065 10115
rect 49099 10112 49111 10115
rect 49326 10112 49332 10124
rect 49099 10084 49332 10112
rect 49099 10081 49111 10084
rect 49053 10075 49111 10081
rect 49326 10072 49332 10084
rect 49384 10112 49390 10124
rect 49789 10115 49847 10121
rect 49789 10112 49801 10115
rect 49384 10084 49801 10112
rect 49384 10072 49390 10084
rect 49789 10081 49801 10084
rect 49835 10081 49847 10115
rect 50356 10112 50384 10152
rect 50525 10115 50583 10121
rect 50525 10112 50537 10115
rect 50356 10084 50537 10112
rect 49789 10075 49847 10081
rect 50525 10081 50537 10084
rect 50571 10081 50583 10115
rect 50525 10075 50583 10081
rect 46400 10016 47164 10044
rect 44637 9979 44695 9985
rect 41472 9948 42012 9976
rect 42536 9948 44588 9976
rect 41472 9936 41478 9948
rect 29086 9908 29092 9920
rect 28644 9880 29092 9908
rect 28445 9871 28503 9877
rect 29086 9868 29092 9880
rect 29144 9908 29150 9920
rect 29457 9911 29515 9917
rect 29457 9908 29469 9911
rect 29144 9880 29469 9908
rect 29144 9868 29150 9880
rect 29457 9877 29469 9880
rect 29503 9877 29515 9911
rect 29457 9871 29515 9877
rect 29917 9911 29975 9917
rect 29917 9877 29929 9911
rect 29963 9908 29975 9911
rect 30098 9908 30104 9920
rect 29963 9880 30104 9908
rect 29963 9877 29975 9880
rect 29917 9871 29975 9877
rect 30098 9868 30104 9880
rect 30156 9868 30162 9920
rect 30282 9868 30288 9920
rect 30340 9908 30346 9920
rect 30561 9911 30619 9917
rect 30561 9908 30573 9911
rect 30340 9880 30573 9908
rect 30340 9868 30346 9880
rect 30561 9877 30573 9880
rect 30607 9877 30619 9911
rect 30561 9871 30619 9877
rect 31021 9911 31079 9917
rect 31021 9877 31033 9911
rect 31067 9908 31079 9911
rect 31202 9908 31208 9920
rect 31067 9880 31208 9908
rect 31067 9877 31079 9880
rect 31021 9871 31079 9877
rect 31202 9868 31208 9880
rect 31260 9868 31266 9920
rect 31754 9868 31760 9920
rect 31812 9908 31818 9920
rect 33045 9911 33103 9917
rect 31812 9880 31857 9908
rect 31812 9868 31818 9880
rect 33045 9877 33057 9911
rect 33091 9908 33103 9911
rect 33870 9908 33876 9920
rect 33091 9880 33876 9908
rect 33091 9877 33103 9880
rect 33045 9871 33103 9877
rect 33870 9868 33876 9880
rect 33928 9868 33934 9920
rect 34330 9868 34336 9920
rect 34388 9908 34394 9920
rect 34517 9911 34575 9917
rect 34517 9908 34529 9911
rect 34388 9880 34529 9908
rect 34388 9868 34394 9880
rect 34517 9877 34529 9880
rect 34563 9877 34575 9911
rect 34517 9871 34575 9877
rect 35253 9911 35311 9917
rect 35253 9877 35265 9911
rect 35299 9908 35311 9911
rect 35526 9908 35532 9920
rect 35299 9880 35532 9908
rect 35299 9877 35311 9880
rect 35253 9871 35311 9877
rect 35526 9868 35532 9880
rect 35584 9868 35590 9920
rect 36170 9868 36176 9920
rect 36228 9908 36234 9920
rect 36906 9908 36912 9920
rect 36228 9880 36912 9908
rect 36228 9868 36234 9880
rect 36906 9868 36912 9880
rect 36964 9868 36970 9920
rect 37918 9908 37924 9920
rect 37879 9880 37924 9908
rect 37918 9868 37924 9880
rect 37976 9908 37982 9920
rect 39485 9911 39543 9917
rect 39485 9908 39497 9911
rect 37976 9880 39497 9908
rect 37976 9868 37982 9880
rect 39485 9877 39497 9880
rect 39531 9877 39543 9911
rect 41506 9908 41512 9920
rect 41467 9880 41512 9908
rect 39485 9871 39543 9877
rect 41506 9868 41512 9880
rect 41564 9868 41570 9920
rect 41984 9917 42012 9948
rect 41969 9911 42027 9917
rect 41969 9877 41981 9911
rect 42015 9877 42027 9911
rect 42886 9908 42892 9920
rect 42847 9880 42892 9908
rect 41969 9871 42027 9877
rect 42886 9868 42892 9880
rect 42944 9868 42950 9920
rect 43070 9868 43076 9920
rect 43128 9908 43134 9920
rect 43530 9908 43536 9920
rect 43128 9880 43536 9908
rect 43128 9868 43134 9880
rect 43530 9868 43536 9880
rect 43588 9868 43594 9920
rect 43898 9908 43904 9920
rect 43859 9880 43904 9908
rect 43898 9868 43904 9880
rect 43956 9868 43962 9920
rect 44560 9908 44588 9948
rect 44637 9945 44649 9979
rect 44683 9976 44695 9979
rect 45462 9976 45468 9988
rect 44683 9948 45468 9976
rect 44683 9945 44695 9948
rect 44637 9939 44695 9945
rect 45462 9936 45468 9948
rect 45520 9936 45526 9988
rect 46400 9908 46428 10016
rect 47210 10004 47216 10056
rect 47268 10044 47274 10056
rect 48961 10047 49019 10053
rect 48961 10044 48973 10047
rect 47268 10016 48973 10044
rect 47268 10004 47274 10016
rect 48961 10013 48973 10016
rect 49007 10013 49019 10047
rect 48961 10007 49019 10013
rect 47118 9936 47124 9988
rect 47176 9976 47182 9988
rect 51092 9976 51120 10152
rect 51534 10140 51540 10192
rect 51592 10180 51598 10192
rect 51721 10183 51779 10189
rect 51721 10180 51733 10183
rect 51592 10152 51733 10180
rect 51592 10140 51598 10152
rect 51721 10149 51733 10152
rect 51767 10149 51779 10183
rect 55398 10180 55404 10192
rect 51721 10143 51779 10149
rect 52656 10152 55404 10180
rect 51258 10112 51264 10124
rect 51219 10084 51264 10112
rect 51258 10072 51264 10084
rect 51316 10112 51322 10124
rect 52656 10112 52684 10152
rect 51316 10084 52684 10112
rect 51316 10072 51322 10084
rect 52730 10072 52736 10124
rect 52788 10112 52794 10124
rect 53009 10115 53067 10121
rect 53009 10112 53021 10115
rect 52788 10084 53021 10112
rect 52788 10072 52794 10084
rect 53009 10081 53021 10084
rect 53055 10081 53067 10115
rect 53009 10075 53067 10081
rect 53377 10115 53435 10121
rect 53377 10081 53389 10115
rect 53423 10081 53435 10115
rect 53377 10075 53435 10081
rect 53469 10115 53527 10121
rect 53469 10081 53481 10115
rect 53515 10112 53527 10115
rect 53558 10112 53564 10124
rect 53515 10084 53564 10112
rect 53515 10081 53527 10084
rect 53469 10075 53527 10081
rect 51169 10047 51227 10053
rect 51169 10013 51181 10047
rect 51215 10044 51227 10047
rect 51534 10044 51540 10056
rect 51215 10016 51540 10044
rect 51215 10013 51227 10016
rect 51169 10007 51227 10013
rect 51534 10004 51540 10016
rect 51592 10004 51598 10056
rect 51626 10004 51632 10056
rect 51684 10044 51690 10056
rect 53392 10044 53420 10075
rect 53558 10072 53564 10084
rect 53616 10112 53622 10124
rect 55048 10121 55076 10152
rect 55398 10140 55404 10152
rect 55456 10140 55462 10192
rect 56244 10180 56272 10220
rect 56321 10217 56333 10251
rect 56367 10248 56379 10251
rect 56410 10248 56416 10260
rect 56367 10220 56416 10248
rect 56367 10217 56379 10220
rect 56321 10211 56379 10217
rect 56410 10208 56416 10220
rect 56468 10208 56474 10260
rect 57238 10248 57244 10260
rect 57199 10220 57244 10248
rect 57238 10208 57244 10220
rect 57296 10208 57302 10260
rect 57330 10208 57336 10260
rect 57388 10248 57394 10260
rect 57609 10251 57667 10257
rect 57609 10248 57621 10251
rect 57388 10220 57621 10248
rect 57388 10208 57394 10220
rect 57609 10217 57621 10220
rect 57655 10217 57667 10251
rect 61838 10248 61844 10260
rect 57609 10211 57667 10217
rect 57716 10220 61844 10248
rect 57716 10180 57744 10220
rect 61838 10208 61844 10220
rect 61896 10208 61902 10260
rect 56244 10152 57744 10180
rect 55033 10115 55091 10121
rect 53616 10084 54708 10112
rect 53616 10072 53622 10084
rect 53834 10044 53840 10056
rect 51684 10016 53840 10044
rect 51684 10004 51690 10016
rect 53834 10004 53840 10016
rect 53892 10004 53898 10056
rect 52365 9979 52423 9985
rect 52365 9976 52377 9979
rect 47176 9948 49280 9976
rect 51092 9948 52377 9976
rect 47176 9936 47182 9948
rect 44560 9880 46428 9908
rect 46474 9868 46480 9920
rect 46532 9908 46538 9920
rect 47210 9908 47216 9920
rect 46532 9880 46577 9908
rect 47171 9880 47216 9908
rect 46532 9868 46538 9880
rect 47210 9868 47216 9880
rect 47268 9868 47274 9920
rect 47673 9911 47731 9917
rect 47673 9877 47685 9911
rect 47719 9908 47731 9911
rect 48406 9908 48412 9920
rect 47719 9880 48412 9908
rect 47719 9877 47731 9880
rect 47673 9871 47731 9877
rect 48406 9868 48412 9880
rect 48464 9868 48470 9920
rect 48682 9908 48688 9920
rect 48643 9880 48688 9908
rect 48682 9868 48688 9880
rect 48740 9868 48746 9920
rect 49252 9917 49280 9948
rect 52365 9945 52377 9948
rect 52411 9945 52423 9979
rect 52822 9976 52828 9988
rect 52783 9948 52828 9976
rect 52365 9939 52423 9945
rect 52822 9936 52828 9948
rect 52880 9936 52886 9988
rect 49237 9911 49295 9917
rect 49237 9877 49249 9911
rect 49283 9877 49295 9911
rect 49237 9871 49295 9877
rect 49602 9868 49608 9920
rect 49660 9908 49666 9920
rect 50157 9911 50215 9917
rect 50157 9908 50169 9911
rect 49660 9880 50169 9908
rect 49660 9868 49666 9880
rect 50157 9877 50169 9880
rect 50203 9877 50215 9911
rect 50157 9871 50215 9877
rect 50246 9868 50252 9920
rect 50304 9908 50310 9920
rect 50341 9911 50399 9917
rect 50341 9908 50353 9911
rect 50304 9880 50353 9908
rect 50304 9868 50310 9880
rect 50341 9877 50353 9880
rect 50387 9877 50399 9911
rect 50341 9871 50399 9877
rect 51810 9868 51816 9920
rect 51868 9908 51874 9920
rect 51997 9911 52055 9917
rect 51997 9908 52009 9911
rect 51868 9880 52009 9908
rect 51868 9868 51874 9880
rect 51997 9877 52009 9880
rect 52043 9877 52055 9911
rect 54680 9908 54708 10084
rect 55033 10081 55045 10115
rect 55079 10081 55091 10115
rect 56502 10112 56508 10124
rect 56463 10084 56508 10112
rect 55033 10075 55091 10081
rect 56502 10072 56508 10084
rect 56560 10072 56566 10124
rect 58434 10112 58440 10124
rect 58395 10084 58440 10112
rect 58434 10072 58440 10084
rect 58492 10072 58498 10124
rect 58805 10115 58863 10121
rect 58805 10081 58817 10115
rect 58851 10112 58863 10115
rect 60185 10115 60243 10121
rect 58851 10084 59768 10112
rect 58851 10081 58863 10084
rect 58805 10075 58863 10081
rect 54754 10004 54760 10056
rect 54812 10044 54818 10056
rect 54941 10047 54999 10053
rect 54941 10044 54953 10047
rect 54812 10016 54953 10044
rect 54812 10004 54818 10016
rect 54941 10013 54953 10016
rect 54987 10013 54999 10047
rect 56410 10044 56416 10056
rect 56371 10016 56416 10044
rect 54941 10007 54999 10013
rect 56410 10004 56416 10016
rect 56468 10004 56474 10056
rect 57790 10004 57796 10056
rect 57848 10044 57854 10056
rect 58345 10047 58403 10053
rect 58345 10044 58357 10047
rect 57848 10016 58357 10044
rect 57848 10004 57854 10016
rect 58345 10013 58357 10016
rect 58391 10013 58403 10047
rect 58345 10007 58403 10013
rect 58897 10047 58955 10053
rect 58897 10013 58909 10047
rect 58943 10044 58955 10047
rect 58943 10016 59400 10044
rect 58943 10013 58955 10016
rect 58897 10007 58955 10013
rect 59078 9976 59084 9988
rect 55048 9948 59084 9976
rect 55048 9908 55076 9948
rect 59078 9936 59084 9948
rect 59136 9936 59142 9988
rect 55214 9908 55220 9920
rect 54680 9880 55076 9908
rect 55175 9880 55220 9908
rect 51997 9871 52055 9877
rect 55214 9868 55220 9880
rect 55272 9868 55278 9920
rect 56594 9868 56600 9920
rect 56652 9908 56658 9920
rect 56689 9911 56747 9917
rect 56689 9908 56701 9911
rect 56652 9880 56701 9908
rect 56652 9868 56658 9880
rect 56689 9877 56701 9880
rect 56735 9877 56747 9911
rect 56689 9871 56747 9877
rect 57885 9911 57943 9917
rect 57885 9877 57897 9911
rect 57931 9908 57943 9911
rect 58158 9908 58164 9920
rect 57931 9880 58164 9908
rect 57931 9877 57943 9880
rect 57885 9871 57943 9877
rect 58158 9868 58164 9880
rect 58216 9868 58222 9920
rect 59372 9917 59400 10016
rect 59357 9911 59415 9917
rect 59357 9877 59369 9911
rect 59403 9908 59415 9911
rect 59446 9908 59452 9920
rect 59403 9880 59452 9908
rect 59403 9877 59415 9880
rect 59357 9871 59415 9877
rect 59446 9868 59452 9880
rect 59504 9868 59510 9920
rect 59740 9917 59768 10084
rect 60185 10081 60197 10115
rect 60231 10112 60243 10115
rect 61286 10112 61292 10124
rect 60231 10084 61292 10112
rect 60231 10081 60243 10084
rect 60185 10075 60243 10081
rect 61286 10072 61292 10084
rect 61344 10072 61350 10124
rect 60458 10044 60464 10056
rect 60419 10016 60464 10044
rect 60458 10004 60464 10016
rect 60516 10004 60522 10056
rect 59725 9911 59783 9917
rect 59725 9877 59737 9911
rect 59771 9908 59783 9911
rect 59814 9908 59820 9920
rect 59771 9880 59820 9908
rect 59771 9877 59783 9880
rect 59725 9871 59783 9877
rect 59814 9868 59820 9880
rect 59872 9868 59878 9920
rect 61749 9911 61807 9917
rect 61749 9877 61761 9911
rect 61795 9908 61807 9911
rect 61838 9908 61844 9920
rect 61795 9880 61844 9908
rect 61795 9877 61807 9880
rect 61749 9871 61807 9877
rect 61838 9868 61844 9880
rect 61896 9868 61902 9920
rect 1104 9818 63480 9840
rect 1104 9766 11378 9818
rect 11430 9766 11442 9818
rect 11494 9766 11506 9818
rect 11558 9766 11570 9818
rect 11622 9766 32170 9818
rect 32222 9766 32234 9818
rect 32286 9766 32298 9818
rect 32350 9766 32362 9818
rect 32414 9766 52962 9818
rect 53014 9766 53026 9818
rect 53078 9766 53090 9818
rect 53142 9766 53154 9818
rect 53206 9766 63480 9818
rect 1104 9744 63480 9766
rect 4798 9664 4804 9716
rect 4856 9704 4862 9716
rect 5905 9707 5963 9713
rect 5905 9704 5917 9707
rect 4856 9676 5917 9704
rect 4856 9664 4862 9676
rect 5905 9673 5917 9676
rect 5951 9704 5963 9707
rect 6273 9707 6331 9713
rect 6273 9704 6285 9707
rect 5951 9676 6285 9704
rect 5951 9673 5963 9676
rect 5905 9667 5963 9673
rect 6273 9673 6285 9676
rect 6319 9704 6331 9707
rect 6362 9704 6368 9716
rect 6319 9676 6368 9704
rect 6319 9673 6331 9676
rect 6273 9667 6331 9673
rect 6362 9664 6368 9676
rect 6420 9704 6426 9716
rect 9950 9704 9956 9716
rect 6420 9676 9956 9704
rect 6420 9664 6426 9676
rect 2958 9636 2964 9648
rect 2919 9608 2964 9636
rect 2958 9596 2964 9608
rect 3016 9596 3022 9648
rect 5261 9639 5319 9645
rect 5261 9605 5273 9639
rect 5307 9636 5319 9639
rect 5350 9636 5356 9648
rect 5307 9608 5356 9636
rect 5307 9605 5319 9608
rect 5261 9599 5319 9605
rect 5350 9596 5356 9608
rect 5408 9596 5414 9648
rect 3789 9571 3847 9577
rect 3789 9537 3801 9571
rect 3835 9568 3847 9571
rect 3881 9571 3939 9577
rect 3881 9568 3893 9571
rect 3835 9540 3893 9568
rect 3835 9537 3847 9540
rect 3789 9531 3847 9537
rect 3881 9537 3893 9540
rect 3927 9568 3939 9571
rect 4246 9568 4252 9580
rect 3927 9540 4252 9568
rect 3927 9537 3939 9540
rect 3881 9531 3939 9537
rect 4246 9528 4252 9540
rect 4304 9528 4310 9580
rect 6840 9577 6868 9676
rect 9950 9664 9956 9676
rect 10008 9664 10014 9716
rect 11790 9704 11796 9716
rect 11751 9676 11796 9704
rect 11790 9664 11796 9676
rect 11848 9664 11854 9716
rect 12250 9704 12256 9716
rect 12211 9676 12256 9704
rect 12250 9664 12256 9676
rect 12308 9664 12314 9716
rect 14185 9707 14243 9713
rect 14185 9673 14197 9707
rect 14231 9704 14243 9707
rect 14274 9704 14280 9716
rect 14231 9676 14280 9704
rect 14231 9673 14243 9676
rect 14185 9667 14243 9673
rect 14274 9664 14280 9676
rect 14332 9664 14338 9716
rect 15013 9707 15071 9713
rect 15013 9673 15025 9707
rect 15059 9704 15071 9707
rect 16022 9704 16028 9716
rect 15059 9676 15240 9704
rect 15983 9676 16028 9704
rect 15059 9673 15071 9676
rect 15013 9667 15071 9673
rect 9217 9639 9275 9645
rect 9217 9605 9229 9639
rect 9263 9636 9275 9639
rect 9674 9636 9680 9648
rect 9263 9608 9680 9636
rect 9263 9605 9275 9608
rect 9217 9599 9275 9605
rect 9674 9596 9680 9608
rect 9732 9596 9738 9648
rect 12713 9639 12771 9645
rect 12713 9605 12725 9639
rect 12759 9636 12771 9639
rect 12802 9636 12808 9648
rect 12759 9608 12808 9636
rect 12759 9605 12771 9608
rect 12713 9599 12771 9605
rect 12802 9596 12808 9608
rect 12860 9596 12866 9648
rect 13538 9596 13544 9648
rect 13596 9636 13602 9648
rect 15105 9639 15163 9645
rect 15105 9636 15117 9639
rect 13596 9608 15117 9636
rect 13596 9596 13602 9608
rect 15105 9605 15117 9608
rect 15151 9605 15163 9639
rect 15212 9636 15240 9676
rect 16022 9664 16028 9676
rect 16080 9664 16086 9716
rect 17954 9664 17960 9716
rect 18012 9704 18018 9716
rect 18012 9676 18552 9704
rect 18012 9664 18018 9676
rect 15381 9639 15439 9645
rect 15381 9636 15393 9639
rect 15212 9608 15393 9636
rect 15105 9599 15163 9605
rect 15381 9605 15393 9608
rect 15427 9605 15439 9639
rect 15381 9599 15439 9605
rect 16485 9639 16543 9645
rect 16485 9605 16497 9639
rect 16531 9636 16543 9639
rect 18322 9636 18328 9648
rect 16531 9608 18328 9636
rect 16531 9605 16543 9608
rect 16485 9599 16543 9605
rect 6825 9571 6883 9577
rect 6825 9537 6837 9571
rect 6871 9537 6883 9571
rect 6825 9531 6883 9537
rect 8481 9571 8539 9577
rect 8481 9537 8493 9571
rect 8527 9568 8539 9571
rect 10502 9568 10508 9580
rect 8527 9540 10508 9568
rect 8527 9537 8539 9540
rect 8481 9531 8539 9537
rect 10502 9528 10508 9540
rect 10560 9528 10566 9580
rect 11517 9571 11575 9577
rect 11517 9537 11529 9571
rect 11563 9568 11575 9571
rect 12158 9568 12164 9580
rect 11563 9540 12164 9568
rect 11563 9537 11575 9540
rect 11517 9531 11575 9537
rect 12158 9528 12164 9540
rect 12216 9528 12222 9580
rect 12618 9528 12624 9580
rect 12676 9568 12682 9580
rect 13725 9571 13783 9577
rect 13725 9568 13737 9571
rect 12676 9540 13737 9568
rect 12676 9528 12682 9540
rect 2777 9503 2835 9509
rect 2777 9469 2789 9503
rect 2823 9500 2835 9503
rect 4154 9500 4160 9512
rect 2823 9472 3096 9500
rect 4115 9472 4160 9500
rect 2823 9469 2835 9472
rect 2777 9463 2835 9469
rect 3068 9376 3096 9472
rect 4154 9460 4160 9472
rect 4212 9460 4218 9512
rect 7098 9500 7104 9512
rect 6932 9472 7104 9500
rect 6641 9435 6699 9441
rect 6641 9401 6653 9435
rect 6687 9432 6699 9435
rect 6932 9432 6960 9472
rect 7098 9460 7104 9472
rect 7156 9460 7162 9512
rect 9306 9500 9312 9512
rect 9267 9472 9312 9500
rect 9306 9460 9312 9472
rect 9364 9460 9370 9512
rect 9401 9503 9459 9509
rect 9401 9469 9413 9503
rect 9447 9500 9459 9503
rect 9447 9472 10272 9500
rect 9447 9469 9459 9472
rect 9401 9463 9459 9469
rect 9858 9432 9864 9444
rect 6687 9404 6960 9432
rect 9819 9404 9864 9432
rect 6687 9401 6699 9404
rect 6641 9395 6699 9401
rect 9858 9392 9864 9404
rect 9916 9392 9922 9444
rect 10244 9441 10272 9472
rect 10686 9460 10692 9512
rect 10744 9500 10750 9512
rect 10965 9503 11023 9509
rect 10965 9500 10977 9503
rect 10744 9472 10977 9500
rect 10744 9460 10750 9472
rect 10965 9469 10977 9472
rect 11011 9469 11023 9503
rect 10965 9463 11023 9469
rect 11057 9503 11115 9509
rect 11057 9469 11069 9503
rect 11103 9469 11115 9503
rect 12894 9500 12900 9512
rect 12855 9472 12900 9500
rect 11057 9463 11115 9469
rect 10229 9435 10287 9441
rect 10229 9401 10241 9435
rect 10275 9432 10287 9435
rect 10870 9432 10876 9444
rect 10275 9404 10876 9432
rect 10275 9401 10287 9404
rect 10229 9395 10287 9401
rect 10870 9392 10876 9404
rect 10928 9432 10934 9444
rect 11072 9432 11100 9463
rect 12894 9460 12900 9472
rect 12952 9460 12958 9512
rect 13096 9509 13124 9540
rect 13725 9537 13737 9540
rect 13771 9537 13783 9571
rect 15120 9568 15148 9599
rect 18322 9596 18328 9608
rect 18380 9596 18386 9648
rect 18524 9636 18552 9676
rect 18782 9664 18788 9716
rect 18840 9704 18846 9716
rect 18969 9707 19027 9713
rect 18969 9704 18981 9707
rect 18840 9676 18981 9704
rect 18840 9664 18846 9676
rect 18969 9673 18981 9676
rect 19015 9673 19027 9707
rect 18969 9667 19027 9673
rect 20806 9664 20812 9716
rect 20864 9704 20870 9716
rect 22557 9707 22615 9713
rect 22557 9704 22569 9707
rect 20864 9676 22569 9704
rect 20864 9664 20870 9676
rect 22557 9673 22569 9676
rect 22603 9673 22615 9707
rect 23198 9704 23204 9716
rect 23159 9676 23204 9704
rect 22557 9667 22615 9673
rect 23198 9664 23204 9676
rect 23256 9664 23262 9716
rect 27430 9704 27436 9716
rect 27391 9676 27436 9704
rect 27430 9664 27436 9676
rect 27488 9704 27494 9716
rect 27614 9704 27620 9716
rect 27488 9676 27620 9704
rect 27488 9664 27494 9676
rect 27614 9664 27620 9676
rect 27672 9664 27678 9716
rect 28902 9704 28908 9716
rect 27724 9676 28908 9704
rect 19150 9636 19156 9648
rect 18524 9608 19156 9636
rect 19150 9596 19156 9608
rect 19208 9636 19214 9648
rect 19337 9639 19395 9645
rect 19337 9636 19349 9639
rect 19208 9608 19349 9636
rect 19208 9596 19214 9608
rect 19337 9605 19349 9608
rect 19383 9605 19395 9639
rect 19794 9636 19800 9648
rect 19755 9608 19800 9636
rect 19337 9599 19395 9605
rect 19794 9596 19800 9608
rect 19852 9596 19858 9648
rect 22005 9639 22063 9645
rect 22005 9636 22017 9639
rect 19904 9608 22017 9636
rect 16390 9568 16396 9580
rect 15120 9540 16396 9568
rect 13725 9531 13783 9537
rect 16390 9528 16396 9540
rect 16448 9528 16454 9580
rect 16577 9571 16635 9577
rect 16577 9537 16589 9571
rect 16623 9568 16635 9571
rect 16623 9540 16896 9568
rect 16623 9537 16635 9540
rect 16577 9531 16635 9537
rect 13081 9503 13139 9509
rect 13081 9469 13093 9503
rect 13127 9469 13139 9503
rect 13081 9463 13139 9469
rect 13265 9503 13323 9509
rect 13265 9469 13277 9503
rect 13311 9500 13323 9503
rect 14274 9500 14280 9512
rect 13311 9472 14280 9500
rect 13311 9469 13323 9472
rect 13265 9463 13323 9469
rect 14274 9460 14280 9472
rect 14332 9460 14338 9512
rect 14645 9503 14703 9509
rect 14645 9469 14657 9503
rect 14691 9500 14703 9503
rect 14734 9500 14740 9512
rect 14691 9472 14740 9500
rect 14691 9469 14703 9472
rect 14645 9463 14703 9469
rect 14734 9460 14740 9472
rect 14792 9460 14798 9512
rect 15194 9460 15200 9512
rect 15252 9500 15258 9512
rect 15289 9503 15347 9509
rect 15289 9500 15301 9503
rect 15252 9472 15301 9500
rect 15252 9460 15258 9472
rect 15289 9469 15301 9472
rect 15335 9469 15347 9503
rect 15289 9463 15347 9469
rect 15381 9503 15439 9509
rect 15381 9469 15393 9503
rect 15427 9500 15439 9503
rect 15473 9503 15531 9509
rect 15473 9500 15485 9503
rect 15427 9472 15485 9500
rect 15427 9469 15439 9472
rect 15381 9463 15439 9469
rect 15473 9469 15485 9472
rect 15519 9500 15531 9503
rect 16022 9500 16028 9512
rect 15519 9472 16028 9500
rect 15519 9469 15531 9472
rect 15473 9463 15531 9469
rect 16022 9460 16028 9472
rect 16080 9460 16086 9512
rect 16209 9503 16267 9509
rect 16209 9469 16221 9503
rect 16255 9500 16267 9503
rect 16666 9500 16672 9512
rect 16255 9472 16672 9500
rect 16255 9469 16267 9472
rect 16209 9463 16267 9469
rect 16666 9460 16672 9472
rect 16724 9460 16730 9512
rect 16868 9500 16896 9540
rect 16942 9528 16948 9580
rect 17000 9568 17006 9580
rect 17129 9571 17187 9577
rect 17129 9568 17141 9571
rect 17000 9540 17141 9568
rect 17000 9528 17006 9540
rect 17129 9537 17141 9540
rect 17175 9537 17187 9571
rect 18506 9568 18512 9580
rect 17129 9531 17187 9537
rect 17420 9540 18512 9568
rect 17420 9509 17448 9540
rect 18506 9528 18512 9540
rect 18564 9528 18570 9580
rect 18693 9571 18751 9577
rect 18693 9537 18705 9571
rect 18739 9568 18751 9571
rect 19058 9568 19064 9580
rect 18739 9540 19064 9568
rect 18739 9537 18751 9540
rect 18693 9531 18751 9537
rect 19058 9528 19064 9540
rect 19116 9528 19122 9580
rect 19242 9528 19248 9580
rect 19300 9568 19306 9580
rect 19904 9568 19932 9608
rect 22005 9605 22017 9608
rect 22051 9605 22063 9639
rect 22005 9599 22063 9605
rect 22741 9639 22799 9645
rect 22741 9605 22753 9639
rect 22787 9605 22799 9639
rect 22741 9599 22799 9605
rect 20714 9568 20720 9580
rect 19300 9540 19932 9568
rect 19996 9540 20720 9568
rect 19300 9528 19306 9540
rect 19996 9512 20024 9540
rect 20714 9528 20720 9540
rect 20772 9528 20778 9580
rect 21361 9571 21419 9577
rect 21361 9537 21373 9571
rect 21407 9568 21419 9571
rect 21910 9568 21916 9580
rect 21407 9540 21588 9568
rect 21871 9540 21916 9568
rect 21407 9537 21419 9540
rect 21361 9531 21419 9537
rect 17405 9503 17463 9509
rect 17405 9500 17417 9503
rect 16868 9472 17417 9500
rect 17405 9469 17417 9472
rect 17451 9469 17463 9503
rect 17405 9463 17463 9469
rect 18046 9460 18052 9512
rect 18104 9500 18110 9512
rect 18141 9503 18199 9509
rect 18141 9500 18153 9503
rect 18104 9472 18153 9500
rect 18104 9460 18110 9472
rect 18141 9469 18153 9472
rect 18187 9469 18199 9503
rect 18141 9463 18199 9469
rect 18230 9460 18236 9512
rect 18288 9500 18294 9512
rect 19978 9500 19984 9512
rect 18288 9472 18333 9500
rect 19939 9472 19984 9500
rect 18288 9460 18294 9472
rect 19978 9460 19984 9472
rect 20036 9460 20042 9512
rect 20165 9503 20223 9509
rect 20165 9469 20177 9503
rect 20211 9469 20223 9503
rect 20165 9463 20223 9469
rect 20349 9503 20407 9509
rect 20349 9469 20361 9503
rect 20395 9500 20407 9503
rect 21082 9500 21088 9512
rect 20395 9472 21088 9500
rect 20395 9469 20407 9472
rect 20349 9463 20407 9469
rect 17218 9432 17224 9444
rect 10928 9404 17224 9432
rect 10928 9392 10934 9404
rect 17218 9392 17224 9404
rect 17276 9392 17282 9444
rect 18690 9392 18696 9444
rect 18748 9432 18754 9444
rect 19242 9432 19248 9444
rect 18748 9404 19248 9432
rect 18748 9392 18754 9404
rect 19242 9392 19248 9404
rect 19300 9432 19306 9444
rect 20180 9432 20208 9463
rect 21082 9460 21088 9472
rect 21140 9460 21146 9512
rect 21453 9503 21511 9509
rect 21453 9500 21465 9503
rect 21284 9472 21465 9500
rect 20254 9432 20260 9444
rect 19300 9404 20260 9432
rect 19300 9392 19306 9404
rect 20254 9392 20260 9404
rect 20312 9432 20318 9444
rect 20806 9432 20812 9444
rect 20312 9404 20812 9432
rect 20312 9392 20318 9404
rect 20806 9392 20812 9404
rect 20864 9392 20870 9444
rect 21284 9376 21312 9472
rect 21453 9469 21465 9472
rect 21499 9469 21511 9503
rect 21453 9463 21511 9469
rect 3050 9324 3056 9376
rect 3108 9364 3114 9376
rect 3329 9367 3387 9373
rect 3329 9364 3341 9367
rect 3108 9336 3341 9364
rect 3108 9324 3114 9336
rect 3329 9333 3341 9336
rect 3375 9333 3387 9367
rect 3329 9327 3387 9333
rect 8849 9367 8907 9373
rect 8849 9333 8861 9367
rect 8895 9364 8907 9367
rect 8938 9364 8944 9376
rect 8895 9336 8944 9364
rect 8895 9333 8907 9336
rect 8849 9327 8907 9333
rect 8938 9324 8944 9336
rect 8996 9324 9002 9376
rect 10686 9324 10692 9376
rect 10744 9364 10750 9376
rect 10781 9367 10839 9373
rect 10781 9364 10793 9367
rect 10744 9336 10793 9364
rect 10744 9324 10750 9336
rect 10781 9333 10793 9336
rect 10827 9333 10839 9367
rect 10781 9327 10839 9333
rect 11054 9324 11060 9376
rect 11112 9364 11118 9376
rect 15657 9367 15715 9373
rect 15657 9364 15669 9367
rect 11112 9336 15669 9364
rect 11112 9324 11118 9336
rect 15657 9333 15669 9336
rect 15703 9364 15715 9367
rect 16209 9367 16267 9373
rect 16209 9364 16221 9367
rect 15703 9336 16221 9364
rect 15703 9333 15715 9336
rect 15657 9327 15715 9333
rect 16209 9333 16221 9336
rect 16255 9333 16267 9367
rect 16209 9327 16267 9333
rect 17586 9324 17592 9376
rect 17644 9364 17650 9376
rect 17773 9367 17831 9373
rect 17773 9364 17785 9367
rect 17644 9336 17785 9364
rect 17644 9324 17650 9336
rect 17773 9333 17785 9336
rect 17819 9333 17831 9367
rect 17773 9327 17831 9333
rect 18138 9324 18144 9376
rect 18196 9364 18202 9376
rect 21082 9364 21088 9376
rect 18196 9336 21088 9364
rect 18196 9324 18202 9336
rect 21082 9324 21088 9336
rect 21140 9324 21146 9376
rect 21266 9364 21272 9376
rect 21227 9336 21272 9364
rect 21266 9324 21272 9336
rect 21324 9324 21330 9376
rect 21560 9364 21588 9540
rect 21910 9528 21916 9540
rect 21968 9528 21974 9580
rect 22097 9571 22155 9577
rect 22097 9537 22109 9571
rect 22143 9568 22155 9571
rect 22756 9568 22784 9599
rect 23382 9596 23388 9648
rect 23440 9636 23446 9648
rect 23845 9639 23903 9645
rect 23845 9636 23857 9639
rect 23440 9608 23857 9636
rect 23440 9596 23446 9608
rect 23845 9605 23857 9608
rect 23891 9605 23903 9639
rect 23845 9599 23903 9605
rect 24581 9639 24639 9645
rect 24581 9605 24593 9639
rect 24627 9636 24639 9639
rect 25038 9636 25044 9648
rect 24627 9608 25044 9636
rect 24627 9605 24639 9608
rect 24581 9599 24639 9605
rect 22143 9540 22784 9568
rect 22143 9537 22155 9540
rect 22097 9531 22155 9537
rect 22925 9503 22983 9509
rect 22925 9469 22937 9503
rect 22971 9500 22983 9503
rect 23106 9500 23112 9512
rect 22971 9472 23112 9500
rect 22971 9469 22983 9472
rect 22925 9463 22983 9469
rect 23106 9460 23112 9472
rect 23164 9460 23170 9512
rect 24029 9503 24087 9509
rect 24029 9469 24041 9503
rect 24075 9500 24087 9503
rect 24596 9500 24624 9599
rect 25038 9596 25044 9608
rect 25096 9596 25102 9648
rect 26786 9596 26792 9648
rect 26844 9636 26850 9648
rect 26973 9639 27031 9645
rect 26973 9636 26985 9639
rect 26844 9608 26985 9636
rect 26844 9596 26850 9608
rect 26973 9605 26985 9608
rect 27019 9636 27031 9639
rect 27246 9636 27252 9648
rect 27019 9608 27252 9636
rect 27019 9605 27031 9608
rect 26973 9599 27031 9605
rect 27246 9596 27252 9608
rect 27304 9596 27310 9648
rect 27724 9636 27752 9676
rect 28902 9664 28908 9676
rect 28960 9664 28966 9716
rect 35894 9664 35900 9716
rect 35952 9704 35958 9716
rect 36357 9707 36415 9713
rect 36357 9704 36369 9707
rect 35952 9676 36369 9704
rect 35952 9664 35958 9676
rect 36357 9673 36369 9676
rect 36403 9704 36415 9707
rect 36538 9704 36544 9716
rect 36403 9676 36544 9704
rect 36403 9673 36415 9676
rect 36357 9667 36415 9673
rect 36538 9664 36544 9676
rect 36596 9704 36602 9716
rect 37090 9704 37096 9716
rect 36596 9676 37096 9704
rect 36596 9664 36602 9676
rect 37090 9664 37096 9676
rect 37148 9664 37154 9716
rect 38304 9676 38608 9704
rect 27540 9608 27752 9636
rect 30101 9639 30159 9645
rect 26142 9568 26148 9580
rect 24075 9472 24624 9500
rect 24780 9540 26148 9568
rect 24075 9469 24087 9472
rect 24029 9463 24087 9469
rect 24121 9435 24179 9441
rect 24121 9401 24133 9435
rect 24167 9432 24179 9435
rect 24780 9432 24808 9540
rect 26142 9528 26148 9540
rect 26200 9528 26206 9580
rect 27062 9528 27068 9580
rect 27120 9568 27126 9580
rect 27540 9577 27568 9608
rect 30101 9605 30113 9639
rect 30147 9636 30159 9639
rect 30282 9636 30288 9648
rect 30147 9608 30288 9636
rect 30147 9605 30159 9608
rect 30101 9599 30159 9605
rect 30282 9596 30288 9608
rect 30340 9596 30346 9648
rect 31573 9639 31631 9645
rect 31573 9605 31585 9639
rect 31619 9636 31631 9639
rect 31938 9636 31944 9648
rect 31619 9608 31944 9636
rect 31619 9605 31631 9608
rect 31573 9599 31631 9605
rect 31938 9596 31944 9608
rect 31996 9636 32002 9648
rect 34330 9636 34336 9648
rect 31996 9608 34336 9636
rect 31996 9596 32002 9608
rect 34330 9596 34336 9608
rect 34388 9596 34394 9648
rect 36722 9636 36728 9648
rect 36683 9608 36728 9636
rect 36722 9596 36728 9608
rect 36780 9596 36786 9648
rect 37108 9636 37136 9664
rect 37737 9639 37795 9645
rect 37737 9636 37749 9639
rect 37108 9608 37749 9636
rect 37737 9605 37749 9608
rect 37783 9605 37795 9639
rect 37737 9599 37795 9605
rect 37826 9596 37832 9648
rect 37884 9636 37890 9648
rect 38304 9636 38332 9676
rect 38470 9636 38476 9648
rect 37884 9608 38332 9636
rect 38431 9608 38476 9636
rect 37884 9596 37890 9608
rect 38470 9596 38476 9608
rect 38528 9596 38534 9648
rect 38580 9636 38608 9676
rect 39022 9664 39028 9716
rect 39080 9704 39086 9716
rect 39577 9707 39635 9713
rect 39577 9704 39589 9707
rect 39080 9676 39589 9704
rect 39080 9664 39086 9676
rect 39577 9673 39589 9676
rect 39623 9673 39635 9707
rect 39577 9667 39635 9673
rect 41598 9664 41604 9716
rect 41656 9704 41662 9716
rect 41656 9676 49556 9704
rect 41656 9664 41662 9676
rect 38838 9636 38844 9648
rect 38580 9608 38844 9636
rect 38838 9596 38844 9608
rect 38896 9596 38902 9648
rect 38930 9596 38936 9648
rect 38988 9636 38994 9648
rect 39209 9639 39267 9645
rect 39209 9636 39221 9639
rect 38988 9608 39221 9636
rect 38988 9596 38994 9608
rect 39209 9605 39221 9608
rect 39255 9605 39267 9639
rect 39209 9599 39267 9605
rect 41049 9639 41107 9645
rect 41049 9605 41061 9639
rect 41095 9605 41107 9639
rect 41049 9599 41107 9605
rect 27525 9571 27583 9577
rect 27525 9568 27537 9571
rect 27120 9540 27537 9568
rect 27120 9528 27126 9540
rect 27525 9537 27537 9540
rect 27571 9537 27583 9571
rect 27525 9531 27583 9537
rect 27982 9528 27988 9580
rect 28040 9568 28046 9580
rect 28077 9571 28135 9577
rect 28077 9568 28089 9571
rect 28040 9540 28089 9568
rect 28040 9528 28046 9540
rect 28077 9537 28089 9540
rect 28123 9537 28135 9571
rect 33502 9568 33508 9580
rect 33463 9540 33508 9568
rect 28077 9531 28135 9537
rect 33502 9528 33508 9540
rect 33560 9528 33566 9580
rect 41064 9568 41092 9599
rect 41414 9596 41420 9648
rect 41472 9636 41478 9648
rect 42337 9639 42395 9645
rect 42337 9636 42349 9639
rect 41472 9608 42349 9636
rect 41472 9596 41478 9608
rect 42337 9605 42349 9608
rect 42383 9636 42395 9639
rect 42429 9639 42487 9645
rect 42429 9636 42441 9639
rect 42383 9608 42441 9636
rect 42383 9605 42395 9608
rect 42337 9599 42395 9605
rect 42429 9605 42441 9608
rect 42475 9605 42487 9639
rect 44174 9636 44180 9648
rect 44135 9608 44180 9636
rect 42429 9599 42487 9605
rect 44174 9596 44180 9608
rect 44232 9596 44238 9648
rect 45278 9636 45284 9648
rect 45239 9608 45284 9636
rect 45278 9596 45284 9608
rect 45336 9596 45342 9648
rect 45554 9636 45560 9648
rect 45515 9608 45560 9636
rect 45554 9596 45560 9608
rect 45612 9596 45618 9648
rect 46658 9636 46664 9648
rect 46619 9608 46664 9636
rect 46658 9596 46664 9608
rect 46716 9596 46722 9648
rect 47026 9636 47032 9648
rect 46987 9608 47032 9636
rect 47026 9596 47032 9608
rect 47084 9596 47090 9648
rect 47489 9639 47547 9645
rect 47489 9605 47501 9639
rect 47535 9636 47547 9639
rect 47854 9636 47860 9648
rect 47535 9608 47860 9636
rect 47535 9605 47547 9608
rect 47489 9599 47547 9605
rect 42886 9568 42892 9580
rect 33612 9540 36308 9568
rect 24946 9460 24952 9512
rect 25004 9500 25010 9512
rect 25041 9503 25099 9509
rect 25041 9500 25053 9503
rect 25004 9472 25053 9500
rect 25004 9460 25010 9472
rect 25041 9469 25053 9472
rect 25087 9469 25099 9503
rect 25317 9503 25375 9509
rect 25317 9500 25329 9503
rect 25041 9463 25099 9469
rect 25148 9472 25329 9500
rect 25148 9432 25176 9472
rect 25317 9469 25329 9472
rect 25363 9469 25375 9503
rect 27614 9500 27620 9512
rect 27575 9472 27620 9500
rect 25317 9463 25375 9469
rect 27614 9460 27620 9472
rect 27672 9500 27678 9512
rect 28353 9503 28411 9509
rect 28353 9500 28365 9503
rect 27672 9472 28365 9500
rect 27672 9460 27678 9472
rect 28353 9469 28365 9472
rect 28399 9500 28411 9503
rect 28442 9500 28448 9512
rect 28399 9472 28448 9500
rect 28399 9469 28411 9472
rect 28353 9463 28411 9469
rect 28442 9460 28448 9472
rect 28500 9500 28506 9512
rect 28718 9500 28724 9512
rect 28500 9472 28724 9500
rect 28500 9460 28506 9472
rect 28718 9460 28724 9472
rect 28776 9460 28782 9512
rect 29917 9503 29975 9509
rect 29917 9469 29929 9503
rect 29963 9500 29975 9503
rect 29963 9472 29997 9500
rect 29963 9469 29975 9472
rect 29917 9463 29975 9469
rect 29086 9432 29092 9444
rect 24167 9404 24808 9432
rect 24872 9404 25176 9432
rect 26436 9404 29092 9432
rect 24167 9401 24179 9404
rect 24121 9395 24179 9401
rect 24872 9376 24900 9404
rect 22281 9367 22339 9373
rect 22281 9364 22293 9367
rect 21560 9336 22293 9364
rect 22281 9333 22293 9336
rect 22327 9364 22339 9367
rect 23014 9364 23020 9376
rect 22327 9336 23020 9364
rect 22327 9333 22339 9336
rect 22281 9327 22339 9333
rect 23014 9324 23020 9336
rect 23072 9324 23078 9376
rect 24854 9364 24860 9376
rect 24815 9336 24860 9364
rect 24854 9324 24860 9336
rect 24912 9324 24918 9376
rect 25314 9324 25320 9376
rect 25372 9364 25378 9376
rect 26436 9373 26464 9404
rect 29086 9392 29092 9404
rect 29144 9392 29150 9444
rect 29825 9435 29883 9441
rect 29825 9401 29837 9435
rect 29871 9432 29883 9435
rect 29932 9432 29960 9463
rect 30282 9460 30288 9512
rect 30340 9500 30346 9512
rect 30561 9503 30619 9509
rect 30561 9500 30573 9503
rect 30340 9472 30573 9500
rect 30340 9460 30346 9472
rect 30561 9469 30573 9472
rect 30607 9500 30619 9503
rect 31205 9503 31263 9509
rect 31205 9500 31217 9503
rect 30607 9472 31217 9500
rect 30607 9469 30619 9472
rect 30561 9463 30619 9469
rect 31205 9469 31217 9472
rect 31251 9500 31263 9503
rect 31251 9472 32168 9500
rect 31251 9469 31263 9472
rect 31205 9463 31263 9469
rect 30650 9432 30656 9444
rect 29871 9404 30656 9432
rect 29871 9401 29883 9404
rect 29825 9395 29883 9401
rect 30650 9392 30656 9404
rect 30708 9392 30714 9444
rect 30834 9392 30840 9444
rect 30892 9432 30898 9444
rect 31665 9435 31723 9441
rect 31665 9432 31677 9435
rect 30892 9404 31677 9432
rect 30892 9392 30898 9404
rect 31665 9401 31677 9404
rect 31711 9432 31723 9435
rect 31754 9432 31760 9444
rect 31711 9404 31760 9432
rect 31711 9401 31723 9404
rect 31665 9395 31723 9401
rect 31754 9392 31760 9404
rect 31812 9392 31818 9444
rect 32140 9432 32168 9472
rect 33318 9460 33324 9512
rect 33376 9500 33382 9512
rect 33413 9503 33471 9509
rect 33413 9500 33425 9503
rect 33376 9472 33425 9500
rect 33376 9460 33382 9472
rect 33413 9469 33425 9472
rect 33459 9500 33471 9503
rect 33612 9500 33640 9540
rect 33962 9500 33968 9512
rect 33459 9472 33640 9500
rect 33923 9472 33968 9500
rect 33459 9469 33471 9472
rect 33413 9463 33471 9469
rect 33962 9460 33968 9472
rect 34020 9460 34026 9512
rect 34146 9500 34152 9512
rect 34107 9472 34152 9500
rect 34146 9460 34152 9472
rect 34204 9460 34210 9512
rect 34330 9500 34336 9512
rect 34291 9472 34336 9500
rect 34330 9460 34336 9472
rect 34388 9460 34394 9512
rect 34977 9503 35035 9509
rect 34977 9469 34989 9503
rect 35023 9500 35035 9503
rect 35069 9503 35127 9509
rect 35069 9500 35081 9503
rect 35023 9472 35081 9500
rect 35023 9469 35035 9472
rect 34977 9463 35035 9469
rect 35069 9469 35081 9472
rect 35115 9469 35127 9503
rect 35069 9463 35127 9469
rect 35161 9503 35219 9509
rect 35161 9469 35173 9503
rect 35207 9500 35219 9503
rect 35526 9500 35532 9512
rect 35207 9472 35532 9500
rect 35207 9469 35219 9472
rect 35161 9463 35219 9469
rect 35526 9460 35532 9472
rect 35584 9460 35590 9512
rect 35621 9503 35679 9509
rect 35621 9469 35633 9503
rect 35667 9500 35679 9503
rect 36170 9500 36176 9512
rect 35667 9472 36176 9500
rect 35667 9469 35679 9472
rect 35621 9463 35679 9469
rect 36170 9460 36176 9472
rect 36228 9460 36234 9512
rect 36280 9500 36308 9540
rect 36648 9540 38792 9568
rect 41064 9540 42892 9568
rect 36648 9500 36676 9540
rect 36906 9500 36912 9512
rect 36280 9472 36676 9500
rect 36867 9472 36912 9500
rect 36906 9460 36912 9472
rect 36964 9460 36970 9512
rect 37090 9500 37096 9512
rect 37051 9472 37096 9500
rect 37090 9460 37096 9472
rect 37148 9460 37154 9512
rect 37277 9503 37335 9509
rect 37277 9469 37289 9503
rect 37323 9500 37335 9503
rect 37918 9500 37924 9512
rect 37323 9472 37924 9500
rect 37323 9469 37335 9472
rect 37277 9463 37335 9469
rect 37918 9460 37924 9472
rect 37976 9460 37982 9512
rect 38289 9503 38347 9509
rect 38289 9500 38301 9503
rect 38120 9472 38301 9500
rect 36538 9432 36544 9444
rect 32140 9404 36544 9432
rect 36538 9392 36544 9404
rect 36596 9392 36602 9444
rect 26421 9367 26479 9373
rect 26421 9364 26433 9367
rect 25372 9336 26433 9364
rect 25372 9324 25378 9336
rect 26421 9333 26433 9336
rect 26467 9333 26479 9367
rect 26421 9327 26479 9333
rect 27430 9324 27436 9376
rect 27488 9364 27494 9376
rect 29914 9364 29920 9376
rect 27488 9336 29920 9364
rect 27488 9324 27494 9336
rect 29914 9324 29920 9336
rect 29972 9324 29978 9376
rect 30006 9324 30012 9376
rect 30064 9364 30070 9376
rect 30745 9367 30803 9373
rect 30745 9364 30757 9367
rect 30064 9336 30757 9364
rect 30064 9324 30070 9336
rect 30745 9333 30757 9336
rect 30791 9333 30803 9367
rect 30745 9327 30803 9333
rect 31110 9324 31116 9376
rect 31168 9364 31174 9376
rect 34977 9367 35035 9373
rect 34977 9364 34989 9367
rect 31168 9336 34989 9364
rect 31168 9324 31174 9336
rect 34977 9333 34989 9336
rect 35023 9364 35035 9367
rect 35897 9367 35955 9373
rect 35897 9364 35909 9367
rect 35023 9336 35909 9364
rect 35023 9333 35035 9336
rect 34977 9327 35035 9333
rect 35897 9333 35909 9336
rect 35943 9364 35955 9367
rect 35986 9364 35992 9376
rect 35943 9336 35992 9364
rect 35943 9333 35955 9336
rect 35897 9327 35955 9333
rect 35986 9324 35992 9336
rect 36044 9324 36050 9376
rect 36170 9324 36176 9376
rect 36228 9364 36234 9376
rect 38120 9364 38148 9472
rect 38289 9469 38301 9472
rect 38335 9469 38347 9503
rect 38289 9463 38347 9469
rect 38197 9435 38255 9441
rect 38197 9401 38209 9435
rect 38243 9432 38255 9435
rect 38654 9432 38660 9444
rect 38243 9404 38660 9432
rect 38243 9401 38255 9404
rect 38197 9395 38255 9401
rect 38654 9392 38660 9404
rect 38712 9392 38718 9444
rect 38764 9432 38792 9540
rect 42886 9528 42892 9540
rect 42944 9528 42950 9580
rect 42978 9528 42984 9580
rect 43036 9568 43042 9580
rect 43036 9540 45600 9568
rect 43036 9528 43042 9540
rect 40313 9503 40371 9509
rect 40313 9469 40325 9503
rect 40359 9500 40371 9503
rect 40402 9500 40408 9512
rect 40359 9472 40408 9500
rect 40359 9469 40371 9472
rect 40313 9463 40371 9469
rect 40402 9460 40408 9472
rect 40460 9460 40466 9512
rect 41230 9500 41236 9512
rect 41191 9472 41236 9500
rect 41230 9460 41236 9472
rect 41288 9460 41294 9512
rect 41414 9460 41420 9512
rect 41472 9500 41478 9512
rect 41598 9500 41604 9512
rect 41472 9472 41517 9500
rect 41559 9472 41604 9500
rect 41472 9460 41478 9472
rect 41598 9460 41604 9472
rect 41656 9460 41662 9512
rect 42334 9460 42340 9512
rect 42392 9500 42398 9512
rect 42613 9503 42671 9509
rect 42613 9500 42625 9503
rect 42392 9472 42625 9500
rect 42392 9460 42398 9472
rect 42613 9469 42625 9472
rect 42659 9469 42671 9503
rect 43898 9500 43904 9512
rect 42613 9463 42671 9469
rect 42720 9472 43904 9500
rect 42720 9432 42748 9472
rect 43898 9460 43904 9472
rect 43956 9460 43962 9512
rect 45572 9500 45600 9540
rect 45646 9528 45652 9580
rect 45704 9568 45710 9580
rect 45704 9540 46888 9568
rect 45704 9528 45710 9540
rect 45925 9503 45983 9509
rect 45572 9472 45876 9500
rect 38764 9404 42748 9432
rect 44082 9392 44088 9444
rect 44140 9432 44146 9444
rect 44140 9404 45784 9432
rect 44140 9392 44146 9404
rect 38841 9367 38899 9373
rect 38841 9364 38853 9367
rect 36228 9336 38853 9364
rect 36228 9324 36234 9336
rect 38841 9333 38853 9336
rect 38887 9333 38899 9367
rect 38841 9327 38899 9333
rect 40034 9324 40040 9376
rect 40092 9364 40098 9376
rect 41598 9364 41604 9376
rect 40092 9336 41604 9364
rect 40092 9324 40098 9336
rect 41598 9324 41604 9336
rect 41656 9324 41662 9376
rect 41690 9324 41696 9376
rect 41748 9364 41754 9376
rect 42061 9367 42119 9373
rect 42061 9364 42073 9367
rect 41748 9336 42073 9364
rect 41748 9324 41754 9336
rect 42061 9333 42073 9336
rect 42107 9333 42119 9367
rect 42061 9327 42119 9333
rect 42337 9367 42395 9373
rect 42337 9333 42349 9367
rect 42383 9364 42395 9367
rect 42978 9364 42984 9376
rect 42383 9336 42984 9364
rect 42383 9333 42395 9336
rect 42337 9327 42395 9333
rect 42978 9324 42984 9336
rect 43036 9324 43042 9376
rect 44818 9364 44824 9376
rect 44779 9336 44824 9364
rect 44818 9324 44824 9336
rect 44876 9324 44882 9376
rect 45756 9373 45784 9404
rect 45741 9367 45799 9373
rect 45741 9333 45753 9367
rect 45787 9333 45799 9367
rect 45848 9364 45876 9472
rect 45925 9469 45937 9503
rect 45971 9500 45983 9503
rect 46014 9500 46020 9512
rect 45971 9472 46020 9500
rect 45971 9469 45983 9472
rect 45925 9463 45983 9469
rect 46014 9460 46020 9472
rect 46072 9460 46078 9512
rect 46860 9509 46888 9540
rect 46845 9503 46903 9509
rect 46845 9469 46857 9503
rect 46891 9500 46903 9503
rect 47504 9500 47532 9599
rect 47854 9596 47860 9608
rect 47912 9596 47918 9648
rect 49528 9636 49556 9676
rect 49602 9664 49608 9716
rect 49660 9704 49666 9716
rect 49660 9676 49705 9704
rect 50264 9676 53328 9704
rect 49660 9664 49666 9676
rect 50264 9636 50292 9676
rect 50430 9636 50436 9648
rect 49528 9608 50292 9636
rect 50391 9608 50436 9636
rect 50430 9596 50436 9608
rect 50488 9596 50494 9648
rect 50709 9639 50767 9645
rect 50709 9605 50721 9639
rect 50755 9636 50767 9639
rect 51258 9636 51264 9648
rect 50755 9608 51264 9636
rect 50755 9605 50767 9608
rect 50709 9599 50767 9605
rect 51258 9596 51264 9608
rect 51316 9636 51322 9648
rect 51445 9639 51503 9645
rect 51445 9636 51457 9639
rect 51316 9608 51457 9636
rect 51316 9596 51322 9608
rect 51445 9605 51457 9608
rect 51491 9605 51503 9639
rect 53300 9636 53328 9676
rect 53834 9664 53840 9716
rect 53892 9704 53898 9716
rect 54021 9707 54079 9713
rect 54021 9704 54033 9707
rect 53892 9676 54033 9704
rect 53892 9664 53898 9676
rect 54021 9673 54033 9676
rect 54067 9704 54079 9707
rect 54386 9704 54392 9716
rect 54067 9676 54392 9704
rect 54067 9673 54079 9676
rect 54021 9667 54079 9673
rect 54386 9664 54392 9676
rect 54444 9664 54450 9716
rect 55398 9704 55404 9716
rect 55359 9676 55404 9704
rect 55398 9664 55404 9676
rect 55456 9664 55462 9716
rect 56042 9664 56048 9716
rect 56100 9704 56106 9716
rect 56410 9704 56416 9716
rect 56100 9676 56416 9704
rect 56100 9664 56106 9676
rect 56410 9664 56416 9676
rect 56468 9664 56474 9716
rect 58158 9704 58164 9716
rect 58119 9676 58164 9704
rect 58158 9664 58164 9676
rect 58216 9664 58222 9716
rect 53653 9639 53711 9645
rect 53653 9636 53665 9639
rect 53300 9608 53665 9636
rect 51445 9599 51503 9605
rect 53576 9580 53604 9608
rect 53653 9605 53665 9608
rect 53699 9605 53711 9639
rect 53653 9599 53711 9605
rect 48314 9568 48320 9580
rect 48275 9540 48320 9568
rect 48314 9528 48320 9540
rect 48372 9528 48378 9580
rect 49234 9528 49240 9580
rect 49292 9568 49298 9580
rect 49292 9540 52132 9568
rect 49292 9528 49298 9540
rect 46891 9472 47532 9500
rect 48041 9503 48099 9509
rect 46891 9469 46903 9472
rect 46845 9463 46903 9469
rect 48041 9469 48053 9503
rect 48087 9500 48099 9503
rect 49694 9500 49700 9512
rect 48087 9472 49700 9500
rect 48087 9469 48099 9472
rect 48041 9463 48099 9469
rect 49694 9460 49700 9472
rect 49752 9500 49758 9512
rect 50246 9500 50252 9512
rect 49752 9472 50252 9500
rect 49752 9460 49758 9472
rect 50246 9460 50252 9472
rect 50304 9460 50310 9512
rect 50522 9500 50528 9512
rect 50435 9472 50528 9500
rect 50522 9460 50528 9472
rect 50580 9500 50586 9512
rect 51718 9500 51724 9512
rect 50580 9472 51120 9500
rect 51679 9472 51724 9500
rect 50580 9460 50586 9472
rect 46385 9435 46443 9441
rect 46385 9401 46397 9435
rect 46431 9432 46443 9435
rect 47210 9432 47216 9444
rect 46431 9404 47216 9432
rect 46431 9401 46443 9404
rect 46385 9395 46443 9401
rect 47210 9392 47216 9404
rect 47268 9392 47274 9444
rect 50062 9432 50068 9444
rect 47688 9404 48176 9432
rect 50023 9404 50068 9432
rect 47688 9364 47716 9404
rect 45848 9336 47716 9364
rect 45741 9327 45799 9333
rect 47762 9324 47768 9376
rect 47820 9364 47826 9376
rect 47857 9367 47915 9373
rect 47857 9364 47869 9367
rect 47820 9336 47869 9364
rect 47820 9324 47826 9336
rect 47857 9333 47869 9336
rect 47903 9364 47915 9367
rect 48038 9364 48044 9376
rect 47903 9336 48044 9364
rect 47903 9333 47915 9336
rect 47857 9327 47915 9333
rect 48038 9324 48044 9336
rect 48096 9324 48102 9376
rect 48148 9364 48176 9404
rect 50062 9392 50068 9404
rect 50120 9432 50126 9444
rect 50338 9432 50344 9444
rect 50120 9404 50344 9432
rect 50120 9392 50126 9404
rect 50338 9392 50344 9404
rect 50396 9392 50402 9444
rect 51092 9432 51120 9472
rect 51718 9460 51724 9472
rect 51776 9460 51782 9512
rect 51810 9460 51816 9512
rect 51868 9500 51874 9512
rect 51997 9503 52055 9509
rect 51997 9500 52009 9503
rect 51868 9472 52009 9500
rect 51868 9460 51874 9472
rect 51997 9469 52009 9472
rect 52043 9469 52055 9503
rect 52104 9500 52132 9540
rect 52362 9528 52368 9580
rect 52420 9568 52426 9580
rect 53101 9571 53159 9577
rect 53101 9568 53113 9571
rect 52420 9540 53113 9568
rect 52420 9528 52426 9540
rect 53101 9537 53113 9540
rect 53147 9568 53159 9571
rect 53282 9568 53288 9580
rect 53147 9540 53288 9568
rect 53147 9537 53159 9540
rect 53101 9531 53159 9537
rect 53282 9528 53288 9540
rect 53340 9528 53346 9580
rect 53558 9528 53564 9580
rect 53616 9528 53622 9580
rect 54404 9568 54432 9664
rect 56502 9596 56508 9648
rect 56560 9636 56566 9648
rect 56781 9639 56839 9645
rect 56781 9636 56793 9639
rect 56560 9608 56793 9636
rect 56560 9596 56566 9608
rect 56781 9605 56793 9608
rect 56827 9605 56839 9639
rect 56781 9599 56839 9605
rect 54573 9571 54631 9577
rect 54573 9568 54585 9571
rect 54404 9540 54585 9568
rect 54573 9537 54585 9540
rect 54619 9537 54631 9571
rect 55122 9568 55128 9580
rect 55083 9540 55128 9568
rect 54573 9531 54631 9537
rect 55122 9528 55128 9540
rect 55180 9528 55186 9580
rect 58176 9568 58204 9664
rect 58621 9571 58679 9577
rect 58621 9568 58633 9571
rect 58176 9540 58633 9568
rect 58621 9537 58633 9540
rect 58667 9537 58679 9571
rect 58621 9531 58679 9537
rect 52638 9500 52644 9512
rect 52104 9472 52644 9500
rect 51997 9463 52055 9469
rect 52638 9460 52644 9472
rect 52696 9460 52702 9512
rect 54665 9503 54723 9509
rect 54665 9469 54677 9503
rect 54711 9500 54723 9503
rect 54938 9500 54944 9512
rect 54711 9472 54944 9500
rect 54711 9469 54723 9472
rect 54665 9463 54723 9469
rect 54938 9460 54944 9472
rect 54996 9460 55002 9512
rect 55953 9503 56011 9509
rect 55953 9500 55965 9503
rect 55784 9472 55965 9500
rect 51092 9404 51212 9432
rect 48774 9364 48780 9376
rect 48148 9336 48780 9364
rect 48774 9324 48780 9336
rect 48832 9364 48838 9376
rect 50890 9364 50896 9376
rect 48832 9336 50896 9364
rect 48832 9324 48838 9336
rect 50890 9324 50896 9336
rect 50948 9324 50954 9376
rect 51184 9373 51212 9404
rect 51169 9367 51227 9373
rect 51169 9333 51181 9367
rect 51215 9364 51227 9367
rect 51442 9364 51448 9376
rect 51215 9336 51448 9364
rect 51215 9333 51227 9336
rect 51169 9327 51227 9333
rect 51442 9324 51448 9336
rect 51500 9324 51506 9376
rect 55674 9324 55680 9376
rect 55732 9364 55738 9376
rect 55784 9373 55812 9472
rect 55953 9469 55965 9472
rect 55999 9469 56011 9503
rect 55953 9463 56011 9469
rect 56134 9460 56140 9512
rect 56192 9500 56198 9512
rect 58342 9500 58348 9512
rect 56192 9472 58348 9500
rect 56192 9460 56198 9472
rect 58342 9460 58348 9472
rect 58400 9460 58406 9512
rect 60550 9500 60556 9512
rect 58452 9472 60556 9500
rect 56045 9435 56103 9441
rect 56045 9401 56057 9435
rect 56091 9432 56103 9435
rect 58452 9432 58480 9472
rect 60550 9460 60556 9472
rect 60608 9460 60614 9512
rect 56091 9404 58480 9432
rect 56091 9401 56103 9404
rect 56045 9395 56103 9401
rect 55769 9367 55827 9373
rect 55769 9364 55781 9367
rect 55732 9336 55781 9364
rect 55732 9324 55738 9336
rect 55769 9333 55781 9336
rect 55815 9333 55827 9367
rect 55769 9327 55827 9333
rect 57330 9324 57336 9376
rect 57388 9364 57394 9376
rect 57790 9364 57796 9376
rect 57388 9336 57796 9364
rect 57388 9324 57394 9336
rect 57790 9324 57796 9336
rect 57848 9324 57854 9376
rect 59725 9367 59783 9373
rect 59725 9333 59737 9367
rect 59771 9364 59783 9367
rect 59814 9364 59820 9376
rect 59771 9336 59820 9364
rect 59771 9333 59783 9336
rect 59725 9327 59783 9333
rect 59814 9324 59820 9336
rect 59872 9324 59878 9376
rect 60458 9364 60464 9376
rect 60419 9336 60464 9364
rect 60458 9324 60464 9336
rect 60516 9324 60522 9376
rect 60921 9367 60979 9373
rect 60921 9333 60933 9367
rect 60967 9364 60979 9367
rect 61286 9364 61292 9376
rect 60967 9336 61292 9364
rect 60967 9333 60979 9336
rect 60921 9327 60979 9333
rect 61286 9324 61292 9336
rect 61344 9324 61350 9376
rect 1104 9274 63480 9296
rect 1104 9222 21774 9274
rect 21826 9222 21838 9274
rect 21890 9222 21902 9274
rect 21954 9222 21966 9274
rect 22018 9222 42566 9274
rect 42618 9222 42630 9274
rect 42682 9222 42694 9274
rect 42746 9222 42758 9274
rect 42810 9222 63480 9274
rect 1104 9200 63480 9222
rect 7837 9163 7895 9169
rect 7837 9160 7849 9163
rect 3160 9132 7849 9160
rect 2590 9024 2596 9036
rect 2551 8996 2596 9024
rect 2590 8984 2596 8996
rect 2648 8984 2654 9036
rect 2866 8984 2872 9036
rect 2924 9024 2930 9036
rect 2961 9027 3019 9033
rect 2961 9024 2973 9027
rect 2924 8996 2973 9024
rect 2924 8984 2930 8996
rect 2961 8993 2973 8996
rect 3007 8993 3019 9027
rect 2961 8987 3019 8993
rect 3050 8984 3056 9036
rect 3108 9024 3114 9036
rect 3160 9024 3188 9132
rect 7837 9129 7849 9132
rect 7883 9129 7895 9163
rect 7837 9123 7895 9129
rect 17218 9120 17224 9172
rect 17276 9160 17282 9172
rect 17276 9132 23060 9160
rect 17276 9120 17282 9132
rect 4706 9052 4712 9104
rect 4764 9092 4770 9104
rect 4801 9095 4859 9101
rect 4801 9092 4813 9095
rect 4764 9064 4813 9092
rect 4764 9052 4770 9064
rect 4801 9061 4813 9064
rect 4847 9092 4859 9095
rect 6733 9095 6791 9101
rect 6733 9092 6745 9095
rect 4847 9064 6745 9092
rect 4847 9061 4859 9064
rect 4801 9055 4859 9061
rect 6733 9061 6745 9064
rect 6779 9061 6791 9095
rect 6733 9055 6791 9061
rect 7098 9052 7104 9104
rect 7156 9092 7162 9104
rect 9677 9095 9735 9101
rect 9677 9092 9689 9095
rect 7156 9064 9689 9092
rect 7156 9052 7162 9064
rect 9677 9061 9689 9064
rect 9723 9061 9735 9095
rect 9677 9055 9735 9061
rect 17773 9095 17831 9101
rect 17773 9061 17785 9095
rect 17819 9092 17831 9095
rect 18414 9092 18420 9104
rect 17819 9064 18420 9092
rect 17819 9061 17831 9064
rect 17773 9055 17831 9061
rect 18414 9052 18420 9064
rect 18472 9052 18478 9104
rect 18598 9092 18604 9104
rect 18559 9064 18604 9092
rect 18598 9052 18604 9064
rect 18656 9052 18662 9104
rect 18690 9052 18696 9104
rect 18748 9092 18754 9104
rect 21634 9092 21640 9104
rect 18748 9064 21640 9092
rect 18748 9052 18754 9064
rect 21634 9052 21640 9064
rect 21692 9052 21698 9104
rect 22833 9095 22891 9101
rect 22833 9092 22845 9095
rect 21744 9064 22845 9092
rect 5721 9027 5779 9033
rect 3108 8996 3201 9024
rect 3108 8984 3114 8996
rect 5721 8993 5733 9027
rect 5767 9024 5779 9027
rect 6546 9024 6552 9036
rect 5767 8996 6552 9024
rect 5767 8993 5779 8996
rect 5721 8987 5779 8993
rect 6546 8984 6552 8996
rect 6604 8984 6610 9036
rect 6641 9027 6699 9033
rect 6641 8993 6653 9027
rect 6687 9024 6699 9027
rect 7190 9024 7196 9036
rect 6687 8996 7196 9024
rect 6687 8993 6699 8996
rect 6641 8987 6699 8993
rect 7190 8984 7196 8996
rect 7248 8984 7254 9036
rect 7282 8984 7288 9036
rect 7340 9024 7346 9036
rect 7561 9027 7619 9033
rect 7561 9024 7573 9027
rect 7340 8996 7573 9024
rect 7340 8984 7346 8996
rect 7561 8993 7573 8996
rect 7607 9024 7619 9027
rect 8018 9024 8024 9036
rect 7607 8996 8024 9024
rect 7607 8993 7619 8996
rect 7561 8987 7619 8993
rect 8018 8984 8024 8996
rect 8076 8984 8082 9036
rect 8754 9024 8760 9036
rect 8715 8996 8760 9024
rect 8754 8984 8760 8996
rect 8812 8984 8818 9036
rect 9493 9027 9551 9033
rect 9493 8993 9505 9027
rect 9539 9024 9551 9027
rect 10134 9024 10140 9036
rect 9539 8996 10140 9024
rect 9539 8993 9551 8996
rect 9493 8987 9551 8993
rect 10134 8984 10140 8996
rect 10192 8984 10198 9036
rect 10502 9024 10508 9036
rect 10463 8996 10508 9024
rect 10502 8984 10508 8996
rect 10560 8984 10566 9036
rect 10870 8984 10876 9036
rect 10928 9024 10934 9036
rect 12342 9024 12348 9036
rect 10928 8996 12204 9024
rect 12303 8996 12348 9024
rect 10928 8984 10934 8996
rect 4338 8916 4344 8968
rect 4396 8956 4402 8968
rect 4893 8959 4951 8965
rect 4893 8956 4905 8959
rect 4396 8928 4905 8956
rect 4396 8916 4402 8928
rect 4893 8925 4905 8928
rect 4939 8925 4951 8959
rect 5442 8956 5448 8968
rect 5403 8928 5448 8956
rect 4893 8919 4951 8925
rect 5442 8916 5448 8928
rect 5500 8916 5506 8968
rect 5905 8959 5963 8965
rect 5905 8925 5917 8959
rect 5951 8956 5963 8959
rect 7653 8959 7711 8965
rect 5951 8928 6316 8956
rect 5951 8925 5963 8928
rect 5905 8919 5963 8925
rect 2409 8891 2467 8897
rect 2409 8857 2421 8891
rect 2455 8888 2467 8891
rect 4154 8888 4160 8900
rect 2455 8860 4160 8888
rect 2455 8857 2467 8860
rect 2409 8851 2467 8857
rect 4154 8848 4160 8860
rect 4212 8848 4218 8900
rect 6288 8832 6316 8928
rect 7653 8925 7665 8959
rect 7699 8956 7711 8959
rect 7837 8959 7895 8965
rect 7837 8956 7849 8959
rect 7699 8928 7849 8956
rect 7699 8925 7711 8928
rect 7653 8919 7711 8925
rect 7837 8925 7849 8928
rect 7883 8956 7895 8959
rect 8113 8959 8171 8965
rect 8113 8956 8125 8959
rect 7883 8928 8125 8956
rect 7883 8925 7895 8928
rect 7837 8919 7895 8925
rect 8113 8925 8125 8928
rect 8159 8956 8171 8959
rect 10594 8956 10600 8968
rect 8159 8928 10600 8956
rect 8159 8925 8171 8928
rect 8113 8919 8171 8925
rect 10594 8916 10600 8928
rect 10652 8916 10658 8968
rect 10778 8916 10784 8968
rect 10836 8956 10842 8968
rect 11517 8959 11575 8965
rect 11517 8956 11529 8959
rect 10836 8928 11529 8956
rect 10836 8916 10842 8928
rect 11517 8925 11529 8928
rect 11563 8925 11575 8959
rect 11517 8919 11575 8925
rect 12069 8959 12127 8965
rect 12069 8925 12081 8959
rect 12115 8925 12127 8959
rect 12176 8956 12204 8996
rect 12342 8984 12348 8996
rect 12400 8984 12406 9036
rect 12986 8984 12992 9036
rect 13044 9024 13050 9036
rect 13538 9024 13544 9036
rect 13044 8996 13544 9024
rect 13044 8984 13050 8996
rect 13538 8984 13544 8996
rect 13596 8984 13602 9036
rect 13722 9024 13728 9036
rect 13683 8996 13728 9024
rect 13722 8984 13728 8996
rect 13780 9024 13786 9036
rect 15381 9027 15439 9033
rect 15381 9024 15393 9027
rect 13780 8996 15393 9024
rect 13780 8984 13786 8996
rect 15381 8993 15393 8996
rect 15427 9024 15439 9027
rect 15930 9024 15936 9036
rect 15427 8996 15936 9024
rect 15427 8993 15439 8996
rect 15381 8987 15439 8993
rect 15930 8984 15936 8996
rect 15988 8984 15994 9036
rect 16022 8984 16028 9036
rect 16080 9024 16086 9036
rect 16758 9024 16764 9036
rect 16080 8996 16764 9024
rect 16080 8984 16086 8996
rect 16758 8984 16764 8996
rect 16816 8984 16822 9036
rect 17013 9027 17071 9033
rect 17013 9024 17025 9027
rect 16868 8996 17025 9024
rect 12526 8956 12532 8968
rect 12176 8928 12532 8956
rect 12069 8919 12127 8925
rect 8202 8848 8208 8900
rect 8260 8888 8266 8900
rect 9033 8891 9091 8897
rect 9033 8888 9045 8891
rect 8260 8860 9045 8888
rect 8260 8848 8266 8860
rect 9033 8857 9045 8860
rect 9079 8857 9091 8891
rect 11146 8888 11152 8900
rect 11107 8860 11152 8888
rect 9033 8851 9091 8857
rect 11146 8848 11152 8860
rect 11204 8848 11210 8900
rect 12084 8888 12112 8919
rect 12526 8916 12532 8928
rect 12584 8916 12590 8968
rect 12897 8959 12955 8965
rect 12897 8956 12909 8959
rect 12636 8928 12909 8956
rect 12636 8888 12664 8928
rect 12897 8925 12909 8928
rect 12943 8956 12955 8959
rect 12943 8928 13584 8956
rect 12943 8925 12955 8928
rect 12897 8919 12955 8925
rect 13357 8891 13415 8897
rect 13357 8888 13369 8891
rect 12084 8860 12664 8888
rect 12728 8860 13369 8888
rect 4062 8780 4068 8832
rect 4120 8820 4126 8832
rect 4249 8823 4307 8829
rect 4249 8820 4261 8823
rect 4120 8792 4261 8820
rect 4120 8780 4126 8792
rect 4249 8789 4261 8792
rect 4295 8820 4307 8823
rect 4798 8820 4804 8832
rect 4295 8792 4804 8820
rect 4295 8789 4307 8792
rect 4249 8783 4307 8789
rect 4798 8780 4804 8792
rect 4856 8780 4862 8832
rect 6270 8820 6276 8832
rect 6231 8792 6276 8820
rect 6270 8780 6276 8792
rect 6328 8780 6334 8832
rect 6362 8780 6368 8832
rect 6420 8820 6426 8832
rect 10502 8820 10508 8832
rect 6420 8792 10508 8820
rect 6420 8780 6426 8792
rect 10502 8780 10508 8792
rect 10560 8780 10566 8832
rect 12250 8780 12256 8832
rect 12308 8820 12314 8832
rect 12728 8820 12756 8860
rect 13357 8857 13369 8860
rect 13403 8857 13415 8891
rect 13556 8888 13584 8928
rect 13630 8916 13636 8968
rect 13688 8956 13694 8968
rect 15289 8959 15347 8965
rect 13688 8928 13733 8956
rect 13688 8916 13694 8928
rect 15289 8925 15301 8959
rect 15335 8956 15347 8959
rect 16114 8956 16120 8968
rect 15335 8928 16120 8956
rect 15335 8925 15347 8928
rect 15289 8919 15347 8925
rect 16114 8916 16120 8928
rect 16172 8916 16178 8968
rect 16390 8916 16396 8968
rect 16448 8956 16454 8968
rect 16868 8956 16896 8996
rect 17013 8993 17025 8996
rect 17059 8993 17071 9027
rect 17013 8987 17071 8993
rect 17310 8984 17316 9036
rect 17368 9024 17374 9036
rect 19061 9027 19119 9033
rect 17368 8996 17413 9024
rect 17368 8984 17374 8996
rect 19061 8993 19073 9027
rect 19107 9024 19119 9027
rect 19150 9024 19156 9036
rect 19107 8996 19156 9024
rect 19107 8993 19119 8996
rect 19061 8987 19119 8993
rect 19150 8984 19156 8996
rect 19208 8984 19214 9036
rect 19242 8984 19248 9036
rect 19300 9024 19306 9036
rect 19429 9027 19487 9033
rect 19300 8996 19345 9024
rect 19300 8984 19306 8996
rect 19429 8993 19441 9027
rect 19475 8993 19487 9027
rect 19429 8987 19487 8993
rect 20993 9027 21051 9033
rect 20993 8993 21005 9027
rect 21039 8993 21051 9027
rect 21450 9024 21456 9036
rect 21411 8996 21456 9024
rect 20993 8987 21051 8993
rect 17218 8956 17224 8968
rect 16448 8928 16896 8956
rect 17179 8928 17224 8956
rect 16448 8916 16454 8928
rect 17218 8916 17224 8928
rect 17276 8916 17282 8968
rect 17494 8916 17500 8968
rect 17552 8956 17558 8968
rect 19334 8956 19340 8968
rect 17552 8928 19340 8956
rect 17552 8916 17558 8928
rect 19334 8916 19340 8928
rect 19392 8916 19398 8968
rect 19444 8956 19472 8987
rect 19702 8956 19708 8968
rect 19444 8928 19708 8956
rect 19702 8916 19708 8928
rect 19760 8956 19766 8968
rect 20625 8959 20683 8965
rect 20625 8956 20637 8959
rect 19760 8928 20637 8956
rect 19760 8916 19766 8928
rect 20625 8925 20637 8928
rect 20671 8925 20683 8959
rect 20898 8956 20904 8968
rect 20859 8928 20904 8956
rect 20625 8919 20683 8925
rect 20898 8916 20904 8928
rect 20956 8916 20962 8968
rect 21008 8956 21036 8987
rect 21450 8984 21456 8996
rect 21508 8984 21514 9036
rect 21542 8984 21548 9036
rect 21600 9024 21606 9036
rect 21744 9024 21772 9064
rect 22833 9061 22845 9064
rect 22879 9061 22891 9095
rect 23032 9092 23060 9132
rect 23106 9120 23112 9172
rect 23164 9160 23170 9172
rect 23569 9163 23627 9169
rect 23569 9160 23581 9163
rect 23164 9132 23581 9160
rect 23164 9120 23170 9132
rect 23569 9129 23581 9132
rect 23615 9160 23627 9163
rect 33318 9160 33324 9172
rect 23615 9132 30972 9160
rect 23615 9129 23627 9132
rect 23569 9123 23627 9129
rect 24581 9095 24639 9101
rect 23032 9064 24072 9092
rect 22833 9055 22891 9061
rect 22370 9024 22376 9036
rect 21600 8996 21772 9024
rect 21836 8996 22376 9024
rect 21600 8984 21606 8996
rect 21266 8956 21272 8968
rect 21008 8928 21272 8956
rect 21266 8916 21272 8928
rect 21324 8956 21330 8968
rect 21836 8956 21864 8996
rect 22370 8984 22376 8996
rect 22428 8984 22434 9036
rect 22278 8956 22284 8968
rect 21324 8928 21864 8956
rect 22239 8928 22284 8956
rect 21324 8916 21330 8928
rect 22278 8916 22284 8928
rect 22336 8916 22342 8968
rect 22554 8916 22560 8968
rect 22612 8956 22618 8968
rect 23201 8959 23259 8965
rect 23201 8956 23213 8959
rect 22612 8928 23213 8956
rect 22612 8916 22618 8928
rect 23201 8925 23213 8928
rect 23247 8956 23259 8959
rect 23934 8956 23940 8968
rect 23247 8928 23940 8956
rect 23247 8925 23259 8928
rect 23201 8919 23259 8925
rect 23934 8916 23940 8928
rect 23992 8916 23998 8968
rect 24044 8956 24072 9064
rect 24581 9061 24593 9095
rect 24627 9092 24639 9095
rect 24854 9092 24860 9104
rect 24627 9064 24860 9092
rect 24627 9061 24639 9064
rect 24581 9055 24639 9061
rect 24854 9052 24860 9064
rect 24912 9052 24918 9104
rect 30282 9092 30288 9104
rect 24964 9064 25268 9092
rect 24394 8984 24400 9036
rect 24452 9024 24458 9036
rect 24964 9024 24992 9064
rect 24452 8996 24992 9024
rect 24452 8984 24458 8996
rect 25038 8984 25044 9036
rect 25096 9024 25102 9036
rect 25240 9033 25268 9064
rect 25516 9064 30288 9092
rect 25225 9027 25283 9033
rect 25096 8996 25141 9024
rect 25096 8984 25102 8996
rect 25225 8993 25237 9027
rect 25271 8993 25283 9027
rect 25406 9024 25412 9036
rect 25367 8996 25412 9024
rect 25225 8987 25283 8993
rect 25406 8984 25412 8996
rect 25464 8984 25470 9036
rect 25516 8956 25544 9064
rect 30282 9052 30288 9064
rect 30340 9052 30346 9104
rect 30374 9052 30380 9104
rect 30432 9092 30438 9104
rect 30469 9095 30527 9101
rect 30469 9092 30481 9095
rect 30432 9064 30481 9092
rect 30432 9052 30438 9064
rect 30469 9061 30481 9064
rect 30515 9061 30527 9095
rect 30944 9092 30972 9132
rect 31588 9132 33324 9160
rect 31588 9092 31616 9132
rect 33318 9120 33324 9132
rect 33376 9120 33382 9172
rect 33502 9160 33508 9172
rect 33463 9132 33508 9160
rect 33502 9120 33508 9132
rect 33560 9120 33566 9172
rect 34514 9120 34520 9172
rect 34572 9160 34578 9172
rect 36446 9160 36452 9172
rect 34572 9132 36452 9160
rect 34572 9120 34578 9132
rect 36446 9120 36452 9132
rect 36504 9120 36510 9172
rect 36538 9120 36544 9172
rect 36596 9160 36602 9172
rect 49145 9163 49203 9169
rect 36596 9132 49004 9160
rect 36596 9120 36602 9132
rect 33686 9092 33692 9104
rect 30944 9064 31616 9092
rect 33647 9064 33692 9092
rect 30469 9055 30527 9061
rect 33686 9052 33692 9064
rect 33744 9052 33750 9104
rect 34606 9092 34612 9104
rect 34164 9064 34612 9092
rect 26142 8984 26148 9036
rect 26200 9024 26206 9036
rect 27341 9027 27399 9033
rect 27341 9024 27353 9027
rect 26200 8996 27353 9024
rect 26200 8984 26206 8996
rect 27341 8993 27353 8996
rect 27387 9024 27399 9027
rect 27801 9027 27859 9033
rect 27801 9024 27813 9027
rect 27387 8996 27813 9024
rect 27387 8993 27399 8996
rect 27341 8987 27399 8993
rect 27801 8993 27813 8996
rect 27847 8993 27859 9027
rect 28442 9024 28448 9036
rect 28403 8996 28448 9024
rect 27801 8987 27859 8993
rect 28442 8984 28448 8996
rect 28500 8984 28506 9036
rect 30006 9024 30012 9036
rect 29967 8996 30012 9024
rect 30006 8984 30012 8996
rect 30064 8984 30070 9036
rect 30098 8984 30104 9036
rect 30156 9024 30162 9036
rect 31113 9027 31171 9033
rect 31113 9024 31125 9027
rect 30156 8996 31125 9024
rect 30156 8984 30162 8996
rect 31113 8993 31125 8996
rect 31159 8993 31171 9027
rect 32398 9024 32404 9036
rect 32359 8996 32404 9024
rect 31113 8987 31171 8993
rect 32398 8984 32404 8996
rect 32456 8984 32462 9036
rect 34164 9033 34192 9064
rect 34606 9052 34612 9064
rect 34664 9052 34670 9104
rect 34882 9052 34888 9104
rect 34940 9092 34946 9104
rect 34940 9064 37228 9092
rect 34940 9052 34946 9064
rect 34149 9027 34207 9033
rect 34149 8993 34161 9027
rect 34195 8993 34207 9027
rect 34514 9024 34520 9036
rect 34475 8996 34520 9024
rect 34149 8987 34207 8993
rect 34514 8984 34520 8996
rect 34572 8984 34578 9036
rect 34698 8984 34704 9036
rect 34756 9024 34762 9036
rect 35621 9027 35679 9033
rect 35621 9024 35633 9027
rect 34756 8996 35633 9024
rect 34756 8984 34762 8996
rect 35621 8993 35633 8996
rect 35667 9024 35679 9027
rect 36357 9027 36415 9033
rect 36357 9024 36369 9027
rect 35667 8996 36369 9024
rect 35667 8993 35679 8996
rect 35621 8987 35679 8993
rect 36357 8993 36369 8996
rect 36403 8993 36415 9027
rect 37200 9024 37228 9064
rect 37274 9052 37280 9104
rect 37332 9092 37338 9104
rect 37921 9095 37979 9101
rect 37921 9092 37933 9095
rect 37332 9064 37933 9092
rect 37332 9052 37338 9064
rect 37921 9061 37933 9064
rect 37967 9061 37979 9095
rect 38286 9092 38292 9104
rect 38247 9064 38292 9092
rect 37921 9055 37979 9061
rect 37936 9024 37964 9055
rect 38286 9052 38292 9064
rect 38344 9052 38350 9104
rect 39482 9052 39488 9104
rect 39540 9092 39546 9104
rect 42337 9095 42395 9101
rect 42337 9092 42349 9095
rect 39540 9064 42349 9092
rect 39540 9052 39546 9064
rect 42337 9061 42349 9064
rect 42383 9061 42395 9095
rect 42337 9055 42395 9061
rect 43901 9095 43959 9101
rect 43901 9061 43913 9095
rect 43947 9092 43959 9095
rect 44818 9092 44824 9104
rect 43947 9064 44824 9092
rect 43947 9061 43959 9064
rect 43901 9055 43959 9061
rect 44818 9052 44824 9064
rect 44876 9052 44882 9104
rect 47765 9095 47823 9101
rect 47765 9061 47777 9095
rect 47811 9092 47823 9095
rect 48682 9092 48688 9104
rect 47811 9064 48688 9092
rect 47811 9061 47823 9064
rect 47765 9055 47823 9061
rect 48682 9052 48688 9064
rect 48740 9052 48746 9104
rect 48976 9092 49004 9132
rect 49145 9129 49157 9163
rect 49191 9160 49203 9163
rect 49326 9160 49332 9172
rect 49191 9132 49332 9160
rect 49191 9129 49203 9132
rect 49145 9123 49203 9129
rect 49326 9120 49332 9132
rect 49384 9120 49390 9172
rect 49970 9120 49976 9172
rect 50028 9160 50034 9172
rect 60642 9160 60648 9172
rect 50028 9132 60648 9160
rect 50028 9120 50034 9132
rect 60642 9120 60648 9132
rect 60700 9160 60706 9172
rect 61841 9163 61899 9169
rect 61841 9160 61853 9163
rect 60700 9132 61853 9160
rect 60700 9120 60706 9132
rect 61841 9129 61853 9132
rect 61887 9129 61899 9163
rect 61841 9123 61899 9129
rect 49605 9095 49663 9101
rect 49605 9092 49617 9095
rect 48976 9064 49617 9092
rect 40034 9024 40040 9036
rect 37200 8996 37872 9024
rect 37936 8996 40040 9024
rect 36357 8987 36415 8993
rect 24044 8928 25544 8956
rect 26513 8959 26571 8965
rect 26513 8925 26525 8959
rect 26559 8925 26571 8959
rect 26513 8919 26571 8925
rect 27065 8959 27123 8965
rect 27065 8925 27077 8959
rect 27111 8956 27123 8959
rect 27154 8956 27160 8968
rect 27111 8928 27160 8956
rect 27111 8925 27123 8928
rect 27065 8919 27123 8925
rect 13998 8888 14004 8900
rect 13556 8860 14004 8888
rect 13357 8851 13415 8857
rect 13998 8848 14004 8860
rect 14056 8888 14062 8900
rect 14553 8891 14611 8897
rect 14553 8888 14565 8891
rect 14056 8860 14565 8888
rect 14056 8848 14062 8860
rect 14553 8857 14565 8860
rect 14599 8888 14611 8891
rect 26528 8888 26556 8919
rect 27154 8916 27160 8928
rect 27212 8916 27218 8968
rect 27525 8959 27583 8965
rect 27525 8925 27537 8959
rect 27571 8925 27583 8959
rect 28350 8956 28356 8968
rect 28263 8928 28356 8956
rect 27525 8919 27583 8925
rect 14599 8860 26556 8888
rect 14599 8857 14611 8860
rect 14553 8851 14611 8857
rect 26602 8848 26608 8900
rect 26660 8888 26666 8900
rect 27430 8888 27436 8900
rect 26660 8860 27436 8888
rect 26660 8848 26666 8860
rect 27430 8848 27436 8860
rect 27488 8888 27494 8900
rect 27540 8888 27568 8919
rect 28350 8916 28356 8928
rect 28408 8956 28414 8968
rect 28810 8956 28816 8968
rect 28408 8928 28816 8956
rect 28408 8916 28414 8928
rect 28810 8916 28816 8928
rect 28868 8916 28874 8968
rect 29454 8916 29460 8968
rect 29512 8956 29518 8968
rect 29917 8959 29975 8965
rect 29917 8956 29929 8959
rect 29512 8928 29929 8956
rect 29512 8916 29518 8928
rect 29917 8925 29929 8928
rect 29963 8956 29975 8959
rect 30742 8956 30748 8968
rect 29963 8928 30748 8956
rect 29963 8925 29975 8928
rect 29917 8919 29975 8925
rect 30742 8916 30748 8928
rect 30800 8916 30806 8968
rect 32309 8959 32367 8965
rect 32309 8925 32321 8959
rect 32355 8956 32367 8959
rect 32766 8956 32772 8968
rect 32355 8928 32772 8956
rect 32355 8925 32367 8928
rect 32309 8919 32367 8925
rect 32766 8916 32772 8928
rect 32824 8916 32830 8968
rect 32861 8959 32919 8965
rect 32861 8925 32873 8959
rect 32907 8925 32919 8959
rect 32861 8919 32919 8925
rect 34609 8959 34667 8965
rect 34609 8925 34621 8959
rect 34655 8956 34667 8959
rect 34790 8956 34796 8968
rect 34655 8928 34796 8956
rect 34655 8925 34667 8928
rect 34609 8919 34667 8925
rect 27488 8860 27568 8888
rect 27488 8848 27494 8860
rect 27614 8848 27620 8900
rect 27672 8888 27678 8900
rect 28169 8891 28227 8897
rect 28169 8888 28181 8891
rect 27672 8860 28181 8888
rect 27672 8848 27678 8860
rect 28169 8857 28181 8860
rect 28215 8857 28227 8891
rect 32876 8888 32904 8919
rect 34790 8916 34796 8928
rect 34848 8916 34854 8968
rect 35526 8956 35532 8968
rect 35487 8928 35532 8956
rect 35526 8916 35532 8928
rect 35584 8916 35590 8968
rect 35710 8916 35716 8968
rect 35768 8956 35774 8968
rect 36081 8959 36139 8965
rect 36081 8956 36093 8959
rect 35768 8928 36093 8956
rect 35768 8916 35774 8928
rect 36081 8925 36093 8928
rect 36127 8956 36139 8959
rect 36127 8928 37228 8956
rect 36127 8925 36139 8928
rect 36081 8919 36139 8925
rect 36262 8888 36268 8900
rect 32876 8860 36268 8888
rect 28169 8851 28227 8857
rect 36262 8848 36268 8860
rect 36320 8848 36326 8900
rect 37200 8832 37228 8928
rect 12308 8792 12756 8820
rect 12308 8780 12314 8792
rect 12986 8780 12992 8832
rect 13044 8820 13050 8832
rect 13173 8823 13231 8829
rect 13173 8820 13185 8823
rect 13044 8792 13185 8820
rect 13044 8780 13050 8792
rect 13173 8789 13185 8792
rect 13219 8789 13231 8823
rect 13173 8783 13231 8789
rect 13814 8780 13820 8832
rect 13872 8820 13878 8832
rect 13909 8823 13967 8829
rect 13909 8820 13921 8823
rect 13872 8792 13921 8820
rect 13872 8780 13878 8792
rect 13909 8789 13921 8792
rect 13955 8789 13967 8823
rect 13909 8783 13967 8789
rect 15105 8823 15163 8829
rect 15105 8789 15117 8823
rect 15151 8820 15163 8823
rect 15194 8820 15200 8832
rect 15151 8792 15200 8820
rect 15151 8789 15163 8792
rect 15105 8783 15163 8789
rect 15194 8780 15200 8792
rect 15252 8780 15258 8832
rect 15470 8780 15476 8832
rect 15528 8820 15534 8832
rect 15565 8823 15623 8829
rect 15565 8820 15577 8823
rect 15528 8792 15577 8820
rect 15528 8780 15534 8792
rect 15565 8789 15577 8792
rect 15611 8789 15623 8823
rect 16114 8820 16120 8832
rect 16075 8792 16120 8820
rect 15565 8783 15623 8789
rect 16114 8780 16120 8792
rect 16172 8780 16178 8832
rect 16758 8820 16764 8832
rect 16719 8792 16764 8820
rect 16758 8780 16764 8792
rect 16816 8780 16822 8832
rect 16850 8780 16856 8832
rect 16908 8820 16914 8832
rect 16908 8792 16953 8820
rect 16908 8780 16914 8792
rect 17402 8780 17408 8832
rect 17460 8820 17466 8832
rect 18138 8820 18144 8832
rect 17460 8792 18144 8820
rect 17460 8780 17466 8792
rect 18138 8780 18144 8792
rect 18196 8820 18202 8832
rect 18233 8823 18291 8829
rect 18233 8820 18245 8823
rect 18196 8792 18245 8820
rect 18196 8780 18202 8792
rect 18233 8789 18245 8792
rect 18279 8789 18291 8823
rect 18233 8783 18291 8789
rect 18506 8780 18512 8832
rect 18564 8820 18570 8832
rect 19886 8820 19892 8832
rect 18564 8792 19892 8820
rect 18564 8780 18570 8792
rect 19886 8780 19892 8792
rect 19944 8780 19950 8832
rect 19981 8823 20039 8829
rect 19981 8789 19993 8823
rect 20027 8820 20039 8823
rect 20254 8820 20260 8832
rect 20027 8792 20260 8820
rect 20027 8789 20039 8792
rect 19981 8783 20039 8789
rect 20254 8780 20260 8792
rect 20312 8780 20318 8832
rect 20346 8780 20352 8832
rect 20404 8820 20410 8832
rect 20404 8792 20449 8820
rect 20404 8780 20410 8792
rect 21542 8780 21548 8832
rect 21600 8820 21606 8832
rect 21729 8823 21787 8829
rect 21729 8820 21741 8823
rect 21600 8792 21741 8820
rect 21600 8780 21606 8792
rect 21729 8789 21741 8792
rect 21775 8789 21787 8823
rect 21729 8783 21787 8789
rect 21818 8780 21824 8832
rect 21876 8820 21882 8832
rect 22097 8823 22155 8829
rect 22097 8820 22109 8823
rect 21876 8792 22109 8820
rect 21876 8780 21882 8792
rect 22097 8789 22109 8792
rect 22143 8789 22155 8823
rect 22097 8783 22155 8789
rect 23474 8780 23480 8832
rect 23532 8820 23538 8832
rect 24029 8823 24087 8829
rect 24029 8820 24041 8823
rect 23532 8792 24041 8820
rect 23532 8780 23538 8792
rect 24029 8789 24041 8792
rect 24075 8789 24087 8823
rect 24394 8820 24400 8832
rect 24355 8792 24400 8820
rect 24029 8783 24087 8789
rect 24394 8780 24400 8792
rect 24452 8780 24458 8832
rect 25866 8820 25872 8832
rect 25827 8792 25872 8820
rect 25866 8780 25872 8792
rect 25924 8780 25930 8832
rect 26234 8820 26240 8832
rect 26195 8792 26240 8820
rect 26234 8780 26240 8792
rect 26292 8820 26298 8832
rect 27706 8820 27712 8832
rect 26292 8792 27712 8820
rect 26292 8780 26298 8792
rect 27706 8780 27712 8792
rect 27764 8780 27770 8832
rect 28626 8820 28632 8832
rect 28587 8792 28632 8820
rect 28626 8780 28632 8792
rect 28684 8780 28690 8832
rect 29270 8820 29276 8832
rect 29231 8792 29276 8820
rect 29270 8780 29276 8792
rect 29328 8780 29334 8832
rect 29362 8780 29368 8832
rect 29420 8820 29426 8832
rect 29641 8823 29699 8829
rect 29641 8820 29653 8823
rect 29420 8792 29653 8820
rect 29420 8780 29426 8792
rect 29641 8789 29653 8792
rect 29687 8789 29699 8823
rect 29641 8783 29699 8789
rect 31202 8780 31208 8832
rect 31260 8820 31266 8832
rect 31573 8823 31631 8829
rect 31573 8820 31585 8823
rect 31260 8792 31585 8820
rect 31260 8780 31266 8792
rect 31573 8789 31585 8792
rect 31619 8820 31631 8823
rect 31941 8823 31999 8829
rect 31941 8820 31953 8823
rect 31619 8792 31953 8820
rect 31619 8789 31631 8792
rect 31573 8783 31631 8789
rect 31941 8789 31953 8792
rect 31987 8820 31999 8823
rect 33410 8820 33416 8832
rect 31987 8792 33416 8820
rect 31987 8789 31999 8792
rect 31941 8783 31999 8789
rect 33410 8780 33416 8792
rect 33468 8780 33474 8832
rect 33870 8780 33876 8832
rect 33928 8820 33934 8832
rect 34882 8820 34888 8832
rect 33928 8792 34888 8820
rect 33928 8780 33934 8792
rect 34882 8780 34888 8792
rect 34940 8780 34946 8832
rect 35066 8820 35072 8832
rect 35027 8792 35072 8820
rect 35066 8780 35072 8792
rect 35124 8780 35130 8832
rect 36722 8820 36728 8832
rect 36683 8792 36728 8820
rect 36722 8780 36728 8792
rect 36780 8780 36786 8832
rect 37182 8820 37188 8832
rect 37143 8792 37188 8820
rect 37182 8780 37188 8792
rect 37240 8780 37246 8832
rect 37844 8820 37872 8996
rect 40034 8984 40040 8996
rect 40092 8984 40098 9036
rect 41690 9024 41696 9036
rect 41524 8996 41696 9024
rect 38470 8956 38476 8968
rect 38431 8928 38476 8956
rect 38470 8916 38476 8928
rect 38528 8916 38534 8968
rect 38746 8956 38752 8968
rect 38707 8928 38752 8956
rect 38746 8916 38752 8928
rect 38804 8916 38810 8968
rect 38838 8916 38844 8968
rect 38896 8956 38902 8968
rect 41524 8956 41552 8996
rect 41690 8984 41696 8996
rect 41748 9024 41754 9036
rect 41877 9027 41935 9033
rect 41877 9024 41889 9027
rect 41748 8996 41889 9024
rect 41748 8984 41754 8996
rect 41877 8993 41889 8996
rect 41923 8993 41935 9027
rect 41877 8987 41935 8993
rect 41966 8984 41972 9036
rect 42024 9024 42030 9036
rect 43441 9027 43499 9033
rect 43441 9024 43453 9027
rect 42024 8996 43453 9024
rect 42024 8984 42030 8996
rect 43441 8993 43453 8996
rect 43487 9024 43499 9027
rect 43530 9024 43536 9036
rect 43487 8996 43536 9024
rect 43487 8993 43499 8996
rect 43441 8987 43499 8993
rect 43530 8984 43536 8996
rect 43588 9024 43594 9036
rect 44358 9024 44364 9036
rect 43588 8996 44364 9024
rect 43588 8984 43594 8996
rect 44358 8984 44364 8996
rect 44416 8984 44422 9036
rect 47394 9033 47400 9036
rect 47346 9027 47400 9033
rect 47346 8993 47358 9027
rect 47392 8993 47400 9027
rect 47346 8987 47400 8993
rect 47394 8984 47400 8987
rect 47452 9024 47458 9036
rect 48976 9033 49004 9064
rect 49605 9061 49617 9064
rect 49651 9092 49663 9095
rect 50522 9092 50528 9104
rect 49651 9064 50528 9092
rect 49651 9061 49663 9064
rect 49605 9055 49663 9061
rect 50522 9052 50528 9064
rect 50580 9052 50586 9104
rect 51166 9092 51172 9104
rect 50724 9064 51172 9092
rect 50724 9033 50752 9064
rect 51166 9052 51172 9064
rect 51224 9052 51230 9104
rect 52362 9092 52368 9104
rect 51368 9064 52368 9092
rect 51368 9036 51396 9064
rect 52362 9052 52368 9064
rect 52420 9052 52426 9104
rect 52454 9052 52460 9104
rect 52512 9092 52518 9104
rect 52641 9095 52699 9101
rect 52641 9092 52653 9095
rect 52512 9064 52653 9092
rect 52512 9052 52518 9064
rect 52641 9061 52653 9064
rect 52687 9061 52699 9095
rect 52641 9055 52699 9061
rect 54202 9052 54208 9104
rect 54260 9092 54266 9104
rect 54297 9095 54355 9101
rect 54297 9092 54309 9095
rect 54260 9064 54309 9092
rect 54260 9052 54266 9064
rect 54297 9061 54309 9064
rect 54343 9092 54355 9095
rect 54343 9064 55996 9092
rect 54343 9061 54355 9064
rect 54297 9055 54355 9061
rect 48041 9027 48099 9033
rect 48041 9024 48053 9027
rect 47452 8996 48053 9024
rect 47452 8984 47458 8996
rect 48041 8993 48053 8996
rect 48087 8993 48099 9027
rect 48041 8987 48099 8993
rect 48961 9027 49019 9033
rect 48961 8993 48973 9027
rect 49007 8993 49019 9027
rect 48961 8987 49019 8993
rect 49329 9027 49387 9033
rect 49329 8993 49341 9027
rect 49375 9024 49387 9027
rect 50709 9027 50767 9033
rect 49375 8996 50292 9024
rect 49375 8993 49387 8996
rect 49329 8987 49387 8993
rect 38896 8928 41552 8956
rect 38896 8916 38902 8928
rect 41598 8916 41604 8968
rect 41656 8956 41662 8968
rect 41785 8959 41843 8965
rect 41656 8928 41701 8956
rect 41656 8916 41662 8928
rect 41785 8925 41797 8959
rect 41831 8956 41843 8959
rect 42242 8956 42248 8968
rect 41831 8928 42248 8956
rect 41831 8925 41843 8928
rect 41785 8919 41843 8925
rect 42242 8916 42248 8928
rect 42300 8916 42306 8968
rect 43346 8916 43352 8968
rect 43404 8956 43410 8968
rect 43404 8928 43449 8956
rect 43404 8916 43410 8928
rect 44082 8916 44088 8968
rect 44140 8956 44146 8968
rect 44729 8959 44787 8965
rect 44729 8956 44741 8959
rect 44140 8928 44741 8956
rect 44140 8916 44146 8928
rect 44729 8925 44741 8928
rect 44775 8925 44787 8959
rect 44729 8919 44787 8925
rect 45005 8959 45063 8965
rect 45005 8925 45017 8959
rect 45051 8956 45063 8959
rect 45094 8956 45100 8968
rect 45051 8928 45100 8956
rect 45051 8925 45063 8928
rect 45005 8919 45063 8925
rect 45094 8916 45100 8928
rect 45152 8916 45158 8968
rect 47213 8959 47271 8965
rect 47213 8925 47225 8959
rect 47259 8956 47271 8959
rect 47762 8956 47768 8968
rect 47259 8928 47768 8956
rect 47259 8925 47271 8928
rect 47213 8919 47271 8925
rect 47762 8916 47768 8928
rect 47820 8916 47826 8968
rect 48056 8956 48084 8987
rect 49786 8956 49792 8968
rect 48056 8928 49792 8956
rect 49786 8916 49792 8928
rect 49844 8916 49850 8968
rect 50264 8956 50292 8996
rect 50709 8993 50721 9027
rect 50755 8993 50767 9027
rect 50890 9024 50896 9036
rect 50851 8996 50896 9024
rect 50709 8987 50767 8993
rect 50890 8984 50896 8996
rect 50948 8984 50954 9036
rect 51077 9027 51135 9033
rect 51077 8993 51089 9027
rect 51123 9024 51135 9027
rect 51350 9024 51356 9036
rect 51123 8996 51356 9024
rect 51123 8993 51135 8996
rect 51077 8987 51135 8993
rect 51350 8984 51356 8996
rect 51408 8984 51414 9036
rect 51442 8984 51448 9036
rect 51500 9024 51506 9036
rect 52181 9027 52239 9033
rect 52181 9024 52193 9027
rect 51500 8996 52193 9024
rect 51500 8984 51506 8996
rect 52181 8993 52193 8996
rect 52227 9024 52239 9027
rect 52730 9024 52736 9036
rect 52227 8996 52736 9024
rect 52227 8993 52239 8996
rect 52181 8987 52239 8993
rect 52730 8984 52736 8996
rect 52788 8984 52794 9036
rect 53469 9027 53527 9033
rect 53469 8993 53481 9027
rect 53515 9024 53527 9027
rect 53558 9024 53564 9036
rect 53515 8996 53564 9024
rect 53515 8993 53527 8996
rect 53469 8987 53527 8993
rect 53558 8984 53564 8996
rect 53616 8984 53622 9036
rect 54665 9027 54723 9033
rect 54665 8993 54677 9027
rect 54711 9024 54723 9027
rect 55214 9024 55220 9036
rect 54711 8996 55220 9024
rect 54711 8993 54723 8996
rect 54665 8987 54723 8993
rect 55214 8984 55220 8996
rect 55272 9024 55278 9036
rect 55398 9024 55404 9036
rect 55272 8996 55404 9024
rect 55272 8984 55278 8996
rect 55398 8984 55404 8996
rect 55456 8984 55462 9036
rect 55968 9024 55996 9064
rect 58713 9027 58771 9033
rect 58713 9024 58725 9027
rect 55968 8996 58725 9024
rect 58713 8993 58725 8996
rect 58759 9024 58771 9027
rect 59262 9024 59268 9036
rect 58759 8996 59268 9024
rect 58759 8993 58771 8996
rect 58713 8987 58771 8993
rect 59262 8984 59268 8996
rect 59320 8984 59326 9036
rect 60645 9027 60703 9033
rect 60645 8993 60657 9027
rect 60691 9024 60703 9027
rect 61013 9027 61071 9033
rect 60691 8996 60964 9024
rect 60691 8993 60703 8996
rect 60645 8987 60703 8993
rect 52089 8959 52147 8965
rect 50264 8928 52040 8956
rect 40037 8891 40095 8897
rect 40037 8857 40049 8891
rect 40083 8888 40095 8891
rect 40310 8888 40316 8900
rect 40083 8860 40316 8888
rect 40083 8857 40095 8860
rect 40037 8851 40095 8857
rect 40310 8848 40316 8860
rect 40368 8848 40374 8900
rect 42334 8848 42340 8900
rect 42392 8888 42398 8900
rect 42981 8891 43039 8897
rect 42981 8888 42993 8891
rect 42392 8860 42993 8888
rect 42392 8848 42398 8860
rect 42981 8857 42993 8860
rect 43027 8888 43039 8891
rect 43070 8888 43076 8900
rect 43027 8860 43076 8888
rect 43027 8857 43039 8860
rect 42981 8851 43039 8857
rect 43070 8848 43076 8860
rect 43128 8848 43134 8900
rect 46106 8848 46112 8900
rect 46164 8888 46170 8900
rect 46661 8891 46719 8897
rect 46661 8888 46673 8891
rect 46164 8860 46673 8888
rect 46164 8848 46170 8860
rect 46661 8857 46673 8860
rect 46707 8857 46719 8891
rect 46661 8851 46719 8857
rect 48777 8891 48835 8897
rect 48777 8857 48789 8891
rect 48823 8888 48835 8891
rect 49970 8888 49976 8900
rect 48823 8860 49976 8888
rect 48823 8857 48835 8860
rect 48777 8851 48835 8857
rect 49970 8848 49976 8860
rect 50028 8848 50034 8900
rect 50525 8891 50583 8897
rect 50525 8857 50537 8891
rect 50571 8888 50583 8891
rect 51810 8888 51816 8900
rect 50571 8860 51816 8888
rect 50571 8857 50583 8860
rect 50525 8851 50583 8857
rect 51810 8848 51816 8860
rect 51868 8848 51874 8900
rect 52012 8888 52040 8928
rect 52089 8925 52101 8959
rect 52135 8956 52147 8959
rect 53282 8956 53288 8968
rect 52135 8928 53288 8956
rect 52135 8925 52147 8928
rect 52089 8919 52147 8925
rect 53282 8916 53288 8928
rect 53340 8916 53346 8968
rect 54294 8916 54300 8968
rect 54352 8956 54358 8968
rect 54573 8959 54631 8965
rect 54573 8956 54585 8959
rect 54352 8928 54585 8956
rect 54352 8916 54358 8928
rect 54573 8925 54585 8928
rect 54619 8925 54631 8959
rect 54573 8919 54631 8925
rect 55122 8916 55128 8968
rect 55180 8956 55186 8968
rect 56134 8956 56140 8968
rect 55180 8928 56140 8956
rect 55180 8916 55186 8928
rect 56134 8916 56140 8928
rect 56192 8916 56198 8968
rect 56410 8956 56416 8968
rect 56371 8928 56416 8956
rect 56410 8916 56416 8928
rect 56468 8916 56474 8968
rect 56502 8916 56508 8968
rect 56560 8956 56566 8968
rect 57054 8956 57060 8968
rect 56560 8928 57060 8956
rect 56560 8916 56566 8928
rect 57054 8916 57060 8928
rect 57112 8956 57118 8968
rect 58618 8956 58624 8968
rect 57112 8928 58624 8956
rect 57112 8916 57118 8928
rect 58618 8916 58624 8928
rect 58676 8916 58682 8968
rect 53561 8891 53619 8897
rect 53561 8888 53573 8891
rect 52012 8860 53573 8888
rect 53561 8857 53573 8860
rect 53607 8857 53619 8891
rect 53561 8851 53619 8857
rect 54754 8848 54760 8900
rect 54812 8888 54818 8900
rect 55401 8891 55459 8897
rect 55401 8888 55413 8891
rect 54812 8860 55413 8888
rect 54812 8848 54818 8860
rect 55401 8857 55413 8860
rect 55447 8857 55459 8891
rect 55401 8851 55459 8857
rect 58161 8891 58219 8897
rect 58161 8857 58173 8891
rect 58207 8888 58219 8891
rect 58250 8888 58256 8900
rect 58207 8860 58256 8888
rect 58207 8857 58219 8860
rect 58161 8851 58219 8857
rect 58250 8848 58256 8860
rect 58308 8888 58314 8900
rect 60458 8888 60464 8900
rect 58308 8860 58940 8888
rect 60419 8860 60464 8888
rect 58308 8848 58314 8860
rect 40586 8820 40592 8832
rect 37844 8792 40592 8820
rect 40586 8780 40592 8792
rect 40644 8820 40650 8832
rect 41046 8820 41052 8832
rect 40644 8792 41052 8820
rect 40644 8780 40650 8792
rect 41046 8780 41052 8792
rect 41104 8780 41110 8832
rect 41230 8820 41236 8832
rect 41191 8792 41236 8820
rect 41230 8780 41236 8792
rect 41288 8780 41294 8832
rect 41966 8780 41972 8832
rect 42024 8820 42030 8832
rect 42613 8823 42671 8829
rect 42613 8820 42625 8823
rect 42024 8792 42625 8820
rect 42024 8780 42030 8792
rect 42613 8789 42625 8792
rect 42659 8789 42671 8823
rect 44266 8820 44272 8832
rect 44227 8792 44272 8820
rect 42613 8783 42671 8789
rect 44266 8780 44272 8792
rect 44324 8780 44330 8832
rect 44634 8820 44640 8832
rect 44595 8792 44640 8820
rect 44634 8780 44640 8792
rect 44692 8780 44698 8832
rect 46290 8820 46296 8832
rect 46251 8792 46296 8820
rect 46290 8780 46296 8792
rect 46348 8780 46354 8832
rect 47026 8820 47032 8832
rect 46987 8792 47032 8820
rect 47026 8780 47032 8792
rect 47084 8780 47090 8832
rect 47394 8780 47400 8832
rect 47452 8820 47458 8832
rect 49329 8823 49387 8829
rect 49329 8820 49341 8823
rect 47452 8792 49341 8820
rect 47452 8780 47458 8792
rect 49329 8789 49341 8792
rect 49375 8789 49387 8823
rect 50062 8820 50068 8832
rect 50023 8792 50068 8820
rect 49329 8783 49387 8789
rect 50062 8780 50068 8792
rect 50120 8780 50126 8832
rect 51534 8820 51540 8832
rect 51495 8792 51540 8820
rect 51534 8780 51540 8792
rect 51592 8780 51598 8832
rect 51718 8780 51724 8832
rect 51776 8820 51782 8832
rect 51997 8823 52055 8829
rect 51997 8820 52009 8823
rect 51776 8792 52009 8820
rect 51776 8780 51782 8792
rect 51997 8789 52009 8792
rect 52043 8820 52055 8823
rect 52270 8820 52276 8832
rect 52043 8792 52276 8820
rect 52043 8789 52055 8792
rect 51997 8783 52055 8789
rect 52270 8780 52276 8792
rect 52328 8780 52334 8832
rect 52822 8780 52828 8832
rect 52880 8820 52886 8832
rect 53009 8823 53067 8829
rect 53009 8820 53021 8823
rect 52880 8792 53021 8820
rect 52880 8780 52886 8792
rect 53009 8789 53021 8792
rect 53055 8789 53067 8823
rect 54846 8820 54852 8832
rect 54807 8792 54852 8820
rect 53009 8783 53067 8789
rect 54846 8780 54852 8792
rect 54904 8780 54910 8832
rect 56045 8823 56103 8829
rect 56045 8789 56057 8823
rect 56091 8820 56103 8823
rect 56318 8820 56324 8832
rect 56091 8792 56324 8820
rect 56091 8789 56103 8792
rect 56045 8783 56103 8789
rect 56318 8780 56324 8792
rect 56376 8780 56382 8832
rect 56502 8780 56508 8832
rect 56560 8820 56566 8832
rect 57517 8823 57575 8829
rect 57517 8820 57529 8823
rect 56560 8792 57529 8820
rect 56560 8780 56566 8792
rect 57517 8789 57529 8792
rect 57563 8789 57575 8823
rect 58434 8820 58440 8832
rect 58395 8792 58440 8820
rect 57517 8783 57575 8789
rect 58434 8780 58440 8792
rect 58492 8780 58498 8832
rect 58912 8829 58940 8860
rect 60458 8848 60464 8860
rect 60516 8848 60522 8900
rect 60936 8888 60964 8996
rect 61013 8993 61025 9027
rect 61059 9024 61071 9027
rect 61838 9024 61844 9036
rect 61059 8996 61844 9024
rect 61059 8993 61071 8996
rect 61013 8987 61071 8993
rect 61838 8984 61844 8996
rect 61896 8984 61902 9036
rect 61102 8956 61108 8968
rect 61063 8928 61108 8956
rect 61102 8916 61108 8928
rect 61160 8916 61166 8968
rect 61378 8916 61384 8968
rect 61436 8956 61442 8968
rect 61473 8959 61531 8965
rect 61473 8956 61485 8959
rect 61436 8928 61485 8956
rect 61436 8916 61442 8928
rect 61473 8925 61485 8928
rect 61519 8925 61531 8959
rect 61473 8919 61531 8925
rect 61396 8888 61424 8916
rect 60936 8860 61424 8888
rect 58897 8823 58955 8829
rect 58897 8789 58909 8823
rect 58943 8789 58955 8823
rect 58897 8783 58955 8789
rect 59078 8780 59084 8832
rect 59136 8820 59142 8832
rect 59449 8823 59507 8829
rect 59449 8820 59461 8823
rect 59136 8792 59461 8820
rect 59136 8780 59142 8792
rect 59449 8789 59461 8792
rect 59495 8789 59507 8823
rect 59814 8820 59820 8832
rect 59775 8792 59820 8820
rect 59449 8783 59507 8789
rect 59814 8780 59820 8792
rect 59872 8780 59878 8832
rect 1104 8730 63480 8752
rect 1104 8678 11378 8730
rect 11430 8678 11442 8730
rect 11494 8678 11506 8730
rect 11558 8678 11570 8730
rect 11622 8678 32170 8730
rect 32222 8678 32234 8730
rect 32286 8678 32298 8730
rect 32350 8678 32362 8730
rect 32414 8678 52962 8730
rect 53014 8678 53026 8730
rect 53078 8678 53090 8730
rect 53142 8678 53154 8730
rect 53206 8678 63480 8730
rect 1104 8656 63480 8678
rect 3050 8616 3056 8628
rect 3011 8588 3056 8616
rect 3050 8576 3056 8588
rect 3108 8576 3114 8628
rect 6362 8616 6368 8628
rect 3436 8588 6368 8616
rect 2866 8508 2872 8560
rect 2924 8548 2930 8560
rect 3329 8551 3387 8557
rect 3329 8548 3341 8551
rect 2924 8520 3341 8548
rect 2924 8508 2930 8520
rect 3329 8517 3341 8520
rect 3375 8517 3387 8551
rect 3329 8511 3387 8517
rect 2590 8440 2596 8492
rect 2648 8480 2654 8492
rect 2685 8483 2743 8489
rect 2685 8480 2697 8483
rect 2648 8452 2697 8480
rect 2648 8440 2654 8452
rect 2685 8449 2697 8452
rect 2731 8480 2743 8483
rect 3436 8480 3464 8588
rect 6362 8576 6368 8588
rect 6420 8576 6426 8628
rect 8665 8619 8723 8625
rect 8665 8585 8677 8619
rect 8711 8616 8723 8619
rect 8754 8616 8760 8628
rect 8711 8588 8760 8616
rect 8711 8585 8723 8588
rect 8665 8579 8723 8585
rect 8754 8576 8760 8588
rect 8812 8616 8818 8628
rect 11146 8616 11152 8628
rect 8812 8588 11152 8616
rect 8812 8576 8818 8588
rect 11146 8576 11152 8588
rect 11204 8576 11210 8628
rect 11882 8616 11888 8628
rect 11843 8588 11888 8616
rect 11882 8576 11888 8588
rect 11940 8576 11946 8628
rect 12253 8619 12311 8625
rect 12253 8585 12265 8619
rect 12299 8616 12311 8619
rect 12342 8616 12348 8628
rect 12299 8588 12348 8616
rect 12299 8585 12311 8588
rect 12253 8579 12311 8585
rect 12342 8576 12348 8588
rect 12400 8576 12406 8628
rect 12526 8576 12532 8628
rect 12584 8616 12590 8628
rect 12621 8619 12679 8625
rect 12621 8616 12633 8619
rect 12584 8588 12633 8616
rect 12584 8576 12590 8588
rect 12621 8585 12633 8588
rect 12667 8585 12679 8619
rect 15102 8616 15108 8628
rect 15063 8588 15108 8616
rect 12621 8579 12679 8585
rect 15102 8576 15108 8588
rect 15160 8576 15166 8628
rect 15930 8576 15936 8628
rect 15988 8616 15994 8628
rect 16025 8619 16083 8625
rect 16025 8616 16037 8619
rect 15988 8588 16037 8616
rect 15988 8576 15994 8588
rect 16025 8585 16037 8588
rect 16071 8585 16083 8619
rect 16025 8579 16083 8585
rect 16853 8619 16911 8625
rect 16853 8585 16865 8619
rect 16899 8616 16911 8619
rect 19978 8616 19984 8628
rect 16899 8588 19984 8616
rect 16899 8585 16911 8588
rect 16853 8579 16911 8585
rect 19978 8576 19984 8588
rect 20036 8576 20042 8628
rect 20165 8619 20223 8625
rect 20165 8585 20177 8619
rect 20211 8616 20223 8619
rect 20254 8616 20260 8628
rect 20211 8588 20260 8616
rect 20211 8585 20223 8588
rect 20165 8579 20223 8585
rect 20254 8576 20260 8588
rect 20312 8576 20318 8628
rect 20898 8576 20904 8628
rect 20956 8616 20962 8628
rect 21177 8619 21235 8625
rect 21177 8616 21189 8619
rect 20956 8588 21189 8616
rect 20956 8576 20962 8588
rect 21177 8585 21189 8588
rect 21223 8616 21235 8619
rect 21634 8616 21640 8628
rect 21223 8588 21640 8616
rect 21223 8585 21235 8588
rect 21177 8579 21235 8585
rect 21634 8576 21640 8588
rect 21692 8576 21698 8628
rect 22370 8576 22376 8628
rect 22428 8616 22434 8628
rect 22833 8619 22891 8625
rect 22833 8616 22845 8619
rect 22428 8588 22845 8616
rect 22428 8576 22434 8588
rect 22833 8585 22845 8588
rect 22879 8585 22891 8619
rect 22833 8579 22891 8585
rect 24029 8619 24087 8625
rect 24029 8585 24041 8619
rect 24075 8616 24087 8619
rect 25406 8616 25412 8628
rect 24075 8588 25412 8616
rect 24075 8585 24087 8588
rect 24029 8579 24087 8585
rect 25406 8576 25412 8588
rect 25464 8616 25470 8628
rect 26510 8616 26516 8628
rect 25464 8588 26516 8616
rect 25464 8576 25470 8588
rect 26510 8576 26516 8588
rect 26568 8576 26574 8628
rect 28442 8616 28448 8628
rect 28403 8588 28448 8616
rect 28442 8576 28448 8588
rect 28500 8576 28506 8628
rect 28534 8576 28540 8628
rect 28592 8616 28598 8628
rect 30837 8619 30895 8625
rect 30837 8616 30849 8619
rect 28592 8588 30849 8616
rect 28592 8576 28598 8588
rect 30837 8585 30849 8588
rect 30883 8585 30895 8619
rect 30837 8579 30895 8585
rect 32490 8576 32496 8628
rect 32548 8616 32554 8628
rect 33045 8619 33103 8625
rect 33045 8616 33057 8619
rect 32548 8588 33057 8616
rect 32548 8576 32554 8588
rect 33045 8585 33057 8588
rect 33091 8585 33103 8619
rect 33045 8579 33103 8585
rect 33321 8619 33379 8625
rect 33321 8585 33333 8619
rect 33367 8616 33379 8619
rect 34609 8619 34667 8625
rect 34609 8616 34621 8619
rect 33367 8588 34621 8616
rect 33367 8585 33379 8588
rect 33321 8579 33379 8585
rect 34609 8585 34621 8588
rect 34655 8616 34667 8619
rect 34790 8616 34796 8628
rect 34655 8588 34796 8616
rect 34655 8585 34667 8588
rect 34609 8579 34667 8585
rect 34790 8576 34796 8588
rect 34848 8616 34854 8628
rect 35894 8616 35900 8628
rect 34848 8588 35900 8616
rect 34848 8576 34854 8588
rect 35894 8576 35900 8588
rect 35952 8576 35958 8628
rect 36446 8576 36452 8628
rect 36504 8616 36510 8628
rect 36633 8619 36691 8625
rect 36633 8616 36645 8619
rect 36504 8588 36645 8616
rect 36504 8576 36510 8588
rect 36633 8585 36645 8588
rect 36679 8585 36691 8619
rect 38746 8616 38752 8628
rect 38707 8588 38752 8616
rect 36633 8579 36691 8585
rect 38746 8576 38752 8588
rect 38804 8576 38810 8628
rect 41414 8616 41420 8628
rect 38948 8588 41420 8616
rect 8021 8551 8079 8557
rect 8021 8517 8033 8551
rect 8067 8548 8079 8551
rect 8573 8551 8631 8557
rect 8573 8548 8585 8551
rect 8067 8520 8585 8548
rect 8067 8517 8079 8520
rect 8021 8511 8079 8517
rect 8573 8517 8585 8520
rect 8619 8548 8631 8551
rect 11054 8548 11060 8560
rect 8619 8520 11060 8548
rect 8619 8517 8631 8520
rect 8573 8511 8631 8517
rect 11054 8508 11060 8520
rect 11112 8508 11118 8560
rect 2731 8452 3464 8480
rect 4157 8483 4215 8489
rect 2731 8449 2743 8452
rect 2685 8443 2743 8449
rect 4157 8449 4169 8483
rect 4203 8480 4215 8483
rect 4203 8452 4568 8480
rect 4203 8449 4215 8452
rect 4157 8443 4215 8449
rect 4062 8372 4068 8424
rect 4120 8412 4126 8424
rect 4540 8421 4568 8452
rect 7282 8440 7288 8492
rect 7340 8480 7346 8492
rect 7837 8483 7895 8489
rect 7837 8480 7849 8483
rect 7340 8452 7849 8480
rect 7340 8440 7346 8452
rect 7837 8449 7849 8452
rect 7883 8449 7895 8483
rect 7837 8443 7895 8449
rect 7929 8483 7987 8489
rect 7929 8449 7941 8483
rect 7975 8480 7987 8483
rect 8205 8483 8263 8489
rect 8205 8480 8217 8483
rect 7975 8452 8217 8480
rect 7975 8449 7987 8452
rect 7929 8443 7987 8449
rect 8205 8449 8217 8452
rect 8251 8480 8263 8483
rect 9401 8483 9459 8489
rect 8251 8452 9076 8480
rect 8251 8449 8263 8452
rect 8205 8443 8263 8449
rect 4249 8415 4307 8421
rect 4249 8412 4261 8415
rect 4120 8384 4261 8412
rect 4120 8372 4126 8384
rect 4249 8381 4261 8384
rect 4295 8381 4307 8415
rect 4249 8375 4307 8381
rect 4525 8415 4583 8421
rect 4525 8381 4537 8415
rect 4571 8412 4583 8415
rect 6825 8415 6883 8421
rect 6825 8412 6837 8415
rect 4571 8384 6837 8412
rect 4571 8381 4583 8384
rect 4525 8375 4583 8381
rect 6825 8381 6837 8384
rect 6871 8381 6883 8415
rect 6825 8375 6883 8381
rect 7377 8415 7435 8421
rect 7377 8381 7389 8415
rect 7423 8381 7435 8415
rect 7377 8375 7435 8381
rect 7653 8415 7711 8421
rect 7653 8381 7665 8415
rect 7699 8412 7711 8415
rect 8021 8415 8079 8421
rect 8021 8412 8033 8415
rect 7699 8384 8033 8412
rect 7699 8381 7711 8384
rect 7653 8375 7711 8381
rect 8021 8381 8033 8384
rect 8067 8381 8079 8415
rect 8941 8415 8999 8421
rect 8941 8412 8953 8415
rect 8021 8375 8079 8381
rect 8772 8384 8953 8412
rect 5442 8304 5448 8356
rect 5500 8344 5506 8356
rect 6638 8344 6644 8356
rect 5500 8316 6132 8344
rect 6599 8316 6644 8344
rect 5500 8304 5506 8316
rect 6104 8288 6132 8316
rect 6638 8304 6644 8316
rect 6696 8304 6702 8356
rect 7392 8344 7420 8375
rect 7929 8347 7987 8353
rect 7929 8344 7941 8347
rect 6748 8316 7941 8344
rect 5810 8276 5816 8288
rect 5771 8248 5816 8276
rect 5810 8236 5816 8248
rect 5868 8236 5874 8288
rect 6086 8236 6092 8288
rect 6144 8276 6150 8288
rect 6273 8279 6331 8285
rect 6273 8276 6285 8279
rect 6144 8248 6285 8276
rect 6144 8236 6150 8248
rect 6273 8245 6285 8248
rect 6319 8276 6331 8279
rect 6748 8276 6776 8316
rect 7929 8313 7941 8316
rect 7975 8313 7987 8347
rect 7929 8307 7987 8313
rect 8202 8304 8208 8356
rect 8260 8344 8266 8356
rect 8772 8344 8800 8384
rect 8941 8381 8953 8384
rect 8987 8381 8999 8415
rect 9048 8412 9076 8452
rect 9401 8449 9413 8483
rect 9447 8480 9459 8483
rect 10870 8480 10876 8492
rect 9447 8452 10876 8480
rect 9447 8449 9459 8452
rect 9401 8443 9459 8449
rect 10870 8440 10876 8452
rect 10928 8440 10934 8492
rect 11900 8480 11928 8576
rect 15657 8551 15715 8557
rect 15657 8517 15669 8551
rect 15703 8548 15715 8551
rect 18046 8548 18052 8560
rect 15703 8520 18052 8548
rect 15703 8517 15715 8520
rect 15657 8511 15715 8517
rect 18046 8508 18052 8520
rect 18104 8508 18110 8560
rect 18322 8508 18328 8560
rect 18380 8557 18386 8560
rect 18380 8551 18429 8557
rect 18380 8517 18383 8551
rect 18417 8517 18429 8551
rect 18380 8511 18429 8517
rect 18380 8508 18386 8511
rect 19334 8508 19340 8560
rect 19392 8548 19398 8560
rect 20346 8548 20352 8560
rect 19392 8520 20352 8548
rect 19392 8508 19398 8520
rect 20346 8508 20352 8520
rect 20404 8548 20410 8560
rect 24121 8551 24179 8557
rect 24121 8548 24133 8551
rect 20404 8520 24133 8548
rect 20404 8508 20410 8520
rect 24121 8517 24133 8520
rect 24167 8517 24179 8551
rect 24121 8511 24179 8517
rect 24946 8508 24952 8560
rect 25004 8548 25010 8560
rect 26694 8548 26700 8560
rect 25004 8520 26700 8548
rect 25004 8508 25010 8520
rect 26694 8508 26700 8520
rect 26752 8548 26758 8560
rect 27338 8548 27344 8560
rect 26752 8520 27344 8548
rect 26752 8508 26758 8520
rect 27338 8508 27344 8520
rect 27396 8508 27402 8560
rect 28902 8508 28908 8560
rect 28960 8548 28966 8560
rect 29917 8551 29975 8557
rect 29917 8548 29929 8551
rect 28960 8520 29929 8548
rect 28960 8508 28966 8520
rect 29917 8517 29929 8520
rect 29963 8517 29975 8551
rect 29917 8511 29975 8517
rect 30006 8508 30012 8560
rect 30064 8548 30070 8560
rect 30193 8551 30251 8557
rect 30193 8548 30205 8551
rect 30064 8520 30205 8548
rect 30064 8508 30070 8520
rect 30193 8517 30205 8520
rect 30239 8548 30251 8551
rect 38838 8548 38844 8560
rect 30239 8520 38844 8548
rect 30239 8517 30251 8520
rect 30193 8511 30251 8517
rect 38838 8508 38844 8520
rect 38896 8508 38902 8560
rect 11164 8452 11928 8480
rect 11164 8421 11192 8452
rect 12066 8440 12072 8492
rect 12124 8480 12130 8492
rect 14737 8483 14795 8489
rect 14737 8480 14749 8483
rect 12124 8452 14749 8480
rect 12124 8440 12130 8452
rect 10597 8415 10655 8421
rect 9048 8384 10272 8412
rect 8941 8375 8999 8381
rect 8260 8316 8800 8344
rect 8260 8304 8266 8316
rect 8846 8304 8852 8356
rect 8904 8344 8910 8356
rect 9677 8347 9735 8353
rect 9677 8344 9689 8347
rect 8904 8316 9689 8344
rect 8904 8304 8910 8316
rect 9677 8313 9689 8316
rect 9723 8313 9735 8347
rect 9677 8307 9735 8313
rect 6319 8248 6776 8276
rect 10244 8276 10272 8384
rect 10597 8381 10609 8415
rect 10643 8381 10655 8415
rect 10597 8375 10655 8381
rect 11149 8415 11207 8421
rect 11149 8381 11161 8415
rect 11195 8381 11207 8415
rect 11149 8375 11207 8381
rect 10321 8347 10379 8353
rect 10321 8313 10333 8347
rect 10367 8344 10379 8347
rect 10612 8344 10640 8375
rect 11238 8372 11244 8424
rect 11296 8412 11302 8424
rect 13998 8412 14004 8424
rect 11296 8384 11341 8412
rect 13959 8384 14004 8412
rect 11296 8372 11302 8384
rect 13998 8372 14004 8384
rect 14056 8372 14062 8424
rect 14292 8421 14320 8452
rect 14737 8449 14749 8452
rect 14783 8449 14795 8483
rect 14737 8443 14795 8449
rect 15010 8440 15016 8492
rect 15068 8480 15074 8492
rect 16114 8480 16120 8492
rect 15068 8452 16120 8480
rect 15068 8440 15074 8452
rect 16114 8440 16120 8452
rect 16172 8440 16178 8492
rect 16577 8483 16635 8489
rect 16577 8449 16589 8483
rect 16623 8480 16635 8483
rect 16623 8452 17448 8480
rect 16623 8449 16635 8452
rect 16577 8443 16635 8449
rect 14277 8415 14335 8421
rect 14277 8381 14289 8415
rect 14323 8381 14335 8415
rect 14277 8375 14335 8381
rect 14461 8415 14519 8421
rect 14461 8381 14473 8415
rect 14507 8412 14519 8415
rect 15102 8412 15108 8424
rect 14507 8384 15108 8412
rect 14507 8381 14519 8384
rect 14461 8375 14519 8381
rect 15102 8372 15108 8384
rect 15160 8372 15166 8424
rect 15194 8372 15200 8424
rect 15252 8412 15258 8424
rect 15473 8415 15531 8421
rect 15473 8412 15485 8415
rect 15252 8384 15485 8412
rect 15252 8372 15258 8384
rect 15473 8381 15485 8384
rect 15519 8412 15531 8415
rect 15746 8412 15752 8424
rect 15519 8384 15752 8412
rect 15519 8381 15531 8384
rect 15473 8375 15531 8381
rect 15746 8372 15752 8384
rect 15804 8372 15810 8424
rect 16669 8415 16727 8421
rect 16669 8381 16681 8415
rect 16715 8412 16727 8415
rect 16758 8412 16764 8424
rect 16715 8384 16764 8412
rect 16715 8381 16727 8384
rect 16669 8375 16727 8381
rect 16758 8372 16764 8384
rect 16816 8412 16822 8424
rect 17218 8412 17224 8424
rect 16816 8384 17224 8412
rect 16816 8372 16822 8384
rect 17218 8372 17224 8384
rect 17276 8372 17282 8424
rect 17420 8356 17448 8452
rect 17494 8440 17500 8492
rect 17552 8480 17558 8492
rect 18601 8483 18659 8489
rect 18601 8480 18613 8483
rect 17552 8452 18613 8480
rect 17552 8440 17558 8452
rect 18601 8449 18613 8452
rect 18647 8480 18659 8483
rect 22002 8480 22008 8492
rect 18647 8452 22008 8480
rect 18647 8449 18659 8452
rect 18601 8443 18659 8449
rect 22002 8440 22008 8452
rect 22060 8440 22066 8492
rect 22094 8440 22100 8492
rect 22152 8480 22158 8492
rect 24305 8483 24363 8489
rect 24305 8480 24317 8483
rect 22152 8452 24317 8480
rect 22152 8440 22158 8452
rect 24305 8449 24317 8452
rect 24351 8480 24363 8483
rect 24581 8483 24639 8489
rect 24581 8480 24593 8483
rect 24351 8452 24593 8480
rect 24351 8449 24363 8452
rect 24305 8443 24363 8449
rect 24581 8449 24593 8452
rect 24627 8480 24639 8483
rect 28534 8480 28540 8492
rect 24627 8452 26372 8480
rect 24627 8449 24639 8452
rect 24581 8443 24639 8449
rect 18049 8415 18107 8421
rect 18049 8381 18061 8415
rect 18095 8412 18107 8415
rect 18463 8415 18521 8421
rect 18463 8412 18475 8415
rect 18095 8384 18475 8412
rect 18095 8381 18107 8384
rect 18049 8375 18107 8381
rect 18463 8381 18475 8384
rect 18509 8412 18521 8415
rect 19245 8415 19303 8421
rect 19245 8412 19257 8415
rect 18509 8384 19257 8412
rect 18509 8381 18521 8384
rect 18463 8375 18521 8381
rect 19245 8381 19257 8384
rect 19291 8381 19303 8415
rect 20346 8412 20352 8424
rect 20307 8384 20352 8412
rect 19245 8375 19303 8381
rect 20346 8372 20352 8384
rect 20404 8372 20410 8424
rect 20714 8412 20720 8424
rect 20675 8384 20720 8412
rect 20714 8372 20720 8384
rect 20772 8412 20778 8424
rect 21361 8415 21419 8421
rect 21361 8412 21373 8415
rect 20772 8384 21373 8412
rect 20772 8372 20778 8384
rect 21361 8381 21373 8384
rect 21407 8412 21419 8415
rect 21453 8415 21511 8421
rect 21453 8412 21465 8415
rect 21407 8384 21465 8412
rect 21407 8381 21419 8384
rect 21361 8375 21419 8381
rect 21453 8381 21465 8384
rect 21499 8381 21511 8415
rect 21453 8375 21511 8381
rect 21542 8372 21548 8424
rect 21600 8412 21606 8424
rect 21637 8415 21695 8421
rect 21637 8412 21649 8415
rect 21600 8384 21649 8412
rect 21600 8372 21606 8384
rect 21637 8381 21649 8384
rect 21683 8381 21695 8415
rect 21637 8375 21695 8381
rect 21726 8372 21732 8424
rect 21784 8412 21790 8424
rect 21784 8384 21829 8412
rect 21784 8372 21790 8384
rect 22186 8372 22192 8424
rect 22244 8412 22250 8424
rect 22244 8384 22289 8412
rect 22244 8372 22250 8384
rect 23474 8372 23480 8424
rect 23532 8412 23538 8424
rect 24489 8415 24547 8421
rect 24489 8412 24501 8415
rect 23532 8384 24501 8412
rect 23532 8372 23538 8384
rect 24489 8381 24501 8384
rect 24535 8412 24547 8415
rect 25222 8412 25228 8424
rect 24535 8384 25228 8412
rect 24535 8381 24547 8384
rect 24489 8375 24547 8381
rect 25222 8372 25228 8384
rect 25280 8372 25286 8424
rect 25685 8415 25743 8421
rect 25685 8381 25697 8415
rect 25731 8412 25743 8415
rect 25866 8412 25872 8424
rect 25731 8384 25872 8412
rect 25731 8381 25743 8384
rect 25685 8375 25743 8381
rect 25866 8372 25872 8384
rect 25924 8372 25930 8424
rect 26053 8415 26111 8421
rect 26053 8381 26065 8415
rect 26099 8412 26111 8415
rect 26234 8412 26240 8424
rect 26099 8384 26240 8412
rect 26099 8381 26111 8384
rect 26053 8375 26111 8381
rect 26234 8372 26240 8384
rect 26292 8372 26298 8424
rect 26344 8421 26372 8452
rect 28276 8452 28540 8480
rect 26329 8415 26387 8421
rect 26329 8381 26341 8415
rect 26375 8381 26387 8415
rect 26329 8375 26387 8381
rect 26510 8372 26516 8424
rect 26568 8412 26574 8424
rect 26605 8415 26663 8421
rect 26605 8412 26617 8415
rect 26568 8384 26617 8412
rect 26568 8372 26574 8384
rect 26605 8381 26617 8384
rect 26651 8381 26663 8415
rect 27154 8412 27160 8424
rect 27067 8384 27160 8412
rect 26605 8375 26663 8381
rect 27154 8372 27160 8384
rect 27212 8412 27218 8424
rect 27338 8412 27344 8424
rect 27212 8384 27344 8412
rect 27212 8372 27218 8384
rect 27338 8372 27344 8384
rect 27396 8372 27402 8424
rect 27614 8412 27620 8424
rect 27575 8384 27620 8412
rect 27614 8372 27620 8384
rect 27672 8372 27678 8424
rect 27890 8412 27896 8424
rect 27851 8384 27896 8412
rect 27890 8372 27896 8384
rect 27948 8412 27954 8424
rect 28276 8412 28304 8452
rect 28534 8440 28540 8452
rect 28592 8480 28598 8492
rect 28813 8483 28871 8489
rect 28813 8480 28825 8483
rect 28592 8452 28825 8480
rect 28592 8440 28598 8452
rect 28813 8449 28825 8452
rect 28859 8449 28871 8483
rect 29270 8480 29276 8492
rect 29183 8452 29276 8480
rect 28813 8443 28871 8449
rect 29270 8440 29276 8452
rect 29328 8480 29334 8492
rect 30558 8480 30564 8492
rect 29328 8452 30564 8480
rect 29328 8440 29334 8452
rect 30558 8440 30564 8452
rect 30616 8440 30622 8492
rect 31757 8483 31815 8489
rect 31757 8449 31769 8483
rect 31803 8480 31815 8483
rect 32401 8483 32459 8489
rect 31803 8452 31984 8480
rect 31803 8449 31815 8452
rect 31757 8443 31815 8449
rect 27948 8384 28304 8412
rect 27948 8372 27954 8384
rect 28718 8372 28724 8424
rect 28776 8412 28782 8424
rect 29362 8412 29368 8424
rect 28776 8384 29368 8412
rect 28776 8372 28782 8384
rect 29362 8372 29368 8384
rect 29420 8372 29426 8424
rect 30650 8412 30656 8424
rect 29472 8384 29960 8412
rect 30563 8384 30656 8412
rect 11514 8344 11520 8356
rect 10367 8316 11520 8344
rect 10367 8313 10379 8316
rect 10321 8307 10379 8313
rect 11514 8304 11520 8316
rect 11572 8304 11578 8356
rect 13446 8344 13452 8356
rect 13407 8316 13452 8344
rect 13446 8304 13452 8316
rect 13504 8304 13510 8356
rect 15930 8304 15936 8356
rect 15988 8344 15994 8356
rect 17402 8344 17408 8356
rect 15988 8316 17264 8344
rect 17363 8316 17408 8344
rect 15988 8304 15994 8316
rect 10505 8279 10563 8285
rect 10505 8276 10517 8279
rect 10244 8248 10517 8276
rect 6319 8245 6331 8248
rect 6273 8239 6331 8245
rect 10505 8245 10517 8248
rect 10551 8245 10563 8279
rect 10505 8239 10563 8245
rect 13170 8236 13176 8288
rect 13228 8276 13234 8288
rect 13265 8279 13323 8285
rect 13265 8276 13277 8279
rect 13228 8248 13277 8276
rect 13228 8236 13234 8248
rect 13265 8245 13277 8248
rect 13311 8276 13323 8279
rect 13722 8276 13728 8288
rect 13311 8248 13728 8276
rect 13311 8245 13323 8248
rect 13265 8239 13323 8245
rect 13722 8236 13728 8248
rect 13780 8236 13786 8288
rect 16485 8279 16543 8285
rect 16485 8245 16497 8279
rect 16531 8276 16543 8279
rect 16574 8276 16580 8288
rect 16531 8248 16580 8276
rect 16531 8245 16543 8248
rect 16485 8239 16543 8245
rect 16574 8236 16580 8248
rect 16632 8236 16638 8288
rect 17236 8276 17264 8316
rect 17402 8304 17408 8316
rect 17460 8304 17466 8356
rect 18233 8347 18291 8353
rect 18233 8313 18245 8347
rect 18279 8313 18291 8347
rect 18233 8307 18291 8313
rect 17773 8279 17831 8285
rect 17773 8276 17785 8279
rect 17236 8248 17785 8276
rect 17773 8245 17785 8248
rect 17819 8276 17831 8279
rect 18138 8276 18144 8288
rect 17819 8248 18144 8276
rect 17819 8245 17831 8248
rect 17773 8239 17831 8245
rect 18138 8236 18144 8248
rect 18196 8236 18202 8288
rect 18248 8276 18276 8307
rect 18874 8304 18880 8356
rect 18932 8344 18938 8356
rect 18969 8347 19027 8353
rect 18969 8344 18981 8347
rect 18932 8316 18981 8344
rect 18932 8304 18938 8316
rect 18969 8313 18981 8316
rect 19015 8313 19027 8347
rect 18969 8307 19027 8313
rect 19702 8304 19708 8356
rect 19760 8344 19766 8356
rect 22002 8344 22008 8356
rect 19760 8316 22008 8344
rect 19760 8304 19766 8316
rect 22002 8304 22008 8316
rect 22060 8304 22066 8356
rect 22278 8304 22284 8356
rect 22336 8344 22342 8356
rect 22557 8347 22615 8353
rect 22557 8344 22569 8347
rect 22336 8316 22569 8344
rect 22336 8304 22342 8316
rect 22557 8313 22569 8316
rect 22603 8344 22615 8347
rect 22738 8344 22744 8356
rect 22603 8316 22744 8344
rect 22603 8313 22615 8316
rect 22557 8307 22615 8313
rect 22738 8304 22744 8316
rect 22796 8304 22802 8356
rect 24121 8347 24179 8353
rect 23216 8316 23520 8344
rect 19613 8279 19671 8285
rect 19613 8276 19625 8279
rect 18248 8248 19625 8276
rect 19613 8245 19625 8248
rect 19659 8276 19671 8279
rect 19794 8276 19800 8288
rect 19659 8248 19800 8276
rect 19659 8245 19671 8248
rect 19613 8239 19671 8245
rect 19794 8236 19800 8248
rect 19852 8236 19858 8288
rect 21361 8279 21419 8285
rect 21361 8245 21373 8279
rect 21407 8276 21419 8279
rect 23216 8276 23244 8316
rect 21407 8248 23244 8276
rect 21407 8245 21419 8248
rect 21361 8239 21419 8245
rect 23290 8236 23296 8288
rect 23348 8276 23354 8288
rect 23385 8279 23443 8285
rect 23385 8276 23397 8279
rect 23348 8248 23397 8276
rect 23348 8236 23354 8248
rect 23385 8245 23397 8248
rect 23431 8245 23443 8279
rect 23492 8276 23520 8316
rect 24121 8313 24133 8347
rect 24167 8344 24179 8347
rect 29472 8344 29500 8384
rect 29825 8347 29883 8353
rect 29825 8344 29837 8347
rect 24167 8316 29500 8344
rect 29564 8316 29837 8344
rect 24167 8313 24179 8316
rect 24121 8307 24179 8313
rect 24946 8276 24952 8288
rect 23492 8248 24952 8276
rect 23385 8239 23443 8245
rect 24946 8236 24952 8248
rect 25004 8236 25010 8288
rect 25038 8236 25044 8288
rect 25096 8276 25102 8288
rect 25096 8248 25141 8276
rect 25096 8236 25102 8248
rect 25314 8236 25320 8288
rect 25372 8276 25378 8288
rect 26970 8276 26976 8288
rect 25372 8248 26976 8276
rect 25372 8236 25378 8248
rect 26970 8236 26976 8248
rect 27028 8236 27034 8288
rect 27522 8276 27528 8288
rect 27483 8248 27528 8276
rect 27522 8236 27528 8248
rect 27580 8236 27586 8288
rect 27706 8236 27712 8288
rect 27764 8276 27770 8288
rect 28166 8276 28172 8288
rect 27764 8248 28172 8276
rect 27764 8236 27770 8248
rect 28166 8236 28172 8248
rect 28224 8276 28230 8288
rect 29564 8276 29592 8316
rect 29825 8313 29837 8316
rect 29871 8313 29883 8347
rect 29932 8344 29960 8384
rect 30650 8372 30656 8384
rect 30708 8412 30714 8424
rect 31294 8412 31300 8424
rect 30708 8384 31300 8412
rect 30708 8372 30714 8384
rect 31294 8372 31300 8384
rect 31352 8372 31358 8424
rect 31846 8412 31852 8424
rect 31807 8384 31852 8412
rect 31846 8372 31852 8384
rect 31904 8372 31910 8424
rect 31956 8421 31984 8452
rect 32401 8449 32413 8483
rect 32447 8480 32459 8483
rect 36078 8480 36084 8492
rect 32447 8452 36084 8480
rect 32447 8449 32459 8452
rect 32401 8443 32459 8449
rect 36078 8440 36084 8452
rect 36136 8480 36142 8492
rect 36722 8480 36728 8492
rect 36136 8452 36728 8480
rect 36136 8440 36142 8452
rect 36722 8440 36728 8452
rect 36780 8440 36786 8492
rect 36814 8440 36820 8492
rect 36872 8480 36878 8492
rect 37093 8483 37151 8489
rect 37093 8480 37105 8483
rect 36872 8452 37105 8480
rect 36872 8440 36878 8452
rect 37093 8449 37105 8452
rect 37139 8480 37151 8483
rect 37645 8483 37703 8489
rect 37139 8452 37320 8480
rect 37139 8449 37151 8452
rect 37093 8443 37151 8449
rect 31941 8415 31999 8421
rect 31941 8381 31953 8415
rect 31987 8412 31999 8415
rect 32030 8412 32036 8424
rect 31987 8384 32036 8412
rect 31987 8381 31999 8384
rect 31941 8375 31999 8381
rect 32030 8372 32036 8384
rect 32088 8372 32094 8424
rect 33229 8415 33287 8421
rect 33229 8412 33241 8415
rect 32324 8384 33241 8412
rect 32324 8356 32352 8384
rect 33229 8381 33241 8384
rect 33275 8381 33287 8415
rect 33229 8375 33287 8381
rect 32306 8344 32312 8356
rect 29932 8316 32312 8344
rect 29825 8307 29883 8313
rect 32306 8304 32312 8316
rect 32364 8304 32370 8356
rect 28224 8248 29592 8276
rect 29917 8279 29975 8285
rect 28224 8236 28230 8248
rect 29917 8245 29929 8279
rect 29963 8276 29975 8279
rect 30561 8279 30619 8285
rect 30561 8276 30573 8279
rect 29963 8248 30573 8276
rect 29963 8245 29975 8248
rect 29917 8239 29975 8245
rect 30561 8245 30573 8248
rect 30607 8276 30619 8279
rect 30650 8276 30656 8288
rect 30607 8248 30656 8276
rect 30607 8245 30619 8248
rect 30561 8239 30619 8245
rect 30650 8236 30656 8248
rect 30708 8236 30714 8288
rect 31294 8276 31300 8288
rect 31255 8248 31300 8276
rect 31294 8236 31300 8248
rect 31352 8236 31358 8288
rect 31846 8236 31852 8288
rect 31904 8276 31910 8288
rect 32769 8279 32827 8285
rect 32769 8276 32781 8279
rect 31904 8248 32781 8276
rect 31904 8236 31910 8248
rect 32769 8245 32781 8248
rect 32815 8276 32827 8279
rect 33042 8276 33048 8288
rect 32815 8248 33048 8276
rect 32815 8245 32827 8248
rect 32769 8239 32827 8245
rect 33042 8236 33048 8248
rect 33100 8236 33106 8288
rect 33244 8276 33272 8375
rect 33686 8372 33692 8424
rect 33744 8412 33750 8424
rect 33781 8415 33839 8421
rect 33781 8412 33793 8415
rect 33744 8384 33793 8412
rect 33744 8372 33750 8384
rect 33781 8381 33793 8384
rect 33827 8412 33839 8415
rect 34241 8415 34299 8421
rect 34241 8412 34253 8415
rect 33827 8384 34253 8412
rect 33827 8381 33839 8384
rect 33781 8375 33839 8381
rect 34241 8381 34253 8384
rect 34287 8412 34299 8415
rect 34517 8415 34575 8421
rect 34517 8412 34529 8415
rect 34287 8384 34529 8412
rect 34287 8381 34299 8384
rect 34241 8375 34299 8381
rect 34517 8381 34529 8384
rect 34563 8381 34575 8415
rect 34517 8375 34575 8381
rect 34885 8415 34943 8421
rect 34885 8381 34897 8415
rect 34931 8412 34943 8415
rect 35066 8412 35072 8424
rect 34931 8384 35072 8412
rect 34931 8381 34943 8384
rect 34885 8375 34943 8381
rect 34900 8344 34928 8375
rect 35066 8372 35072 8384
rect 35124 8372 35130 8424
rect 35158 8372 35164 8424
rect 35216 8412 35222 8424
rect 35253 8415 35311 8421
rect 35253 8412 35265 8415
rect 35216 8384 35265 8412
rect 35216 8372 35222 8384
rect 35253 8381 35265 8384
rect 35299 8381 35311 8415
rect 35434 8412 35440 8424
rect 35395 8384 35440 8412
rect 35253 8375 35311 8381
rect 34440 8316 34928 8344
rect 35268 8344 35296 8375
rect 35434 8372 35440 8384
rect 35492 8372 35498 8424
rect 37182 8412 37188 8424
rect 35728 8384 37044 8412
rect 37143 8384 37188 8412
rect 35728 8344 35756 8384
rect 35897 8347 35955 8353
rect 35897 8344 35909 8347
rect 35268 8316 35756 8344
rect 35820 8316 35909 8344
rect 34440 8276 34468 8316
rect 33244 8248 34468 8276
rect 34517 8279 34575 8285
rect 34517 8245 34529 8279
rect 34563 8276 34575 8279
rect 35526 8276 35532 8288
rect 34563 8248 35532 8276
rect 34563 8245 34575 8248
rect 34517 8239 34575 8245
rect 35526 8236 35532 8248
rect 35584 8276 35590 8288
rect 35820 8276 35848 8316
rect 35897 8313 35909 8316
rect 35943 8313 35955 8347
rect 37016 8344 37044 8384
rect 37182 8372 37188 8384
rect 37240 8372 37246 8424
rect 37292 8412 37320 8452
rect 37645 8449 37657 8483
rect 37691 8480 37703 8483
rect 38654 8480 38660 8492
rect 37691 8452 38660 8480
rect 37691 8449 37703 8452
rect 37645 8443 37703 8449
rect 38654 8440 38660 8452
rect 38712 8440 38718 8492
rect 38948 8480 38976 8588
rect 41414 8576 41420 8588
rect 41472 8576 41478 8628
rect 41874 8576 41880 8628
rect 41932 8616 41938 8628
rect 42245 8619 42303 8625
rect 42245 8616 42257 8619
rect 41932 8588 42257 8616
rect 41932 8576 41938 8588
rect 42245 8585 42257 8588
rect 42291 8585 42303 8619
rect 42245 8579 42303 8585
rect 42705 8619 42763 8625
rect 42705 8585 42717 8619
rect 42751 8616 42763 8619
rect 45554 8616 45560 8628
rect 42751 8588 45560 8616
rect 42751 8585 42763 8588
rect 42705 8579 42763 8585
rect 45554 8576 45560 8588
rect 45612 8576 45618 8628
rect 46290 8576 46296 8628
rect 46348 8616 46354 8628
rect 48961 8619 49019 8625
rect 46348 8588 48636 8616
rect 46348 8576 46354 8588
rect 40129 8551 40187 8557
rect 40129 8517 40141 8551
rect 40175 8548 40187 8551
rect 47302 8548 47308 8560
rect 40175 8520 47308 8548
rect 40175 8517 40187 8520
rect 40129 8511 40187 8517
rect 47302 8508 47308 8520
rect 47360 8548 47366 8560
rect 48498 8548 48504 8560
rect 47360 8520 48504 8548
rect 47360 8508 47366 8520
rect 48498 8508 48504 8520
rect 48556 8508 48562 8560
rect 48608 8548 48636 8588
rect 48961 8585 48973 8619
rect 49007 8616 49019 8619
rect 52730 8616 52736 8628
rect 49007 8588 52132 8616
rect 52691 8588 52736 8616
rect 49007 8585 49019 8588
rect 48961 8579 49019 8585
rect 48608 8520 50200 8548
rect 50172 8492 50200 8520
rect 50246 8508 50252 8560
rect 50304 8548 50310 8560
rect 51353 8551 51411 8557
rect 51353 8548 51365 8551
rect 50304 8520 51365 8548
rect 50304 8508 50310 8520
rect 51353 8517 51365 8520
rect 51399 8517 51411 8551
rect 51997 8551 52055 8557
rect 51997 8548 52009 8551
rect 51353 8511 51411 8517
rect 51460 8520 52009 8548
rect 38856 8452 38976 8480
rect 39025 8483 39083 8489
rect 37829 8415 37887 8421
rect 37829 8412 37841 8415
rect 37292 8384 37841 8412
rect 37829 8381 37841 8384
rect 37875 8412 37887 8415
rect 37921 8415 37979 8421
rect 37921 8412 37933 8415
rect 37875 8384 37933 8412
rect 37875 8381 37887 8384
rect 37829 8375 37887 8381
rect 37921 8381 37933 8384
rect 37967 8381 37979 8415
rect 38856 8412 38884 8452
rect 39025 8449 39037 8483
rect 39071 8480 39083 8483
rect 39577 8483 39635 8489
rect 39071 8452 39344 8480
rect 39071 8449 39083 8452
rect 39025 8443 39083 8449
rect 37921 8375 37979 8381
rect 38212 8384 38884 8412
rect 39117 8415 39175 8421
rect 38212 8344 38240 8384
rect 39117 8381 39129 8415
rect 39163 8381 39175 8415
rect 39316 8412 39344 8452
rect 39577 8449 39589 8483
rect 39623 8480 39635 8483
rect 41230 8480 41236 8492
rect 39623 8452 41236 8480
rect 39623 8449 39635 8452
rect 39577 8443 39635 8449
rect 41230 8440 41236 8452
rect 41288 8440 41294 8492
rect 41966 8480 41972 8492
rect 41927 8452 41972 8480
rect 41966 8440 41972 8452
rect 42024 8480 42030 8492
rect 42705 8483 42763 8489
rect 42705 8480 42717 8483
rect 42024 8452 42717 8480
rect 42024 8440 42030 8452
rect 42705 8449 42717 8452
rect 42751 8449 42763 8483
rect 42705 8443 42763 8449
rect 44266 8440 44272 8492
rect 44324 8480 44330 8492
rect 44361 8483 44419 8489
rect 44361 8480 44373 8483
rect 44324 8452 44373 8480
rect 44324 8440 44330 8452
rect 44361 8449 44373 8452
rect 44407 8480 44419 8483
rect 46290 8480 46296 8492
rect 44407 8452 46296 8480
rect 44407 8449 44419 8452
rect 44361 8443 44419 8449
rect 46290 8440 46296 8452
rect 46348 8440 46354 8492
rect 48685 8483 48743 8489
rect 48685 8449 48697 8483
rect 48731 8449 48743 8483
rect 50062 8480 50068 8492
rect 50023 8452 50068 8480
rect 48685 8443 48743 8449
rect 39853 8415 39911 8421
rect 39853 8412 39865 8415
rect 39316 8384 39865 8412
rect 39117 8375 39175 8381
rect 39853 8381 39865 8384
rect 39899 8412 39911 8415
rect 39942 8412 39948 8424
rect 39899 8384 39948 8412
rect 39899 8381 39911 8384
rect 39853 8375 39911 8381
rect 38378 8344 38384 8356
rect 37016 8316 38240 8344
rect 38339 8316 38384 8344
rect 35897 8307 35955 8313
rect 38378 8304 38384 8316
rect 38436 8344 38442 8356
rect 39132 8344 39160 8375
rect 39942 8372 39948 8384
rect 40000 8372 40006 8424
rect 40310 8412 40316 8424
rect 40271 8384 40316 8412
rect 40310 8372 40316 8384
rect 40368 8372 40374 8424
rect 40494 8412 40500 8424
rect 40455 8384 40500 8412
rect 40494 8372 40500 8384
rect 40552 8372 40558 8424
rect 40586 8372 40592 8424
rect 40644 8412 40650 8424
rect 41049 8415 41107 8421
rect 40644 8384 40689 8412
rect 40644 8372 40650 8384
rect 41049 8381 41061 8415
rect 41095 8412 41107 8415
rect 41506 8412 41512 8424
rect 41095 8384 41512 8412
rect 41095 8381 41107 8384
rect 41049 8375 41107 8381
rect 41506 8372 41512 8384
rect 41564 8372 41570 8424
rect 42061 8415 42119 8421
rect 42061 8412 42073 8415
rect 41800 8384 42073 8412
rect 40129 8347 40187 8353
rect 40129 8344 40141 8347
rect 38436 8316 40141 8344
rect 38436 8304 38442 8316
rect 40129 8313 40141 8316
rect 40175 8313 40187 8347
rect 40512 8344 40540 8372
rect 41325 8347 41383 8353
rect 41325 8344 41337 8347
rect 40512 8316 41337 8344
rect 40129 8307 40187 8313
rect 41325 8313 41337 8316
rect 41371 8313 41383 8347
rect 41325 8307 41383 8313
rect 36262 8276 36268 8288
rect 35584 8248 35848 8276
rect 36223 8248 36268 8276
rect 35584 8236 35590 8248
rect 36262 8236 36268 8248
rect 36320 8236 36326 8288
rect 37829 8279 37887 8285
rect 37829 8245 37841 8279
rect 37875 8276 37887 8279
rect 41598 8276 41604 8288
rect 37875 8248 41604 8276
rect 37875 8245 37887 8248
rect 37829 8239 37887 8245
rect 41598 8236 41604 8248
rect 41656 8236 41662 8288
rect 41690 8236 41696 8288
rect 41748 8276 41754 8288
rect 41800 8285 41828 8384
rect 42061 8381 42073 8384
rect 42107 8412 42119 8415
rect 42797 8415 42855 8421
rect 42797 8412 42809 8415
rect 42107 8384 42809 8412
rect 42107 8381 42119 8384
rect 42061 8375 42119 8381
rect 42797 8381 42809 8384
rect 42843 8381 42855 8415
rect 42797 8375 42855 8381
rect 43254 8372 43260 8424
rect 43312 8412 43318 8424
rect 43349 8415 43407 8421
rect 43349 8412 43361 8415
rect 43312 8384 43361 8412
rect 43312 8372 43318 8384
rect 43349 8381 43361 8384
rect 43395 8381 43407 8415
rect 43349 8375 43407 8381
rect 44450 8372 44456 8424
rect 44508 8421 44514 8424
rect 44508 8415 44557 8421
rect 44508 8381 44511 8415
rect 44545 8381 44557 8415
rect 44634 8412 44640 8424
rect 44595 8384 44640 8412
rect 44508 8375 44557 8381
rect 44508 8372 44514 8375
rect 44634 8372 44640 8384
rect 44692 8372 44698 8424
rect 45925 8415 45983 8421
rect 45925 8381 45937 8415
rect 45971 8412 45983 8415
rect 46201 8415 46259 8421
rect 46201 8412 46213 8415
rect 45971 8384 46213 8412
rect 45971 8381 45983 8384
rect 45925 8375 45983 8381
rect 46201 8381 46213 8384
rect 46247 8412 46259 8415
rect 46842 8412 46848 8424
rect 46247 8384 46848 8412
rect 46247 8381 46259 8384
rect 46201 8375 46259 8381
rect 46842 8372 46848 8384
rect 46900 8372 46906 8424
rect 47029 8415 47087 8421
rect 47029 8412 47041 8415
rect 46952 8384 47041 8412
rect 43809 8347 43867 8353
rect 43809 8313 43821 8347
rect 43855 8344 43867 8347
rect 44726 8344 44732 8356
rect 43855 8316 44732 8344
rect 43855 8313 43867 8316
rect 43809 8307 43867 8313
rect 44726 8304 44732 8316
rect 44784 8304 44790 8356
rect 45462 8344 45468 8356
rect 44836 8316 45232 8344
rect 45423 8316 45468 8344
rect 41785 8279 41843 8285
rect 41785 8276 41797 8279
rect 41748 8248 41797 8276
rect 41748 8236 41754 8248
rect 41785 8245 41797 8248
rect 41831 8245 41843 8279
rect 41785 8239 41843 8245
rect 41874 8236 41880 8288
rect 41932 8276 41938 8288
rect 44836 8276 44864 8316
rect 45094 8276 45100 8288
rect 41932 8248 44864 8276
rect 45055 8248 45100 8276
rect 41932 8236 41938 8248
rect 45094 8236 45100 8248
rect 45152 8236 45158 8288
rect 45204 8276 45232 8316
rect 45462 8304 45468 8316
rect 45520 8304 45526 8356
rect 45738 8304 45744 8356
rect 45796 8344 45802 8356
rect 46293 8347 46351 8353
rect 46293 8344 46305 8347
rect 45796 8316 46305 8344
rect 45796 8304 45802 8316
rect 46293 8313 46305 8316
rect 46339 8313 46351 8347
rect 46952 8344 46980 8384
rect 47029 8381 47041 8384
rect 47075 8381 47087 8415
rect 47029 8375 47087 8381
rect 47167 8415 47225 8421
rect 47167 8381 47179 8415
rect 47213 8412 47225 8415
rect 47302 8412 47308 8424
rect 47213 8384 47308 8412
rect 47213 8381 47225 8384
rect 47167 8375 47225 8381
rect 47302 8372 47308 8384
rect 47360 8372 47366 8424
rect 47486 8412 47492 8424
rect 47447 8384 47492 8412
rect 47486 8372 47492 8384
rect 47544 8372 47550 8424
rect 47762 8372 47768 8424
rect 47820 8412 47826 8424
rect 47857 8415 47915 8421
rect 47857 8412 47869 8415
rect 47820 8384 47869 8412
rect 47820 8372 47826 8384
rect 47857 8381 47869 8384
rect 47903 8381 47915 8415
rect 47857 8375 47915 8381
rect 48498 8372 48504 8424
rect 48556 8412 48562 8424
rect 48700 8412 48728 8443
rect 50062 8440 50068 8452
rect 50120 8440 50126 8492
rect 50154 8440 50160 8492
rect 50212 8480 50218 8492
rect 50614 8480 50620 8492
rect 50212 8452 50620 8480
rect 50212 8440 50218 8452
rect 50614 8440 50620 8452
rect 50672 8440 50678 8492
rect 50890 8440 50896 8492
rect 50948 8480 50954 8492
rect 51077 8483 51135 8489
rect 51077 8480 51089 8483
rect 50948 8452 51089 8480
rect 50948 8440 50954 8452
rect 51077 8449 51089 8452
rect 51123 8449 51135 8483
rect 51077 8443 51135 8449
rect 51258 8440 51264 8492
rect 51316 8480 51322 8492
rect 51460 8489 51488 8520
rect 51997 8517 52009 8520
rect 52043 8517 52055 8551
rect 52104 8548 52132 8588
rect 52730 8576 52736 8588
rect 52788 8576 52794 8628
rect 53558 8616 53564 8628
rect 53471 8588 53564 8616
rect 53558 8576 53564 8588
rect 53616 8616 53622 8628
rect 55309 8619 55367 8625
rect 55309 8616 55321 8619
rect 53616 8588 55321 8616
rect 53616 8576 53622 8588
rect 55309 8585 55321 8588
rect 55355 8616 55367 8619
rect 55858 8616 55864 8628
rect 55355 8588 55864 8616
rect 55355 8585 55367 8588
rect 55309 8579 55367 8585
rect 55858 8576 55864 8588
rect 55916 8576 55922 8628
rect 56134 8576 56140 8628
rect 56192 8616 56198 8628
rect 56594 8616 56600 8628
rect 56192 8588 56600 8616
rect 56192 8576 56198 8588
rect 56594 8576 56600 8588
rect 56652 8616 56658 8628
rect 57149 8619 57207 8625
rect 57149 8616 57161 8619
rect 56652 8588 57161 8616
rect 56652 8576 56658 8588
rect 57149 8585 57161 8588
rect 57195 8616 57207 8619
rect 57698 8616 57704 8628
rect 57195 8588 57704 8616
rect 57195 8585 57207 8588
rect 57149 8579 57207 8585
rect 57698 8576 57704 8588
rect 57756 8576 57762 8628
rect 58618 8616 58624 8628
rect 58579 8588 58624 8616
rect 58618 8576 58624 8588
rect 58676 8616 58682 8628
rect 61473 8619 61531 8625
rect 61473 8616 61485 8619
rect 58676 8588 61485 8616
rect 58676 8576 58682 8588
rect 61473 8585 61485 8588
rect 61519 8585 61531 8619
rect 61838 8616 61844 8628
rect 61799 8588 61844 8616
rect 61473 8579 61531 8585
rect 61838 8576 61844 8588
rect 61896 8576 61902 8628
rect 52822 8548 52828 8560
rect 52104 8520 52828 8548
rect 51997 8511 52055 8517
rect 52822 8508 52828 8520
rect 52880 8508 52886 8560
rect 52917 8551 52975 8557
rect 52917 8517 52929 8551
rect 52963 8548 52975 8551
rect 53193 8551 53251 8557
rect 53193 8548 53205 8551
rect 52963 8520 53205 8548
rect 52963 8517 52975 8520
rect 52917 8511 52975 8517
rect 53193 8517 53205 8520
rect 53239 8548 53251 8551
rect 61102 8548 61108 8560
rect 53239 8520 57560 8548
rect 61063 8520 61108 8548
rect 53239 8517 53251 8520
rect 53193 8511 53251 8517
rect 51445 8483 51503 8489
rect 51445 8480 51457 8483
rect 51316 8452 51457 8480
rect 51316 8440 51322 8452
rect 51445 8449 51457 8452
rect 51491 8449 51503 8483
rect 51445 8443 51503 8449
rect 52089 8483 52147 8489
rect 52089 8449 52101 8483
rect 52135 8480 52147 8483
rect 52178 8480 52184 8492
rect 52135 8452 52184 8480
rect 52135 8449 52147 8452
rect 52089 8443 52147 8449
rect 52178 8440 52184 8452
rect 52236 8440 52242 8492
rect 52270 8440 52276 8492
rect 52328 8480 52334 8492
rect 56502 8480 56508 8492
rect 52328 8452 55812 8480
rect 52328 8440 52334 8452
rect 48866 8421 48872 8424
rect 48556 8384 48728 8412
rect 48818 8415 48872 8421
rect 48556 8372 48562 8384
rect 48818 8381 48830 8415
rect 48864 8381 48872 8415
rect 48818 8375 48872 8381
rect 48866 8372 48872 8375
rect 48924 8372 48930 8424
rect 49973 8415 50031 8421
rect 49973 8381 49985 8415
rect 50019 8412 50031 8415
rect 51166 8412 51172 8424
rect 50019 8384 51172 8412
rect 50019 8381 50031 8384
rect 49973 8375 50031 8381
rect 51166 8372 51172 8384
rect 51224 8372 51230 8424
rect 51353 8415 51411 8421
rect 51353 8381 51365 8415
rect 51399 8412 51411 8415
rect 51868 8415 51926 8421
rect 51868 8412 51880 8415
rect 51399 8384 51880 8412
rect 51399 8381 51411 8384
rect 51353 8375 51411 8381
rect 51868 8381 51880 8384
rect 51914 8412 51926 8415
rect 52917 8415 52975 8421
rect 52917 8412 52929 8415
rect 51914 8384 52929 8412
rect 51914 8381 51926 8384
rect 51868 8375 51926 8381
rect 52917 8381 52929 8384
rect 52963 8381 52975 8415
rect 54202 8412 54208 8424
rect 54163 8384 54208 8412
rect 52917 8375 52975 8381
rect 54202 8372 54208 8384
rect 54260 8372 54266 8424
rect 54941 8415 54999 8421
rect 54941 8381 54953 8415
rect 54987 8412 54999 8415
rect 55214 8412 55220 8424
rect 54987 8384 55220 8412
rect 54987 8381 54999 8384
rect 54941 8375 54999 8381
rect 55214 8372 55220 8384
rect 55272 8372 55278 8424
rect 47504 8344 47532 8372
rect 46952 8316 47532 8344
rect 46293 8307 46351 8313
rect 48038 8304 48044 8356
rect 48096 8344 48102 8356
rect 49234 8344 49240 8356
rect 48096 8316 49240 8344
rect 48096 8304 48102 8316
rect 49234 8304 49240 8316
rect 49292 8304 49298 8356
rect 50246 8344 50252 8356
rect 49344 8316 49648 8344
rect 50207 8316 50252 8344
rect 49344 8276 49372 8316
rect 49510 8276 49516 8288
rect 45204 8248 49372 8276
rect 49471 8248 49516 8276
rect 49510 8236 49516 8248
rect 49568 8236 49574 8288
rect 49620 8276 49648 8316
rect 50246 8304 50252 8316
rect 50304 8304 50310 8356
rect 50433 8347 50491 8353
rect 50433 8313 50445 8347
rect 50479 8344 50491 8347
rect 50614 8344 50620 8356
rect 50479 8316 50620 8344
rect 50479 8313 50491 8316
rect 50433 8307 50491 8313
rect 50614 8304 50620 8316
rect 50672 8304 50678 8356
rect 50798 8344 50804 8356
rect 50759 8316 50804 8344
rect 50798 8304 50804 8316
rect 50856 8304 50862 8356
rect 51074 8304 51080 8356
rect 51132 8344 51138 8356
rect 51626 8344 51632 8356
rect 51132 8316 51632 8344
rect 51132 8304 51138 8316
rect 51626 8304 51632 8316
rect 51684 8344 51690 8356
rect 51721 8347 51779 8353
rect 51721 8344 51733 8347
rect 51684 8316 51733 8344
rect 51684 8304 51690 8316
rect 51721 8313 51733 8316
rect 51767 8313 51779 8347
rect 52454 8344 52460 8356
rect 52415 8316 52460 8344
rect 51721 8307 51779 8313
rect 52454 8304 52460 8316
rect 52512 8304 52518 8356
rect 53834 8344 53840 8356
rect 53795 8316 53840 8344
rect 53834 8304 53840 8316
rect 53892 8344 53898 8356
rect 54021 8347 54079 8353
rect 54021 8344 54033 8347
rect 53892 8316 54033 8344
rect 53892 8304 53898 8316
rect 54021 8313 54033 8316
rect 54067 8313 54079 8347
rect 54021 8307 54079 8313
rect 54573 8347 54631 8353
rect 54573 8313 54585 8347
rect 54619 8344 54631 8347
rect 55306 8344 55312 8356
rect 54619 8316 55312 8344
rect 54619 8313 54631 8316
rect 54573 8307 54631 8313
rect 55306 8304 55312 8316
rect 55364 8304 55370 8356
rect 55398 8304 55404 8356
rect 55456 8344 55462 8356
rect 55456 8316 55501 8344
rect 55456 8304 55462 8316
rect 55784 8288 55812 8452
rect 55968 8452 56508 8480
rect 55858 8372 55864 8424
rect 55916 8412 55922 8424
rect 55968 8412 55996 8452
rect 56502 8440 56508 8452
rect 56560 8440 56566 8492
rect 57532 8480 57560 8520
rect 61102 8508 61108 8520
rect 61160 8508 61166 8560
rect 61286 8508 61292 8560
rect 61344 8548 61350 8560
rect 62209 8551 62267 8557
rect 62209 8548 62221 8551
rect 61344 8520 62221 8548
rect 61344 8508 61350 8520
rect 62209 8517 62221 8520
rect 62255 8517 62267 8551
rect 62209 8511 62267 8517
rect 59814 8480 59820 8492
rect 57532 8452 59820 8480
rect 55916 8384 56009 8412
rect 55916 8372 55922 8384
rect 56134 8372 56140 8424
rect 56192 8421 56198 8424
rect 56192 8415 56241 8421
rect 56192 8381 56195 8415
rect 56229 8381 56241 8415
rect 56318 8412 56324 8424
rect 56279 8384 56324 8412
rect 56192 8375 56241 8381
rect 56192 8372 56198 8375
rect 56318 8372 56324 8384
rect 56376 8372 56382 8424
rect 57532 8421 57560 8452
rect 59814 8440 59820 8452
rect 59872 8440 59878 8492
rect 57517 8415 57575 8421
rect 57517 8381 57529 8415
rect 57563 8381 57575 8415
rect 57517 8375 57575 8381
rect 58342 8372 58348 8424
rect 58400 8412 58406 8424
rect 58526 8412 58532 8424
rect 58400 8384 58532 8412
rect 58400 8372 58406 8384
rect 58526 8372 58532 8384
rect 58584 8412 58590 8424
rect 58805 8415 58863 8421
rect 58805 8412 58817 8415
rect 58584 8384 58817 8412
rect 58584 8372 58590 8384
rect 58805 8381 58817 8384
rect 58851 8381 58863 8415
rect 59078 8412 59084 8424
rect 59039 8384 59084 8412
rect 58805 8375 58863 8381
rect 59078 8372 59084 8384
rect 59136 8372 59142 8424
rect 60461 8415 60519 8421
rect 60461 8381 60473 8415
rect 60507 8412 60519 8415
rect 60642 8412 60648 8424
rect 60507 8384 60648 8412
rect 60507 8381 60519 8384
rect 60461 8375 60519 8381
rect 60642 8372 60648 8384
rect 60700 8412 60706 8424
rect 61289 8415 61347 8421
rect 61289 8412 61301 8415
rect 60700 8384 61301 8412
rect 60700 8372 60706 8384
rect 61289 8381 61301 8384
rect 61335 8381 61347 8415
rect 61289 8375 61347 8381
rect 55950 8304 55956 8356
rect 56008 8344 56014 8356
rect 56410 8344 56416 8356
rect 56008 8316 56416 8344
rect 56008 8304 56014 8316
rect 56410 8304 56416 8316
rect 56468 8344 56474 8356
rect 56689 8347 56747 8353
rect 56689 8344 56701 8347
rect 56468 8316 56701 8344
rect 56468 8304 56474 8316
rect 56689 8313 56701 8316
rect 56735 8313 56747 8347
rect 57333 8347 57391 8353
rect 57333 8344 57345 8347
rect 56689 8307 56747 8313
rect 56796 8316 57345 8344
rect 49878 8276 49884 8288
rect 49620 8248 49884 8276
rect 49878 8236 49884 8248
rect 49936 8236 49942 8288
rect 50341 8279 50399 8285
rect 50341 8245 50353 8279
rect 50387 8276 50399 8279
rect 50706 8276 50712 8288
rect 50387 8248 50712 8276
rect 50387 8245 50399 8248
rect 50341 8239 50399 8245
rect 50706 8236 50712 8248
rect 50764 8236 50770 8288
rect 51994 8236 52000 8288
rect 52052 8276 52058 8288
rect 52178 8276 52184 8288
rect 52052 8248 52184 8276
rect 52052 8236 52058 8248
rect 52178 8236 52184 8248
rect 52236 8236 52242 8288
rect 55766 8236 55772 8288
rect 55824 8276 55830 8288
rect 56796 8276 56824 8316
rect 57333 8313 57345 8316
rect 57379 8344 57391 8347
rect 58161 8347 58219 8353
rect 58161 8344 58173 8347
rect 57379 8316 58173 8344
rect 57379 8313 57391 8316
rect 57333 8307 57391 8313
rect 58161 8313 58173 8316
rect 58207 8313 58219 8347
rect 58161 8307 58219 8313
rect 58544 8316 58756 8344
rect 57606 8276 57612 8288
rect 55824 8248 56824 8276
rect 57567 8248 57612 8276
rect 55824 8236 55830 8248
rect 57606 8236 57612 8248
rect 57664 8236 57670 8288
rect 57698 8236 57704 8288
rect 57756 8276 57762 8288
rect 58544 8276 58572 8316
rect 57756 8248 58572 8276
rect 58728 8276 58756 8316
rect 60918 8276 60924 8288
rect 58728 8248 60924 8276
rect 57756 8236 57762 8248
rect 60918 8236 60924 8248
rect 60976 8236 60982 8288
rect 1104 8186 63480 8208
rect 1104 8134 21774 8186
rect 21826 8134 21838 8186
rect 21890 8134 21902 8186
rect 21954 8134 21966 8186
rect 22018 8134 42566 8186
rect 42618 8134 42630 8186
rect 42682 8134 42694 8186
rect 42746 8134 42758 8186
rect 42810 8134 63480 8186
rect 1104 8112 63480 8134
rect 5810 8032 5816 8084
rect 5868 8072 5874 8084
rect 6365 8075 6423 8081
rect 6365 8072 6377 8075
rect 5868 8044 6377 8072
rect 5868 8032 5874 8044
rect 6365 8041 6377 8044
rect 6411 8041 6423 8075
rect 6365 8035 6423 8041
rect 6825 8075 6883 8081
rect 6825 8041 6837 8075
rect 6871 8072 6883 8075
rect 8202 8072 8208 8084
rect 6871 8044 8208 8072
rect 6871 8041 6883 8044
rect 6825 8035 6883 8041
rect 6086 8004 6092 8016
rect 6047 7976 6092 8004
rect 6086 7964 6092 7976
rect 6144 7964 6150 8016
rect 4338 7936 4344 7948
rect 4299 7908 4344 7936
rect 4338 7896 4344 7908
rect 4396 7896 4402 7948
rect 6380 7936 6408 8035
rect 8202 8032 8208 8044
rect 8260 8032 8266 8084
rect 11514 8072 11520 8084
rect 11475 8044 11520 8072
rect 11514 8032 11520 8044
rect 11572 8032 11578 8084
rect 17218 8072 17224 8084
rect 12176 8044 17224 8072
rect 8757 8007 8815 8013
rect 8757 8004 8769 8007
rect 7300 7976 8769 8004
rect 7300 7948 7328 7976
rect 8757 7973 8769 7976
rect 8803 7973 8815 8007
rect 8757 7967 8815 7973
rect 7193 7939 7251 7945
rect 7193 7936 7205 7939
rect 6380 7908 7205 7936
rect 7193 7905 7205 7908
rect 7239 7936 7251 7939
rect 7282 7936 7288 7948
rect 7239 7908 7288 7936
rect 7239 7905 7251 7908
rect 7193 7899 7251 7905
rect 7282 7896 7288 7908
rect 7340 7896 7346 7948
rect 7558 7936 7564 7948
rect 7519 7908 7564 7936
rect 7558 7896 7564 7908
rect 7616 7896 7622 7948
rect 7745 7939 7803 7945
rect 7745 7905 7757 7939
rect 7791 7936 7803 7939
rect 9125 7939 9183 7945
rect 9125 7936 9137 7939
rect 7791 7908 9137 7936
rect 7791 7905 7803 7908
rect 7745 7899 7803 7905
rect 9125 7905 9137 7908
rect 9171 7905 9183 7939
rect 9950 7936 9956 7948
rect 9911 7908 9956 7936
rect 9125 7899 9183 7905
rect 4062 7868 4068 7880
rect 4023 7840 4068 7868
rect 4062 7828 4068 7840
rect 4120 7828 4126 7880
rect 6822 7828 6828 7880
rect 6880 7868 6886 7880
rect 7009 7871 7067 7877
rect 7009 7868 7021 7871
rect 6880 7840 7021 7868
rect 6880 7828 6886 7840
rect 7009 7837 7021 7840
rect 7055 7837 7067 7871
rect 7009 7831 7067 7837
rect 6546 7760 6552 7812
rect 6604 7800 6610 7812
rect 7760 7800 7788 7899
rect 9950 7896 9956 7908
rect 10008 7896 10014 7948
rect 10413 7939 10471 7945
rect 10413 7905 10425 7939
rect 10459 7936 10471 7939
rect 10505 7939 10563 7945
rect 10505 7936 10517 7939
rect 10459 7908 10517 7936
rect 10459 7905 10471 7908
rect 10413 7899 10471 7905
rect 10505 7905 10517 7908
rect 10551 7905 10563 7939
rect 11238 7936 11244 7948
rect 11199 7908 11244 7936
rect 10505 7899 10563 7905
rect 11238 7896 11244 7908
rect 11296 7896 11302 7948
rect 11425 7939 11483 7945
rect 11425 7905 11437 7939
rect 11471 7936 11483 7939
rect 11882 7936 11888 7948
rect 11471 7908 11888 7936
rect 11471 7905 11483 7908
rect 11425 7899 11483 7905
rect 11882 7896 11888 7908
rect 11940 7896 11946 7948
rect 8018 7828 8024 7880
rect 8076 7868 8082 7880
rect 8389 7871 8447 7877
rect 8389 7868 8401 7871
rect 8076 7840 8401 7868
rect 8076 7828 8082 7840
rect 8389 7837 8401 7840
rect 8435 7837 8447 7871
rect 8389 7831 8447 7837
rect 10045 7871 10103 7877
rect 10045 7837 10057 7871
rect 10091 7868 10103 7871
rect 10594 7868 10600 7880
rect 10091 7840 10600 7868
rect 10091 7837 10103 7840
rect 10045 7831 10103 7837
rect 10594 7828 10600 7840
rect 10652 7868 10658 7880
rect 11057 7871 11115 7877
rect 11057 7868 11069 7871
rect 10652 7840 11069 7868
rect 10652 7828 10658 7840
rect 11057 7837 11069 7840
rect 11103 7837 11115 7871
rect 11256 7868 11284 7896
rect 12066 7868 12072 7880
rect 11256 7840 12072 7868
rect 11057 7831 11115 7837
rect 12066 7828 12072 7840
rect 12124 7828 12130 7880
rect 6604 7772 7788 7800
rect 6604 7760 6610 7772
rect 8202 7760 8208 7812
rect 8260 7800 8266 7812
rect 12176 7800 12204 8044
rect 17218 8032 17224 8044
rect 17276 8032 17282 8084
rect 17310 8032 17316 8084
rect 17368 8072 17374 8084
rect 17954 8072 17960 8084
rect 17368 8044 17960 8072
rect 17368 8032 17374 8044
rect 17954 8032 17960 8044
rect 18012 8032 18018 8084
rect 18322 8032 18328 8084
rect 18380 8072 18386 8084
rect 18969 8075 19027 8081
rect 18969 8072 18981 8075
rect 18380 8044 18981 8072
rect 18380 8032 18386 8044
rect 18969 8041 18981 8044
rect 19015 8041 19027 8075
rect 18969 8035 19027 8041
rect 12526 7964 12532 8016
rect 12584 8004 12590 8016
rect 14093 8007 14151 8013
rect 14093 8004 14105 8007
rect 12584 7976 14105 8004
rect 12584 7964 12590 7976
rect 14093 7973 14105 7976
rect 14139 8004 14151 8007
rect 17494 8004 17500 8016
rect 14139 7976 17500 8004
rect 14139 7973 14151 7976
rect 14093 7967 14151 7973
rect 12897 7939 12955 7945
rect 12897 7905 12909 7939
rect 12943 7936 12955 7939
rect 13170 7936 13176 7948
rect 12943 7908 13176 7936
rect 12943 7905 12955 7908
rect 12897 7899 12955 7905
rect 13170 7896 13176 7908
rect 13228 7896 13234 7948
rect 14182 7896 14188 7948
rect 14240 7936 14246 7948
rect 15010 7936 15016 7948
rect 14240 7908 15016 7936
rect 14240 7896 14246 7908
rect 15010 7896 15016 7908
rect 15068 7896 15074 7948
rect 15856 7945 15884 7976
rect 17494 7964 17500 7976
rect 17552 7964 17558 8016
rect 18984 8004 19012 8035
rect 19518 8032 19524 8084
rect 19576 8072 19582 8084
rect 20717 8075 20775 8081
rect 20717 8072 20729 8075
rect 19576 8044 20729 8072
rect 19576 8032 19582 8044
rect 20717 8041 20729 8044
rect 20763 8072 20775 8075
rect 21082 8072 21088 8084
rect 20763 8044 21088 8072
rect 20763 8041 20775 8044
rect 20717 8035 20775 8041
rect 21082 8032 21088 8044
rect 21140 8072 21146 8084
rect 24765 8075 24823 8081
rect 21140 8044 24532 8072
rect 21140 8032 21146 8044
rect 24504 8016 24532 8044
rect 24765 8041 24777 8075
rect 24811 8072 24823 8075
rect 29638 8072 29644 8084
rect 24811 8044 29644 8072
rect 24811 8041 24823 8044
rect 24765 8035 24823 8041
rect 29638 8032 29644 8044
rect 29696 8072 29702 8084
rect 30009 8075 30067 8081
rect 30009 8072 30021 8075
rect 29696 8044 30021 8072
rect 29696 8032 29702 8044
rect 30009 8041 30021 8044
rect 30055 8041 30067 8075
rect 30009 8035 30067 8041
rect 30742 8032 30748 8084
rect 30800 8072 30806 8084
rect 31849 8075 31907 8081
rect 31849 8072 31861 8075
rect 30800 8044 31861 8072
rect 30800 8032 30806 8044
rect 31849 8041 31861 8044
rect 31895 8041 31907 8075
rect 31849 8035 31907 8041
rect 32306 8032 32312 8084
rect 32364 8072 32370 8084
rect 32585 8075 32643 8081
rect 32585 8072 32597 8075
rect 32364 8044 32597 8072
rect 32364 8032 32370 8044
rect 32585 8041 32597 8044
rect 32631 8072 32643 8075
rect 33413 8075 33471 8081
rect 33413 8072 33425 8075
rect 32631 8044 33425 8072
rect 32631 8041 32643 8044
rect 32585 8035 32643 8041
rect 33413 8041 33425 8044
rect 33459 8041 33471 8075
rect 34606 8072 34612 8084
rect 34567 8044 34612 8072
rect 33413 8035 33471 8041
rect 34606 8032 34612 8044
rect 34664 8032 34670 8084
rect 35250 8072 35256 8084
rect 35211 8044 35256 8072
rect 35250 8032 35256 8044
rect 35308 8032 35314 8084
rect 35434 8032 35440 8084
rect 35492 8072 35498 8084
rect 35802 8072 35808 8084
rect 35492 8044 35808 8072
rect 35492 8032 35498 8044
rect 35802 8032 35808 8044
rect 35860 8072 35866 8084
rect 36262 8072 36268 8084
rect 35860 8044 36268 8072
rect 35860 8032 35866 8044
rect 36262 8032 36268 8044
rect 36320 8032 36326 8084
rect 39114 8032 39120 8084
rect 39172 8072 39178 8084
rect 43530 8072 43536 8084
rect 39172 8044 39712 8072
rect 43491 8044 43536 8072
rect 39172 8032 39178 8044
rect 21453 8007 21511 8013
rect 18984 7976 21414 8004
rect 15841 7939 15899 7945
rect 15841 7905 15853 7939
rect 15887 7905 15899 7939
rect 15841 7899 15899 7905
rect 16117 7939 16175 7945
rect 16117 7905 16129 7939
rect 16163 7936 16175 7939
rect 16574 7936 16580 7948
rect 16163 7908 16580 7936
rect 16163 7905 16175 7908
rect 16117 7899 16175 7905
rect 16574 7896 16580 7908
rect 16632 7896 16638 7948
rect 16942 7896 16948 7948
rect 17000 7936 17006 7948
rect 20162 7936 20168 7948
rect 17000 7908 20168 7936
rect 17000 7896 17006 7908
rect 20162 7896 20168 7908
rect 20220 7896 20226 7948
rect 20898 7936 20904 7948
rect 20859 7908 20904 7936
rect 20898 7896 20904 7908
rect 20956 7896 20962 7948
rect 21082 7936 21088 7948
rect 21043 7908 21088 7936
rect 21082 7896 21088 7908
rect 21140 7896 21146 7948
rect 21386 7936 21414 7976
rect 21453 7973 21465 8007
rect 21499 8004 21511 8007
rect 24394 8004 24400 8016
rect 21499 7976 24400 8004
rect 21499 7973 21511 7976
rect 21453 7967 21511 7973
rect 24394 7964 24400 7976
rect 24452 7964 24458 8016
rect 24486 7964 24492 8016
rect 24544 8004 24550 8016
rect 24581 8007 24639 8013
rect 24581 8004 24593 8007
rect 24544 7976 24593 8004
rect 24544 7964 24550 7976
rect 24581 7973 24593 7976
rect 24627 8004 24639 8007
rect 25866 8004 25872 8016
rect 24627 7976 25872 8004
rect 24627 7973 24639 7976
rect 24581 7967 24639 7973
rect 25866 7964 25872 7976
rect 25924 7964 25930 8016
rect 26510 7964 26516 8016
rect 26568 7964 26574 8016
rect 27890 7964 27896 8016
rect 27948 8004 27954 8016
rect 28902 8004 28908 8016
rect 27948 7976 28908 8004
rect 27948 7964 27954 7976
rect 28902 7964 28908 7976
rect 28960 8004 28966 8016
rect 29181 8007 29239 8013
rect 29181 8004 29193 8007
rect 28960 7976 29193 8004
rect 28960 7964 28966 7976
rect 29181 7973 29193 7976
rect 29227 7973 29239 8007
rect 29181 7967 29239 7973
rect 29362 7964 29368 8016
rect 29420 8004 29426 8016
rect 30190 8004 30196 8016
rect 29420 7976 30196 8004
rect 29420 7964 29426 7976
rect 30190 7964 30196 7976
rect 30248 7964 30254 8016
rect 32766 7964 32772 8016
rect 32824 8004 32830 8016
rect 32953 8007 33011 8013
rect 32953 8004 32965 8007
rect 32824 7976 32965 8004
rect 32824 7964 32830 7976
rect 32953 7973 32965 7976
rect 32999 8004 33011 8007
rect 34238 8004 34244 8016
rect 32999 7976 34244 8004
rect 32999 7973 33011 7976
rect 32953 7967 33011 7973
rect 34238 7964 34244 7976
rect 34296 7964 34302 8016
rect 34333 8007 34391 8013
rect 34333 7973 34345 8007
rect 34379 8004 34391 8007
rect 35618 8004 35624 8016
rect 34379 7976 35624 8004
rect 34379 7973 34391 7976
rect 34333 7967 34391 7973
rect 35618 7964 35624 7976
rect 35676 7964 35682 8016
rect 37921 8007 37979 8013
rect 37921 8004 37933 8007
rect 35728 7976 37933 8004
rect 22281 7939 22339 7945
rect 22281 7936 22293 7939
rect 21386 7908 22293 7936
rect 22281 7905 22293 7908
rect 22327 7936 22339 7939
rect 22925 7939 22983 7945
rect 22925 7936 22937 7939
rect 22327 7908 22937 7936
rect 22327 7905 22339 7908
rect 22281 7899 22339 7905
rect 22925 7905 22937 7908
rect 22971 7936 22983 7939
rect 24302 7936 24308 7948
rect 22971 7908 24308 7936
rect 22971 7905 22983 7908
rect 22925 7899 22983 7905
rect 24302 7896 24308 7908
rect 24360 7936 24366 7948
rect 24857 7939 24915 7945
rect 24857 7936 24869 7939
rect 24360 7908 24869 7936
rect 24360 7896 24366 7908
rect 24857 7905 24869 7908
rect 24903 7905 24915 7939
rect 24857 7899 24915 7905
rect 25961 7939 26019 7945
rect 25961 7905 25973 7939
rect 26007 7936 26019 7939
rect 26326 7936 26332 7948
rect 26007 7908 26332 7936
rect 26007 7905 26019 7908
rect 25961 7899 26019 7905
rect 26326 7896 26332 7908
rect 26384 7896 26390 7948
rect 26528 7936 26556 7964
rect 26789 7939 26847 7945
rect 26789 7936 26801 7939
rect 26528 7908 26801 7936
rect 26789 7905 26801 7908
rect 26835 7905 26847 7939
rect 26789 7899 26847 7905
rect 27430 7896 27436 7948
rect 27488 7936 27494 7948
rect 28810 7936 28816 7948
rect 27488 7908 28816 7936
rect 27488 7896 27494 7908
rect 28810 7896 28816 7908
rect 28868 7896 28874 7948
rect 29086 7896 29092 7948
rect 29144 7936 29150 7948
rect 29273 7939 29331 7945
rect 29273 7936 29285 7939
rect 29144 7908 29285 7936
rect 29144 7896 29150 7908
rect 29273 7905 29285 7908
rect 29319 7905 29331 7939
rect 29273 7899 29331 7905
rect 12805 7871 12863 7877
rect 12805 7837 12817 7871
rect 12851 7868 12863 7871
rect 13354 7868 13360 7880
rect 12851 7840 13360 7868
rect 12851 7837 12863 7840
rect 12805 7831 12863 7837
rect 13354 7828 13360 7840
rect 13412 7828 13418 7880
rect 13906 7828 13912 7880
rect 13964 7868 13970 7880
rect 15289 7871 15347 7877
rect 15289 7868 15301 7871
rect 13964 7840 15301 7868
rect 13964 7828 13970 7840
rect 15289 7837 15301 7840
rect 15335 7837 15347 7871
rect 15289 7831 15347 7837
rect 16206 7828 16212 7880
rect 16264 7868 16270 7880
rect 16301 7871 16359 7877
rect 16301 7868 16313 7871
rect 16264 7840 16313 7868
rect 16264 7828 16270 7840
rect 16301 7837 16313 7840
rect 16347 7837 16359 7871
rect 16301 7831 16359 7837
rect 17494 7828 17500 7880
rect 17552 7868 17558 7880
rect 17589 7871 17647 7877
rect 17589 7868 17601 7871
rect 17552 7840 17601 7868
rect 17552 7828 17558 7840
rect 17589 7837 17601 7840
rect 17635 7837 17647 7871
rect 17589 7831 17647 7837
rect 17865 7871 17923 7877
rect 17865 7837 17877 7871
rect 17911 7868 17923 7871
rect 18230 7868 18236 7880
rect 17911 7840 18236 7868
rect 17911 7837 17923 7840
rect 17865 7831 17923 7837
rect 18230 7828 18236 7840
rect 18288 7828 18294 7880
rect 19702 7868 19708 7880
rect 19663 7840 19708 7868
rect 19702 7828 19708 7840
rect 19760 7828 19766 7880
rect 20916 7868 20944 7896
rect 22097 7871 22155 7877
rect 22097 7868 22109 7871
rect 20916 7840 22109 7868
rect 22097 7837 22109 7840
rect 22143 7837 22155 7871
rect 25222 7868 25228 7880
rect 25183 7840 25228 7868
rect 22097 7831 22155 7837
rect 25222 7828 25228 7840
rect 25280 7828 25286 7880
rect 26513 7871 26571 7877
rect 26513 7837 26525 7871
rect 26559 7868 26571 7871
rect 26694 7868 26700 7880
rect 26559 7840 26700 7868
rect 26559 7837 26571 7840
rect 26513 7831 26571 7837
rect 26694 7828 26700 7840
rect 26752 7828 26758 7880
rect 26970 7828 26976 7880
rect 27028 7868 27034 7880
rect 28169 7871 28227 7877
rect 27028 7840 27476 7868
rect 27028 7828 27034 7840
rect 8260 7772 12204 7800
rect 8260 7760 8266 7772
rect 12434 7760 12440 7812
rect 12492 7800 12498 7812
rect 12529 7803 12587 7809
rect 12529 7800 12541 7803
rect 12492 7772 12541 7800
rect 12492 7760 12498 7772
rect 12529 7769 12541 7772
rect 12575 7800 12587 7803
rect 12575 7772 15516 7800
rect 12575 7769 12587 7772
rect 12529 7763 12587 7769
rect 5629 7735 5687 7741
rect 5629 7701 5641 7735
rect 5675 7732 5687 7735
rect 6270 7732 6276 7744
rect 5675 7704 6276 7732
rect 5675 7701 5687 7704
rect 5629 7695 5687 7701
rect 6270 7692 6276 7704
rect 6328 7732 6334 7744
rect 6730 7732 6736 7744
rect 6328 7704 6736 7732
rect 6328 7692 6334 7704
rect 6730 7692 6736 7704
rect 6788 7692 6794 7744
rect 7558 7692 7564 7744
rect 7616 7732 7622 7744
rect 8021 7735 8079 7741
rect 8021 7732 8033 7735
rect 7616 7704 8033 7732
rect 7616 7692 7622 7704
rect 8021 7701 8033 7704
rect 8067 7701 8079 7735
rect 8021 7695 8079 7701
rect 8754 7692 8760 7744
rect 8812 7732 8818 7744
rect 10505 7735 10563 7741
rect 10505 7732 10517 7735
rect 8812 7704 10517 7732
rect 8812 7692 8818 7704
rect 10505 7701 10517 7704
rect 10551 7732 10563 7735
rect 10781 7735 10839 7741
rect 10781 7732 10793 7735
rect 10551 7704 10793 7732
rect 10551 7701 10563 7704
rect 10505 7695 10563 7701
rect 10781 7701 10793 7704
rect 10827 7732 10839 7735
rect 10962 7732 10968 7744
rect 10827 7704 10968 7732
rect 10827 7701 10839 7704
rect 10781 7695 10839 7701
rect 10962 7692 10968 7704
rect 11020 7692 11026 7744
rect 13078 7732 13084 7744
rect 13039 7704 13084 7732
rect 13078 7692 13084 7704
rect 13136 7692 13142 7744
rect 13262 7692 13268 7744
rect 13320 7732 13326 7744
rect 13630 7732 13636 7744
rect 13320 7704 13636 7732
rect 13320 7692 13326 7704
rect 13630 7692 13636 7704
rect 13688 7692 13694 7744
rect 14458 7732 14464 7744
rect 14419 7704 14464 7732
rect 14458 7692 14464 7704
rect 14516 7692 14522 7744
rect 15488 7732 15516 7772
rect 15746 7760 15752 7812
rect 15804 7800 15810 7812
rect 15804 7772 17356 7800
rect 15804 7760 15810 7772
rect 16666 7732 16672 7744
rect 15488 7704 16672 7732
rect 16666 7692 16672 7704
rect 16724 7692 16730 7744
rect 17328 7732 17356 7772
rect 18874 7760 18880 7812
rect 18932 7800 18938 7812
rect 19981 7803 20039 7809
rect 19981 7800 19993 7803
rect 18932 7772 19993 7800
rect 18932 7760 18938 7772
rect 19981 7769 19993 7772
rect 20027 7769 20039 7803
rect 24121 7803 24179 7809
rect 24121 7800 24133 7803
rect 19981 7763 20039 7769
rect 20088 7772 24133 7800
rect 20088 7732 20116 7772
rect 24121 7769 24133 7772
rect 24167 7769 24179 7803
rect 24121 7763 24179 7769
rect 17328 7704 20116 7732
rect 21821 7735 21879 7741
rect 21821 7701 21833 7735
rect 21867 7732 21879 7735
rect 22278 7732 22284 7744
rect 21867 7704 22284 7732
rect 21867 7701 21879 7704
rect 21821 7695 21879 7701
rect 22278 7692 22284 7704
rect 22336 7692 22342 7744
rect 22462 7732 22468 7744
rect 22423 7704 22468 7732
rect 22462 7692 22468 7704
rect 22520 7692 22526 7744
rect 23290 7732 23296 7744
rect 23251 7704 23296 7732
rect 23290 7692 23296 7704
rect 23348 7732 23354 7744
rect 23753 7735 23811 7741
rect 23753 7732 23765 7735
rect 23348 7704 23765 7732
rect 23348 7692 23354 7704
rect 23753 7701 23765 7704
rect 23799 7701 23811 7735
rect 24136 7732 24164 7763
rect 24854 7760 24860 7812
rect 24912 7800 24918 7812
rect 26234 7800 26240 7812
rect 24912 7772 26240 7800
rect 24912 7760 24918 7772
rect 26234 7760 26240 7772
rect 26292 7760 26298 7812
rect 27448 7800 27476 7840
rect 28169 7837 28181 7871
rect 28215 7868 28227 7871
rect 28997 7871 29055 7877
rect 28997 7868 29009 7871
rect 28215 7840 29009 7868
rect 28215 7837 28227 7840
rect 28169 7831 28227 7837
rect 28997 7837 29009 7840
rect 29043 7837 29055 7871
rect 28997 7831 29055 7837
rect 29012 7800 29040 7831
rect 29086 7800 29092 7812
rect 27448 7772 28580 7800
rect 29012 7772 29092 7800
rect 24765 7735 24823 7741
rect 24765 7732 24777 7735
rect 24136 7704 24777 7732
rect 23753 7695 23811 7701
rect 24765 7701 24777 7704
rect 24811 7732 24823 7735
rect 24995 7735 25053 7741
rect 24995 7732 25007 7735
rect 24811 7704 25007 7732
rect 24811 7701 24823 7704
rect 24765 7695 24823 7701
rect 24995 7701 25007 7704
rect 25041 7701 25053 7735
rect 24995 7695 25053 7701
rect 25133 7735 25191 7741
rect 25133 7701 25145 7735
rect 25179 7732 25191 7735
rect 25314 7732 25320 7744
rect 25179 7704 25320 7732
rect 25179 7701 25191 7704
rect 25133 7695 25191 7701
rect 25314 7692 25320 7704
rect 25372 7692 25378 7744
rect 25501 7735 25559 7741
rect 25501 7701 25513 7735
rect 25547 7732 25559 7735
rect 25774 7732 25780 7744
rect 25547 7704 25780 7732
rect 25547 7701 25559 7704
rect 25501 7695 25559 7701
rect 25774 7692 25780 7704
rect 25832 7692 25838 7744
rect 25866 7692 25872 7744
rect 25924 7732 25930 7744
rect 27982 7732 27988 7744
rect 25924 7704 27988 7732
rect 25924 7692 25930 7704
rect 27982 7692 27988 7704
rect 28040 7692 28046 7744
rect 28442 7732 28448 7744
rect 28403 7704 28448 7732
rect 28442 7692 28448 7704
rect 28500 7692 28506 7744
rect 28552 7732 28580 7772
rect 29086 7760 29092 7772
rect 29144 7760 29150 7812
rect 29288 7800 29316 7899
rect 29914 7896 29920 7948
rect 29972 7936 29978 7948
rect 30561 7939 30619 7945
rect 30561 7936 30573 7939
rect 29972 7908 30573 7936
rect 29972 7896 29978 7908
rect 30561 7905 30573 7908
rect 30607 7936 30619 7939
rect 31202 7936 31208 7948
rect 30607 7908 31208 7936
rect 30607 7905 30619 7908
rect 30561 7899 30619 7905
rect 31202 7896 31208 7908
rect 31260 7896 31266 7948
rect 32401 7939 32459 7945
rect 32401 7905 32413 7939
rect 32447 7936 32459 7939
rect 32490 7936 32496 7948
rect 32447 7908 32496 7936
rect 32447 7905 32459 7908
rect 32401 7899 32459 7905
rect 32490 7896 32496 7908
rect 32548 7936 32554 7948
rect 33873 7939 33931 7945
rect 33873 7936 33885 7939
rect 32548 7908 33885 7936
rect 32548 7896 32554 7908
rect 33873 7905 33885 7908
rect 33919 7936 33931 7939
rect 34698 7936 34704 7948
rect 33919 7908 34704 7936
rect 33919 7905 33931 7908
rect 33873 7899 33931 7905
rect 34698 7896 34704 7908
rect 34756 7896 34762 7948
rect 35161 7939 35219 7945
rect 35161 7936 35173 7939
rect 34900 7908 35173 7936
rect 29454 7828 29460 7880
rect 29512 7868 29518 7880
rect 29733 7871 29791 7877
rect 29733 7868 29745 7871
rect 29512 7840 29745 7868
rect 29512 7828 29518 7840
rect 29733 7837 29745 7840
rect 29779 7837 29791 7871
rect 29733 7831 29791 7837
rect 29822 7828 29828 7880
rect 29880 7868 29886 7880
rect 33686 7868 33692 7880
rect 29880 7840 33692 7868
rect 29880 7828 29886 7840
rect 33686 7828 33692 7840
rect 33744 7828 33750 7880
rect 33778 7828 33784 7880
rect 33836 7868 33842 7880
rect 33836 7840 33881 7868
rect 33836 7828 33842 7840
rect 34238 7828 34244 7880
rect 34296 7868 34302 7880
rect 34900 7868 34928 7908
rect 35161 7905 35173 7908
rect 35207 7936 35219 7939
rect 35728 7936 35756 7976
rect 37921 7973 37933 7976
rect 37967 8004 37979 8007
rect 38010 8004 38016 8016
rect 37967 7976 38016 8004
rect 37967 7973 37979 7976
rect 37921 7967 37979 7973
rect 38010 7964 38016 7976
rect 38068 7964 38074 8016
rect 38470 7964 38476 8016
rect 38528 8004 38534 8016
rect 39684 8004 39712 8044
rect 43530 8032 43536 8044
rect 43588 8032 43594 8084
rect 44085 8075 44143 8081
rect 44085 8041 44097 8075
rect 44131 8072 44143 8075
rect 44266 8072 44272 8084
rect 44131 8044 44272 8072
rect 44131 8041 44143 8044
rect 44085 8035 44143 8041
rect 44266 8032 44272 8044
rect 44324 8032 44330 8084
rect 44450 8032 44456 8084
rect 44508 8072 44514 8084
rect 45462 8072 45468 8084
rect 44508 8044 45468 8072
rect 44508 8032 44514 8044
rect 45462 8032 45468 8044
rect 45520 8032 45526 8084
rect 45738 8072 45744 8084
rect 45699 8044 45744 8072
rect 45738 8032 45744 8044
rect 45796 8032 45802 8084
rect 46937 8075 46995 8081
rect 46937 8041 46949 8075
rect 46983 8041 46995 8075
rect 46937 8035 46995 8041
rect 41877 8007 41935 8013
rect 38528 7976 39620 8004
rect 39684 7976 41828 8004
rect 38528 7964 38534 7976
rect 35207 7908 35756 7936
rect 35989 7939 36047 7945
rect 35207 7905 35219 7908
rect 35161 7899 35219 7905
rect 35989 7905 36001 7939
rect 36035 7936 36047 7939
rect 36357 7939 36415 7945
rect 36357 7936 36369 7939
rect 36035 7908 36369 7936
rect 36035 7905 36047 7908
rect 35989 7899 36047 7905
rect 36357 7905 36369 7908
rect 36403 7905 36415 7939
rect 36357 7899 36415 7905
rect 39114 7896 39120 7948
rect 39172 7936 39178 7948
rect 39592 7945 39620 7976
rect 39209 7939 39267 7945
rect 39209 7936 39221 7939
rect 39172 7908 39221 7936
rect 39172 7896 39178 7908
rect 39209 7905 39221 7908
rect 39255 7905 39267 7939
rect 39209 7899 39267 7905
rect 39577 7939 39635 7945
rect 39577 7905 39589 7939
rect 39623 7936 39635 7939
rect 40310 7936 40316 7948
rect 39623 7908 40316 7936
rect 39623 7905 39635 7908
rect 39577 7899 39635 7905
rect 40310 7896 40316 7908
rect 40368 7896 40374 7948
rect 41417 7939 41475 7945
rect 41417 7905 41429 7939
rect 41463 7936 41475 7939
rect 41690 7936 41696 7948
rect 41463 7908 41696 7936
rect 41463 7905 41475 7908
rect 41417 7899 41475 7905
rect 41690 7896 41696 7908
rect 41748 7896 41754 7948
rect 41800 7936 41828 7976
rect 41877 7973 41889 8007
rect 41923 8004 41935 8007
rect 43622 8004 43628 8016
rect 41923 7976 43628 8004
rect 41923 7973 41935 7976
rect 41877 7967 41935 7973
rect 43622 7964 43628 7976
rect 43680 7964 43686 8016
rect 44177 8007 44235 8013
rect 44177 7973 44189 8007
rect 44223 8004 44235 8007
rect 45094 8004 45100 8016
rect 44223 7976 45100 8004
rect 44223 7973 44235 7976
rect 44177 7967 44235 7973
rect 45094 7964 45100 7976
rect 45152 7964 45158 8016
rect 45480 8004 45508 8032
rect 45646 8004 45652 8016
rect 45480 7976 45652 8004
rect 45646 7964 45652 7976
rect 45704 7964 45710 8016
rect 44818 7936 44824 7948
rect 41800 7908 44824 7936
rect 44818 7896 44824 7908
rect 44876 7896 44882 7948
rect 45186 7936 45192 7948
rect 45147 7908 45192 7936
rect 45186 7896 45192 7908
rect 45244 7896 45250 7948
rect 45373 7939 45431 7945
rect 45373 7905 45385 7939
rect 45419 7936 45431 7939
rect 45756 7936 45784 8032
rect 46952 8004 46980 8035
rect 47026 8032 47032 8084
rect 47084 8072 47090 8084
rect 47302 8072 47308 8084
rect 47084 8044 47308 8072
rect 47084 8032 47090 8044
rect 47302 8032 47308 8044
rect 47360 8032 47366 8084
rect 48041 8075 48099 8081
rect 48041 8041 48053 8075
rect 48087 8072 48099 8075
rect 50338 8072 50344 8084
rect 48087 8044 50344 8072
rect 48087 8041 48099 8044
rect 48041 8035 48099 8041
rect 50338 8032 50344 8044
rect 50396 8032 50402 8084
rect 50985 8075 51043 8081
rect 50985 8041 50997 8075
rect 51031 8072 51043 8075
rect 51074 8072 51080 8084
rect 51031 8044 51080 8072
rect 51031 8041 51043 8044
rect 50985 8035 51043 8041
rect 51074 8032 51080 8044
rect 51132 8032 51138 8084
rect 51350 8072 51356 8084
rect 51311 8044 51356 8072
rect 51350 8032 51356 8044
rect 51408 8032 51414 8084
rect 52178 8032 52184 8084
rect 52236 8072 52242 8084
rect 52825 8075 52883 8081
rect 52825 8072 52837 8075
rect 52236 8044 52837 8072
rect 52236 8032 52242 8044
rect 52825 8041 52837 8044
rect 52871 8072 52883 8075
rect 53374 8072 53380 8084
rect 52871 8044 53380 8072
rect 52871 8041 52883 8044
rect 52825 8035 52883 8041
rect 53374 8032 53380 8044
rect 53432 8032 53438 8084
rect 53926 8072 53932 8084
rect 53839 8044 53932 8072
rect 53926 8032 53932 8044
rect 53984 8072 53990 8084
rect 54297 8075 54355 8081
rect 54297 8072 54309 8075
rect 53984 8044 54309 8072
rect 53984 8032 53990 8044
rect 54297 8041 54309 8044
rect 54343 8072 54355 8075
rect 55122 8072 55128 8084
rect 54343 8044 55128 8072
rect 54343 8041 54355 8044
rect 54297 8035 54355 8041
rect 55122 8032 55128 8044
rect 55180 8032 55186 8084
rect 55306 8032 55312 8084
rect 55364 8072 55370 8084
rect 55493 8075 55551 8081
rect 55493 8072 55505 8075
rect 55364 8044 55505 8072
rect 55364 8032 55370 8044
rect 55493 8041 55505 8044
rect 55539 8041 55551 8075
rect 55493 8035 55551 8041
rect 57425 8075 57483 8081
rect 57425 8041 57437 8075
rect 57471 8072 57483 8075
rect 57606 8072 57612 8084
rect 57471 8044 57612 8072
rect 57471 8041 57483 8044
rect 57425 8035 57483 8041
rect 53834 8004 53840 8016
rect 46952 7976 53840 8004
rect 53834 7964 53840 7976
rect 53892 7964 53898 8016
rect 55508 8004 55536 8035
rect 57606 8032 57612 8044
rect 57664 8032 57670 8084
rect 58158 8032 58164 8084
rect 58216 8072 58222 8084
rect 58434 8072 58440 8084
rect 58216 8044 58440 8072
rect 58216 8032 58222 8044
rect 58434 8032 58440 8044
rect 58492 8072 58498 8084
rect 58989 8075 59047 8081
rect 58989 8072 59001 8075
rect 58492 8044 59001 8072
rect 58492 8032 58498 8044
rect 58989 8041 59001 8044
rect 59035 8041 59047 8075
rect 58989 8035 59047 8041
rect 59262 8032 59268 8084
rect 59320 8072 59326 8084
rect 59357 8075 59415 8081
rect 59357 8072 59369 8075
rect 59320 8044 59369 8072
rect 59320 8032 59326 8044
rect 59357 8041 59369 8044
rect 59403 8041 59415 8075
rect 59357 8035 59415 8041
rect 57517 8007 57575 8013
rect 55508 7976 56364 8004
rect 45419 7908 45784 7936
rect 47305 7939 47363 7945
rect 45419 7905 45431 7908
rect 45373 7899 45431 7905
rect 47305 7905 47317 7939
rect 47351 7936 47363 7939
rect 47394 7936 47400 7948
rect 47351 7908 47400 7936
rect 47351 7905 47363 7908
rect 47305 7899 47363 7905
rect 47394 7896 47400 7908
rect 47452 7896 47458 7948
rect 47670 7936 47676 7948
rect 47631 7908 47676 7936
rect 47670 7896 47676 7908
rect 47728 7896 47734 7948
rect 47765 7939 47823 7945
rect 47765 7905 47777 7939
rect 47811 7905 47823 7939
rect 47765 7899 47823 7905
rect 34296 7840 34928 7868
rect 34296 7828 34302 7840
rect 34974 7828 34980 7880
rect 35032 7868 35038 7880
rect 35069 7871 35127 7877
rect 35069 7868 35081 7871
rect 35032 7840 35081 7868
rect 35032 7828 35038 7840
rect 35069 7837 35081 7840
rect 35115 7868 35127 7871
rect 35710 7868 35716 7880
rect 35115 7840 35716 7868
rect 35115 7837 35127 7840
rect 35069 7831 35127 7837
rect 35710 7828 35716 7840
rect 35768 7828 35774 7880
rect 35894 7868 35900 7880
rect 35855 7840 35900 7868
rect 35894 7828 35900 7840
rect 35952 7868 35958 7880
rect 36909 7871 36967 7877
rect 36909 7868 36921 7871
rect 35952 7840 36921 7868
rect 35952 7828 35958 7840
rect 36909 7837 36921 7840
rect 36955 7868 36967 7871
rect 37369 7871 37427 7877
rect 37369 7868 37381 7871
rect 36955 7840 37381 7868
rect 36955 7837 36967 7840
rect 36909 7831 36967 7837
rect 37369 7837 37381 7840
rect 37415 7837 37427 7871
rect 37369 7831 37427 7837
rect 38473 7871 38531 7877
rect 38473 7837 38485 7871
rect 38519 7868 38531 7871
rect 39298 7868 39304 7880
rect 38519 7840 39304 7868
rect 38519 7837 38531 7840
rect 38473 7831 38531 7837
rect 39298 7828 39304 7840
rect 39356 7828 39362 7880
rect 39666 7868 39672 7880
rect 39627 7840 39672 7868
rect 39666 7828 39672 7840
rect 39724 7828 39730 7880
rect 41325 7871 41383 7877
rect 41325 7837 41337 7871
rect 41371 7868 41383 7871
rect 41966 7868 41972 7880
rect 41371 7840 41972 7868
rect 41371 7837 41383 7840
rect 41325 7831 41383 7837
rect 41966 7828 41972 7840
rect 42024 7828 42030 7880
rect 42242 7868 42248 7880
rect 42155 7840 42248 7868
rect 42242 7828 42248 7840
rect 42300 7868 42306 7880
rect 44266 7868 44272 7880
rect 42300 7840 44272 7868
rect 42300 7828 42306 7840
rect 44266 7828 44272 7840
rect 44324 7828 44330 7880
rect 44726 7868 44732 7880
rect 44687 7840 44732 7868
rect 44726 7828 44732 7840
rect 44784 7828 44790 7880
rect 46934 7828 46940 7880
rect 46992 7868 46998 7880
rect 47121 7871 47179 7877
rect 47121 7868 47133 7871
rect 46992 7840 47133 7868
rect 46992 7828 46998 7840
rect 47121 7837 47133 7840
rect 47167 7837 47179 7871
rect 47780 7868 47808 7899
rect 48774 7896 48780 7948
rect 48832 7936 48838 7948
rect 48961 7939 49019 7945
rect 48961 7936 48973 7939
rect 48832 7908 48973 7936
rect 48832 7896 48838 7908
rect 48961 7905 48973 7908
rect 49007 7905 49019 7939
rect 49142 7936 49148 7948
rect 49103 7908 49148 7936
rect 48961 7899 49019 7905
rect 49142 7896 49148 7908
rect 49200 7896 49206 7948
rect 50341 7939 50399 7945
rect 50341 7936 50353 7939
rect 49436 7908 50353 7936
rect 47121 7831 47179 7837
rect 47688 7840 47808 7868
rect 47688 7812 47716 7840
rect 48130 7828 48136 7880
rect 48188 7868 48194 7880
rect 48501 7871 48559 7877
rect 48501 7868 48513 7871
rect 48188 7840 48513 7868
rect 48188 7828 48194 7840
rect 48501 7837 48513 7840
rect 48547 7868 48559 7871
rect 49436 7868 49464 7908
rect 50341 7905 50353 7908
rect 50387 7936 50399 7939
rect 51994 7936 52000 7948
rect 50387 7908 50936 7936
rect 51955 7908 52000 7936
rect 50387 7905 50399 7908
rect 50341 7899 50399 7905
rect 48547 7840 49464 7868
rect 49513 7871 49571 7877
rect 48547 7837 48559 7840
rect 48501 7831 48559 7837
rect 49513 7837 49525 7871
rect 49559 7868 49571 7871
rect 49786 7868 49792 7880
rect 49559 7840 49792 7868
rect 49559 7837 49571 7840
rect 49513 7831 49571 7837
rect 49786 7828 49792 7840
rect 49844 7828 49850 7880
rect 49878 7828 49884 7880
rect 49936 7868 49942 7880
rect 50246 7868 50252 7880
rect 49936 7840 50252 7868
rect 49936 7828 49942 7840
rect 50246 7828 50252 7840
rect 50304 7868 50310 7880
rect 50304 7840 50660 7868
rect 50304 7828 50310 7840
rect 30377 7803 30435 7809
rect 30377 7800 30389 7803
rect 29288 7772 30389 7800
rect 30377 7769 30389 7772
rect 30423 7769 30435 7803
rect 30377 7763 30435 7769
rect 36357 7803 36415 7809
rect 36357 7769 36369 7803
rect 36403 7800 36415 7803
rect 36633 7803 36691 7809
rect 36633 7800 36645 7803
rect 36403 7772 36645 7800
rect 36403 7769 36415 7772
rect 36357 7763 36415 7769
rect 36633 7769 36645 7772
rect 36679 7800 36691 7803
rect 38286 7800 38292 7812
rect 36679 7772 38292 7800
rect 36679 7769 36691 7772
rect 36633 7763 36691 7769
rect 38286 7760 38292 7772
rect 38344 7760 38350 7812
rect 38657 7803 38715 7809
rect 38657 7769 38669 7803
rect 38703 7800 38715 7803
rect 38746 7800 38752 7812
rect 38703 7772 38752 7800
rect 38703 7769 38715 7772
rect 38657 7763 38715 7769
rect 38746 7760 38752 7772
rect 38804 7760 38810 7812
rect 39206 7760 39212 7812
rect 39264 7800 39270 7812
rect 40129 7803 40187 7809
rect 40129 7800 40141 7803
rect 39264 7772 40141 7800
rect 39264 7760 39270 7772
rect 40129 7769 40141 7772
rect 40175 7800 40187 7803
rect 40175 7772 41460 7800
rect 40175 7769 40187 7772
rect 40129 7763 40187 7769
rect 29362 7732 29368 7744
rect 28552 7704 29368 7732
rect 29362 7692 29368 7704
rect 29420 7692 29426 7744
rect 29914 7692 29920 7744
rect 29972 7732 29978 7744
rect 30745 7735 30803 7741
rect 30745 7732 30757 7735
rect 29972 7704 30757 7732
rect 29972 7692 29978 7704
rect 30745 7701 30757 7704
rect 30791 7701 30803 7735
rect 31202 7732 31208 7744
rect 31163 7704 31208 7732
rect 30745 7695 30803 7701
rect 31202 7692 31208 7704
rect 31260 7692 31266 7744
rect 31478 7732 31484 7744
rect 31439 7704 31484 7732
rect 31478 7692 31484 7704
rect 31536 7692 31542 7744
rect 33962 7692 33968 7744
rect 34020 7732 34026 7744
rect 34514 7732 34520 7744
rect 34020 7704 34520 7732
rect 34020 7692 34026 7704
rect 34514 7692 34520 7704
rect 34572 7692 34578 7744
rect 39758 7692 39764 7744
rect 39816 7732 39822 7744
rect 40497 7735 40555 7741
rect 40497 7732 40509 7735
rect 39816 7704 40509 7732
rect 39816 7692 39822 7704
rect 40497 7701 40509 7704
rect 40543 7701 40555 7735
rect 40862 7732 40868 7744
rect 40823 7704 40868 7732
rect 40497 7695 40555 7701
rect 40862 7692 40868 7704
rect 40920 7692 40926 7744
rect 41432 7732 41460 7772
rect 41598 7760 41604 7812
rect 41656 7800 41662 7812
rect 47486 7800 47492 7812
rect 41656 7772 47492 7800
rect 41656 7760 41662 7772
rect 47486 7760 47492 7772
rect 47544 7760 47550 7812
rect 47670 7760 47676 7812
rect 47728 7760 47734 7812
rect 47946 7760 47952 7812
rect 48004 7800 48010 7812
rect 48406 7800 48412 7812
rect 48004 7772 48412 7800
rect 48004 7760 48010 7772
rect 48406 7760 48412 7772
rect 48464 7760 48470 7812
rect 48590 7760 48596 7812
rect 48648 7800 48654 7812
rect 50479 7803 50537 7809
rect 50479 7800 50491 7803
rect 48648 7772 50491 7800
rect 48648 7760 48654 7772
rect 50479 7769 50491 7772
rect 50525 7769 50537 7803
rect 50632 7800 50660 7840
rect 50706 7828 50712 7880
rect 50764 7868 50770 7880
rect 50908 7868 50936 7908
rect 51994 7896 52000 7908
rect 52052 7896 52058 7948
rect 52454 7896 52460 7948
rect 52512 7936 52518 7948
rect 53285 7939 53343 7945
rect 53285 7936 53297 7939
rect 52512 7908 53297 7936
rect 52512 7896 52518 7908
rect 53285 7905 53297 7908
rect 53331 7936 53343 7939
rect 53742 7936 53748 7948
rect 53331 7908 53748 7936
rect 53331 7905 53343 7908
rect 53285 7899 53343 7905
rect 53742 7896 53748 7908
rect 53800 7896 53806 7948
rect 56134 7936 56140 7948
rect 56095 7908 56140 7936
rect 56134 7896 56140 7908
rect 56192 7896 56198 7948
rect 56336 7945 56364 7976
rect 57517 7973 57529 8007
rect 57563 8004 57575 8007
rect 59078 8004 59084 8016
rect 57563 7976 59084 8004
rect 57563 7973 57575 7976
rect 57517 7967 57575 7973
rect 59078 7964 59084 7976
rect 59136 7964 59142 8016
rect 61197 8007 61255 8013
rect 61197 8004 61209 8007
rect 60476 7976 61209 8004
rect 56321 7939 56379 7945
rect 56321 7905 56333 7939
rect 56367 7905 56379 7939
rect 56321 7899 56379 7905
rect 56505 7939 56563 7945
rect 56505 7905 56517 7939
rect 56551 7905 56563 7939
rect 56505 7899 56563 7905
rect 51721 7871 51779 7877
rect 51721 7868 51733 7871
rect 50764 7840 50809 7868
rect 50908 7840 51733 7868
rect 50764 7828 50770 7840
rect 51721 7837 51733 7840
rect 51767 7837 51779 7871
rect 51902 7868 51908 7880
rect 51863 7840 51908 7868
rect 51721 7831 51779 7837
rect 51902 7828 51908 7840
rect 51960 7828 51966 7880
rect 55398 7828 55404 7880
rect 55456 7868 55462 7880
rect 56520 7868 56548 7899
rect 56686 7896 56692 7948
rect 56744 7936 56750 7948
rect 58158 7936 58164 7948
rect 56744 7908 58164 7936
rect 56744 7896 56750 7908
rect 58158 7896 58164 7908
rect 58216 7896 58222 7948
rect 58250 7896 58256 7948
rect 58308 7936 58314 7948
rect 58529 7939 58587 7945
rect 58308 7908 58353 7936
rect 58308 7896 58314 7908
rect 58529 7905 58541 7939
rect 58575 7905 58587 7939
rect 58710 7936 58716 7948
rect 58671 7908 58716 7936
rect 58529 7899 58587 7905
rect 55456 7840 56548 7868
rect 55456 7828 55462 7840
rect 57514 7828 57520 7880
rect 57572 7868 57578 7880
rect 58544 7868 58572 7899
rect 58710 7896 58716 7908
rect 58768 7896 58774 7948
rect 60476 7945 60504 7976
rect 61197 7973 61209 7976
rect 61243 7973 61255 8007
rect 61197 7967 61255 7973
rect 60461 7939 60519 7945
rect 60461 7905 60473 7939
rect 60507 7905 60519 7939
rect 60918 7936 60924 7948
rect 60879 7908 60924 7936
rect 60461 7899 60519 7905
rect 60476 7868 60504 7899
rect 60918 7896 60924 7908
rect 60976 7896 60982 7948
rect 57572 7840 58572 7868
rect 58636 7840 60504 7868
rect 57572 7828 57578 7840
rect 53469 7803 53527 7809
rect 53469 7800 53481 7803
rect 50632 7772 53481 7800
rect 50479 7763 50537 7769
rect 53469 7769 53481 7772
rect 53515 7769 53527 7803
rect 55950 7800 55956 7812
rect 55911 7772 55956 7800
rect 53469 7763 53527 7769
rect 55950 7760 55956 7772
rect 56008 7760 56014 7812
rect 56318 7760 56324 7812
rect 56376 7800 56382 7812
rect 58636 7800 58664 7840
rect 56376 7772 58664 7800
rect 56376 7760 56382 7772
rect 59446 7760 59452 7812
rect 59504 7800 59510 7812
rect 60277 7803 60335 7809
rect 60277 7800 60289 7803
rect 59504 7772 60289 7800
rect 59504 7760 59510 7772
rect 60277 7769 60289 7772
rect 60323 7769 60335 7803
rect 60277 7763 60335 7769
rect 41874 7732 41880 7744
rect 41432 7704 41880 7732
rect 41874 7692 41880 7704
rect 41932 7692 41938 7744
rect 42426 7692 42432 7744
rect 42484 7732 42490 7744
rect 42613 7735 42671 7741
rect 42613 7732 42625 7735
rect 42484 7704 42625 7732
rect 42484 7692 42490 7704
rect 42613 7701 42625 7704
rect 42659 7701 42671 7735
rect 43070 7732 43076 7744
rect 43031 7704 43076 7732
rect 42613 7695 42671 7701
rect 43070 7692 43076 7704
rect 43128 7692 43134 7744
rect 46198 7732 46204 7744
rect 46159 7704 46204 7732
rect 46198 7692 46204 7704
rect 46256 7692 46262 7744
rect 46658 7692 46664 7744
rect 46716 7732 46722 7744
rect 48041 7735 48099 7741
rect 48041 7732 48053 7735
rect 46716 7704 48053 7732
rect 46716 7692 46722 7704
rect 48041 7701 48053 7704
rect 48087 7701 48099 7735
rect 48222 7732 48228 7744
rect 48183 7704 48228 7732
rect 48041 7695 48099 7701
rect 48222 7692 48228 7704
rect 48280 7692 48286 7744
rect 49602 7692 49608 7744
rect 49660 7732 49666 7744
rect 49881 7735 49939 7741
rect 49881 7732 49893 7735
rect 49660 7704 49893 7732
rect 49660 7692 49666 7704
rect 49881 7701 49893 7704
rect 49927 7701 49939 7735
rect 50614 7732 50620 7744
rect 50575 7704 50620 7732
rect 49881 7695 49939 7701
rect 50614 7692 50620 7704
rect 50672 7692 50678 7744
rect 51166 7692 51172 7744
rect 51224 7732 51230 7744
rect 52181 7735 52239 7741
rect 52181 7732 52193 7735
rect 51224 7704 52193 7732
rect 51224 7692 51230 7704
rect 52181 7701 52193 7704
rect 52227 7701 52239 7735
rect 52181 7695 52239 7701
rect 53193 7735 53251 7741
rect 53193 7701 53205 7735
rect 53239 7732 53251 7735
rect 53282 7732 53288 7744
rect 53239 7704 53288 7732
rect 53239 7701 53251 7704
rect 53193 7695 53251 7701
rect 53282 7692 53288 7704
rect 53340 7692 53346 7744
rect 54294 7692 54300 7744
rect 54352 7732 54358 7744
rect 54757 7735 54815 7741
rect 54757 7732 54769 7735
rect 54352 7704 54769 7732
rect 54352 7692 54358 7704
rect 54757 7701 54769 7704
rect 54803 7701 54815 7735
rect 54757 7695 54815 7701
rect 55858 7692 55864 7744
rect 55916 7732 55922 7744
rect 56965 7735 57023 7741
rect 56965 7732 56977 7735
rect 55916 7704 56977 7732
rect 55916 7692 55922 7704
rect 56965 7701 56977 7704
rect 57011 7701 57023 7735
rect 56965 7695 57023 7701
rect 59630 7692 59636 7744
rect 59688 7732 59694 7744
rect 59817 7735 59875 7741
rect 59817 7732 59829 7735
rect 59688 7704 59829 7732
rect 59688 7692 59694 7704
rect 59817 7701 59829 7704
rect 59863 7701 59875 7735
rect 59817 7695 59875 7701
rect 1104 7642 63480 7664
rect 1104 7590 11378 7642
rect 11430 7590 11442 7642
rect 11494 7590 11506 7642
rect 11558 7590 11570 7642
rect 11622 7590 32170 7642
rect 32222 7590 32234 7642
rect 32286 7590 32298 7642
rect 32350 7590 32362 7642
rect 32414 7590 52962 7642
rect 53014 7590 53026 7642
rect 53078 7590 53090 7642
rect 53142 7590 53154 7642
rect 53206 7590 63480 7642
rect 1104 7568 63480 7590
rect 4338 7528 4344 7540
rect 4299 7500 4344 7528
rect 4338 7488 4344 7500
rect 4396 7488 4402 7540
rect 7101 7531 7159 7537
rect 7101 7497 7113 7531
rect 7147 7528 7159 7531
rect 8846 7528 8852 7540
rect 7147 7500 8852 7528
rect 7147 7497 7159 7500
rect 7101 7491 7159 7497
rect 8846 7488 8852 7500
rect 8904 7488 8910 7540
rect 11425 7531 11483 7537
rect 9140 7500 10824 7528
rect 7742 7420 7748 7472
rect 7800 7460 7806 7472
rect 8754 7460 8760 7472
rect 7800 7432 8760 7460
rect 7800 7420 7806 7432
rect 8754 7420 8760 7432
rect 8812 7420 8818 7472
rect 5442 7392 5448 7404
rect 5403 7364 5448 7392
rect 5442 7352 5448 7364
rect 5500 7352 5506 7404
rect 6270 7392 6276 7404
rect 5736 7364 6276 7392
rect 5736 7333 5764 7364
rect 6270 7352 6276 7364
rect 6328 7352 6334 7404
rect 6730 7352 6736 7404
rect 6788 7392 6794 7404
rect 9033 7395 9091 7401
rect 9033 7392 9045 7395
rect 6788 7364 9045 7392
rect 6788 7352 6794 7364
rect 5721 7327 5779 7333
rect 5721 7293 5733 7327
rect 5767 7293 5779 7327
rect 5721 7287 5779 7293
rect 5905 7327 5963 7333
rect 5905 7293 5917 7327
rect 5951 7324 5963 7327
rect 6546 7324 6552 7336
rect 5951 7296 6552 7324
rect 5951 7293 5963 7296
rect 5905 7287 5963 7293
rect 6546 7284 6552 7296
rect 6604 7284 6610 7336
rect 7098 7284 7104 7336
rect 7156 7324 7162 7336
rect 7484 7333 7512 7364
rect 9033 7361 9045 7364
rect 9079 7361 9091 7395
rect 9033 7355 9091 7361
rect 7285 7327 7343 7333
rect 7285 7324 7297 7327
rect 7156 7296 7297 7324
rect 7156 7284 7162 7296
rect 7285 7293 7297 7296
rect 7331 7293 7343 7327
rect 7285 7287 7343 7293
rect 7469 7327 7527 7333
rect 7469 7293 7481 7327
rect 7515 7293 7527 7327
rect 7469 7287 7527 7293
rect 4890 7256 4896 7268
rect 4851 7228 4896 7256
rect 4890 7216 4896 7228
rect 4948 7216 4954 7268
rect 7300 7256 7328 7287
rect 7742 7284 7748 7336
rect 7800 7333 7806 7336
rect 7800 7327 7849 7333
rect 7800 7293 7803 7327
rect 7837 7293 7849 7327
rect 7926 7324 7932 7336
rect 7887 7296 7932 7324
rect 7800 7287 7849 7293
rect 7800 7284 7806 7287
rect 7926 7284 7932 7296
rect 7984 7284 7990 7336
rect 8202 7256 8208 7268
rect 7300 7228 8208 7256
rect 8202 7216 8208 7228
rect 8260 7256 8266 7268
rect 8297 7259 8355 7265
rect 8297 7256 8309 7259
rect 8260 7228 8309 7256
rect 8260 7216 8266 7228
rect 8297 7225 8309 7228
rect 8343 7225 8355 7259
rect 8297 7219 8355 7225
rect 3694 7188 3700 7200
rect 3655 7160 3700 7188
rect 3694 7148 3700 7160
rect 3752 7188 3758 7200
rect 3973 7191 4031 7197
rect 3973 7188 3985 7191
rect 3752 7160 3985 7188
rect 3752 7148 3758 7160
rect 3973 7157 3985 7160
rect 4019 7188 4031 7191
rect 4062 7188 4068 7200
rect 4019 7160 4068 7188
rect 4019 7157 4031 7160
rect 3973 7151 4031 7157
rect 4062 7148 4068 7160
rect 4120 7188 4126 7200
rect 4709 7191 4767 7197
rect 4709 7188 4721 7191
rect 4120 7160 4721 7188
rect 4120 7148 4126 7160
rect 4709 7157 4721 7160
rect 4755 7157 4767 7191
rect 4709 7151 4767 7157
rect 5534 7148 5540 7200
rect 5592 7188 5598 7200
rect 6549 7191 6607 7197
rect 6549 7188 6561 7191
rect 5592 7160 6561 7188
rect 5592 7148 5598 7160
rect 6549 7157 6561 7160
rect 6595 7188 6607 7191
rect 6822 7188 6828 7200
rect 6595 7160 6828 7188
rect 6595 7157 6607 7160
rect 6549 7151 6607 7157
rect 6822 7148 6828 7160
rect 6880 7188 6886 7200
rect 9140 7188 9168 7500
rect 10796 7460 10824 7500
rect 11425 7497 11437 7531
rect 11471 7528 11483 7531
rect 12526 7528 12532 7540
rect 11471 7500 12532 7528
rect 11471 7497 11483 7500
rect 11425 7491 11483 7497
rect 12526 7488 12532 7500
rect 12584 7488 12590 7540
rect 12621 7531 12679 7537
rect 12621 7497 12633 7531
rect 12667 7528 12679 7531
rect 12897 7531 12955 7537
rect 12897 7528 12909 7531
rect 12667 7500 12909 7528
rect 12667 7497 12679 7500
rect 12621 7491 12679 7497
rect 12897 7497 12909 7500
rect 12943 7528 12955 7531
rect 12943 7500 15700 7528
rect 12943 7497 12955 7500
rect 12897 7491 12955 7497
rect 13354 7460 13360 7472
rect 10796 7432 13216 7460
rect 13315 7432 13360 7460
rect 9769 7395 9827 7401
rect 9769 7361 9781 7395
rect 9815 7392 9827 7395
rect 10137 7395 10195 7401
rect 10137 7392 10149 7395
rect 9815 7364 10149 7392
rect 9815 7361 9827 7364
rect 9769 7355 9827 7361
rect 10137 7361 10149 7364
rect 10183 7392 10195 7395
rect 12526 7392 12532 7404
rect 10183 7364 12532 7392
rect 10183 7361 10195 7364
rect 10137 7355 10195 7361
rect 12526 7352 12532 7364
rect 12584 7352 12590 7404
rect 13078 7392 13084 7404
rect 13039 7364 13084 7392
rect 13078 7352 13084 7364
rect 13136 7352 13142 7404
rect 9861 7327 9919 7333
rect 9861 7293 9873 7327
rect 9907 7324 9919 7327
rect 10226 7324 10232 7336
rect 9907 7296 10232 7324
rect 9907 7293 9919 7296
rect 9861 7287 9919 7293
rect 10226 7284 10232 7296
rect 10284 7324 10290 7336
rect 12342 7324 12348 7336
rect 10284 7296 12348 7324
rect 10284 7284 10290 7296
rect 12342 7284 12348 7296
rect 12400 7284 12406 7336
rect 12434 7284 12440 7336
rect 12492 7324 12498 7336
rect 12492 7296 12537 7324
rect 12492 7284 12498 7296
rect 12897 7259 12955 7265
rect 12897 7256 12909 7259
rect 10796 7228 12909 7256
rect 6880 7160 9168 7188
rect 6880 7148 6886 7160
rect 9950 7148 9956 7200
rect 10008 7188 10014 7200
rect 10796 7188 10824 7228
rect 12897 7225 12909 7228
rect 12943 7225 12955 7259
rect 13188 7256 13216 7432
rect 13354 7420 13360 7432
rect 13412 7420 13418 7472
rect 15672 7460 15700 7500
rect 16758 7488 16764 7540
rect 16816 7528 16822 7540
rect 16853 7531 16911 7537
rect 16853 7528 16865 7531
rect 16816 7500 16865 7528
rect 16816 7488 16822 7500
rect 16853 7497 16865 7500
rect 16899 7497 16911 7531
rect 18230 7528 18236 7540
rect 18191 7500 18236 7528
rect 16853 7491 16911 7497
rect 18230 7488 18236 7500
rect 18288 7488 18294 7540
rect 19245 7531 19303 7537
rect 19245 7497 19257 7531
rect 19291 7528 19303 7531
rect 20898 7528 20904 7540
rect 19291 7500 20904 7528
rect 19291 7497 19303 7500
rect 19245 7491 19303 7497
rect 20898 7488 20904 7500
rect 20956 7488 20962 7540
rect 23474 7528 23480 7540
rect 23435 7500 23480 7528
rect 23474 7488 23480 7500
rect 23532 7488 23538 7540
rect 25041 7531 25099 7537
rect 25041 7497 25053 7531
rect 25087 7528 25099 7531
rect 25314 7528 25320 7540
rect 25087 7500 25320 7528
rect 25087 7497 25099 7500
rect 25041 7491 25099 7497
rect 25314 7488 25320 7500
rect 25372 7488 25378 7540
rect 25869 7531 25927 7537
rect 25869 7497 25881 7531
rect 25915 7528 25927 7531
rect 26510 7528 26516 7540
rect 25915 7500 26516 7528
rect 25915 7497 25927 7500
rect 25869 7491 25927 7497
rect 26510 7488 26516 7500
rect 26568 7528 26574 7540
rect 27249 7531 27307 7537
rect 27249 7528 27261 7531
rect 26568 7500 27261 7528
rect 26568 7488 26574 7500
rect 27249 7497 27261 7500
rect 27295 7497 27307 7531
rect 27249 7491 27307 7497
rect 28445 7531 28503 7537
rect 28445 7497 28457 7531
rect 28491 7528 28503 7531
rect 28718 7528 28724 7540
rect 28491 7500 28724 7528
rect 28491 7497 28503 7500
rect 28445 7491 28503 7497
rect 28718 7488 28724 7500
rect 28776 7488 28782 7540
rect 28810 7488 28816 7540
rect 28868 7528 28874 7540
rect 28868 7500 29960 7528
rect 28868 7488 28874 7500
rect 24762 7460 24768 7472
rect 15672 7432 24768 7460
rect 24762 7420 24768 7432
rect 24820 7420 24826 7472
rect 29822 7460 29828 7472
rect 24872 7432 29828 7460
rect 13538 7352 13544 7404
rect 13596 7392 13602 7404
rect 14093 7395 14151 7401
rect 14093 7392 14105 7395
rect 13596 7364 14105 7392
rect 13596 7352 13602 7364
rect 14093 7361 14105 7364
rect 14139 7392 14151 7395
rect 15286 7392 15292 7404
rect 14139 7364 15292 7392
rect 14139 7361 14151 7364
rect 14093 7355 14151 7361
rect 15286 7352 15292 7364
rect 15344 7352 15350 7404
rect 15746 7392 15752 7404
rect 15707 7364 15752 7392
rect 15746 7352 15752 7364
rect 15804 7352 15810 7404
rect 17218 7352 17224 7404
rect 17276 7392 17282 7404
rect 24872 7392 24900 7432
rect 29822 7420 29828 7432
rect 29880 7420 29886 7472
rect 29932 7460 29960 7500
rect 30190 7488 30196 7540
rect 30248 7528 30254 7540
rect 30653 7531 30711 7537
rect 30653 7528 30665 7531
rect 30248 7500 30665 7528
rect 30248 7488 30254 7500
rect 30653 7497 30665 7500
rect 30699 7497 30711 7531
rect 31018 7528 31024 7540
rect 30979 7500 31024 7528
rect 30653 7491 30711 7497
rect 31018 7488 31024 7500
rect 31076 7488 31082 7540
rect 33870 7528 33876 7540
rect 33831 7500 33876 7528
rect 33870 7488 33876 7500
rect 33928 7488 33934 7540
rect 34606 7488 34612 7540
rect 34664 7528 34670 7540
rect 35161 7531 35219 7537
rect 35161 7528 35173 7531
rect 34664 7500 35173 7528
rect 34664 7488 34670 7500
rect 35161 7497 35173 7500
rect 35207 7497 35219 7531
rect 41690 7528 41696 7540
rect 41651 7500 41696 7528
rect 35161 7491 35219 7497
rect 41690 7488 41696 7500
rect 41748 7488 41754 7540
rect 41966 7488 41972 7540
rect 42024 7528 42030 7540
rect 42061 7531 42119 7537
rect 42061 7528 42073 7531
rect 42024 7500 42073 7528
rect 42024 7488 42030 7500
rect 42061 7497 42073 7500
rect 42107 7528 42119 7531
rect 42794 7528 42800 7540
rect 42107 7500 42800 7528
rect 42107 7497 42119 7500
rect 42061 7491 42119 7497
rect 42794 7488 42800 7500
rect 42852 7488 42858 7540
rect 44726 7528 44732 7540
rect 44687 7500 44732 7528
rect 44726 7488 44732 7500
rect 44784 7488 44790 7540
rect 44818 7488 44824 7540
rect 44876 7528 44882 7540
rect 45465 7531 45523 7537
rect 45465 7528 45477 7531
rect 44876 7500 45477 7528
rect 44876 7488 44882 7500
rect 45465 7497 45477 7500
rect 45511 7528 45523 7531
rect 45511 7500 46612 7528
rect 45511 7497 45523 7500
rect 45465 7491 45523 7497
rect 32769 7463 32827 7469
rect 32769 7460 32781 7463
rect 29932 7432 32781 7460
rect 32769 7429 32781 7432
rect 32815 7460 32827 7463
rect 35894 7460 35900 7472
rect 32815 7432 35900 7460
rect 32815 7429 32827 7432
rect 32769 7423 32827 7429
rect 35894 7420 35900 7432
rect 35952 7420 35958 7472
rect 38841 7463 38899 7469
rect 38841 7429 38853 7463
rect 38887 7460 38899 7463
rect 39666 7460 39672 7472
rect 38887 7432 39672 7460
rect 38887 7429 38899 7432
rect 38841 7423 38899 7429
rect 39666 7420 39672 7432
rect 39724 7420 39730 7472
rect 45554 7420 45560 7472
rect 45612 7460 45618 7472
rect 46474 7460 46480 7472
rect 45612 7432 46480 7460
rect 45612 7420 45618 7432
rect 46474 7420 46480 7432
rect 46532 7420 46538 7472
rect 46584 7460 46612 7500
rect 46658 7488 46664 7540
rect 46716 7528 46722 7540
rect 47213 7531 47271 7537
rect 47213 7528 47225 7531
rect 46716 7500 47225 7528
rect 46716 7488 46722 7500
rect 47213 7497 47225 7500
rect 47259 7497 47271 7531
rect 47213 7491 47271 7497
rect 47486 7488 47492 7540
rect 47544 7528 47550 7540
rect 47581 7531 47639 7537
rect 47581 7528 47593 7531
rect 47544 7500 47593 7528
rect 47544 7488 47550 7500
rect 47581 7497 47593 7500
rect 47627 7497 47639 7531
rect 47581 7491 47639 7497
rect 47670 7488 47676 7540
rect 47728 7528 47734 7540
rect 50617 7531 50675 7537
rect 50617 7528 50629 7531
rect 47728 7500 50629 7528
rect 47728 7488 47734 7500
rect 50617 7497 50629 7500
rect 50663 7528 50675 7531
rect 51626 7528 51632 7540
rect 50663 7500 51632 7528
rect 50663 7497 50675 7500
rect 50617 7491 50675 7497
rect 51626 7488 51632 7500
rect 51684 7488 51690 7540
rect 51994 7488 52000 7540
rect 52052 7528 52058 7540
rect 52641 7531 52699 7537
rect 52641 7528 52653 7531
rect 52052 7500 52653 7528
rect 52052 7488 52058 7500
rect 52641 7497 52653 7500
rect 52687 7497 52699 7531
rect 53742 7528 53748 7540
rect 53703 7500 53748 7528
rect 52641 7491 52699 7497
rect 52546 7460 52552 7472
rect 46584 7432 52552 7460
rect 52546 7420 52552 7432
rect 52604 7420 52610 7472
rect 17276 7364 24900 7392
rect 24949 7395 25007 7401
rect 17276 7352 17282 7364
rect 24949 7361 24961 7395
rect 24995 7392 25007 7395
rect 26513 7395 26571 7401
rect 26513 7392 26525 7395
rect 24995 7364 26525 7392
rect 24995 7361 25007 7364
rect 24949 7355 25007 7361
rect 26513 7361 26525 7364
rect 26559 7392 26571 7395
rect 28442 7392 28448 7404
rect 26559 7364 28448 7392
rect 26559 7361 26571 7364
rect 26513 7355 26571 7361
rect 28442 7352 28448 7364
rect 28500 7352 28506 7404
rect 28994 7352 29000 7404
rect 29052 7392 29058 7404
rect 31478 7392 31484 7404
rect 29052 7364 31484 7392
rect 29052 7352 29058 7364
rect 14001 7327 14059 7333
rect 14001 7293 14013 7327
rect 14047 7324 14059 7327
rect 14182 7324 14188 7336
rect 14047 7296 14188 7324
rect 14047 7293 14059 7296
rect 14001 7287 14059 7293
rect 14182 7284 14188 7296
rect 14240 7284 14246 7336
rect 14369 7327 14427 7333
rect 14369 7293 14381 7327
rect 14415 7324 14427 7327
rect 14458 7324 14464 7336
rect 14415 7296 14464 7324
rect 14415 7293 14427 7296
rect 14369 7287 14427 7293
rect 14458 7284 14464 7296
rect 14516 7324 14522 7336
rect 16298 7324 16304 7336
rect 14516 7296 16304 7324
rect 14516 7284 14522 7296
rect 16298 7284 16304 7296
rect 16356 7284 16362 7336
rect 16577 7327 16635 7333
rect 16577 7293 16589 7327
rect 16623 7293 16635 7327
rect 16577 7287 16635 7293
rect 16592 7256 16620 7287
rect 16666 7284 16672 7336
rect 16724 7324 16730 7336
rect 17678 7324 17684 7336
rect 16724 7296 17684 7324
rect 16724 7284 16730 7296
rect 17678 7284 17684 7296
rect 17736 7284 17742 7336
rect 18138 7284 18144 7336
rect 18196 7324 18202 7336
rect 18874 7324 18880 7336
rect 18196 7296 18880 7324
rect 18196 7284 18202 7296
rect 18874 7284 18880 7296
rect 18932 7324 18938 7336
rect 19429 7327 19487 7333
rect 19429 7324 19441 7327
rect 18932 7296 19441 7324
rect 18932 7284 18938 7296
rect 19429 7293 19441 7296
rect 19475 7293 19487 7327
rect 19429 7287 19487 7293
rect 19613 7327 19671 7333
rect 19613 7293 19625 7327
rect 19659 7324 19671 7327
rect 19702 7324 19708 7336
rect 19659 7296 19708 7324
rect 19659 7293 19671 7296
rect 19613 7287 19671 7293
rect 19702 7284 19708 7296
rect 19760 7284 19766 7336
rect 19981 7327 20039 7333
rect 19981 7293 19993 7327
rect 20027 7293 20039 7327
rect 19981 7287 20039 7293
rect 13188 7228 14228 7256
rect 12897 7219 12955 7225
rect 10008 7160 10824 7188
rect 10008 7148 10014 7160
rect 10870 7148 10876 7200
rect 10928 7188 10934 7200
rect 11882 7188 11888 7200
rect 10928 7160 11888 7188
rect 10928 7148 10934 7160
rect 11882 7148 11888 7160
rect 11940 7148 11946 7200
rect 12250 7188 12256 7200
rect 12211 7160 12256 7188
rect 12250 7148 12256 7160
rect 12308 7148 12314 7200
rect 14200 7188 14228 7228
rect 16040 7228 16620 7256
rect 16040 7188 16068 7228
rect 16206 7188 16212 7200
rect 14200 7160 16068 7188
rect 16167 7160 16212 7188
rect 16206 7148 16212 7160
rect 16264 7148 16270 7200
rect 16592 7188 16620 7228
rect 17494 7216 17500 7268
rect 17552 7256 17558 7268
rect 17865 7259 17923 7265
rect 17865 7256 17877 7259
rect 17552 7228 17877 7256
rect 17552 7216 17558 7228
rect 17865 7225 17877 7228
rect 17911 7256 17923 7259
rect 19518 7256 19524 7268
rect 17911 7228 19524 7256
rect 17911 7225 17923 7228
rect 17865 7219 17923 7225
rect 19518 7216 19524 7228
rect 19576 7216 19582 7268
rect 19996 7256 20024 7287
rect 20070 7284 20076 7336
rect 20128 7324 20134 7336
rect 20165 7327 20223 7333
rect 20165 7324 20177 7327
rect 20128 7296 20177 7324
rect 20128 7284 20134 7296
rect 20165 7293 20177 7296
rect 20211 7324 20223 7327
rect 20441 7327 20499 7333
rect 20441 7324 20453 7327
rect 20211 7296 20453 7324
rect 20211 7293 20223 7296
rect 20165 7287 20223 7293
rect 20441 7293 20453 7296
rect 20487 7293 20499 7327
rect 21174 7324 21180 7336
rect 21135 7296 21180 7324
rect 20441 7287 20499 7293
rect 21174 7284 21180 7296
rect 21232 7324 21238 7336
rect 21542 7324 21548 7336
rect 21232 7296 21548 7324
rect 21232 7284 21238 7296
rect 21542 7284 21548 7296
rect 21600 7324 21606 7336
rect 21821 7327 21879 7333
rect 21821 7324 21833 7327
rect 21600 7296 21833 7324
rect 21600 7284 21606 7296
rect 21821 7293 21833 7296
rect 21867 7293 21879 7327
rect 21821 7287 21879 7293
rect 22094 7284 22100 7336
rect 22152 7324 22158 7336
rect 22465 7327 22523 7333
rect 22465 7324 22477 7327
rect 22152 7296 22477 7324
rect 22152 7284 22158 7296
rect 22465 7293 22477 7296
rect 22511 7324 22523 7327
rect 23017 7327 23075 7333
rect 23017 7324 23029 7327
rect 22511 7296 23029 7324
rect 22511 7293 22523 7296
rect 22465 7287 22523 7293
rect 23017 7293 23029 7296
rect 23063 7324 23075 7327
rect 23842 7324 23848 7336
rect 23063 7296 23848 7324
rect 23063 7293 23075 7296
rect 23017 7287 23075 7293
rect 23842 7284 23848 7296
rect 23900 7284 23906 7336
rect 24302 7324 24308 7336
rect 24263 7296 24308 7324
rect 24302 7284 24308 7296
rect 24360 7284 24366 7336
rect 24397 7327 24455 7333
rect 24397 7293 24409 7327
rect 24443 7293 24455 7327
rect 24397 7287 24455 7293
rect 19996 7228 20208 7256
rect 17405 7191 17463 7197
rect 17405 7188 17417 7191
rect 16592 7160 17417 7188
rect 17405 7157 17417 7160
rect 17451 7188 17463 7191
rect 18598 7188 18604 7200
rect 17451 7160 18604 7188
rect 17451 7157 17463 7160
rect 17405 7151 17463 7157
rect 18598 7148 18604 7160
rect 18656 7148 18662 7200
rect 18782 7188 18788 7200
rect 18743 7160 18788 7188
rect 18782 7148 18788 7160
rect 18840 7148 18846 7200
rect 18874 7148 18880 7200
rect 18932 7188 18938 7200
rect 20070 7188 20076 7200
rect 18932 7160 20076 7188
rect 18932 7148 18938 7160
rect 20070 7148 20076 7160
rect 20128 7148 20134 7200
rect 20180 7188 20208 7228
rect 20254 7216 20260 7268
rect 20312 7256 20318 7268
rect 20993 7259 21051 7265
rect 20312 7228 20944 7256
rect 20312 7216 20318 7228
rect 20806 7188 20812 7200
rect 20180 7160 20812 7188
rect 20806 7148 20812 7160
rect 20864 7148 20870 7200
rect 20916 7188 20944 7228
rect 20993 7225 21005 7259
rect 21039 7256 21051 7259
rect 22189 7259 22247 7265
rect 22189 7256 22201 7259
rect 21039 7228 22201 7256
rect 21039 7225 21051 7228
rect 20993 7219 21051 7225
rect 22189 7225 22201 7228
rect 22235 7256 22247 7259
rect 22278 7256 22284 7268
rect 22235 7228 22284 7256
rect 22235 7225 22247 7228
rect 22189 7219 22247 7225
rect 22278 7216 22284 7228
rect 22336 7216 22342 7268
rect 24412 7256 24440 7287
rect 24486 7284 24492 7336
rect 24544 7324 24550 7336
rect 25314 7324 25320 7336
rect 24544 7296 24589 7324
rect 24688 7296 25320 7324
rect 24544 7284 24550 7296
rect 24688 7256 24716 7296
rect 25314 7284 25320 7296
rect 25372 7284 25378 7336
rect 25958 7284 25964 7336
rect 26016 7324 26022 7336
rect 26421 7327 26479 7333
rect 26421 7324 26433 7327
rect 26016 7296 26433 7324
rect 26016 7284 26022 7296
rect 26421 7293 26433 7296
rect 26467 7293 26479 7327
rect 26421 7287 26479 7293
rect 26789 7327 26847 7333
rect 26789 7293 26801 7327
rect 26835 7293 26847 7327
rect 26789 7287 26847 7293
rect 24412 7228 24716 7256
rect 26234 7216 26240 7268
rect 26292 7256 26298 7268
rect 26804 7256 26832 7287
rect 26878 7284 26884 7336
rect 26936 7324 26942 7336
rect 26936 7296 26981 7324
rect 26936 7284 26942 7296
rect 27154 7284 27160 7336
rect 27212 7324 27218 7336
rect 27617 7327 27675 7333
rect 27617 7324 27629 7327
rect 27212 7296 27629 7324
rect 27212 7284 27218 7296
rect 27617 7293 27629 7296
rect 27663 7293 27675 7327
rect 27617 7287 27675 7293
rect 27890 7284 27896 7336
rect 27948 7324 27954 7336
rect 27985 7327 28043 7333
rect 27985 7324 27997 7327
rect 27948 7296 27997 7324
rect 27948 7284 27954 7296
rect 27985 7293 27997 7296
rect 28031 7293 28043 7327
rect 27985 7287 28043 7293
rect 28074 7284 28080 7336
rect 28132 7324 28138 7336
rect 29472 7333 29500 7364
rect 31478 7352 31484 7364
rect 31536 7352 31542 7404
rect 32030 7352 32036 7404
rect 32088 7392 32094 7404
rect 32088 7364 33640 7392
rect 32088 7352 32094 7364
rect 29457 7327 29515 7333
rect 28132 7296 29408 7324
rect 28132 7284 28138 7296
rect 26292 7228 26832 7256
rect 26292 7216 26298 7228
rect 27062 7216 27068 7268
rect 27120 7256 27126 7268
rect 27120 7228 27752 7256
rect 27120 7216 27126 7228
rect 21269 7191 21327 7197
rect 21269 7188 21281 7191
rect 20916 7160 21281 7188
rect 21269 7157 21281 7160
rect 21315 7157 21327 7191
rect 21269 7151 21327 7157
rect 22649 7191 22707 7197
rect 22649 7157 22661 7191
rect 22695 7188 22707 7191
rect 23106 7188 23112 7200
rect 22695 7160 23112 7188
rect 22695 7157 22707 7160
rect 22649 7151 22707 7157
rect 23106 7148 23112 7160
rect 23164 7148 23170 7200
rect 23934 7188 23940 7200
rect 23847 7160 23940 7188
rect 23934 7148 23940 7160
rect 23992 7188 23998 7200
rect 25041 7191 25099 7197
rect 25041 7188 25053 7191
rect 23992 7160 25053 7188
rect 23992 7148 23998 7160
rect 25041 7157 25053 7160
rect 25087 7157 25099 7191
rect 25314 7188 25320 7200
rect 25275 7160 25320 7188
rect 25041 7151 25099 7157
rect 25314 7148 25320 7160
rect 25372 7148 25378 7200
rect 25685 7191 25743 7197
rect 25685 7157 25697 7191
rect 25731 7188 25743 7191
rect 25958 7188 25964 7200
rect 25731 7160 25964 7188
rect 25731 7157 25743 7160
rect 25685 7151 25743 7157
rect 25958 7148 25964 7160
rect 26016 7148 26022 7200
rect 27724 7188 27752 7228
rect 27798 7216 27804 7268
rect 27856 7256 27862 7268
rect 28445 7259 28503 7265
rect 28445 7256 28457 7259
rect 27856 7228 28457 7256
rect 27856 7216 27862 7228
rect 28445 7225 28457 7228
rect 28491 7225 28503 7259
rect 29270 7256 29276 7268
rect 29231 7228 29276 7256
rect 28445 7219 28503 7225
rect 29270 7216 29276 7228
rect 29328 7216 29334 7268
rect 28077 7191 28135 7197
rect 28077 7188 28089 7191
rect 27724 7160 28089 7188
rect 28077 7157 28089 7160
rect 28123 7157 28135 7191
rect 28077 7151 28135 7157
rect 28258 7148 28264 7200
rect 28316 7188 28322 7200
rect 28997 7191 29055 7197
rect 28997 7188 29009 7191
rect 28316 7160 29009 7188
rect 28316 7148 28322 7160
rect 28997 7157 29009 7160
rect 29043 7157 29055 7191
rect 29380 7188 29408 7296
rect 29457 7293 29469 7327
rect 29503 7293 29515 7327
rect 30285 7327 30343 7333
rect 30285 7324 30297 7327
rect 29457 7287 29515 7293
rect 29656 7296 30297 7324
rect 29546 7256 29552 7268
rect 29507 7228 29552 7256
rect 29546 7216 29552 7228
rect 29604 7216 29610 7268
rect 29656 7265 29684 7296
rect 30285 7293 30297 7296
rect 30331 7293 30343 7327
rect 30285 7287 30343 7293
rect 30742 7284 30748 7336
rect 30800 7324 30806 7336
rect 30837 7327 30895 7333
rect 30837 7324 30849 7327
rect 30800 7296 30849 7324
rect 30800 7284 30806 7296
rect 30837 7293 30849 7296
rect 30883 7324 30895 7327
rect 31294 7324 31300 7336
rect 30883 7296 31300 7324
rect 30883 7293 30895 7296
rect 30837 7287 30895 7293
rect 31294 7284 31300 7296
rect 31352 7324 31358 7336
rect 33612 7333 33640 7364
rect 33778 7352 33784 7404
rect 33836 7392 33842 7404
rect 34241 7395 34299 7401
rect 34241 7392 34253 7395
rect 33836 7364 34253 7392
rect 33836 7352 33842 7364
rect 34241 7361 34253 7364
rect 34287 7361 34299 7395
rect 34698 7392 34704 7404
rect 34659 7364 34704 7392
rect 34241 7355 34299 7361
rect 34698 7352 34704 7364
rect 34756 7352 34762 7404
rect 35713 7395 35771 7401
rect 35713 7392 35725 7395
rect 34900 7364 35725 7392
rect 31389 7327 31447 7333
rect 31389 7324 31401 7327
rect 31352 7296 31401 7324
rect 31352 7284 31358 7296
rect 31389 7293 31401 7296
rect 31435 7293 31447 7327
rect 31389 7287 31447 7293
rect 32585 7327 32643 7333
rect 32585 7293 32597 7327
rect 32631 7324 32643 7327
rect 33597 7327 33655 7333
rect 32631 7296 33272 7324
rect 32631 7293 32643 7296
rect 32585 7287 32643 7293
rect 29641 7259 29699 7265
rect 29641 7225 29653 7259
rect 29687 7225 29699 7259
rect 30006 7256 30012 7268
rect 29967 7228 30012 7256
rect 29641 7219 29699 7225
rect 29656 7188 29684 7219
rect 30006 7216 30012 7228
rect 30064 7216 30070 7268
rect 29380 7160 29684 7188
rect 28997 7151 29055 7157
rect 30650 7148 30656 7200
rect 30708 7188 30714 7200
rect 31754 7188 31760 7200
rect 30708 7160 31760 7188
rect 30708 7148 30714 7160
rect 31754 7148 31760 7160
rect 31812 7148 31818 7200
rect 32398 7188 32404 7200
rect 32359 7160 32404 7188
rect 32398 7148 32404 7160
rect 32456 7148 32462 7200
rect 33244 7197 33272 7296
rect 33597 7293 33609 7327
rect 33643 7324 33655 7327
rect 33689 7327 33747 7333
rect 33689 7324 33701 7327
rect 33643 7296 33701 7324
rect 33643 7293 33655 7296
rect 33597 7287 33655 7293
rect 33689 7293 33701 7296
rect 33735 7293 33747 7327
rect 33689 7287 33747 7293
rect 33704 7256 33732 7287
rect 34606 7284 34612 7336
rect 34664 7324 34670 7336
rect 34900 7333 34928 7364
rect 35713 7361 35725 7364
rect 35759 7361 35771 7395
rect 35912 7392 35940 7420
rect 43993 7395 44051 7401
rect 35912 7364 37044 7392
rect 35713 7355 35771 7361
rect 34885 7327 34943 7333
rect 34885 7324 34897 7327
rect 34664 7296 34897 7324
rect 34664 7284 34670 7296
rect 34885 7293 34897 7296
rect 34931 7293 34943 7327
rect 34885 7287 34943 7293
rect 34974 7284 34980 7336
rect 35032 7324 35038 7336
rect 37016 7333 37044 7364
rect 39040 7364 43392 7392
rect 39040 7333 39068 7364
rect 36817 7327 36875 7333
rect 35032 7296 35077 7324
rect 35032 7284 35038 7296
rect 36817 7293 36829 7327
rect 36863 7293 36875 7327
rect 36817 7287 36875 7293
rect 37001 7327 37059 7333
rect 37001 7293 37013 7327
rect 37047 7293 37059 7327
rect 37001 7287 37059 7293
rect 37369 7327 37427 7333
rect 37369 7293 37381 7327
rect 37415 7293 37427 7327
rect 37369 7287 37427 7293
rect 38473 7327 38531 7333
rect 38473 7293 38485 7327
rect 38519 7324 38531 7327
rect 39025 7327 39083 7333
rect 39025 7324 39037 7327
rect 38519 7296 39037 7324
rect 38519 7293 38531 7296
rect 38473 7287 38531 7293
rect 39025 7293 39037 7296
rect 39071 7293 39083 7327
rect 39206 7324 39212 7336
rect 39167 7296 39212 7324
rect 39025 7287 39083 7293
rect 34992 7256 35020 7284
rect 33704 7228 35020 7256
rect 33229 7191 33287 7197
rect 33229 7157 33241 7191
rect 33275 7188 33287 7191
rect 33502 7188 33508 7200
rect 33275 7160 33508 7188
rect 33275 7157 33287 7160
rect 33229 7151 33287 7157
rect 33502 7148 33508 7160
rect 33560 7148 33566 7200
rect 35986 7148 35992 7200
rect 36044 7188 36050 7200
rect 36081 7191 36139 7197
rect 36081 7188 36093 7191
rect 36044 7160 36093 7188
rect 36044 7148 36050 7160
rect 36081 7157 36093 7160
rect 36127 7157 36139 7191
rect 36630 7188 36636 7200
rect 36591 7160 36636 7188
rect 36081 7151 36139 7157
rect 36630 7148 36636 7160
rect 36688 7148 36694 7200
rect 36832 7188 36860 7287
rect 37384 7256 37412 7287
rect 39206 7284 39212 7296
rect 39264 7284 39270 7336
rect 39390 7324 39396 7336
rect 39351 7296 39396 7324
rect 39390 7284 39396 7296
rect 39448 7324 39454 7336
rect 40221 7327 40279 7333
rect 40221 7324 40233 7327
rect 39448 7296 40233 7324
rect 39448 7284 39454 7296
rect 40221 7293 40233 7296
rect 40267 7293 40279 7327
rect 40221 7287 40279 7293
rect 40402 7284 40408 7336
rect 40460 7324 40466 7336
rect 40681 7327 40739 7333
rect 40681 7324 40693 7327
rect 40460 7296 40693 7324
rect 40460 7284 40466 7296
rect 40681 7293 40693 7296
rect 40727 7324 40739 7327
rect 41325 7327 41383 7333
rect 41325 7324 41337 7327
rect 40727 7296 41337 7324
rect 40727 7293 40739 7296
rect 40681 7287 40739 7293
rect 41325 7293 41337 7296
rect 41371 7293 41383 7327
rect 42334 7324 42340 7336
rect 42247 7296 42340 7324
rect 41325 7287 41383 7293
rect 42334 7284 42340 7296
rect 42392 7284 42398 7336
rect 42426 7284 42432 7336
rect 42484 7324 42490 7336
rect 42613 7327 42671 7333
rect 42613 7324 42625 7327
rect 42484 7296 42625 7324
rect 42484 7284 42490 7296
rect 42613 7293 42625 7296
rect 42659 7293 42671 7327
rect 42613 7287 42671 7293
rect 38013 7259 38071 7265
rect 38013 7256 38025 7259
rect 37384 7228 38025 7256
rect 38013 7225 38025 7228
rect 38059 7256 38071 7259
rect 38378 7256 38384 7268
rect 38059 7228 38384 7256
rect 38059 7225 38071 7228
rect 38013 7219 38071 7225
rect 38378 7216 38384 7228
rect 38436 7256 38442 7268
rect 39224 7256 39252 7284
rect 38436 7228 39252 7256
rect 38436 7216 38442 7228
rect 39758 7216 39764 7268
rect 39816 7256 39822 7268
rect 40497 7259 40555 7265
rect 40497 7256 40509 7259
rect 39816 7228 40509 7256
rect 39816 7216 39822 7228
rect 40497 7225 40509 7228
rect 40543 7225 40555 7259
rect 41046 7256 41052 7268
rect 41007 7228 41052 7256
rect 40497 7219 40555 7225
rect 41046 7216 41052 7228
rect 41104 7216 41110 7268
rect 42352 7256 42380 7284
rect 43364 7268 43392 7364
rect 43993 7361 44005 7395
rect 44039 7392 44051 7395
rect 44361 7395 44419 7401
rect 44361 7392 44373 7395
rect 44039 7364 44373 7392
rect 44039 7361 44051 7364
rect 43993 7355 44051 7361
rect 44361 7361 44373 7364
rect 44407 7392 44419 7395
rect 46106 7392 46112 7404
rect 44407 7364 46112 7392
rect 44407 7361 44419 7364
rect 44361 7355 44419 7361
rect 44836 7333 44864 7364
rect 46106 7352 46112 7364
rect 46164 7392 46170 7404
rect 46348 7395 46406 7401
rect 46348 7392 46360 7395
rect 46164 7364 46360 7392
rect 46164 7352 46170 7364
rect 46348 7361 46360 7364
rect 46394 7361 46406 7395
rect 46348 7355 46406 7361
rect 46569 7395 46627 7401
rect 46569 7361 46581 7395
rect 46615 7361 46627 7395
rect 46569 7355 46627 7361
rect 44821 7327 44879 7333
rect 44821 7293 44833 7327
rect 44867 7293 44879 7327
rect 46474 7324 46480 7336
rect 44821 7287 44879 7293
rect 45756 7296 46480 7324
rect 41248 7228 42380 7256
rect 37274 7188 37280 7200
rect 36832 7160 37280 7188
rect 37274 7148 37280 7160
rect 37332 7148 37338 7200
rect 38654 7148 38660 7200
rect 38712 7188 38718 7200
rect 39114 7188 39120 7200
rect 38712 7160 39120 7188
rect 38712 7148 38718 7160
rect 39114 7148 39120 7160
rect 39172 7188 39178 7200
rect 39853 7191 39911 7197
rect 39853 7188 39865 7191
rect 39172 7160 39865 7188
rect 39172 7148 39178 7160
rect 39853 7157 39865 7160
rect 39899 7157 39911 7191
rect 39853 7151 39911 7157
rect 40586 7148 40592 7200
rect 40644 7188 40650 7200
rect 41248 7188 41276 7228
rect 43346 7216 43352 7268
rect 43404 7256 43410 7268
rect 43404 7228 45140 7256
rect 43404 7216 43410 7228
rect 40644 7160 41276 7188
rect 40644 7148 40650 7160
rect 41322 7148 41328 7200
rect 41380 7188 41386 7200
rect 44450 7188 44456 7200
rect 41380 7160 44456 7188
rect 41380 7148 41386 7160
rect 44450 7148 44456 7160
rect 44508 7148 44514 7200
rect 44726 7148 44732 7200
rect 44784 7188 44790 7200
rect 45005 7191 45063 7197
rect 45005 7188 45017 7191
rect 44784 7160 45017 7188
rect 44784 7148 44790 7160
rect 45005 7157 45017 7160
rect 45051 7157 45063 7191
rect 45112 7188 45140 7228
rect 45186 7216 45192 7268
rect 45244 7256 45250 7268
rect 45756 7265 45784 7296
rect 46474 7284 46480 7296
rect 46532 7284 46538 7336
rect 45741 7259 45799 7265
rect 45741 7256 45753 7259
rect 45244 7228 45753 7256
rect 45244 7216 45250 7228
rect 45741 7225 45753 7228
rect 45787 7225 45799 7259
rect 46198 7256 46204 7268
rect 46159 7228 46204 7256
rect 45741 7219 45799 7225
rect 46198 7216 46204 7228
rect 46256 7216 46262 7268
rect 46290 7216 46296 7268
rect 46348 7256 46354 7268
rect 46584 7256 46612 7355
rect 48682 7352 48688 7404
rect 48740 7392 48746 7404
rect 49602 7392 49608 7404
rect 48740 7364 49608 7392
rect 48740 7352 48746 7364
rect 49602 7352 49608 7364
rect 49660 7392 49666 7404
rect 49881 7395 49939 7401
rect 49881 7392 49893 7395
rect 49660 7364 49893 7392
rect 49660 7352 49666 7364
rect 49881 7361 49893 7364
rect 49927 7361 49939 7395
rect 49881 7355 49939 7361
rect 50154 7352 50160 7404
rect 50212 7392 50218 7404
rect 51902 7392 51908 7404
rect 50212 7364 51908 7392
rect 50212 7352 50218 7364
rect 51902 7352 51908 7364
rect 51960 7392 51966 7404
rect 52273 7395 52331 7401
rect 52273 7392 52285 7395
rect 51960 7364 52285 7392
rect 51960 7352 51966 7364
rect 52273 7361 52285 7364
rect 52319 7361 52331 7395
rect 52273 7355 52331 7361
rect 46658 7284 46664 7336
rect 46716 7324 46722 7336
rect 49973 7327 50031 7333
rect 46716 7296 48912 7324
rect 46716 7284 46722 7296
rect 46934 7256 46940 7268
rect 46348 7228 46612 7256
rect 46895 7228 46940 7256
rect 46348 7216 46354 7228
rect 46934 7216 46940 7228
rect 46992 7216 46998 7268
rect 47670 7256 47676 7268
rect 47044 7228 47676 7256
rect 47044 7188 47072 7228
rect 47670 7216 47676 7228
rect 47728 7216 47734 7268
rect 47765 7259 47823 7265
rect 47765 7225 47777 7259
rect 47811 7225 47823 7259
rect 47946 7256 47952 7268
rect 47907 7228 47952 7256
rect 47765 7219 47823 7225
rect 45112 7160 47072 7188
rect 45005 7151 45063 7157
rect 47210 7148 47216 7200
rect 47268 7188 47274 7200
rect 47780 7188 47808 7219
rect 47946 7216 47952 7228
rect 48004 7216 48010 7268
rect 48130 7256 48136 7268
rect 48091 7228 48136 7256
rect 48130 7216 48136 7228
rect 48188 7216 48194 7268
rect 48498 7256 48504 7268
rect 48459 7228 48504 7256
rect 48498 7216 48504 7228
rect 48556 7216 48562 7268
rect 48774 7256 48780 7268
rect 48735 7228 48780 7256
rect 48774 7216 48780 7228
rect 48832 7216 48838 7268
rect 47268 7160 47808 7188
rect 48041 7191 48099 7197
rect 47268 7148 47274 7160
rect 48041 7157 48053 7191
rect 48087 7188 48099 7191
rect 48590 7188 48596 7200
rect 48087 7160 48596 7188
rect 48087 7157 48099 7160
rect 48041 7151 48099 7157
rect 48590 7148 48596 7160
rect 48648 7148 48654 7200
rect 48884 7188 48912 7296
rect 49973 7293 49985 7327
rect 50019 7324 50031 7327
rect 50062 7324 50068 7336
rect 50019 7296 50068 7324
rect 50019 7293 50031 7296
rect 49973 7287 50031 7293
rect 50062 7284 50068 7296
rect 50120 7284 50126 7336
rect 50338 7324 50344 7336
rect 50299 7296 50344 7324
rect 50338 7284 50344 7296
rect 50396 7284 50402 7336
rect 50525 7327 50583 7333
rect 50525 7293 50537 7327
rect 50571 7324 50583 7327
rect 50617 7327 50675 7333
rect 50617 7324 50629 7327
rect 50571 7296 50629 7324
rect 50571 7293 50583 7296
rect 50525 7287 50583 7293
rect 50617 7293 50629 7296
rect 50663 7293 50675 7327
rect 50617 7287 50675 7293
rect 50982 7284 50988 7336
rect 51040 7324 51046 7336
rect 51721 7327 51779 7333
rect 51721 7324 51733 7327
rect 51040 7296 51733 7324
rect 51040 7284 51046 7296
rect 51721 7293 51733 7296
rect 51767 7293 51779 7327
rect 52656 7324 52684 7491
rect 53742 7488 53748 7500
rect 53800 7488 53806 7540
rect 55217 7531 55275 7537
rect 55217 7497 55229 7531
rect 55263 7528 55275 7531
rect 55398 7528 55404 7540
rect 55263 7500 55404 7528
rect 55263 7497 55275 7500
rect 55217 7491 55275 7497
rect 55398 7488 55404 7500
rect 55456 7488 55462 7540
rect 56134 7488 56140 7540
rect 56192 7528 56198 7540
rect 56689 7531 56747 7537
rect 56689 7528 56701 7531
rect 56192 7500 56701 7528
rect 56192 7488 56198 7500
rect 56689 7497 56701 7500
rect 56735 7497 56747 7531
rect 57054 7528 57060 7540
rect 57015 7500 57060 7528
rect 56689 7491 56747 7497
rect 57054 7488 57060 7500
rect 57112 7488 57118 7540
rect 59906 7528 59912 7540
rect 57532 7500 59912 7528
rect 53006 7460 53012 7472
rect 52967 7432 53012 7460
rect 53006 7420 53012 7432
rect 53064 7460 53070 7472
rect 57532 7460 57560 7500
rect 59906 7488 59912 7500
rect 59964 7488 59970 7540
rect 60918 7488 60924 7540
rect 60976 7528 60982 7540
rect 61013 7531 61071 7537
rect 61013 7528 61025 7531
rect 60976 7500 61025 7528
rect 60976 7488 60982 7500
rect 61013 7497 61025 7500
rect 61059 7497 61071 7531
rect 61013 7491 61071 7497
rect 53064 7432 57560 7460
rect 53064 7420 53070 7432
rect 57606 7420 57612 7472
rect 57664 7420 57670 7472
rect 57698 7420 57704 7472
rect 57756 7460 57762 7472
rect 59725 7463 59783 7469
rect 59725 7460 59737 7463
rect 57756 7432 59737 7460
rect 57756 7420 57762 7432
rect 59725 7429 59737 7432
rect 59771 7429 59783 7463
rect 59725 7423 59783 7429
rect 56045 7395 56103 7401
rect 56045 7361 56057 7395
rect 56091 7392 56103 7395
rect 56318 7392 56324 7404
rect 56091 7364 56324 7392
rect 56091 7361 56103 7364
rect 56045 7355 56103 7361
rect 56318 7352 56324 7364
rect 56376 7352 56382 7404
rect 57517 7395 57575 7401
rect 57517 7361 57529 7395
rect 57563 7392 57575 7395
rect 57624 7392 57652 7420
rect 57563 7364 57652 7392
rect 57563 7361 57575 7364
rect 57517 7355 57575 7361
rect 52825 7327 52883 7333
rect 52825 7324 52837 7327
rect 52656 7296 52837 7324
rect 51721 7287 51779 7293
rect 52825 7293 52837 7296
rect 52871 7324 52883 7327
rect 53377 7327 53435 7333
rect 53377 7324 53389 7327
rect 52871 7296 53389 7324
rect 52871 7293 52883 7296
rect 52825 7287 52883 7293
rect 53377 7293 53389 7296
rect 53423 7293 53435 7327
rect 53377 7287 53435 7293
rect 53929 7327 53987 7333
rect 53929 7293 53941 7327
rect 53975 7293 53987 7327
rect 53929 7287 53987 7293
rect 55585 7327 55643 7333
rect 55585 7293 55597 7327
rect 55631 7324 55643 7327
rect 55766 7324 55772 7336
rect 55631 7296 55772 7324
rect 55631 7293 55643 7296
rect 55585 7287 55643 7293
rect 49142 7256 49148 7268
rect 49103 7228 49148 7256
rect 49142 7216 49148 7228
rect 49200 7216 49206 7268
rect 49329 7259 49387 7265
rect 49329 7225 49341 7259
rect 49375 7256 49387 7259
rect 49878 7256 49884 7268
rect 49375 7228 49884 7256
rect 49375 7225 49387 7228
rect 49329 7219 49387 7225
rect 49878 7216 49884 7228
rect 49936 7216 49942 7268
rect 50356 7256 50384 7284
rect 50801 7259 50859 7265
rect 50801 7256 50813 7259
rect 50356 7228 50813 7256
rect 50801 7225 50813 7228
rect 50847 7256 50859 7259
rect 50847 7228 51948 7256
rect 50847 7225 50859 7228
rect 50801 7219 50859 7225
rect 50706 7188 50712 7200
rect 48884 7160 50712 7188
rect 50706 7148 50712 7160
rect 50764 7148 50770 7200
rect 51261 7191 51319 7197
rect 51261 7157 51273 7191
rect 51307 7188 51319 7191
rect 51626 7188 51632 7200
rect 51307 7160 51632 7188
rect 51307 7157 51319 7160
rect 51261 7151 51319 7157
rect 51626 7148 51632 7160
rect 51684 7148 51690 7200
rect 51920 7197 51948 7228
rect 52730 7216 52736 7268
rect 52788 7256 52794 7268
rect 53944 7256 53972 7287
rect 55766 7284 55772 7296
rect 55824 7284 55830 7336
rect 55858 7284 55864 7336
rect 55916 7324 55922 7336
rect 56229 7327 56287 7333
rect 56229 7324 56241 7327
rect 55916 7296 56241 7324
rect 55916 7284 55922 7296
rect 56229 7293 56241 7296
rect 56275 7293 56287 7327
rect 56229 7287 56287 7293
rect 57054 7284 57060 7336
rect 57112 7324 57118 7336
rect 57609 7327 57667 7333
rect 57609 7324 57621 7327
rect 57112 7296 57621 7324
rect 57112 7284 57118 7296
rect 57609 7293 57621 7296
rect 57655 7324 57667 7327
rect 57790 7324 57796 7336
rect 57655 7296 57796 7324
rect 57655 7293 57667 7296
rect 57609 7287 57667 7293
rect 57790 7284 57796 7296
rect 57848 7284 57854 7336
rect 58066 7324 58072 7336
rect 58027 7296 58072 7324
rect 58066 7284 58072 7296
rect 58124 7284 58130 7336
rect 58161 7327 58219 7333
rect 58161 7293 58173 7327
rect 58207 7324 58219 7327
rect 59449 7327 59507 7333
rect 59449 7324 59461 7327
rect 58207 7296 59461 7324
rect 58207 7293 58219 7296
rect 58161 7287 58219 7293
rect 59449 7293 59461 7296
rect 59495 7293 59507 7327
rect 59630 7324 59636 7336
rect 59591 7296 59636 7324
rect 59449 7287 59507 7293
rect 54481 7259 54539 7265
rect 54481 7256 54493 7259
rect 52788 7228 54493 7256
rect 52788 7216 52794 7228
rect 54481 7225 54493 7228
rect 54527 7225 54539 7259
rect 54481 7219 54539 7225
rect 57974 7216 57980 7268
rect 58032 7256 58038 7268
rect 58176 7256 58204 7287
rect 59630 7284 59636 7296
rect 59688 7284 59694 7336
rect 59814 7284 59820 7336
rect 59872 7324 59878 7336
rect 60185 7327 60243 7333
rect 60185 7324 60197 7327
rect 59872 7296 60197 7324
rect 59872 7284 59878 7296
rect 60185 7293 60197 7296
rect 60231 7324 60243 7327
rect 60645 7327 60703 7333
rect 60645 7324 60657 7327
rect 60231 7296 60657 7324
rect 60231 7293 60243 7296
rect 60185 7287 60243 7293
rect 60645 7293 60657 7296
rect 60691 7293 60703 7327
rect 60645 7287 60703 7293
rect 58710 7256 58716 7268
rect 58032 7228 58204 7256
rect 58671 7228 58716 7256
rect 58032 7216 58038 7228
rect 58710 7216 58716 7228
rect 58768 7216 58774 7268
rect 51905 7191 51963 7197
rect 51905 7157 51917 7191
rect 51951 7157 51963 7191
rect 51905 7151 51963 7157
rect 52178 7148 52184 7200
rect 52236 7188 52242 7200
rect 53558 7188 53564 7200
rect 52236 7160 53564 7188
rect 52236 7148 52242 7160
rect 53558 7148 53564 7160
rect 53616 7148 53622 7200
rect 54110 7188 54116 7200
rect 54023 7160 54116 7188
rect 54110 7148 54116 7160
rect 54168 7188 54174 7200
rect 56594 7188 56600 7200
rect 54168 7160 56600 7188
rect 54168 7148 54174 7160
rect 56594 7148 56600 7160
rect 56652 7148 56658 7200
rect 58066 7148 58072 7200
rect 58124 7188 58130 7200
rect 59081 7191 59139 7197
rect 59081 7188 59093 7191
rect 58124 7160 59093 7188
rect 58124 7148 58130 7160
rect 59081 7157 59093 7160
rect 59127 7157 59139 7191
rect 59081 7151 59139 7157
rect 1104 7098 63480 7120
rect 1104 7046 21774 7098
rect 21826 7046 21838 7098
rect 21890 7046 21902 7098
rect 21954 7046 21966 7098
rect 22018 7046 42566 7098
rect 42618 7046 42630 7098
rect 42682 7046 42694 7098
rect 42746 7046 42758 7098
rect 42810 7046 63480 7098
rect 1104 7024 63480 7046
rect 6457 6987 6515 6993
rect 6457 6953 6469 6987
rect 6503 6984 6515 6987
rect 6825 6987 6883 6993
rect 6825 6984 6837 6987
rect 6503 6956 6837 6984
rect 6503 6953 6515 6956
rect 6457 6947 6515 6953
rect 6825 6953 6837 6956
rect 6871 6984 6883 6987
rect 7282 6984 7288 6996
rect 6871 6956 7288 6984
rect 6871 6953 6883 6956
rect 6825 6947 6883 6953
rect 7282 6944 7288 6956
rect 7340 6944 7346 6996
rect 7926 6984 7932 6996
rect 7887 6956 7932 6984
rect 7926 6944 7932 6956
rect 7984 6944 7990 6996
rect 9950 6984 9956 6996
rect 9911 6956 9956 6984
rect 9950 6944 9956 6956
rect 10008 6944 10014 6996
rect 12250 6944 12256 6996
rect 12308 6984 12314 6996
rect 12345 6987 12403 6993
rect 12345 6984 12357 6987
rect 12308 6956 12357 6984
rect 12308 6944 12314 6956
rect 12345 6953 12357 6956
rect 12391 6984 12403 6987
rect 12713 6987 12771 6993
rect 12713 6984 12725 6987
rect 12391 6956 12725 6984
rect 12391 6953 12403 6956
rect 12345 6947 12403 6953
rect 12713 6953 12725 6956
rect 12759 6984 12771 6987
rect 13630 6984 13636 6996
rect 12759 6956 13636 6984
rect 12759 6953 12771 6956
rect 12713 6947 12771 6953
rect 13630 6944 13636 6956
rect 13688 6944 13694 6996
rect 17589 6987 17647 6993
rect 17589 6953 17601 6987
rect 17635 6984 17647 6987
rect 17865 6987 17923 6993
rect 17865 6984 17877 6987
rect 17635 6956 17877 6984
rect 17635 6953 17647 6956
rect 17589 6947 17647 6953
rect 17865 6953 17877 6956
rect 17911 6984 17923 6987
rect 18506 6984 18512 6996
rect 17911 6956 18512 6984
rect 17911 6953 17923 6956
rect 17865 6947 17923 6953
rect 18506 6944 18512 6956
rect 18564 6944 18570 6996
rect 18598 6944 18604 6996
rect 18656 6984 18662 6996
rect 20714 6984 20720 6996
rect 18656 6956 20720 6984
rect 18656 6944 18662 6956
rect 20714 6944 20720 6956
rect 20772 6944 20778 6996
rect 21266 6984 21272 6996
rect 20916 6956 21272 6984
rect 5721 6919 5779 6925
rect 5721 6885 5733 6919
rect 5767 6916 5779 6919
rect 6089 6919 6147 6925
rect 6089 6916 6101 6919
rect 5767 6888 6101 6916
rect 5767 6885 5779 6888
rect 5721 6879 5779 6885
rect 6089 6885 6101 6888
rect 6135 6916 6147 6919
rect 6546 6916 6552 6928
rect 6135 6888 6552 6916
rect 6135 6885 6147 6888
rect 6089 6879 6147 6885
rect 6546 6876 6552 6888
rect 6604 6876 6610 6928
rect 6730 6916 6736 6928
rect 6691 6888 6736 6916
rect 6730 6876 6736 6888
rect 6788 6876 6794 6928
rect 6914 6916 6920 6928
rect 6827 6888 6920 6916
rect 6914 6876 6920 6888
rect 6972 6916 6978 6928
rect 7944 6916 7972 6944
rect 6972 6888 7972 6916
rect 8128 6888 8432 6916
rect 6972 6876 6978 6888
rect 7285 6851 7343 6857
rect 7285 6817 7297 6851
rect 7331 6848 7343 6851
rect 8128 6848 8156 6888
rect 7331 6820 8156 6848
rect 7331 6817 7343 6820
rect 7285 6811 7343 6817
rect 8202 6808 8208 6860
rect 8260 6848 8266 6860
rect 8404 6848 8432 6888
rect 12526 6876 12532 6928
rect 12584 6916 12590 6928
rect 13173 6919 13231 6925
rect 13173 6916 13185 6919
rect 12584 6888 13185 6916
rect 12584 6876 12590 6888
rect 13173 6885 13185 6888
rect 13219 6885 13231 6919
rect 14734 6916 14740 6928
rect 13173 6879 13231 6885
rect 13648 6888 14740 6916
rect 9493 6851 9551 6857
rect 8260 6820 8305 6848
rect 8404 6820 9444 6848
rect 8260 6808 8266 6820
rect 3694 6780 3700 6792
rect 3252 6752 3700 6780
rect 3252 6656 3280 6752
rect 3694 6740 3700 6752
rect 3752 6780 3758 6792
rect 4065 6783 4123 6789
rect 4065 6780 4077 6783
rect 3752 6752 4077 6780
rect 3752 6740 3758 6752
rect 4065 6749 4077 6752
rect 4111 6749 4123 6783
rect 4065 6743 4123 6749
rect 4341 6783 4399 6789
rect 4341 6749 4353 6783
rect 4387 6780 4399 6783
rect 4798 6780 4804 6792
rect 4387 6752 4804 6780
rect 4387 6749 4399 6752
rect 4341 6743 4399 6749
rect 4798 6740 4804 6752
rect 4856 6740 4862 6792
rect 8113 6783 8171 6789
rect 8113 6749 8125 6783
rect 8159 6780 8171 6783
rect 8294 6780 8300 6792
rect 8159 6752 8300 6780
rect 8159 6749 8171 6752
rect 8113 6743 8171 6749
rect 8294 6740 8300 6752
rect 8352 6740 8358 6792
rect 8665 6783 8723 6789
rect 8665 6749 8677 6783
rect 8711 6749 8723 6783
rect 8665 6743 8723 6749
rect 7190 6672 7196 6724
rect 7248 6712 7254 6724
rect 8680 6712 8708 6743
rect 7248 6684 8708 6712
rect 7248 6672 7254 6684
rect 3234 6644 3240 6656
rect 3195 6616 3240 6644
rect 3234 6604 3240 6616
rect 3292 6604 3298 6656
rect 3510 6644 3516 6656
rect 3471 6616 3516 6644
rect 3510 6604 3516 6616
rect 3568 6604 3574 6656
rect 8202 6604 8208 6656
rect 8260 6644 8266 6656
rect 8941 6647 8999 6653
rect 8941 6644 8953 6647
rect 8260 6616 8953 6644
rect 8260 6604 8266 6616
rect 8941 6613 8953 6616
rect 8987 6613 8999 6647
rect 9416 6644 9444 6820
rect 9493 6817 9505 6851
rect 9539 6848 9551 6851
rect 12986 6848 12992 6860
rect 9539 6820 12992 6848
rect 9539 6817 9551 6820
rect 9493 6811 9551 6817
rect 12986 6808 12992 6820
rect 13044 6808 13050 6860
rect 10045 6783 10103 6789
rect 10045 6749 10057 6783
rect 10091 6780 10103 6783
rect 10226 6780 10232 6792
rect 10091 6752 10232 6780
rect 10091 6749 10103 6752
rect 10045 6743 10103 6749
rect 10226 6740 10232 6752
rect 10284 6740 10290 6792
rect 10321 6783 10379 6789
rect 10321 6749 10333 6783
rect 10367 6780 10379 6783
rect 10778 6780 10784 6792
rect 10367 6752 10784 6780
rect 10367 6749 10379 6752
rect 10321 6743 10379 6749
rect 10778 6740 10784 6752
rect 10836 6740 10842 6792
rect 11701 6783 11759 6789
rect 11701 6749 11713 6783
rect 11747 6780 11759 6783
rect 13648 6780 13676 6888
rect 14734 6876 14740 6888
rect 14792 6876 14798 6928
rect 16298 6916 16304 6928
rect 16259 6888 16304 6916
rect 16298 6876 16304 6888
rect 16356 6876 16362 6928
rect 17328 6888 17632 6916
rect 13814 6848 13820 6860
rect 13775 6820 13820 6848
rect 13814 6808 13820 6820
rect 13872 6808 13878 6860
rect 14185 6851 14243 6857
rect 14185 6817 14197 6851
rect 14231 6817 14243 6851
rect 14366 6848 14372 6860
rect 14327 6820 14372 6848
rect 14185 6811 14243 6817
rect 11747 6752 13676 6780
rect 13725 6783 13783 6789
rect 11747 6749 11759 6752
rect 11701 6743 11759 6749
rect 13725 6749 13737 6783
rect 13771 6780 13783 6783
rect 13906 6780 13912 6792
rect 13771 6752 13912 6780
rect 13771 6749 13783 6752
rect 13725 6743 13783 6749
rect 13906 6740 13912 6752
rect 13964 6740 13970 6792
rect 14200 6780 14228 6811
rect 14366 6808 14372 6820
rect 14424 6808 14430 6860
rect 15013 6851 15071 6857
rect 15013 6848 15025 6851
rect 14660 6820 15025 6848
rect 14660 6780 14688 6820
rect 15013 6817 15025 6820
rect 15059 6848 15071 6851
rect 15654 6848 15660 6860
rect 15059 6820 15660 6848
rect 15059 6817 15071 6820
rect 15013 6811 15071 6817
rect 15654 6808 15660 6820
rect 15712 6808 15718 6860
rect 16206 6848 16212 6860
rect 15764 6820 16212 6848
rect 14200 6752 14688 6780
rect 14737 6783 14795 6789
rect 14737 6749 14749 6783
rect 14783 6780 14795 6783
rect 15194 6780 15200 6792
rect 14783 6752 15200 6780
rect 14783 6749 14795 6752
rect 14737 6743 14795 6749
rect 15194 6740 15200 6752
rect 15252 6780 15258 6792
rect 15764 6780 15792 6820
rect 16206 6808 16212 6820
rect 16264 6808 16270 6860
rect 16945 6851 17003 6857
rect 16945 6817 16957 6851
rect 16991 6848 17003 6851
rect 17218 6848 17224 6860
rect 16991 6820 17224 6848
rect 16991 6817 17003 6820
rect 16945 6811 17003 6817
rect 17218 6808 17224 6820
rect 17276 6808 17282 6860
rect 17328 6857 17356 6888
rect 17313 6851 17371 6857
rect 17313 6817 17325 6851
rect 17359 6817 17371 6851
rect 17494 6848 17500 6860
rect 17455 6820 17500 6848
rect 17313 6811 17371 6817
rect 17494 6808 17500 6820
rect 17552 6808 17558 6860
rect 17604 6848 17632 6888
rect 18230 6876 18236 6928
rect 18288 6916 18294 6928
rect 20916 6925 20944 6956
rect 21266 6944 21272 6956
rect 21324 6944 21330 6996
rect 21358 6944 21364 6996
rect 21416 6984 21422 6996
rect 23201 6987 23259 6993
rect 23201 6984 23213 6987
rect 21416 6956 23213 6984
rect 21416 6944 21422 6956
rect 23201 6953 23213 6956
rect 23247 6984 23259 6987
rect 23290 6984 23296 6996
rect 23247 6956 23296 6984
rect 23247 6953 23259 6956
rect 23201 6947 23259 6953
rect 23290 6944 23296 6956
rect 23348 6984 23354 6996
rect 23569 6987 23627 6993
rect 23569 6984 23581 6987
rect 23348 6956 23581 6984
rect 23348 6944 23354 6956
rect 23569 6953 23581 6956
rect 23615 6984 23627 6987
rect 24118 6984 24124 6996
rect 23615 6956 24124 6984
rect 23615 6953 23627 6956
rect 23569 6947 23627 6953
rect 24118 6944 24124 6956
rect 24176 6944 24182 6996
rect 24302 6944 24308 6996
rect 24360 6984 24366 6996
rect 28074 6984 28080 6996
rect 24360 6956 28080 6984
rect 24360 6944 24366 6956
rect 28074 6944 28080 6956
rect 28132 6944 28138 6996
rect 28442 6944 28448 6996
rect 28500 6984 28506 6996
rect 29914 6984 29920 6996
rect 28500 6956 29920 6984
rect 28500 6944 28506 6956
rect 29914 6944 29920 6956
rect 29972 6944 29978 6996
rect 31202 6984 31208 6996
rect 31163 6956 31208 6984
rect 31202 6944 31208 6956
rect 31260 6944 31266 6996
rect 32309 6987 32367 6993
rect 32309 6953 32321 6987
rect 32355 6953 32367 6987
rect 32309 6947 32367 6953
rect 18325 6919 18383 6925
rect 18325 6916 18337 6919
rect 18288 6888 18337 6916
rect 18288 6876 18294 6888
rect 18325 6885 18337 6888
rect 18371 6885 18383 6919
rect 20901 6919 20959 6925
rect 18325 6879 18383 6885
rect 19076 6888 20024 6916
rect 19076 6860 19104 6888
rect 18046 6848 18052 6860
rect 17604 6820 18052 6848
rect 18046 6808 18052 6820
rect 18104 6808 18110 6860
rect 18969 6851 19027 6857
rect 18969 6848 18981 6851
rect 18616 6820 18981 6848
rect 15252 6752 15792 6780
rect 15841 6783 15899 6789
rect 15252 6740 15258 6752
rect 15841 6749 15853 6783
rect 15887 6780 15899 6783
rect 17034 6780 17040 6792
rect 15887 6752 17040 6780
rect 15887 6749 15899 6752
rect 15841 6743 15899 6749
rect 17034 6740 17040 6752
rect 17092 6740 17098 6792
rect 17126 6740 17132 6792
rect 17184 6780 17190 6792
rect 17184 6752 18368 6780
rect 17184 6740 17190 6752
rect 15930 6712 15936 6724
rect 13004 6684 15936 6712
rect 11238 6644 11244 6656
rect 9416 6616 11244 6644
rect 8941 6607 8999 6613
rect 11238 6604 11244 6616
rect 11296 6604 11302 6656
rect 11698 6604 11704 6656
rect 11756 6644 11762 6656
rect 13004 6644 13032 6684
rect 15930 6672 15936 6684
rect 15988 6672 15994 6724
rect 18138 6712 18144 6724
rect 16132 6684 18144 6712
rect 16132 6656 16160 6684
rect 18138 6672 18144 6684
rect 18196 6672 18202 6724
rect 11756 6616 13032 6644
rect 13081 6647 13139 6653
rect 11756 6604 11762 6616
rect 13081 6613 13093 6647
rect 13127 6644 13139 6647
rect 14182 6644 14188 6656
rect 13127 6616 14188 6644
rect 13127 6613 13139 6616
rect 13081 6607 13139 6613
rect 14182 6604 14188 6616
rect 14240 6604 14246 6656
rect 16114 6644 16120 6656
rect 16075 6616 16120 6644
rect 16114 6604 16120 6616
rect 16172 6604 16178 6656
rect 16206 6604 16212 6656
rect 16264 6644 16270 6656
rect 17126 6644 17132 6656
rect 16264 6616 17132 6644
rect 16264 6604 16270 6616
rect 17126 6604 17132 6616
rect 17184 6604 17190 6656
rect 17218 6604 17224 6656
rect 17276 6644 17282 6656
rect 17589 6647 17647 6653
rect 17589 6644 17601 6647
rect 17276 6616 17601 6644
rect 17276 6604 17282 6616
rect 17589 6613 17601 6616
rect 17635 6613 17647 6647
rect 18230 6644 18236 6656
rect 18191 6616 18236 6644
rect 17589 6607 17647 6613
rect 18230 6604 18236 6616
rect 18288 6604 18294 6656
rect 18340 6644 18368 6752
rect 18616 6712 18644 6820
rect 18969 6817 18981 6820
rect 19015 6817 19027 6851
rect 18969 6811 19027 6817
rect 19058 6808 19064 6860
rect 19116 6848 19122 6860
rect 19116 6820 19209 6848
rect 19116 6808 19122 6820
rect 19242 6808 19248 6860
rect 19300 6857 19306 6860
rect 19300 6851 19361 6857
rect 19300 6817 19315 6851
rect 19349 6817 19361 6851
rect 19518 6848 19524 6860
rect 19479 6820 19524 6848
rect 19300 6811 19361 6817
rect 19300 6808 19306 6811
rect 19518 6808 19524 6820
rect 19576 6808 19582 6860
rect 19996 6780 20024 6888
rect 20901 6885 20913 6919
rect 20947 6885 20959 6919
rect 20901 6879 20959 6885
rect 24964 6888 25176 6916
rect 20070 6808 20076 6860
rect 20128 6848 20134 6860
rect 20622 6848 20628 6860
rect 20128 6820 20628 6848
rect 20128 6808 20134 6820
rect 20622 6808 20628 6820
rect 20680 6848 20686 6860
rect 21085 6851 21143 6857
rect 21085 6848 21097 6851
rect 20680 6820 21097 6848
rect 20680 6808 20686 6820
rect 21085 6817 21097 6820
rect 21131 6817 21143 6851
rect 22097 6851 22155 6857
rect 22097 6848 22109 6851
rect 21085 6811 21143 6817
rect 21192 6820 22109 6848
rect 21192 6780 21220 6820
rect 22097 6817 22109 6820
rect 22143 6817 22155 6851
rect 22554 6848 22560 6860
rect 22515 6820 22560 6848
rect 22097 6811 22155 6817
rect 22554 6808 22560 6820
rect 22612 6808 22618 6860
rect 22646 6808 22652 6860
rect 22704 6848 22710 6860
rect 23753 6851 23811 6857
rect 22704 6820 22749 6848
rect 22704 6808 22710 6820
rect 23753 6817 23765 6851
rect 23799 6848 23811 6851
rect 24026 6848 24032 6860
rect 23799 6820 24032 6848
rect 23799 6817 23811 6820
rect 23753 6811 23811 6817
rect 24026 6808 24032 6820
rect 24084 6808 24090 6860
rect 24302 6808 24308 6860
rect 24360 6848 24366 6860
rect 24964 6848 24992 6888
rect 25148 6857 25176 6888
rect 26510 6876 26516 6928
rect 26568 6916 26574 6928
rect 28258 6916 28264 6928
rect 26568 6888 28264 6916
rect 26568 6876 26574 6888
rect 24360 6820 24992 6848
rect 25041 6851 25099 6857
rect 24360 6808 24366 6820
rect 25041 6817 25053 6851
rect 25087 6817 25099 6851
rect 25041 6811 25099 6817
rect 25133 6851 25191 6857
rect 25133 6817 25145 6851
rect 25179 6817 25191 6851
rect 25133 6811 25191 6817
rect 19996 6752 21220 6780
rect 21453 6783 21511 6789
rect 21453 6749 21465 6783
rect 21499 6749 21511 6783
rect 21818 6780 21824 6792
rect 21779 6752 21824 6780
rect 21453 6743 21511 6749
rect 19334 6712 19340 6724
rect 18616 6684 19340 6712
rect 19334 6672 19340 6684
rect 19392 6672 19398 6724
rect 21468 6712 21496 6743
rect 21818 6740 21824 6752
rect 21876 6740 21882 6792
rect 24854 6780 24860 6792
rect 23676 6752 24860 6780
rect 23676 6712 23704 6752
rect 24854 6740 24860 6752
rect 24912 6740 24918 6792
rect 25056 6780 25084 6811
rect 25314 6808 25320 6860
rect 25372 6848 25378 6860
rect 26694 6848 26700 6860
rect 25372 6820 26700 6848
rect 25372 6808 25378 6820
rect 26694 6808 26700 6820
rect 26752 6808 26758 6860
rect 26789 6851 26847 6857
rect 26789 6817 26801 6851
rect 26835 6848 26847 6851
rect 27062 6848 27068 6860
rect 26835 6820 27068 6848
rect 26835 6817 26847 6820
rect 26789 6811 26847 6817
rect 25406 6780 25412 6792
rect 25056 6752 25412 6780
rect 21468 6684 23704 6712
rect 23750 6672 23756 6724
rect 23808 6712 23814 6724
rect 24670 6712 24676 6724
rect 23808 6684 24676 6712
rect 23808 6672 23814 6684
rect 24670 6672 24676 6684
rect 24728 6672 24734 6724
rect 24765 6715 24823 6721
rect 24765 6681 24777 6715
rect 24811 6712 24823 6715
rect 25056 6712 25084 6752
rect 25406 6740 25412 6752
rect 25464 6740 25470 6792
rect 25593 6783 25651 6789
rect 25593 6749 25605 6783
rect 25639 6780 25651 6783
rect 25774 6780 25780 6792
rect 25639 6752 25780 6780
rect 25639 6749 25651 6752
rect 25593 6743 25651 6749
rect 25774 6740 25780 6752
rect 25832 6740 25838 6792
rect 25961 6783 26019 6789
rect 25961 6749 25973 6783
rect 26007 6780 26019 6783
rect 26326 6780 26332 6792
rect 26007 6752 26332 6780
rect 26007 6749 26019 6752
rect 25961 6743 26019 6749
rect 26326 6740 26332 6752
rect 26384 6780 26390 6792
rect 26804 6780 26832 6811
rect 27062 6808 27068 6820
rect 27120 6808 27126 6860
rect 27154 6808 27160 6860
rect 27212 6848 27218 6860
rect 27356 6857 27384 6888
rect 28258 6876 28264 6888
rect 28316 6876 28322 6928
rect 28534 6876 28540 6928
rect 28592 6916 28598 6928
rect 28994 6916 29000 6928
rect 28592 6888 29000 6916
rect 28592 6876 28598 6888
rect 28994 6876 29000 6888
rect 29052 6876 29058 6928
rect 29086 6876 29092 6928
rect 29144 6916 29150 6928
rect 32324 6916 32352 6947
rect 33410 6944 33416 6996
rect 33468 6984 33474 6996
rect 38746 6984 38752 6996
rect 33468 6956 38752 6984
rect 33468 6944 33474 6956
rect 38746 6944 38752 6956
rect 38804 6984 38810 6996
rect 39022 6984 39028 6996
rect 38804 6956 39028 6984
rect 38804 6944 38810 6956
rect 39022 6944 39028 6956
rect 39080 6944 39086 6996
rect 39666 6984 39672 6996
rect 39627 6956 39672 6984
rect 39666 6944 39672 6956
rect 39724 6944 39730 6996
rect 39850 6944 39856 6996
rect 39908 6984 39914 6996
rect 45186 6984 45192 6996
rect 39908 6956 45192 6984
rect 39908 6944 39914 6956
rect 45186 6944 45192 6956
rect 45244 6944 45250 6996
rect 46385 6987 46443 6993
rect 46385 6984 46397 6987
rect 45296 6956 46397 6984
rect 29144 6888 32352 6916
rect 29144 6876 29150 6888
rect 34514 6876 34520 6928
rect 34572 6916 34578 6928
rect 36541 6919 36599 6925
rect 36541 6916 36553 6919
rect 34572 6888 36553 6916
rect 34572 6876 34578 6888
rect 36541 6885 36553 6888
rect 36587 6885 36599 6919
rect 39758 6916 39764 6928
rect 36541 6879 36599 6885
rect 38856 6888 39764 6916
rect 27337 6851 27395 6857
rect 27212 6820 27257 6848
rect 27212 6808 27218 6820
rect 27337 6817 27349 6851
rect 27383 6817 27395 6851
rect 27337 6811 27395 6817
rect 27430 6808 27436 6860
rect 27488 6848 27494 6860
rect 28629 6851 28687 6857
rect 27488 6820 28304 6848
rect 27488 6808 27494 6820
rect 28276 6792 28304 6820
rect 28629 6817 28641 6851
rect 28675 6848 28687 6851
rect 28718 6848 28724 6860
rect 28675 6820 28724 6848
rect 28675 6817 28687 6820
rect 28629 6811 28687 6817
rect 28718 6808 28724 6820
rect 28776 6808 28782 6860
rect 28813 6851 28871 6857
rect 28813 6817 28825 6851
rect 28859 6817 28871 6851
rect 29454 6848 29460 6860
rect 29415 6820 29460 6848
rect 28813 6811 28871 6817
rect 26384 6752 26832 6780
rect 26384 6740 26390 6752
rect 28258 6740 28264 6792
rect 28316 6740 28322 6792
rect 28828 6724 28856 6811
rect 29454 6808 29460 6820
rect 29512 6808 29518 6860
rect 29733 6851 29791 6857
rect 29733 6817 29745 6851
rect 29779 6848 29791 6851
rect 30006 6848 30012 6860
rect 29779 6820 30012 6848
rect 29779 6817 29791 6820
rect 29733 6811 29791 6817
rect 30006 6808 30012 6820
rect 30064 6848 30070 6860
rect 30469 6851 30527 6857
rect 30469 6848 30481 6851
rect 30064 6820 30481 6848
rect 30064 6808 30070 6820
rect 30469 6817 30481 6820
rect 30515 6817 30527 6851
rect 30469 6811 30527 6817
rect 30558 6808 30564 6860
rect 30616 6848 30622 6860
rect 30653 6851 30711 6857
rect 30653 6848 30665 6851
rect 30616 6820 30665 6848
rect 30616 6808 30622 6820
rect 30653 6817 30665 6820
rect 30699 6848 30711 6851
rect 31294 6848 31300 6860
rect 30699 6820 31300 6848
rect 30699 6817 30711 6820
rect 30653 6811 30711 6817
rect 31294 6808 31300 6820
rect 31352 6808 31358 6860
rect 32125 6851 32183 6857
rect 32125 6817 32137 6851
rect 32171 6848 32183 6851
rect 32171 6820 32536 6848
rect 32171 6817 32183 6820
rect 32125 6811 32183 6817
rect 29086 6740 29092 6792
rect 29144 6780 29150 6792
rect 29472 6780 29500 6808
rect 32508 6792 32536 6820
rect 32950 6808 32956 6860
rect 33008 6848 33014 6860
rect 36122 6851 36180 6857
rect 33008 6820 34928 6848
rect 33008 6808 33014 6820
rect 29144 6752 29500 6780
rect 29144 6740 29150 6752
rect 32490 6740 32496 6792
rect 32548 6740 32554 6792
rect 33410 6740 33416 6792
rect 33468 6780 33474 6792
rect 33505 6783 33563 6789
rect 33505 6780 33517 6783
rect 33468 6752 33517 6780
rect 33468 6740 33474 6752
rect 33505 6749 33517 6752
rect 33551 6780 33563 6783
rect 33686 6780 33692 6792
rect 33551 6752 33692 6780
rect 33551 6749 33563 6752
rect 33505 6743 33563 6749
rect 33686 6740 33692 6752
rect 33744 6740 33750 6792
rect 33781 6783 33839 6789
rect 33781 6749 33793 6783
rect 33827 6780 33839 6783
rect 34238 6780 34244 6792
rect 33827 6752 34244 6780
rect 33827 6749 33839 6752
rect 33781 6743 33839 6749
rect 34238 6740 34244 6752
rect 34296 6740 34302 6792
rect 34900 6789 34928 6820
rect 36122 6817 36134 6851
rect 36168 6848 36180 6851
rect 36906 6848 36912 6860
rect 36168 6820 36912 6848
rect 36168 6817 36180 6820
rect 36122 6811 36180 6817
rect 36906 6808 36912 6820
rect 36964 6808 36970 6860
rect 38378 6848 38384 6860
rect 38339 6820 38384 6848
rect 38378 6808 38384 6820
rect 38436 6808 38442 6860
rect 38746 6848 38752 6860
rect 38707 6820 38752 6848
rect 38746 6808 38752 6820
rect 38804 6808 38810 6860
rect 34885 6783 34943 6789
rect 34885 6749 34897 6783
rect 34931 6749 34943 6783
rect 34885 6743 34943 6749
rect 24811 6684 25084 6712
rect 24811 6681 24823 6684
rect 24765 6675 24823 6681
rect 25130 6672 25136 6724
rect 25188 6712 25194 6724
rect 26234 6712 26240 6724
rect 25188 6684 26240 6712
rect 25188 6672 25194 6684
rect 26234 6672 26240 6684
rect 26292 6672 26298 6724
rect 26878 6672 26884 6724
rect 26936 6712 26942 6724
rect 27617 6715 27675 6721
rect 27617 6712 27629 6715
rect 26936 6684 27629 6712
rect 26936 6672 26942 6684
rect 27617 6681 27629 6684
rect 27663 6681 27675 6715
rect 27617 6675 27675 6681
rect 28810 6672 28816 6724
rect 28868 6672 28874 6724
rect 28905 6715 28963 6721
rect 28905 6681 28917 6715
rect 28951 6681 28963 6715
rect 28905 6675 28963 6681
rect 19886 6644 19892 6656
rect 18340 6616 19892 6644
rect 19886 6604 19892 6616
rect 19944 6604 19950 6656
rect 20162 6644 20168 6656
rect 20123 6616 20168 6644
rect 20162 6604 20168 6616
rect 20220 6604 20226 6656
rect 20530 6604 20536 6656
rect 20588 6644 20594 6656
rect 20625 6647 20683 6653
rect 20625 6644 20637 6647
rect 20588 6616 20637 6644
rect 20588 6604 20594 6616
rect 20625 6613 20637 6616
rect 20671 6644 20683 6647
rect 22462 6644 22468 6656
rect 20671 6616 22468 6644
rect 20671 6613 20683 6616
rect 20625 6607 20683 6613
rect 22462 6604 22468 6616
rect 22520 6604 22526 6656
rect 22830 6644 22836 6656
rect 22791 6616 22836 6644
rect 22830 6604 22836 6616
rect 22888 6604 22894 6656
rect 22922 6604 22928 6656
rect 22980 6644 22986 6656
rect 23937 6647 23995 6653
rect 23937 6644 23949 6647
rect 22980 6616 23949 6644
rect 22980 6604 22986 6616
rect 23937 6613 23949 6616
rect 23983 6613 23995 6647
rect 24302 6644 24308 6656
rect 24263 6616 24308 6644
rect 23937 6607 23995 6613
rect 24302 6604 24308 6616
rect 24360 6604 24366 6656
rect 24854 6644 24860 6656
rect 24815 6616 24860 6644
rect 24854 6604 24860 6616
rect 24912 6604 24918 6656
rect 28261 6647 28319 6653
rect 28261 6613 28273 6647
rect 28307 6644 28319 6647
rect 28626 6644 28632 6656
rect 28307 6616 28632 6644
rect 28307 6613 28319 6616
rect 28261 6607 28319 6613
rect 28626 6604 28632 6616
rect 28684 6644 28690 6656
rect 28920 6644 28948 6675
rect 29546 6672 29552 6724
rect 29604 6712 29610 6724
rect 30193 6715 30251 6721
rect 30193 6712 30205 6715
rect 29604 6684 30205 6712
rect 29604 6672 29610 6684
rect 30193 6681 30205 6684
rect 30239 6712 30251 6715
rect 31662 6712 31668 6724
rect 30239 6684 31668 6712
rect 30239 6681 30251 6684
rect 30193 6675 30251 6681
rect 31662 6672 31668 6684
rect 31720 6672 31726 6724
rect 34900 6712 34928 6743
rect 35894 6740 35900 6792
rect 35952 6780 35958 6792
rect 35989 6783 36047 6789
rect 35989 6780 36001 6783
rect 35952 6752 36001 6780
rect 35952 6740 35958 6752
rect 35989 6749 36001 6752
rect 36035 6749 36047 6783
rect 37274 6780 37280 6792
rect 37187 6752 37280 6780
rect 35989 6743 36047 6749
rect 37274 6740 37280 6752
rect 37332 6780 37338 6792
rect 38013 6783 38071 6789
rect 38013 6780 38025 6783
rect 37332 6752 38025 6780
rect 37332 6740 37338 6752
rect 38013 6749 38025 6752
rect 38059 6780 38071 6783
rect 38470 6780 38476 6792
rect 38059 6752 38476 6780
rect 38059 6749 38071 6752
rect 38013 6743 38071 6749
rect 38470 6740 38476 6752
rect 38528 6740 38534 6792
rect 38856 6780 38884 6888
rect 39758 6876 39764 6888
rect 39816 6876 39822 6928
rect 40773 6919 40831 6925
rect 40773 6916 40785 6919
rect 39960 6888 40785 6916
rect 39390 6808 39396 6860
rect 39448 6848 39454 6860
rect 39960 6857 39988 6888
rect 40773 6885 40785 6888
rect 40819 6885 40831 6919
rect 40773 6879 40831 6885
rect 43070 6876 43076 6928
rect 43128 6916 43134 6928
rect 43717 6919 43775 6925
rect 43717 6916 43729 6919
rect 43128 6888 43729 6916
rect 43128 6876 43134 6888
rect 43717 6885 43729 6888
rect 43763 6916 43775 6919
rect 45296 6916 45324 6956
rect 46385 6953 46397 6956
rect 46431 6953 46443 6987
rect 46385 6947 46443 6953
rect 46934 6944 46940 6996
rect 46992 6984 46998 6996
rect 47489 6987 47547 6993
rect 47489 6984 47501 6987
rect 46992 6956 47501 6984
rect 46992 6944 46998 6956
rect 47489 6953 47501 6956
rect 47535 6953 47547 6987
rect 47489 6947 47547 6953
rect 48590 6944 48596 6996
rect 48648 6984 48654 6996
rect 50982 6984 50988 6996
rect 48648 6956 50988 6984
rect 48648 6944 48654 6956
rect 50982 6944 50988 6956
rect 51040 6984 51046 6996
rect 51537 6987 51595 6993
rect 51537 6984 51549 6987
rect 51040 6956 51549 6984
rect 51040 6944 51046 6956
rect 51537 6953 51549 6956
rect 51583 6953 51595 6987
rect 51537 6947 51595 6953
rect 51626 6944 51632 6996
rect 51684 6984 51690 6996
rect 54202 6984 54208 6996
rect 51684 6956 54208 6984
rect 51684 6944 51690 6956
rect 54202 6944 54208 6956
rect 54260 6984 54266 6996
rect 55125 6987 55183 6993
rect 55125 6984 55137 6987
rect 54260 6956 55137 6984
rect 54260 6944 54266 6956
rect 55125 6953 55137 6956
rect 55171 6953 55183 6987
rect 56594 6984 56600 6996
rect 55125 6947 55183 6953
rect 56152 6956 56600 6984
rect 43763 6888 45324 6916
rect 43763 6885 43775 6888
rect 43717 6879 43775 6885
rect 45554 6876 45560 6928
rect 45612 6876 45618 6928
rect 45646 6876 45652 6928
rect 45704 6916 45710 6928
rect 45704 6888 46980 6916
rect 45704 6876 45710 6888
rect 39945 6851 40003 6857
rect 39945 6848 39957 6851
rect 39448 6820 39957 6848
rect 39448 6808 39454 6820
rect 39945 6817 39957 6820
rect 39991 6817 40003 6851
rect 39945 6811 40003 6817
rect 40037 6851 40095 6857
rect 40037 6817 40049 6851
rect 40083 6848 40095 6851
rect 41141 6851 41199 6857
rect 41141 6848 41153 6851
rect 40083 6820 41153 6848
rect 40083 6817 40095 6820
rect 40037 6811 40095 6817
rect 41141 6817 41153 6820
rect 41187 6817 41199 6851
rect 41598 6848 41604 6860
rect 41559 6820 41604 6848
rect 41141 6811 41199 6817
rect 38672 6752 38884 6780
rect 38933 6783 38991 6789
rect 38672 6724 38700 6752
rect 38933 6749 38945 6783
rect 38979 6780 38991 6783
rect 40052 6780 40080 6811
rect 41598 6808 41604 6820
rect 41656 6808 41662 6860
rect 41693 6851 41751 6857
rect 41693 6817 41705 6851
rect 41739 6848 41751 6851
rect 41782 6848 41788 6860
rect 41739 6820 41788 6848
rect 41739 6817 41751 6820
rect 41693 6811 41751 6817
rect 41782 6808 41788 6820
rect 41840 6808 41846 6860
rect 42889 6851 42947 6857
rect 42889 6817 42901 6851
rect 42935 6848 42947 6851
rect 43346 6848 43352 6860
rect 42935 6820 43352 6848
rect 42935 6817 42947 6820
rect 42889 6811 42947 6817
rect 43346 6808 43352 6820
rect 43404 6808 43410 6860
rect 44269 6851 44327 6857
rect 44269 6817 44281 6851
rect 44315 6848 44327 6851
rect 44634 6848 44640 6860
rect 44315 6820 44640 6848
rect 44315 6817 44327 6820
rect 44269 6811 44327 6817
rect 44634 6808 44640 6820
rect 44692 6808 44698 6860
rect 45097 6851 45155 6857
rect 45097 6817 45109 6851
rect 45143 6848 45155 6851
rect 45572 6848 45600 6876
rect 45143 6820 45600 6848
rect 45143 6817 45155 6820
rect 45097 6811 45155 6817
rect 46198 6808 46204 6860
rect 46256 6848 46262 6860
rect 46477 6851 46535 6857
rect 46477 6848 46489 6851
rect 46256 6820 46489 6848
rect 46256 6808 46262 6820
rect 46477 6817 46489 6820
rect 46523 6817 46535 6851
rect 46952 6848 46980 6888
rect 47394 6876 47400 6928
rect 47452 6916 47458 6928
rect 47857 6919 47915 6925
rect 47857 6916 47869 6919
rect 47452 6888 47869 6916
rect 47452 6876 47458 6888
rect 47857 6885 47869 6888
rect 47903 6885 47915 6919
rect 54110 6916 54116 6928
rect 47857 6879 47915 6885
rect 50724 6888 54116 6916
rect 50724 6860 50752 6888
rect 54110 6876 54116 6888
rect 54168 6876 54174 6928
rect 54849 6919 54907 6925
rect 54849 6885 54861 6919
rect 54895 6916 54907 6919
rect 55030 6916 55036 6928
rect 54895 6888 55036 6916
rect 54895 6885 54907 6888
rect 54849 6879 54907 6885
rect 55030 6876 55036 6888
rect 55088 6876 55094 6928
rect 48406 6848 48412 6860
rect 46477 6811 46535 6817
rect 46584 6820 46888 6848
rect 46952 6820 48412 6848
rect 38979 6752 40080 6780
rect 42153 6783 42211 6789
rect 38979 6749 38991 6752
rect 38933 6743 38991 6749
rect 42153 6749 42165 6783
rect 42199 6780 42211 6783
rect 42978 6780 42984 6792
rect 42199 6752 42984 6780
rect 42199 6749 42211 6752
rect 42153 6743 42211 6749
rect 42978 6740 42984 6752
rect 43036 6740 43042 6792
rect 44361 6783 44419 6789
rect 44361 6749 44373 6783
rect 44407 6749 44419 6783
rect 44361 6743 44419 6749
rect 36446 6712 36452 6724
rect 34900 6684 36452 6712
rect 36446 6672 36452 6684
rect 36504 6672 36510 6724
rect 36538 6672 36544 6724
rect 36596 6712 36602 6724
rect 38654 6712 38660 6724
rect 36596 6684 38660 6712
rect 36596 6672 36602 6684
rect 38654 6672 38660 6684
rect 38712 6672 38718 6724
rect 38746 6672 38752 6724
rect 38804 6712 38810 6724
rect 39206 6712 39212 6724
rect 38804 6684 39212 6712
rect 38804 6672 38810 6684
rect 39206 6672 39212 6684
rect 39264 6672 39270 6724
rect 39298 6672 39304 6724
rect 39356 6712 39362 6724
rect 44376 6712 44404 6743
rect 44726 6740 44732 6792
rect 44784 6780 44790 6792
rect 45189 6783 45247 6789
rect 45189 6780 45201 6783
rect 44784 6752 45201 6780
rect 44784 6740 44790 6752
rect 45189 6749 45201 6752
rect 45235 6780 45247 6783
rect 45557 6783 45615 6789
rect 45557 6780 45569 6783
rect 45235 6752 45569 6780
rect 45235 6749 45247 6752
rect 45189 6743 45247 6749
rect 45557 6749 45569 6752
rect 45603 6749 45615 6783
rect 45557 6743 45615 6749
rect 46382 6740 46388 6792
rect 46440 6780 46446 6792
rect 46584 6780 46612 6820
rect 46440 6752 46612 6780
rect 46440 6740 46446 6752
rect 46658 6740 46664 6792
rect 46716 6780 46722 6792
rect 46860 6789 46888 6820
rect 48406 6808 48412 6820
rect 48464 6808 48470 6860
rect 48590 6848 48596 6860
rect 48551 6820 48596 6848
rect 48590 6808 48596 6820
rect 48648 6808 48654 6860
rect 49694 6808 49700 6860
rect 49752 6848 49758 6860
rect 49789 6851 49847 6857
rect 49789 6848 49801 6851
rect 49752 6820 49801 6848
rect 49752 6808 49758 6820
rect 49789 6817 49801 6820
rect 49835 6817 49847 6851
rect 49789 6811 49847 6817
rect 49878 6808 49884 6860
rect 49936 6848 49942 6860
rect 50065 6851 50123 6857
rect 50065 6848 50077 6851
rect 49936 6820 50077 6848
rect 49936 6808 49942 6820
rect 50065 6817 50077 6820
rect 50111 6848 50123 6851
rect 50338 6848 50344 6860
rect 50111 6820 50344 6848
rect 50111 6817 50123 6820
rect 50065 6811 50123 6817
rect 50338 6808 50344 6820
rect 50396 6808 50402 6860
rect 50706 6808 50712 6860
rect 50764 6808 50770 6860
rect 50982 6808 50988 6860
rect 51040 6848 51046 6860
rect 52273 6851 52331 6857
rect 52273 6848 52285 6851
rect 51040 6820 52285 6848
rect 51040 6808 51046 6820
rect 52273 6817 52285 6820
rect 52319 6817 52331 6851
rect 52454 6848 52460 6860
rect 52415 6820 52460 6848
rect 52273 6811 52331 6817
rect 52454 6808 52460 6820
rect 52512 6808 52518 6860
rect 53282 6848 53288 6860
rect 52748 6820 53288 6848
rect 46845 6783 46903 6789
rect 46716 6752 46796 6780
rect 46716 6740 46722 6752
rect 45094 6712 45100 6724
rect 39356 6684 40264 6712
rect 44376 6684 45100 6712
rect 39356 6672 39362 6684
rect 28684 6616 28948 6644
rect 28684 6604 28690 6616
rect 30374 6604 30380 6656
rect 30432 6644 30438 6656
rect 30837 6647 30895 6653
rect 30837 6644 30849 6647
rect 30432 6616 30849 6644
rect 30432 6604 30438 6616
rect 30837 6613 30849 6616
rect 30883 6644 30895 6647
rect 30926 6644 30932 6656
rect 30883 6616 30932 6644
rect 30883 6613 30895 6616
rect 30837 6607 30895 6613
rect 30926 6604 30932 6616
rect 30984 6604 30990 6656
rect 31938 6644 31944 6656
rect 31899 6616 31944 6644
rect 31938 6604 31944 6616
rect 31996 6604 32002 6656
rect 32582 6604 32588 6656
rect 32640 6644 32646 6656
rect 32677 6647 32735 6653
rect 32677 6644 32689 6647
rect 32640 6616 32689 6644
rect 32640 6604 32646 6616
rect 32677 6613 32689 6616
rect 32723 6644 32735 6647
rect 33045 6647 33103 6653
rect 33045 6644 33057 6647
rect 32723 6616 33057 6644
rect 32723 6613 32735 6616
rect 32677 6607 32735 6613
rect 33045 6613 33057 6616
rect 33091 6613 33103 6647
rect 35618 6644 35624 6656
rect 35579 6616 35624 6644
rect 33045 6607 33103 6613
rect 35618 6604 35624 6616
rect 35676 6604 35682 6656
rect 39758 6644 39764 6656
rect 39719 6616 39764 6644
rect 39758 6604 39764 6616
rect 39816 6604 39822 6656
rect 40236 6653 40264 6684
rect 45094 6672 45100 6684
rect 45152 6672 45158 6724
rect 46768 6721 46796 6752
rect 46845 6749 46857 6783
rect 46891 6749 46903 6783
rect 47210 6780 47216 6792
rect 47171 6752 47216 6780
rect 46845 6743 46903 6749
rect 47210 6740 47216 6752
rect 47268 6740 47274 6792
rect 47394 6740 47400 6792
rect 47452 6780 47458 6792
rect 48225 6783 48283 6789
rect 48225 6780 48237 6783
rect 47452 6752 48237 6780
rect 47452 6740 47458 6752
rect 48225 6749 48237 6752
rect 48271 6749 48283 6783
rect 48225 6743 48283 6749
rect 51445 6783 51503 6789
rect 51445 6749 51457 6783
rect 51491 6780 51503 6783
rect 51537 6783 51595 6789
rect 51537 6780 51549 6783
rect 51491 6752 51549 6780
rect 51491 6749 51503 6752
rect 51445 6743 51503 6749
rect 51537 6749 51549 6752
rect 51583 6780 51595 6783
rect 51721 6783 51779 6789
rect 51721 6780 51733 6783
rect 51583 6752 51733 6780
rect 51583 6749 51595 6752
rect 51537 6743 51595 6749
rect 51721 6749 51733 6752
rect 51767 6749 51779 6783
rect 52178 6780 52184 6792
rect 52139 6752 52184 6780
rect 51721 6743 51779 6749
rect 52178 6740 52184 6752
rect 52236 6740 52242 6792
rect 46753 6715 46811 6721
rect 46753 6681 46765 6715
rect 46799 6681 46811 6715
rect 46753 6675 46811 6681
rect 46934 6672 46940 6724
rect 46992 6712 46998 6724
rect 46992 6684 49832 6712
rect 46992 6672 46998 6684
rect 40221 6647 40279 6653
rect 40221 6613 40233 6647
rect 40267 6613 40279 6647
rect 40221 6607 40279 6613
rect 41417 6647 41475 6653
rect 41417 6613 41429 6647
rect 41463 6644 41475 6647
rect 41874 6644 41880 6656
rect 41463 6616 41880 6644
rect 41463 6613 41475 6616
rect 41417 6607 41475 6613
rect 41874 6604 41880 6616
rect 41932 6604 41938 6656
rect 42518 6644 42524 6656
rect 42479 6616 42524 6644
rect 42518 6604 42524 6616
rect 42576 6604 42582 6656
rect 44085 6647 44143 6653
rect 44085 6613 44097 6647
rect 44131 6644 44143 6647
rect 44174 6644 44180 6656
rect 44131 6616 44180 6644
rect 44131 6613 44143 6616
rect 44085 6607 44143 6613
rect 44174 6604 44180 6616
rect 44232 6604 44238 6656
rect 46106 6604 46112 6656
rect 46164 6644 46170 6656
rect 46201 6647 46259 6653
rect 46201 6644 46213 6647
rect 46164 6616 46213 6644
rect 46164 6604 46170 6616
rect 46201 6613 46213 6616
rect 46247 6613 46259 6647
rect 46201 6607 46259 6613
rect 46385 6647 46443 6653
rect 46385 6613 46397 6647
rect 46431 6644 46443 6647
rect 46642 6647 46700 6653
rect 46642 6644 46654 6647
rect 46431 6616 46654 6644
rect 46431 6613 46443 6616
rect 46385 6607 46443 6613
rect 46642 6613 46654 6616
rect 46688 6644 46700 6647
rect 47486 6644 47492 6656
rect 46688 6616 47492 6644
rect 46688 6613 46700 6616
rect 46642 6607 46700 6613
rect 47486 6604 47492 6616
rect 47544 6604 47550 6656
rect 47946 6604 47952 6656
rect 48004 6644 48010 6656
rect 49145 6647 49203 6653
rect 49145 6644 49157 6647
rect 48004 6616 49157 6644
rect 48004 6604 48010 6616
rect 49145 6613 49157 6616
rect 49191 6613 49203 6647
rect 49602 6644 49608 6656
rect 49563 6616 49608 6644
rect 49145 6607 49203 6613
rect 49602 6604 49608 6616
rect 49660 6604 49666 6656
rect 49804 6644 49832 6684
rect 51166 6672 51172 6724
rect 51224 6712 51230 6724
rect 52748 6712 52776 6820
rect 53282 6808 53288 6820
rect 53340 6848 53346 6860
rect 53653 6851 53711 6857
rect 53653 6848 53665 6851
rect 53340 6820 53665 6848
rect 53340 6808 53346 6820
rect 53653 6817 53665 6820
rect 53699 6848 53711 6851
rect 54938 6848 54944 6860
rect 53699 6820 53972 6848
rect 54899 6820 54944 6848
rect 53699 6817 53711 6820
rect 53653 6811 53711 6817
rect 52825 6783 52883 6789
rect 52825 6749 52837 6783
rect 52871 6780 52883 6783
rect 53834 6780 53840 6792
rect 52871 6752 53840 6780
rect 52871 6749 52883 6752
rect 52825 6743 52883 6749
rect 53834 6740 53840 6752
rect 53892 6740 53898 6792
rect 53944 6780 53972 6820
rect 54938 6808 54944 6820
rect 54996 6808 55002 6860
rect 56152 6857 56180 6956
rect 56594 6944 56600 6956
rect 56652 6944 56658 6996
rect 57698 6984 57704 6996
rect 57532 6956 57704 6984
rect 57532 6916 57560 6956
rect 57698 6944 57704 6956
rect 57756 6944 57762 6996
rect 56244 6888 57560 6916
rect 56244 6857 56272 6888
rect 57606 6876 57612 6928
rect 57664 6916 57670 6928
rect 57664 6888 58480 6916
rect 57664 6876 57670 6888
rect 56137 6851 56195 6857
rect 56137 6817 56149 6851
rect 56183 6817 56195 6851
rect 56137 6811 56195 6817
rect 56229 6851 56287 6857
rect 56229 6817 56241 6851
rect 56275 6817 56287 6851
rect 56229 6811 56287 6817
rect 56321 6851 56379 6857
rect 56321 6817 56333 6851
rect 56367 6817 56379 6851
rect 56321 6811 56379 6817
rect 56781 6851 56839 6857
rect 56781 6817 56793 6851
rect 56827 6848 56839 6851
rect 57330 6848 57336 6860
rect 56827 6820 57336 6848
rect 56827 6817 56839 6820
rect 56781 6811 56839 6817
rect 55493 6783 55551 6789
rect 55493 6780 55505 6783
rect 53944 6752 55505 6780
rect 55493 6749 55505 6752
rect 55539 6780 55551 6783
rect 55950 6780 55956 6792
rect 55539 6752 55956 6780
rect 55539 6749 55551 6752
rect 55493 6743 55551 6749
rect 55950 6740 55956 6752
rect 56008 6740 56014 6792
rect 56336 6780 56364 6811
rect 57330 6808 57336 6820
rect 57388 6808 57394 6860
rect 57514 6848 57520 6860
rect 57475 6820 57520 6848
rect 57514 6808 57520 6820
rect 57572 6808 57578 6860
rect 57790 6808 57796 6860
rect 57848 6848 57854 6860
rect 58452 6857 58480 6888
rect 59722 6876 59728 6928
rect 59780 6916 59786 6928
rect 60737 6919 60795 6925
rect 60737 6916 60749 6919
rect 59780 6888 60749 6916
rect 59780 6876 59786 6888
rect 60737 6885 60749 6888
rect 60783 6885 60795 6919
rect 60737 6879 60795 6885
rect 58437 6851 58495 6857
rect 57848 6820 58388 6848
rect 57848 6808 57854 6820
rect 57057 6783 57115 6789
rect 57057 6780 57069 6783
rect 56244 6752 57069 6780
rect 56244 6712 56272 6752
rect 57057 6749 57069 6752
rect 57103 6749 57115 6783
rect 57057 6743 57115 6749
rect 57609 6783 57667 6789
rect 57609 6749 57621 6783
rect 57655 6780 57667 6783
rect 57974 6780 57980 6792
rect 57655 6752 57980 6780
rect 57655 6749 57667 6752
rect 57609 6743 57667 6749
rect 57974 6740 57980 6752
rect 58032 6740 58038 6792
rect 58161 6783 58219 6789
rect 58161 6749 58173 6783
rect 58207 6780 58219 6783
rect 58250 6780 58256 6792
rect 58207 6752 58256 6780
rect 58207 6749 58219 6752
rect 58161 6743 58219 6749
rect 58250 6740 58256 6752
rect 58308 6740 58314 6792
rect 58360 6780 58388 6820
rect 58437 6817 58449 6851
rect 58483 6848 58495 6851
rect 59265 6851 59323 6857
rect 59265 6848 59277 6851
rect 58483 6820 59277 6848
rect 58483 6817 58495 6820
rect 58437 6811 58495 6817
rect 59265 6817 59277 6820
rect 59311 6848 59323 6851
rect 59630 6848 59636 6860
rect 59311 6820 59636 6848
rect 59311 6817 59323 6820
rect 59265 6811 59323 6817
rect 59630 6808 59636 6820
rect 59688 6808 59694 6860
rect 59906 6848 59912 6860
rect 59867 6820 59912 6848
rect 59906 6808 59912 6820
rect 59964 6848 59970 6860
rect 60277 6851 60335 6857
rect 60277 6848 60289 6851
rect 59964 6820 60289 6848
rect 59964 6808 59970 6820
rect 60277 6817 60289 6820
rect 60323 6848 60335 6851
rect 60642 6848 60648 6860
rect 60323 6820 60648 6848
rect 60323 6817 60335 6820
rect 60277 6811 60335 6817
rect 60642 6808 60648 6820
rect 60700 6848 60706 6860
rect 61105 6851 61163 6857
rect 61105 6848 61117 6851
rect 60700 6820 61117 6848
rect 60700 6808 60706 6820
rect 61105 6817 61117 6820
rect 61151 6848 61163 6851
rect 61657 6851 61715 6857
rect 61657 6848 61669 6851
rect 61151 6820 61669 6848
rect 61151 6817 61163 6820
rect 61105 6811 61163 6817
rect 61657 6817 61669 6820
rect 61703 6817 61715 6851
rect 61657 6811 61715 6817
rect 58621 6783 58679 6789
rect 58621 6780 58633 6783
rect 58360 6752 58633 6780
rect 58621 6749 58633 6752
rect 58667 6780 58679 6783
rect 58897 6783 58955 6789
rect 58897 6780 58909 6783
rect 58667 6752 58909 6780
rect 58667 6749 58679 6752
rect 58621 6743 58679 6749
rect 58897 6749 58909 6752
rect 58943 6749 58955 6783
rect 58897 6743 58955 6749
rect 59998 6740 60004 6792
rect 60056 6780 60062 6792
rect 60185 6783 60243 6789
rect 60185 6780 60197 6783
rect 60056 6752 60197 6780
rect 60056 6740 60062 6752
rect 60185 6749 60197 6752
rect 60231 6749 60243 6783
rect 60185 6743 60243 6749
rect 61286 6740 61292 6792
rect 61344 6780 61350 6792
rect 61381 6783 61439 6789
rect 61381 6780 61393 6783
rect 61344 6752 61393 6780
rect 61344 6740 61350 6752
rect 61381 6749 61393 6752
rect 61427 6749 61439 6783
rect 61562 6780 61568 6792
rect 61523 6752 61568 6780
rect 61381 6743 61439 6749
rect 61562 6740 61568 6752
rect 61620 6740 61626 6792
rect 51224 6684 52776 6712
rect 53116 6684 56272 6712
rect 51224 6672 51230 6684
rect 53116 6644 53144 6684
rect 58526 6672 58532 6724
rect 58584 6712 58590 6724
rect 61304 6712 61332 6740
rect 58584 6684 61332 6712
rect 58584 6672 58590 6684
rect 53282 6644 53288 6656
rect 49804 6616 53144 6644
rect 53243 6616 53288 6644
rect 53282 6604 53288 6616
rect 53340 6604 53346 6656
rect 54018 6644 54024 6656
rect 53979 6616 54024 6644
rect 54018 6604 54024 6616
rect 54076 6604 54082 6656
rect 55582 6604 55588 6656
rect 55640 6644 55646 6656
rect 55858 6644 55864 6656
rect 55640 6616 55864 6644
rect 55640 6604 55646 6616
rect 55858 6604 55864 6616
rect 55916 6604 55922 6656
rect 55950 6604 55956 6656
rect 56008 6644 56014 6656
rect 56134 6644 56140 6656
rect 56008 6616 56140 6644
rect 56008 6604 56014 6616
rect 56134 6604 56140 6616
rect 56192 6644 56198 6656
rect 57606 6644 57612 6656
rect 56192 6616 57612 6644
rect 56192 6604 56198 6616
rect 57606 6604 57612 6616
rect 57664 6604 57670 6656
rect 58802 6604 58808 6656
rect 58860 6644 58866 6656
rect 61841 6647 61899 6653
rect 61841 6644 61853 6647
rect 58860 6616 61853 6644
rect 58860 6604 58866 6616
rect 61841 6613 61853 6616
rect 61887 6613 61899 6647
rect 61841 6607 61899 6613
rect 1104 6554 63480 6576
rect 1104 6502 11378 6554
rect 11430 6502 11442 6554
rect 11494 6502 11506 6554
rect 11558 6502 11570 6554
rect 11622 6502 32170 6554
rect 32222 6502 32234 6554
rect 32286 6502 32298 6554
rect 32350 6502 32362 6554
rect 32414 6502 52962 6554
rect 53014 6502 53026 6554
rect 53078 6502 53090 6554
rect 53142 6502 53154 6554
rect 53206 6502 63480 6554
rect 1104 6480 63480 6502
rect 4890 6400 4896 6452
rect 4948 6440 4954 6452
rect 5169 6443 5227 6449
rect 5169 6440 5181 6443
rect 4948 6412 5181 6440
rect 4948 6400 4954 6412
rect 5169 6409 5181 6412
rect 5215 6409 5227 6443
rect 5169 6403 5227 6409
rect 6273 6443 6331 6449
rect 6273 6409 6285 6443
rect 6319 6440 6331 6443
rect 6914 6440 6920 6452
rect 6319 6412 6920 6440
rect 6319 6409 6331 6412
rect 6273 6403 6331 6409
rect 4801 6375 4859 6381
rect 4801 6341 4813 6375
rect 4847 6372 4859 6375
rect 6288 6372 6316 6403
rect 6914 6400 6920 6412
rect 6972 6400 6978 6452
rect 7374 6400 7380 6452
rect 7432 6440 7438 6452
rect 8481 6443 8539 6449
rect 8481 6440 8493 6443
rect 7432 6412 8493 6440
rect 7432 6400 7438 6412
rect 8481 6409 8493 6412
rect 8527 6409 8539 6443
rect 8481 6403 8539 6409
rect 9306 6400 9312 6452
rect 9364 6440 9370 6452
rect 11701 6443 11759 6449
rect 11701 6440 11713 6443
rect 9364 6412 11713 6440
rect 9364 6400 9370 6412
rect 11701 6409 11713 6412
rect 11747 6409 11759 6443
rect 11701 6403 11759 6409
rect 13173 6443 13231 6449
rect 13173 6409 13185 6443
rect 13219 6440 13231 6443
rect 13906 6440 13912 6452
rect 13219 6412 13912 6440
rect 13219 6409 13231 6412
rect 13173 6403 13231 6409
rect 13906 6400 13912 6412
rect 13964 6400 13970 6452
rect 20162 6440 20168 6452
rect 17788 6412 20168 6440
rect 9125 6375 9183 6381
rect 9125 6372 9137 6375
rect 4847 6344 6316 6372
rect 8220 6344 9137 6372
rect 4847 6341 4859 6344
rect 4801 6335 4859 6341
rect 3510 6304 3516 6316
rect 3471 6276 3516 6304
rect 3510 6264 3516 6276
rect 3568 6264 3574 6316
rect 5905 6307 5963 6313
rect 5905 6273 5917 6307
rect 5951 6304 5963 6307
rect 6730 6304 6736 6316
rect 5951 6276 6736 6304
rect 5951 6273 5963 6276
rect 5905 6267 5963 6273
rect 6730 6264 6736 6276
rect 6788 6264 6794 6316
rect 8220 6313 8248 6344
rect 9125 6341 9137 6344
rect 9171 6372 9183 6375
rect 12710 6372 12716 6384
rect 9171 6344 12716 6372
rect 9171 6341 9183 6344
rect 9125 6335 9183 6341
rect 12710 6332 12716 6344
rect 12768 6332 12774 6384
rect 14461 6375 14519 6381
rect 14461 6341 14473 6375
rect 14507 6372 14519 6375
rect 16022 6372 16028 6384
rect 14507 6344 16028 6372
rect 14507 6341 14519 6344
rect 14461 6335 14519 6341
rect 16022 6332 16028 6344
rect 16080 6332 16086 6384
rect 16298 6332 16304 6384
rect 16356 6372 16362 6384
rect 17788 6372 17816 6412
rect 20162 6400 20168 6412
rect 20220 6400 20226 6452
rect 20714 6400 20720 6452
rect 20772 6440 20778 6452
rect 20772 6412 22048 6440
rect 20772 6400 20778 6412
rect 16356 6344 17816 6372
rect 17865 6375 17923 6381
rect 16356 6332 16362 6344
rect 17865 6341 17877 6375
rect 17911 6372 17923 6375
rect 18046 6372 18052 6384
rect 17911 6344 18052 6372
rect 17911 6341 17923 6344
rect 17865 6335 17923 6341
rect 18046 6332 18052 6344
rect 18104 6372 18110 6384
rect 19153 6375 19211 6381
rect 19153 6372 19165 6375
rect 18104 6344 19165 6372
rect 18104 6332 18110 6344
rect 19153 6341 19165 6344
rect 19199 6372 19211 6375
rect 19337 6375 19395 6381
rect 19337 6372 19349 6375
rect 19199 6344 19349 6372
rect 19199 6341 19211 6344
rect 19153 6335 19211 6341
rect 19337 6341 19349 6344
rect 19383 6341 19395 6375
rect 19978 6372 19984 6384
rect 19939 6344 19984 6372
rect 19337 6335 19395 6341
rect 19978 6332 19984 6344
rect 20036 6332 20042 6384
rect 20530 6372 20536 6384
rect 20088 6344 20536 6372
rect 7745 6307 7803 6313
rect 7745 6304 7757 6307
rect 7024 6276 7757 6304
rect 3234 6236 3240 6248
rect 2976 6208 3240 6236
rect 2314 6060 2320 6112
rect 2372 6100 2378 6112
rect 2976 6109 3004 6208
rect 3234 6196 3240 6208
rect 3292 6196 3298 6248
rect 7024 6245 7052 6276
rect 7745 6273 7757 6276
rect 7791 6304 7803 6307
rect 8205 6307 8263 6313
rect 8205 6304 8217 6307
rect 7791 6276 8217 6304
rect 7791 6273 7803 6276
rect 7745 6267 7803 6273
rect 8205 6273 8217 6276
rect 8251 6273 8263 6307
rect 10134 6304 10140 6316
rect 8205 6267 8263 6273
rect 9140 6276 9720 6304
rect 10095 6276 10140 6304
rect 7009 6239 7067 6245
rect 7009 6205 7021 6239
rect 7055 6205 7067 6239
rect 7009 6199 7067 6205
rect 8110 6196 8116 6248
rect 8168 6236 8174 6248
rect 8297 6239 8355 6245
rect 8297 6236 8309 6239
rect 8168 6208 8309 6236
rect 8168 6196 8174 6208
rect 8297 6205 8309 6208
rect 8343 6205 8355 6239
rect 8297 6199 8355 6205
rect 6549 6171 6607 6177
rect 6549 6137 6561 6171
rect 6595 6168 6607 6171
rect 6825 6171 6883 6177
rect 6825 6168 6837 6171
rect 6595 6140 6837 6168
rect 6595 6137 6607 6140
rect 6549 6131 6607 6137
rect 6825 6137 6837 6140
rect 6871 6168 6883 6171
rect 7190 6168 7196 6180
rect 6871 6140 7196 6168
rect 6871 6137 6883 6140
rect 6825 6131 6883 6137
rect 7190 6128 7196 6140
rect 7248 6128 7254 6180
rect 8202 6128 8208 6180
rect 8260 6168 8266 6180
rect 9140 6168 9168 6276
rect 9214 6196 9220 6248
rect 9272 6236 9278 6248
rect 9692 6245 9720 6276
rect 10134 6264 10140 6276
rect 10192 6264 10198 6316
rect 10778 6304 10784 6316
rect 10739 6276 10784 6304
rect 10778 6264 10784 6276
rect 10836 6264 10842 6316
rect 10965 6307 11023 6313
rect 10965 6273 10977 6307
rect 11011 6304 11023 6307
rect 11793 6307 11851 6313
rect 11793 6304 11805 6307
rect 11011 6276 11805 6304
rect 11011 6273 11023 6276
rect 10965 6267 11023 6273
rect 11793 6273 11805 6276
rect 11839 6304 11851 6307
rect 13541 6307 13599 6313
rect 11839 6276 13492 6304
rect 11839 6273 11851 6276
rect 11793 6267 11851 6273
rect 9585 6239 9643 6245
rect 9585 6236 9597 6239
rect 9272 6208 9597 6236
rect 9272 6196 9278 6208
rect 9401 6171 9459 6177
rect 9401 6168 9413 6171
rect 8260 6140 9413 6168
rect 8260 6128 8266 6140
rect 9401 6137 9413 6140
rect 9447 6137 9459 6171
rect 9508 6168 9536 6208
rect 9585 6205 9597 6208
rect 9631 6205 9643 6239
rect 9585 6199 9643 6205
rect 9677 6239 9735 6245
rect 9677 6205 9689 6239
rect 9723 6236 9735 6239
rect 9766 6236 9772 6248
rect 9723 6208 9772 6236
rect 9723 6205 9735 6208
rect 9677 6199 9735 6205
rect 9766 6196 9772 6208
rect 9824 6196 9830 6248
rect 11054 6236 11060 6248
rect 11015 6208 11060 6236
rect 11054 6196 11060 6208
rect 11112 6196 11118 6248
rect 11517 6239 11575 6245
rect 11517 6205 11529 6239
rect 11563 6236 11575 6239
rect 11974 6236 11980 6248
rect 11563 6208 11980 6236
rect 11563 6205 11575 6208
rect 11517 6199 11575 6205
rect 11974 6196 11980 6208
rect 12032 6196 12038 6248
rect 10413 6171 10471 6177
rect 10413 6168 10425 6171
rect 9508 6140 10425 6168
rect 9401 6131 9459 6137
rect 10413 6137 10425 6140
rect 10459 6137 10471 6171
rect 12434 6168 12440 6180
rect 10413 6131 10471 6137
rect 11624 6140 12440 6168
rect 2593 6103 2651 6109
rect 2593 6100 2605 6103
rect 2372 6072 2605 6100
rect 2372 6060 2378 6072
rect 2593 6069 2605 6072
rect 2639 6100 2651 6103
rect 2961 6103 3019 6109
rect 2961 6100 2973 6103
rect 2639 6072 2973 6100
rect 2639 6069 2651 6072
rect 2593 6063 2651 6069
rect 2961 6069 2973 6072
rect 3007 6069 3019 6103
rect 2961 6063 3019 6069
rect 6638 6060 6644 6112
rect 6696 6100 6702 6112
rect 7101 6103 7159 6109
rect 7101 6100 7113 6103
rect 6696 6072 7113 6100
rect 6696 6060 6702 6072
rect 7101 6069 7113 6072
rect 7147 6069 7159 6103
rect 7101 6063 7159 6069
rect 8113 6103 8171 6109
rect 8113 6069 8125 6103
rect 8159 6100 8171 6103
rect 8294 6100 8300 6112
rect 8159 6072 8300 6100
rect 8159 6069 8171 6072
rect 8113 6063 8171 6069
rect 8294 6060 8300 6072
rect 8352 6100 8358 6112
rect 9306 6100 9312 6112
rect 8352 6072 9312 6100
rect 8352 6060 8358 6072
rect 9306 6060 9312 6072
rect 9364 6060 9370 6112
rect 9490 6060 9496 6112
rect 9548 6100 9554 6112
rect 11624 6100 11652 6140
rect 12434 6128 12440 6140
rect 12492 6128 12498 6180
rect 13464 6168 13492 6276
rect 13541 6273 13553 6307
rect 13587 6304 13599 6307
rect 14366 6304 14372 6316
rect 13587 6276 14372 6304
rect 13587 6273 13599 6276
rect 13541 6267 13599 6273
rect 14366 6264 14372 6276
rect 14424 6304 14430 6316
rect 16209 6307 16267 6313
rect 16209 6304 16221 6307
rect 14424 6276 16221 6304
rect 14424 6264 14430 6276
rect 16209 6273 16221 6276
rect 16255 6273 16267 6307
rect 16209 6267 16267 6273
rect 16684 6276 17080 6304
rect 14645 6239 14703 6245
rect 14645 6205 14657 6239
rect 14691 6205 14703 6239
rect 15010 6236 15016 6248
rect 14971 6208 15016 6236
rect 14645 6199 14703 6205
rect 13538 6168 13544 6180
rect 13464 6140 13544 6168
rect 13538 6128 13544 6140
rect 13596 6128 13602 6180
rect 14660 6168 14688 6199
rect 15010 6196 15016 6208
rect 15068 6196 15074 6248
rect 15105 6239 15163 6245
rect 15105 6205 15117 6239
rect 15151 6236 15163 6239
rect 15746 6236 15752 6248
rect 15151 6208 15752 6236
rect 15151 6205 15163 6208
rect 15105 6199 15163 6205
rect 15746 6196 15752 6208
rect 15804 6236 15810 6248
rect 15841 6239 15899 6245
rect 15841 6236 15853 6239
rect 15804 6208 15853 6236
rect 15804 6196 15810 6208
rect 15841 6205 15853 6208
rect 15887 6205 15899 6239
rect 16114 6236 16120 6248
rect 16075 6208 16120 6236
rect 15841 6199 15899 6205
rect 16114 6196 16120 6208
rect 16172 6196 16178 6248
rect 15194 6168 15200 6180
rect 14660 6140 15200 6168
rect 15194 6128 15200 6140
rect 15252 6128 15258 6180
rect 15930 6128 15936 6180
rect 15988 6168 15994 6180
rect 16684 6168 16712 6276
rect 16758 6196 16764 6248
rect 16816 6245 16822 6248
rect 16816 6239 16865 6245
rect 16816 6205 16819 6239
rect 16853 6205 16865 6239
rect 16816 6199 16865 6205
rect 16945 6239 17003 6245
rect 16945 6205 16957 6239
rect 16991 6205 17003 6239
rect 17052 6236 17080 6276
rect 18230 6264 18236 6316
rect 18288 6304 18294 6316
rect 18601 6307 18659 6313
rect 18601 6304 18613 6307
rect 18288 6276 18613 6304
rect 18288 6264 18294 6276
rect 18601 6273 18613 6276
rect 18647 6304 18659 6307
rect 19426 6304 19432 6316
rect 18647 6276 19432 6304
rect 18647 6273 18659 6276
rect 18601 6267 18659 6273
rect 19426 6264 19432 6276
rect 19484 6264 19490 6316
rect 19797 6307 19855 6313
rect 19797 6273 19809 6307
rect 19843 6304 19855 6307
rect 20088 6304 20116 6344
rect 20530 6332 20536 6344
rect 20588 6332 20594 6384
rect 22020 6372 22048 6412
rect 25774 6400 25780 6452
rect 25832 6440 25838 6452
rect 31938 6440 31944 6452
rect 25832 6412 31944 6440
rect 25832 6400 25838 6412
rect 31938 6400 31944 6412
rect 31996 6400 32002 6452
rect 33870 6440 33876 6452
rect 33831 6412 33876 6440
rect 33870 6400 33876 6412
rect 33928 6400 33934 6452
rect 34425 6443 34483 6449
rect 34425 6409 34437 6443
rect 34471 6440 34483 6443
rect 34701 6443 34759 6449
rect 34701 6440 34713 6443
rect 34471 6412 34713 6440
rect 34471 6409 34483 6412
rect 34425 6403 34483 6409
rect 34701 6409 34713 6412
rect 34747 6440 34759 6443
rect 41969 6443 42027 6449
rect 34747 6412 41000 6440
rect 34747 6409 34759 6412
rect 34701 6403 34759 6409
rect 34900 6384 34928 6412
rect 22922 6372 22928 6384
rect 22020 6344 22928 6372
rect 22922 6332 22928 6344
rect 22980 6332 22986 6384
rect 23937 6375 23995 6381
rect 23937 6341 23949 6375
rect 23983 6372 23995 6375
rect 24026 6372 24032 6384
rect 23983 6344 24032 6372
rect 23983 6341 23995 6344
rect 23937 6335 23995 6341
rect 24026 6332 24032 6344
rect 24084 6332 24090 6384
rect 24397 6375 24455 6381
rect 24397 6341 24409 6375
rect 24443 6372 24455 6375
rect 24854 6372 24860 6384
rect 24443 6344 24860 6372
rect 24443 6341 24455 6344
rect 24397 6335 24455 6341
rect 19843 6276 20116 6304
rect 19843 6273 19855 6276
rect 19797 6267 19855 6273
rect 17052 6208 17632 6236
rect 16945 6199 17003 6205
rect 16816 6196 16822 6199
rect 15988 6140 16712 6168
rect 16960 6168 16988 6199
rect 16960 6140 17172 6168
rect 15988 6128 15994 6140
rect 17144 6112 17172 6140
rect 9548 6072 11652 6100
rect 11701 6103 11759 6109
rect 9548 6060 9554 6072
rect 11701 6069 11713 6103
rect 11747 6100 11759 6103
rect 12253 6103 12311 6109
rect 12253 6100 12265 6103
rect 11747 6072 12265 6100
rect 11747 6069 11759 6072
rect 11701 6063 11759 6069
rect 12253 6069 12265 6072
rect 12299 6100 12311 6103
rect 12526 6100 12532 6112
rect 12299 6072 12532 6100
rect 12299 6069 12311 6072
rect 12253 6063 12311 6069
rect 12526 6060 12532 6072
rect 12584 6060 12590 6112
rect 12805 6103 12863 6109
rect 12805 6069 12817 6103
rect 12851 6100 12863 6103
rect 13170 6100 13176 6112
rect 12851 6072 13176 6100
rect 12851 6069 12863 6072
rect 12805 6063 12863 6069
rect 13170 6060 13176 6072
rect 13228 6060 13234 6112
rect 13814 6060 13820 6112
rect 13872 6100 13878 6112
rect 13909 6103 13967 6109
rect 13909 6100 13921 6103
rect 13872 6072 13921 6100
rect 13872 6060 13878 6072
rect 13909 6069 13921 6072
rect 13955 6100 13967 6103
rect 14642 6100 14648 6112
rect 13955 6072 14648 6100
rect 13955 6069 13967 6072
rect 13909 6063 13967 6069
rect 14642 6060 14648 6072
rect 14700 6060 14706 6112
rect 15010 6060 15016 6112
rect 15068 6100 15074 6112
rect 15565 6103 15623 6109
rect 15565 6100 15577 6103
rect 15068 6072 15577 6100
rect 15068 6060 15074 6072
rect 15565 6069 15577 6072
rect 15611 6100 15623 6103
rect 16114 6100 16120 6112
rect 15611 6072 16120 6100
rect 15611 6069 15623 6072
rect 15565 6063 15623 6069
rect 16114 6060 16120 6072
rect 16172 6060 16178 6112
rect 17126 6060 17132 6112
rect 17184 6100 17190 6112
rect 17402 6100 17408 6112
rect 17184 6072 17408 6100
rect 17184 6060 17190 6072
rect 17402 6060 17408 6072
rect 17460 6060 17466 6112
rect 17604 6100 17632 6208
rect 17954 6196 17960 6248
rect 18012 6236 18018 6248
rect 18690 6236 18696 6248
rect 18012 6208 18696 6236
rect 18012 6196 18018 6208
rect 18690 6196 18696 6208
rect 18748 6236 18754 6248
rect 18877 6239 18935 6245
rect 18877 6236 18889 6239
rect 18748 6208 18889 6236
rect 18748 6196 18754 6208
rect 18877 6205 18889 6208
rect 18923 6205 18935 6239
rect 19058 6236 19064 6248
rect 18971 6208 19064 6236
rect 18877 6199 18935 6205
rect 19058 6196 19064 6208
rect 19116 6236 19122 6248
rect 19153 6239 19211 6245
rect 19153 6236 19165 6239
rect 19116 6208 19165 6236
rect 19116 6196 19122 6208
rect 19153 6205 19165 6208
rect 19199 6205 19211 6239
rect 19153 6199 19211 6205
rect 19334 6196 19340 6248
rect 19392 6236 19398 6248
rect 19812 6236 19840 6267
rect 22646 6264 22652 6316
rect 22704 6304 22710 6316
rect 22741 6307 22799 6313
rect 22741 6304 22753 6307
rect 22704 6276 22753 6304
rect 22704 6264 22710 6276
rect 22741 6273 22753 6276
rect 22787 6304 22799 6307
rect 24412 6304 24440 6335
rect 24854 6332 24860 6344
rect 24912 6372 24918 6384
rect 28350 6372 28356 6384
rect 24912 6344 28356 6372
rect 24912 6332 24918 6344
rect 28350 6332 28356 6344
rect 28408 6332 28414 6384
rect 31478 6332 31484 6384
rect 31536 6372 31542 6384
rect 31536 6344 34836 6372
rect 31536 6332 31542 6344
rect 22787 6276 24440 6304
rect 24489 6307 24547 6313
rect 22787 6273 22799 6276
rect 22741 6267 22799 6273
rect 24489 6273 24501 6307
rect 24535 6273 24547 6307
rect 24489 6267 24547 6273
rect 19392 6208 19840 6236
rect 20073 6239 20131 6245
rect 19392 6196 19398 6208
rect 20073 6205 20085 6239
rect 20119 6236 20131 6239
rect 20162 6236 20168 6248
rect 20119 6208 20168 6236
rect 20119 6205 20131 6208
rect 20073 6199 20131 6205
rect 20162 6196 20168 6208
rect 20220 6196 20226 6248
rect 20530 6236 20536 6248
rect 20491 6208 20536 6236
rect 20530 6196 20536 6208
rect 20588 6196 20594 6248
rect 20622 6196 20628 6248
rect 20680 6236 20686 6248
rect 21085 6239 21143 6245
rect 21085 6236 21097 6239
rect 20680 6208 21097 6236
rect 20680 6196 20686 6208
rect 21085 6205 21097 6208
rect 21131 6205 21143 6239
rect 21634 6236 21640 6248
rect 21595 6208 21640 6236
rect 21085 6199 21143 6205
rect 21634 6196 21640 6208
rect 21692 6236 21698 6248
rect 22281 6239 22339 6245
rect 22281 6236 22293 6239
rect 21692 6208 22293 6236
rect 21692 6196 21698 6208
rect 22281 6205 22293 6208
rect 22327 6205 22339 6239
rect 22281 6199 22339 6205
rect 23109 6239 23167 6245
rect 23109 6205 23121 6239
rect 23155 6236 23167 6239
rect 23750 6236 23756 6248
rect 23155 6208 23756 6236
rect 23155 6205 23167 6208
rect 23109 6199 23167 6205
rect 23750 6196 23756 6208
rect 23808 6196 23814 6248
rect 18046 6168 18052 6180
rect 18007 6140 18052 6168
rect 18046 6128 18052 6140
rect 18104 6128 18110 6180
rect 18230 6128 18236 6180
rect 18288 6168 18294 6180
rect 21453 6171 21511 6177
rect 18288 6140 21036 6168
rect 18288 6128 18294 6140
rect 20898 6100 20904 6112
rect 17604 6072 20904 6100
rect 20898 6060 20904 6072
rect 20956 6060 20962 6112
rect 21008 6100 21036 6140
rect 21453 6137 21465 6171
rect 21499 6168 21511 6171
rect 21818 6168 21824 6180
rect 21499 6140 21824 6168
rect 21499 6137 21511 6140
rect 21453 6131 21511 6137
rect 21818 6128 21824 6140
rect 21876 6128 21882 6180
rect 24504 6168 24532 6267
rect 24578 6264 24584 6316
rect 24636 6304 24642 6316
rect 25041 6307 25099 6313
rect 25041 6304 25053 6307
rect 24636 6276 25053 6304
rect 24636 6264 24642 6276
rect 25041 6273 25053 6276
rect 25087 6304 25099 6307
rect 25130 6304 25136 6316
rect 25087 6276 25136 6304
rect 25087 6273 25099 6276
rect 25041 6267 25099 6273
rect 25130 6264 25136 6276
rect 25188 6264 25194 6316
rect 26329 6307 26387 6313
rect 26329 6304 26341 6307
rect 25332 6276 26341 6304
rect 25332 6248 25360 6276
rect 26329 6273 26341 6276
rect 26375 6304 26387 6307
rect 26510 6304 26516 6316
rect 26375 6276 26516 6304
rect 26375 6273 26387 6276
rect 26329 6267 26387 6273
rect 26510 6264 26516 6276
rect 26568 6264 26574 6316
rect 27614 6304 27620 6316
rect 26896 6276 27620 6304
rect 25314 6236 25320 6248
rect 25227 6208 25320 6236
rect 25314 6196 25320 6208
rect 25372 6196 25378 6248
rect 25501 6239 25559 6245
rect 25501 6205 25513 6239
rect 25547 6236 25559 6239
rect 25590 6236 25596 6248
rect 25547 6208 25596 6236
rect 25547 6205 25559 6208
rect 25501 6199 25559 6205
rect 25590 6196 25596 6208
rect 25648 6236 25654 6248
rect 25777 6239 25835 6245
rect 25777 6236 25789 6239
rect 25648 6208 25789 6236
rect 25648 6196 25654 6208
rect 25777 6205 25789 6208
rect 25823 6205 25835 6239
rect 25777 6199 25835 6205
rect 25866 6196 25872 6248
rect 25924 6236 25930 6248
rect 26896 6245 26924 6276
rect 27614 6264 27620 6276
rect 27672 6264 27678 6316
rect 28442 6304 28448 6316
rect 27724 6276 28448 6304
rect 26881 6239 26939 6245
rect 26881 6236 26893 6239
rect 25924 6208 26893 6236
rect 25924 6196 25930 6208
rect 26881 6205 26893 6208
rect 26927 6205 26939 6239
rect 26881 6199 26939 6205
rect 27062 6196 27068 6248
rect 27120 6236 27126 6248
rect 27157 6239 27215 6245
rect 27157 6236 27169 6239
rect 27120 6208 27169 6236
rect 27120 6196 27126 6208
rect 27157 6205 27169 6208
rect 27203 6205 27215 6239
rect 27157 6199 27215 6205
rect 27341 6239 27399 6245
rect 27341 6205 27353 6239
rect 27387 6236 27399 6239
rect 27433 6239 27491 6245
rect 27433 6236 27445 6239
rect 27387 6208 27445 6236
rect 27387 6205 27399 6208
rect 27341 6199 27399 6205
rect 27433 6205 27445 6208
rect 27479 6236 27491 6239
rect 27724 6236 27752 6276
rect 28442 6264 28448 6276
rect 28500 6264 28506 6316
rect 28718 6304 28724 6316
rect 28679 6276 28724 6304
rect 28718 6264 28724 6276
rect 28776 6264 28782 6316
rect 29546 6304 29552 6316
rect 29507 6276 29552 6304
rect 29546 6264 29552 6276
rect 29604 6264 29610 6316
rect 31662 6264 31668 6316
rect 31720 6304 31726 6316
rect 32217 6307 32275 6313
rect 32217 6304 32229 6307
rect 31720 6276 32229 6304
rect 31720 6264 31726 6276
rect 32217 6273 32229 6276
rect 32263 6273 32275 6307
rect 32217 6267 32275 6273
rect 33229 6307 33287 6313
rect 33229 6273 33241 6307
rect 33275 6304 33287 6307
rect 34425 6307 34483 6313
rect 34425 6304 34437 6307
rect 33275 6276 34437 6304
rect 33275 6273 33287 6276
rect 33229 6267 33287 6273
rect 34425 6273 34437 6276
rect 34471 6273 34483 6307
rect 34808 6304 34836 6344
rect 34882 6332 34888 6384
rect 34940 6372 34946 6384
rect 37918 6372 37924 6384
rect 34940 6344 35033 6372
rect 35452 6344 37780 6372
rect 37879 6344 37924 6372
rect 34940 6332 34946 6344
rect 35452 6304 35480 6344
rect 34808 6276 35480 6304
rect 34425 6267 34483 6273
rect 35526 6264 35532 6316
rect 35584 6304 35590 6316
rect 37093 6307 37151 6313
rect 37093 6304 37105 6307
rect 35584 6276 37105 6304
rect 35584 6264 35590 6276
rect 27479 6208 27752 6236
rect 27479 6205 27491 6208
rect 27433 6199 27491 6205
rect 27798 6196 27804 6248
rect 27856 6236 27862 6248
rect 28169 6239 28227 6245
rect 28169 6236 28181 6239
rect 27856 6208 28181 6236
rect 27856 6196 27862 6208
rect 28169 6205 28181 6208
rect 28215 6236 28227 6239
rect 28736 6236 28764 6264
rect 28215 6208 28764 6236
rect 29273 6239 29331 6245
rect 28215 6205 28227 6208
rect 28169 6199 28227 6205
rect 29273 6205 29285 6239
rect 29319 6236 29331 6239
rect 30006 6236 30012 6248
rect 29319 6208 30012 6236
rect 29319 6205 29331 6208
rect 29273 6199 29331 6205
rect 30006 6196 30012 6208
rect 30064 6196 30070 6248
rect 31294 6236 31300 6248
rect 31255 6208 31300 6236
rect 31294 6196 31300 6208
rect 31352 6196 31358 6248
rect 31757 6239 31815 6245
rect 31757 6205 31769 6239
rect 31803 6205 31815 6239
rect 31757 6199 31815 6205
rect 31849 6239 31907 6245
rect 31849 6205 31861 6239
rect 31895 6205 31907 6239
rect 32030 6236 32036 6248
rect 31991 6208 32036 6236
rect 31849 6199 31907 6205
rect 24854 6168 24860 6180
rect 24504 6140 24860 6168
rect 24854 6128 24860 6140
rect 24912 6128 24918 6180
rect 28258 6168 28264 6180
rect 28171 6140 28264 6168
rect 28258 6128 28264 6140
rect 28316 6168 28322 6180
rect 28810 6168 28816 6180
rect 28316 6140 28816 6168
rect 28316 6128 28322 6140
rect 28810 6128 28816 6140
rect 28868 6128 28874 6180
rect 29086 6168 29092 6180
rect 29047 6140 29092 6168
rect 29086 6128 29092 6140
rect 29144 6128 29150 6180
rect 30929 6171 30987 6177
rect 30929 6137 30941 6171
rect 30975 6168 30987 6171
rect 31662 6168 31668 6180
rect 30975 6140 31668 6168
rect 30975 6137 30987 6140
rect 30929 6131 30987 6137
rect 31662 6128 31668 6140
rect 31720 6128 31726 6180
rect 21729 6103 21787 6109
rect 21729 6100 21741 6103
rect 21008 6072 21741 6100
rect 21729 6069 21741 6072
rect 21775 6069 21787 6103
rect 21729 6063 21787 6069
rect 23477 6103 23535 6109
rect 23477 6069 23489 6103
rect 23523 6100 23535 6103
rect 23658 6100 23664 6112
rect 23523 6072 23664 6100
rect 23523 6069 23535 6072
rect 23477 6063 23535 6069
rect 23658 6060 23664 6072
rect 23716 6100 23722 6112
rect 24486 6100 24492 6112
rect 23716 6072 24492 6100
rect 23716 6060 23722 6072
rect 24486 6060 24492 6072
rect 24544 6060 24550 6112
rect 26237 6103 26295 6109
rect 26237 6069 26249 6103
rect 26283 6100 26295 6103
rect 26786 6100 26792 6112
rect 26283 6072 26792 6100
rect 26283 6069 26295 6072
rect 26237 6063 26295 6069
rect 26786 6060 26792 6072
rect 26844 6100 26850 6112
rect 27433 6103 27491 6109
rect 27433 6100 27445 6103
rect 26844 6072 27445 6100
rect 26844 6060 26850 6072
rect 27433 6069 27445 6072
rect 27479 6100 27491 6103
rect 27617 6103 27675 6109
rect 27617 6100 27629 6103
rect 27479 6072 27629 6100
rect 27479 6069 27491 6072
rect 27433 6063 27491 6069
rect 27617 6069 27629 6072
rect 27663 6069 27675 6103
rect 27617 6063 27675 6069
rect 27706 6060 27712 6112
rect 27764 6100 27770 6112
rect 27985 6103 28043 6109
rect 27985 6100 27997 6103
rect 27764 6072 27997 6100
rect 27764 6060 27770 6072
rect 27985 6069 27997 6072
rect 28031 6100 28043 6103
rect 31386 6100 31392 6112
rect 28031 6072 31392 6100
rect 28031 6069 28043 6072
rect 27985 6063 28043 6069
rect 31386 6060 31392 6072
rect 31444 6060 31450 6112
rect 31478 6060 31484 6112
rect 31536 6100 31542 6112
rect 31573 6103 31631 6109
rect 31573 6100 31585 6103
rect 31536 6072 31585 6100
rect 31536 6060 31542 6072
rect 31573 6069 31585 6072
rect 31619 6069 31631 6103
rect 31772 6100 31800 6199
rect 31864 6168 31892 6199
rect 32030 6196 32036 6208
rect 32088 6196 32094 6248
rect 33689 6239 33747 6245
rect 33689 6236 33701 6239
rect 33520 6208 33701 6236
rect 31938 6168 31944 6180
rect 31864 6140 31944 6168
rect 31938 6128 31944 6140
rect 31996 6128 32002 6180
rect 33520 6112 33548 6208
rect 33689 6205 33701 6208
rect 33735 6205 33747 6239
rect 34238 6236 34244 6248
rect 34199 6208 34244 6236
rect 33689 6199 33747 6205
rect 34238 6196 34244 6208
rect 34296 6196 34302 6248
rect 35618 6236 35624 6248
rect 35579 6208 35624 6236
rect 35618 6196 35624 6208
rect 35676 6196 35682 6248
rect 35986 6236 35992 6248
rect 35947 6208 35992 6236
rect 35986 6196 35992 6208
rect 36044 6196 36050 6248
rect 36188 6245 36216 6276
rect 37093 6273 37105 6276
rect 37139 6273 37151 6307
rect 37093 6267 37151 6273
rect 37752 6245 37780 6344
rect 37918 6332 37924 6344
rect 37976 6332 37982 6384
rect 39577 6375 39635 6381
rect 38304 6344 39528 6372
rect 38304 6245 38332 6344
rect 39390 6304 39396 6316
rect 38396 6276 39252 6304
rect 39351 6276 39396 6304
rect 36173 6239 36231 6245
rect 36173 6205 36185 6239
rect 36219 6205 36231 6239
rect 36173 6199 36231 6205
rect 36541 6239 36599 6245
rect 36541 6205 36553 6239
rect 36587 6205 36599 6239
rect 36541 6199 36599 6205
rect 37737 6239 37795 6245
rect 37737 6205 37749 6239
rect 37783 6236 37795 6239
rect 38289 6239 38347 6245
rect 38289 6236 38301 6239
rect 37783 6208 38301 6236
rect 37783 6205 37795 6208
rect 37737 6199 37795 6205
rect 38289 6205 38301 6208
rect 38335 6205 38347 6239
rect 38289 6199 38347 6205
rect 35250 6168 35256 6180
rect 35211 6140 35256 6168
rect 35250 6128 35256 6140
rect 35308 6128 35314 6180
rect 35710 6128 35716 6180
rect 35768 6168 35774 6180
rect 36556 6168 36584 6199
rect 37461 6171 37519 6177
rect 37461 6168 37473 6171
rect 35768 6140 37473 6168
rect 35768 6128 35774 6140
rect 37461 6137 37473 6140
rect 37507 6137 37519 6171
rect 37461 6131 37519 6137
rect 31846 6100 31852 6112
rect 31772 6072 31852 6100
rect 31573 6063 31631 6069
rect 31846 6060 31852 6072
rect 31904 6060 31910 6112
rect 32490 6060 32496 6112
rect 32548 6100 32554 6112
rect 32769 6103 32827 6109
rect 32769 6100 32781 6103
rect 32548 6072 32781 6100
rect 32548 6060 32554 6072
rect 32769 6069 32781 6072
rect 32815 6069 32827 6103
rect 33502 6100 33508 6112
rect 33463 6072 33508 6100
rect 32769 6063 32827 6069
rect 33502 6060 33508 6072
rect 33560 6060 33566 6112
rect 34606 6060 34612 6112
rect 34664 6100 34670 6112
rect 38396 6100 38424 6276
rect 38654 6236 38660 6248
rect 38615 6208 38660 6236
rect 38654 6196 38660 6208
rect 38712 6236 38718 6248
rect 38841 6239 38899 6245
rect 38841 6236 38853 6239
rect 38712 6208 38853 6236
rect 38712 6196 38718 6208
rect 38841 6205 38853 6208
rect 38887 6205 38899 6239
rect 38841 6199 38899 6205
rect 38930 6196 38936 6248
rect 38988 6236 38994 6248
rect 39025 6239 39083 6245
rect 39025 6236 39037 6239
rect 38988 6208 39037 6236
rect 38988 6196 38994 6208
rect 39025 6205 39037 6208
rect 39071 6205 39083 6239
rect 39224 6236 39252 6276
rect 39390 6264 39396 6276
rect 39448 6264 39454 6316
rect 39500 6304 39528 6344
rect 39577 6341 39589 6375
rect 39623 6372 39635 6375
rect 40494 6372 40500 6384
rect 39623 6344 40500 6372
rect 39623 6341 39635 6344
rect 39577 6335 39635 6341
rect 40494 6332 40500 6344
rect 40552 6332 40558 6384
rect 40972 6372 41000 6412
rect 41969 6409 41981 6443
rect 42015 6440 42027 6443
rect 42426 6440 42432 6452
rect 42015 6412 42432 6440
rect 42015 6409 42027 6412
rect 41969 6403 42027 6409
rect 42426 6400 42432 6412
rect 42484 6400 42490 6452
rect 42886 6400 42892 6452
rect 42944 6440 42950 6452
rect 43349 6443 43407 6449
rect 43349 6440 43361 6443
rect 42944 6412 43361 6440
rect 42944 6400 42950 6412
rect 43349 6409 43361 6412
rect 43395 6409 43407 6443
rect 43349 6403 43407 6409
rect 45005 6443 45063 6449
rect 45005 6409 45017 6443
rect 45051 6440 45063 6443
rect 45281 6443 45339 6449
rect 45281 6440 45293 6443
rect 45051 6412 45293 6440
rect 45051 6409 45063 6412
rect 45005 6403 45063 6409
rect 45281 6409 45293 6412
rect 45327 6440 45339 6443
rect 45554 6440 45560 6452
rect 45327 6412 45560 6440
rect 45327 6409 45339 6412
rect 45281 6403 45339 6409
rect 45554 6400 45560 6412
rect 45612 6400 45618 6452
rect 46198 6400 46204 6452
rect 46256 6440 46262 6452
rect 46256 6412 47164 6440
rect 46256 6400 46262 6412
rect 47029 6375 47087 6381
rect 47029 6372 47041 6375
rect 40972 6344 47041 6372
rect 47029 6341 47041 6344
rect 47075 6341 47087 6375
rect 47136 6372 47164 6412
rect 47302 6400 47308 6452
rect 47360 6440 47366 6452
rect 47946 6440 47952 6452
rect 47360 6412 47952 6440
rect 47360 6400 47366 6412
rect 47946 6400 47952 6412
rect 48004 6400 48010 6452
rect 48498 6400 48504 6452
rect 48556 6440 48562 6452
rect 48869 6443 48927 6449
rect 48869 6440 48881 6443
rect 48556 6412 48881 6440
rect 48556 6400 48562 6412
rect 48869 6409 48881 6412
rect 48915 6409 48927 6443
rect 48869 6403 48927 6409
rect 48976 6412 50292 6440
rect 47489 6375 47547 6381
rect 47489 6372 47501 6375
rect 47136 6344 47501 6372
rect 47029 6335 47087 6341
rect 47489 6341 47501 6344
rect 47535 6372 47547 6375
rect 47581 6375 47639 6381
rect 47581 6372 47593 6375
rect 47535 6344 47593 6372
rect 47535 6341 47547 6344
rect 47489 6335 47547 6341
rect 47581 6341 47593 6344
rect 47627 6341 47639 6375
rect 48976 6372 49004 6412
rect 47581 6335 47639 6341
rect 47688 6344 49004 6372
rect 50264 6372 50292 6412
rect 50338 6400 50344 6452
rect 50396 6440 50402 6452
rect 50433 6443 50491 6449
rect 50433 6440 50445 6443
rect 50396 6412 50445 6440
rect 50396 6400 50402 6412
rect 50433 6409 50445 6412
rect 50479 6409 50491 6443
rect 50985 6443 51043 6449
rect 50985 6440 50997 6443
rect 50433 6403 50491 6409
rect 50540 6412 50997 6440
rect 50540 6372 50568 6412
rect 50985 6409 50997 6412
rect 51031 6409 51043 6443
rect 50985 6403 51043 6409
rect 52178 6400 52184 6452
rect 52236 6440 52242 6452
rect 54573 6443 54631 6449
rect 52236 6412 54524 6440
rect 52236 6400 52242 6412
rect 50264 6344 50568 6372
rect 42058 6304 42064 6316
rect 39500 6276 42064 6304
rect 42058 6264 42064 6276
rect 42116 6264 42122 6316
rect 43901 6307 43959 6313
rect 42536 6276 43852 6304
rect 40681 6239 40739 6245
rect 40681 6236 40693 6239
rect 39224 6208 40693 6236
rect 39025 6199 39083 6205
rect 40681 6205 40693 6208
rect 40727 6236 40739 6239
rect 41325 6239 41383 6245
rect 41325 6236 41337 6239
rect 40727 6208 41337 6236
rect 40727 6205 40739 6208
rect 40681 6199 40739 6205
rect 41325 6205 41337 6208
rect 41371 6205 41383 6239
rect 41325 6199 41383 6205
rect 41785 6239 41843 6245
rect 41785 6205 41797 6239
rect 41831 6236 41843 6239
rect 41874 6236 41880 6248
rect 41831 6208 41880 6236
rect 41831 6205 41843 6208
rect 41785 6199 41843 6205
rect 39040 6168 39068 6199
rect 41874 6196 41880 6208
rect 41932 6196 41938 6248
rect 42426 6196 42432 6248
rect 42484 6245 42490 6248
rect 42484 6239 42501 6245
rect 42489 6205 42501 6239
rect 42484 6199 42501 6205
rect 42484 6196 42490 6199
rect 39577 6171 39635 6177
rect 39577 6168 39589 6171
rect 39040 6140 39589 6168
rect 39577 6137 39589 6140
rect 39623 6168 39635 6171
rect 39669 6171 39727 6177
rect 39669 6168 39681 6171
rect 39623 6140 39681 6168
rect 39623 6137 39635 6140
rect 39577 6131 39635 6137
rect 39669 6137 39681 6140
rect 39715 6137 39727 6171
rect 40494 6168 40500 6180
rect 39669 6131 39727 6137
rect 40236 6140 40500 6168
rect 34664 6072 38424 6100
rect 34664 6060 34670 6072
rect 39482 6060 39488 6112
rect 39540 6100 39546 6112
rect 40236 6109 40264 6140
rect 40494 6128 40500 6140
rect 40552 6128 40558 6180
rect 41049 6171 41107 6177
rect 41049 6137 41061 6171
rect 41095 6168 41107 6171
rect 42536 6168 42564 6276
rect 42613 6239 42671 6245
rect 42613 6205 42625 6239
rect 42659 6205 42671 6239
rect 42886 6236 42892 6248
rect 42847 6208 42892 6236
rect 42613 6199 42671 6205
rect 41095 6140 42564 6168
rect 42628 6168 42656 6199
rect 42886 6196 42892 6208
rect 42944 6196 42950 6248
rect 43073 6239 43131 6245
rect 43073 6205 43085 6239
rect 43119 6236 43131 6239
rect 43346 6236 43352 6248
rect 43119 6208 43352 6236
rect 43119 6205 43131 6208
rect 43073 6199 43131 6205
rect 43346 6196 43352 6208
rect 43404 6196 43410 6248
rect 43824 6236 43852 6276
rect 43901 6273 43913 6307
rect 43947 6304 43959 6307
rect 44082 6304 44088 6316
rect 43947 6276 44088 6304
rect 43947 6273 43959 6276
rect 43901 6267 43959 6273
rect 44082 6264 44088 6276
rect 44140 6304 44146 6316
rect 44634 6304 44640 6316
rect 44140 6276 44640 6304
rect 44140 6264 44146 6276
rect 44634 6264 44640 6276
rect 44692 6264 44698 6316
rect 44913 6307 44971 6313
rect 44913 6273 44925 6307
rect 44959 6304 44971 6307
rect 45005 6307 45063 6313
rect 45005 6304 45017 6307
rect 44959 6276 45017 6304
rect 44959 6273 44971 6276
rect 44913 6267 44971 6273
rect 45005 6273 45017 6276
rect 45051 6273 45063 6307
rect 47688 6304 47716 6344
rect 50614 6332 50620 6384
rect 50672 6372 50678 6384
rect 51169 6375 51227 6381
rect 51169 6372 51181 6375
rect 50672 6344 51181 6372
rect 50672 6332 50678 6344
rect 51169 6341 51181 6344
rect 51215 6341 51227 6375
rect 54496 6372 54524 6412
rect 54573 6409 54585 6443
rect 54619 6440 54631 6443
rect 54754 6440 54760 6452
rect 54619 6412 54760 6440
rect 54619 6409 54631 6412
rect 54573 6403 54631 6409
rect 54754 6400 54760 6412
rect 54812 6400 54818 6452
rect 54938 6440 54944 6452
rect 54899 6412 54944 6440
rect 54938 6400 54944 6412
rect 54996 6400 55002 6452
rect 55401 6443 55459 6449
rect 55401 6409 55413 6443
rect 55447 6440 55459 6443
rect 55490 6440 55496 6452
rect 55447 6412 55496 6440
rect 55447 6409 55459 6412
rect 55401 6403 55459 6409
rect 55490 6400 55496 6412
rect 55548 6440 55554 6452
rect 55766 6440 55772 6452
rect 55548 6412 55772 6440
rect 55548 6400 55554 6412
rect 55766 6400 55772 6412
rect 55824 6400 55830 6452
rect 57149 6443 57207 6449
rect 57149 6409 57161 6443
rect 57195 6440 57207 6443
rect 57698 6440 57704 6452
rect 57195 6412 57704 6440
rect 57195 6409 57207 6412
rect 57149 6403 57207 6409
rect 57698 6400 57704 6412
rect 57756 6400 57762 6452
rect 57790 6400 57796 6452
rect 57848 6440 57854 6452
rect 59449 6443 59507 6449
rect 59449 6440 59461 6443
rect 57848 6412 59461 6440
rect 57848 6400 57854 6412
rect 59449 6409 59461 6412
rect 59495 6409 59507 6443
rect 59449 6403 59507 6409
rect 55217 6375 55275 6381
rect 55217 6372 55229 6375
rect 54496 6344 55229 6372
rect 51169 6335 51227 6341
rect 55217 6341 55229 6344
rect 55263 6341 55275 6375
rect 55217 6335 55275 6341
rect 55677 6375 55735 6381
rect 55677 6341 55689 6375
rect 55723 6372 55735 6375
rect 56594 6372 56600 6384
rect 55723 6344 56600 6372
rect 55723 6341 55735 6344
rect 55677 6335 55735 6341
rect 56594 6332 56600 6344
rect 56652 6332 56658 6384
rect 48317 6307 48375 6313
rect 48317 6304 48329 6307
rect 45005 6267 45063 6273
rect 45480 6276 47716 6304
rect 47780 6276 48329 6304
rect 44358 6236 44364 6248
rect 43824 6208 44364 6236
rect 44358 6196 44364 6208
rect 44416 6196 44422 6248
rect 44453 6239 44511 6245
rect 44453 6205 44465 6239
rect 44499 6205 44511 6239
rect 44726 6236 44732 6248
rect 44687 6208 44732 6236
rect 44453 6199 44511 6205
rect 42978 6168 42984 6180
rect 42628 6140 42984 6168
rect 41095 6137 41107 6140
rect 41049 6131 41107 6137
rect 42978 6128 42984 6140
rect 43036 6128 43042 6180
rect 43714 6168 43720 6180
rect 43675 6140 43720 6168
rect 43714 6128 43720 6140
rect 43772 6168 43778 6180
rect 44468 6168 44496 6199
rect 44726 6196 44732 6208
rect 44784 6196 44790 6248
rect 45480 6236 45508 6276
rect 44928 6208 45508 6236
rect 44928 6180 44956 6208
rect 46106 6196 46112 6248
rect 46164 6236 46170 6248
rect 46201 6239 46259 6245
rect 46201 6236 46213 6239
rect 46164 6208 46213 6236
rect 46164 6196 46170 6208
rect 46201 6205 46213 6208
rect 46247 6205 46259 6239
rect 46201 6199 46259 6205
rect 46290 6196 46296 6248
rect 46348 6236 46354 6248
rect 46477 6239 46535 6245
rect 46477 6236 46489 6239
rect 46348 6208 46489 6236
rect 46348 6196 46354 6208
rect 46477 6205 46489 6208
rect 46523 6236 46535 6239
rect 47394 6236 47400 6248
rect 46523 6208 47400 6236
rect 46523 6205 46535 6208
rect 46477 6199 46535 6205
rect 47394 6196 47400 6208
rect 47452 6196 47458 6248
rect 47780 6245 47808 6276
rect 48317 6273 48329 6276
rect 48363 6273 48375 6307
rect 48317 6267 48375 6273
rect 48498 6264 48504 6316
rect 48556 6304 48562 6316
rect 49881 6307 49939 6313
rect 49881 6304 49893 6307
rect 48556 6276 49893 6304
rect 48556 6264 48562 6276
rect 49881 6273 49893 6276
rect 49927 6273 49939 6307
rect 49881 6267 49939 6273
rect 50985 6307 51043 6313
rect 50985 6273 50997 6307
rect 51031 6304 51043 6307
rect 53282 6304 53288 6316
rect 51031 6276 53144 6304
rect 53243 6276 53288 6304
rect 51031 6273 51043 6276
rect 50985 6267 51043 6273
rect 47489 6239 47547 6245
rect 47489 6205 47501 6239
rect 47535 6236 47547 6239
rect 47765 6239 47823 6245
rect 47765 6236 47777 6239
rect 47535 6208 47777 6236
rect 47535 6205 47547 6208
rect 47489 6199 47547 6205
rect 47765 6205 47777 6208
rect 47811 6205 47823 6239
rect 47765 6199 47823 6205
rect 47946 6196 47952 6248
rect 48004 6236 48010 6248
rect 49053 6239 49111 6245
rect 49053 6236 49065 6239
rect 48004 6208 49065 6236
rect 48004 6196 48010 6208
rect 49053 6205 49065 6208
rect 49099 6205 49111 6239
rect 49053 6199 49111 6205
rect 49789 6239 49847 6245
rect 49789 6205 49801 6239
rect 49835 6236 49847 6239
rect 49970 6236 49976 6248
rect 49835 6208 49976 6236
rect 49835 6205 49847 6208
rect 49789 6199 49847 6205
rect 49970 6196 49976 6208
rect 50028 6236 50034 6248
rect 50430 6236 50436 6248
rect 50028 6208 50436 6236
rect 50028 6196 50034 6208
rect 50430 6196 50436 6208
rect 50488 6196 50494 6248
rect 51902 6236 51908 6248
rect 51863 6208 51908 6236
rect 51902 6196 51908 6208
rect 51960 6196 51966 6248
rect 53006 6236 53012 6248
rect 52967 6208 53012 6236
rect 53006 6196 53012 6208
rect 53064 6196 53070 6248
rect 53116 6236 53144 6276
rect 53282 6264 53288 6276
rect 53340 6264 53346 6316
rect 53374 6264 53380 6316
rect 53432 6304 53438 6316
rect 55858 6304 55864 6316
rect 53432 6276 55864 6304
rect 53432 6264 53438 6276
rect 55858 6264 55864 6276
rect 55916 6264 55922 6316
rect 56413 6307 56471 6313
rect 56413 6273 56425 6307
rect 56459 6304 56471 6307
rect 57514 6304 57520 6316
rect 56459 6276 57520 6304
rect 56459 6273 56471 6276
rect 56413 6267 56471 6273
rect 57514 6264 57520 6276
rect 57572 6264 57578 6316
rect 58250 6304 58256 6316
rect 57992 6276 58256 6304
rect 56045 6239 56103 6245
rect 56045 6236 56057 6239
rect 53116 6208 56057 6236
rect 56045 6205 56057 6208
rect 56091 6236 56103 6239
rect 56689 6239 56747 6245
rect 56689 6236 56701 6239
rect 56091 6208 56701 6236
rect 56091 6205 56103 6208
rect 56045 6199 56103 6205
rect 56689 6205 56701 6208
rect 56735 6205 56747 6239
rect 57992 6236 58020 6276
rect 58250 6264 58256 6276
rect 58308 6264 58314 6316
rect 60553 6307 60611 6313
rect 60553 6304 60565 6307
rect 60384 6276 60565 6304
rect 56689 6199 56747 6205
rect 57532 6208 58020 6236
rect 58069 6239 58127 6245
rect 43772 6140 44496 6168
rect 43772 6128 43778 6140
rect 44910 6128 44916 6180
rect 44968 6128 44974 6180
rect 46385 6171 46443 6177
rect 46385 6137 46397 6171
rect 46431 6168 46443 6171
rect 46750 6168 46756 6180
rect 46431 6140 46756 6168
rect 46431 6137 46443 6140
rect 46385 6131 46443 6137
rect 46750 6128 46756 6140
rect 46808 6128 46814 6180
rect 46842 6128 46848 6180
rect 46900 6168 46906 6180
rect 46937 6171 46995 6177
rect 46937 6168 46949 6171
rect 46900 6140 46949 6168
rect 46900 6128 46906 6140
rect 46937 6137 46949 6140
rect 46983 6137 46995 6171
rect 46937 6131 46995 6137
rect 47029 6171 47087 6177
rect 47029 6137 47041 6171
rect 47075 6168 47087 6171
rect 51920 6168 51948 6196
rect 52457 6171 52515 6177
rect 52457 6168 52469 6171
rect 47075 6140 49188 6168
rect 51920 6140 52469 6168
rect 47075 6137 47087 6140
rect 47029 6131 47087 6137
rect 40221 6103 40279 6109
rect 40221 6100 40233 6103
rect 39540 6072 40233 6100
rect 39540 6060 39546 6072
rect 40221 6069 40233 6072
rect 40267 6069 40279 6103
rect 40221 6063 40279 6069
rect 46658 6060 46664 6112
rect 46716 6100 46722 6112
rect 47213 6103 47271 6109
rect 47213 6100 47225 6103
rect 46716 6072 47225 6100
rect 46716 6060 46722 6072
rect 47213 6069 47225 6072
rect 47259 6100 47271 6103
rect 49050 6100 49056 6112
rect 47259 6072 49056 6100
rect 47259 6069 47271 6072
rect 47213 6063 47271 6069
rect 49050 6060 49056 6072
rect 49108 6060 49114 6112
rect 49160 6109 49188 6140
rect 52457 6137 52469 6140
rect 52503 6137 52515 6171
rect 52457 6131 52515 6137
rect 55582 6128 55588 6180
rect 55640 6168 55646 6180
rect 55861 6171 55919 6177
rect 55861 6168 55873 6171
rect 55640 6140 55873 6168
rect 55640 6128 55646 6140
rect 55861 6137 55873 6140
rect 55907 6137 55919 6171
rect 55861 6131 55919 6137
rect 49145 6103 49203 6109
rect 49145 6069 49157 6103
rect 49191 6069 49203 6103
rect 49145 6063 49203 6069
rect 49694 6060 49700 6112
rect 49752 6100 49758 6112
rect 50062 6100 50068 6112
rect 49752 6072 50068 6100
rect 49752 6060 49758 6072
rect 50062 6060 50068 6072
rect 50120 6060 50126 6112
rect 50798 6100 50804 6112
rect 50759 6072 50804 6100
rect 50798 6060 50804 6072
rect 50856 6060 50862 6112
rect 50890 6060 50896 6112
rect 50948 6100 50954 6112
rect 52089 6103 52147 6109
rect 52089 6100 52101 6103
rect 50948 6072 52101 6100
rect 50948 6060 50954 6072
rect 52089 6069 52101 6072
rect 52135 6100 52147 6103
rect 52362 6100 52368 6112
rect 52135 6072 52368 6100
rect 52135 6069 52147 6072
rect 52089 6063 52147 6069
rect 52362 6060 52368 6072
rect 52420 6060 52426 6112
rect 52546 6060 52552 6112
rect 52604 6100 52610 6112
rect 57532 6109 57560 6208
rect 58069 6205 58081 6239
rect 58115 6205 58127 6239
rect 58342 6236 58348 6248
rect 58303 6208 58348 6236
rect 58069 6199 58127 6205
rect 52825 6103 52883 6109
rect 52825 6100 52837 6103
rect 52604 6072 52837 6100
rect 52604 6060 52610 6072
rect 52825 6069 52837 6072
rect 52871 6069 52883 6103
rect 52825 6063 52883 6069
rect 55217 6103 55275 6109
rect 55217 6069 55229 6103
rect 55263 6100 55275 6103
rect 57517 6103 57575 6109
rect 57517 6100 57529 6103
rect 55263 6072 57529 6100
rect 55263 6069 55275 6072
rect 55217 6063 55275 6069
rect 57517 6069 57529 6072
rect 57563 6069 57575 6103
rect 57974 6100 57980 6112
rect 57935 6072 57980 6100
rect 57517 6063 57575 6069
rect 57974 6060 57980 6072
rect 58032 6060 58038 6112
rect 58084 6100 58112 6199
rect 58342 6196 58348 6208
rect 58400 6196 58406 6248
rect 58434 6100 58440 6112
rect 58084 6072 58440 6100
rect 58434 6060 58440 6072
rect 58492 6060 58498 6112
rect 59998 6100 60004 6112
rect 59959 6072 60004 6100
rect 59998 6060 60004 6072
rect 60056 6060 60062 6112
rect 60274 6060 60280 6112
rect 60332 6100 60338 6112
rect 60384 6109 60412 6276
rect 60553 6273 60565 6276
rect 60599 6273 60611 6307
rect 60553 6267 60611 6273
rect 61105 6307 61163 6313
rect 61105 6273 61117 6307
rect 61151 6304 61163 6307
rect 61378 6304 61384 6316
rect 61151 6276 61384 6304
rect 61151 6273 61163 6276
rect 61105 6267 61163 6273
rect 61378 6264 61384 6276
rect 61436 6264 61442 6316
rect 60642 6236 60648 6248
rect 60603 6208 60648 6236
rect 60642 6196 60648 6208
rect 60700 6236 60706 6248
rect 61933 6239 61991 6245
rect 61933 6236 61945 6239
rect 60700 6208 61945 6236
rect 60700 6196 60706 6208
rect 61933 6205 61945 6208
rect 61979 6205 61991 6239
rect 61933 6199 61991 6205
rect 60369 6103 60427 6109
rect 60369 6100 60381 6103
rect 60332 6072 60381 6100
rect 60332 6060 60338 6072
rect 60369 6069 60381 6072
rect 60415 6069 60427 6103
rect 61562 6100 61568 6112
rect 61523 6072 61568 6100
rect 60369 6063 60427 6069
rect 61562 6060 61568 6072
rect 61620 6060 61626 6112
rect 1104 6010 63480 6032
rect 1104 5958 21774 6010
rect 21826 5958 21838 6010
rect 21890 5958 21902 6010
rect 21954 5958 21966 6010
rect 22018 5958 42566 6010
rect 42618 5958 42630 6010
rect 42682 5958 42694 6010
rect 42746 5958 42758 6010
rect 42810 5958 63480 6010
rect 1104 5936 63480 5958
rect 5629 5899 5687 5905
rect 5629 5865 5641 5899
rect 5675 5896 5687 5899
rect 6914 5896 6920 5908
rect 5675 5868 6920 5896
rect 5675 5865 5687 5868
rect 5629 5859 5687 5865
rect 3510 5788 3516 5840
rect 3568 5828 3574 5840
rect 4249 5831 4307 5837
rect 4249 5828 4261 5831
rect 3568 5800 4261 5828
rect 3568 5788 3574 5800
rect 4249 5797 4261 5800
rect 4295 5797 4307 5831
rect 4249 5791 4307 5797
rect 2682 5760 2688 5772
rect 2643 5732 2688 5760
rect 2682 5720 2688 5732
rect 2740 5720 2746 5772
rect 3145 5763 3203 5769
rect 3145 5729 3157 5763
rect 3191 5760 3203 5763
rect 4614 5760 4620 5772
rect 3191 5732 4620 5760
rect 3191 5729 3203 5732
rect 3145 5723 3203 5729
rect 4614 5720 4620 5732
rect 4672 5720 4678 5772
rect 5077 5763 5135 5769
rect 5077 5760 5089 5763
rect 4724 5732 5089 5760
rect 2590 5692 2596 5704
rect 2551 5664 2596 5692
rect 2590 5652 2596 5664
rect 2648 5652 2654 5704
rect 2700 5692 2728 5720
rect 4724 5692 4752 5732
rect 5077 5729 5089 5732
rect 5123 5760 5135 5763
rect 5166 5760 5172 5772
rect 5123 5732 5172 5760
rect 5123 5729 5135 5732
rect 5077 5723 5135 5729
rect 5166 5720 5172 5732
rect 5224 5720 5230 5772
rect 5261 5763 5319 5769
rect 5261 5729 5273 5763
rect 5307 5760 5319 5763
rect 5644 5760 5672 5859
rect 6914 5856 6920 5868
rect 6972 5856 6978 5908
rect 7190 5856 7196 5908
rect 7248 5896 7254 5908
rect 9398 5896 9404 5908
rect 7248 5868 8340 5896
rect 9311 5868 9404 5896
rect 7248 5856 7254 5868
rect 6546 5788 6552 5840
rect 6604 5828 6610 5840
rect 6641 5831 6699 5837
rect 6641 5828 6653 5831
rect 6604 5800 6653 5828
rect 6604 5788 6610 5800
rect 6641 5797 6653 5800
rect 6687 5797 6699 5831
rect 7837 5831 7895 5837
rect 7837 5828 7849 5831
rect 6641 5791 6699 5797
rect 7300 5800 7849 5828
rect 5307 5732 5672 5760
rect 6089 5763 6147 5769
rect 5307 5729 5319 5732
rect 5261 5723 5319 5729
rect 6089 5729 6101 5763
rect 6135 5760 6147 5763
rect 6178 5760 6184 5772
rect 6135 5732 6184 5760
rect 6135 5729 6147 5732
rect 6089 5723 6147 5729
rect 6178 5720 6184 5732
rect 6236 5760 6242 5772
rect 7300 5760 7328 5800
rect 7837 5797 7849 5800
rect 7883 5828 7895 5831
rect 8202 5828 8208 5840
rect 7883 5800 8208 5828
rect 7883 5797 7895 5800
rect 7837 5791 7895 5797
rect 8202 5788 8208 5800
rect 8260 5788 8266 5840
rect 8312 5828 8340 5868
rect 9398 5856 9404 5868
rect 9456 5896 9462 5908
rect 16758 5896 16764 5908
rect 9456 5868 16764 5896
rect 9456 5856 9462 5868
rect 16758 5856 16764 5868
rect 16816 5896 16822 5908
rect 16945 5899 17003 5905
rect 16945 5896 16957 5899
rect 16816 5868 16957 5896
rect 16816 5856 16822 5868
rect 16945 5865 16957 5868
rect 16991 5865 17003 5899
rect 16945 5859 17003 5865
rect 17034 5856 17040 5908
rect 17092 5896 17098 5908
rect 20714 5896 20720 5908
rect 17092 5868 20024 5896
rect 20675 5868 20720 5896
rect 17092 5856 17098 5868
rect 8386 5828 8392 5840
rect 8299 5800 8392 5828
rect 8386 5788 8392 5800
rect 8444 5828 8450 5840
rect 11698 5828 11704 5840
rect 8444 5800 11704 5828
rect 8444 5788 8450 5800
rect 11698 5788 11704 5800
rect 11756 5788 11762 5840
rect 12069 5831 12127 5837
rect 12069 5797 12081 5831
rect 12115 5828 12127 5831
rect 12894 5828 12900 5840
rect 12115 5800 12900 5828
rect 12115 5797 12127 5800
rect 12069 5791 12127 5797
rect 12894 5788 12900 5800
rect 12952 5788 12958 5840
rect 17497 5831 17555 5837
rect 17497 5797 17509 5831
rect 17543 5828 17555 5831
rect 18782 5828 18788 5840
rect 17543 5800 18788 5828
rect 17543 5797 17555 5800
rect 17497 5791 17555 5797
rect 18782 5788 18788 5800
rect 18840 5828 18846 5840
rect 18969 5831 19027 5837
rect 18840 5800 18920 5828
rect 18840 5788 18846 5800
rect 6236 5732 7328 5760
rect 7377 5763 7435 5769
rect 6236 5720 6242 5732
rect 7377 5729 7389 5763
rect 7423 5760 7435 5763
rect 8294 5760 8300 5772
rect 7423 5732 8300 5760
rect 7423 5729 7435 5732
rect 7377 5723 7435 5729
rect 8294 5720 8300 5732
rect 8352 5720 8358 5772
rect 9766 5760 9772 5772
rect 9727 5732 9772 5760
rect 9766 5720 9772 5732
rect 9824 5760 9830 5772
rect 10505 5763 10563 5769
rect 10505 5760 10517 5763
rect 9824 5732 10517 5760
rect 9824 5720 9830 5732
rect 10505 5729 10517 5732
rect 10551 5729 10563 5763
rect 10505 5723 10563 5729
rect 11054 5720 11060 5772
rect 11112 5760 11118 5772
rect 11609 5763 11667 5769
rect 11609 5760 11621 5763
rect 11112 5732 11621 5760
rect 11112 5720 11118 5732
rect 11609 5729 11621 5732
rect 11655 5760 11667 5763
rect 11882 5760 11888 5772
rect 11655 5732 11888 5760
rect 11655 5729 11667 5732
rect 11609 5723 11667 5729
rect 11882 5720 11888 5732
rect 11940 5720 11946 5772
rect 13541 5763 13599 5769
rect 13541 5729 13553 5763
rect 13587 5760 13599 5763
rect 13630 5760 13636 5772
rect 13587 5732 13636 5760
rect 13587 5729 13599 5732
rect 13541 5723 13599 5729
rect 13630 5720 13636 5732
rect 13688 5720 13694 5772
rect 14093 5763 14151 5769
rect 14093 5729 14105 5763
rect 14139 5760 14151 5763
rect 15010 5760 15016 5772
rect 14139 5732 15016 5760
rect 14139 5729 14151 5732
rect 14093 5723 14151 5729
rect 15010 5720 15016 5732
rect 15068 5720 15074 5772
rect 15933 5763 15991 5769
rect 15933 5729 15945 5763
rect 15979 5760 15991 5763
rect 16114 5760 16120 5772
rect 15979 5732 16120 5760
rect 15979 5729 15991 5732
rect 15933 5723 15991 5729
rect 16114 5720 16120 5732
rect 16172 5720 16178 5772
rect 16298 5760 16304 5772
rect 16259 5732 16304 5760
rect 16298 5720 16304 5732
rect 16356 5720 16362 5772
rect 16485 5763 16543 5769
rect 16485 5729 16497 5763
rect 16531 5760 16543 5763
rect 17770 5760 17776 5772
rect 16531 5732 17776 5760
rect 16531 5729 16543 5732
rect 16485 5723 16543 5729
rect 17770 5720 17776 5732
rect 17828 5720 17834 5772
rect 18138 5720 18144 5772
rect 18196 5760 18202 5772
rect 18233 5763 18291 5769
rect 18233 5760 18245 5763
rect 18196 5732 18245 5760
rect 18196 5720 18202 5732
rect 18233 5729 18245 5732
rect 18279 5729 18291 5763
rect 18233 5723 18291 5729
rect 18325 5763 18383 5769
rect 18325 5729 18337 5763
rect 18371 5760 18383 5763
rect 18690 5760 18696 5772
rect 18371 5732 18696 5760
rect 18371 5729 18383 5732
rect 18325 5723 18383 5729
rect 18690 5720 18696 5732
rect 18748 5720 18754 5772
rect 18892 5760 18920 5800
rect 18969 5797 18981 5831
rect 19015 5828 19027 5831
rect 19153 5831 19211 5837
rect 19153 5828 19165 5831
rect 19015 5800 19165 5828
rect 19015 5797 19027 5800
rect 18969 5791 19027 5797
rect 19153 5797 19165 5800
rect 19199 5828 19211 5831
rect 19334 5828 19340 5840
rect 19199 5800 19340 5828
rect 19199 5797 19211 5800
rect 19153 5791 19211 5797
rect 19334 5788 19340 5800
rect 19392 5788 19398 5840
rect 19429 5831 19487 5837
rect 19429 5797 19441 5831
rect 19475 5828 19487 5831
rect 19794 5828 19800 5840
rect 19475 5800 19800 5828
rect 19475 5797 19487 5800
rect 19429 5791 19487 5797
rect 19794 5788 19800 5800
rect 19852 5788 19858 5840
rect 19996 5837 20024 5868
rect 20714 5856 20720 5868
rect 20772 5856 20778 5908
rect 22094 5856 22100 5908
rect 22152 5896 22158 5908
rect 22465 5899 22523 5905
rect 22465 5896 22477 5899
rect 22152 5868 22477 5896
rect 22152 5856 22158 5868
rect 22465 5865 22477 5868
rect 22511 5896 22523 5899
rect 22830 5896 22836 5908
rect 22511 5868 22836 5896
rect 22511 5865 22523 5868
rect 22465 5859 22523 5865
rect 22830 5856 22836 5868
rect 22888 5856 22894 5908
rect 23106 5896 23112 5908
rect 23067 5868 23112 5896
rect 23106 5856 23112 5868
rect 23164 5856 23170 5908
rect 23658 5896 23664 5908
rect 23619 5868 23664 5896
rect 23658 5856 23664 5868
rect 23716 5856 23722 5908
rect 24026 5856 24032 5908
rect 24084 5896 24090 5908
rect 27249 5899 27307 5905
rect 27249 5896 27261 5899
rect 24084 5868 27261 5896
rect 24084 5856 24090 5868
rect 27249 5865 27261 5868
rect 27295 5865 27307 5899
rect 27249 5859 27307 5865
rect 28258 5856 28264 5908
rect 28316 5896 28322 5908
rect 31297 5899 31355 5905
rect 31297 5896 31309 5899
rect 28316 5868 31309 5896
rect 28316 5856 28322 5868
rect 31297 5865 31309 5868
rect 31343 5865 31355 5899
rect 31297 5859 31355 5865
rect 31386 5856 31392 5908
rect 31444 5896 31450 5908
rect 31444 5868 33272 5896
rect 31444 5856 31450 5868
rect 19981 5831 20039 5837
rect 19981 5797 19993 5831
rect 20027 5797 20039 5831
rect 19981 5791 20039 5797
rect 20898 5788 20904 5840
rect 20956 5828 20962 5840
rect 21177 5831 21235 5837
rect 21177 5828 21189 5831
rect 20956 5800 21189 5828
rect 20956 5788 20962 5800
rect 21177 5797 21189 5800
rect 21223 5828 21235 5831
rect 21266 5828 21272 5840
rect 21223 5800 21272 5828
rect 21223 5797 21235 5800
rect 21177 5791 21235 5797
rect 21266 5788 21272 5800
rect 21324 5788 21330 5840
rect 22741 5831 22799 5837
rect 22741 5828 22753 5831
rect 21560 5800 22753 5828
rect 21560 5772 21588 5800
rect 22741 5797 22753 5800
rect 22787 5797 22799 5831
rect 24854 5828 24860 5840
rect 22741 5791 22799 5797
rect 24136 5800 24860 5828
rect 19521 5763 19579 5769
rect 19521 5760 19533 5763
rect 18892 5732 19533 5760
rect 19521 5729 19533 5732
rect 19567 5729 19579 5763
rect 19521 5723 19579 5729
rect 19610 5720 19616 5772
rect 19668 5760 19674 5772
rect 20257 5763 20315 5769
rect 20257 5760 20269 5763
rect 19668 5732 20269 5760
rect 19668 5720 19674 5732
rect 20257 5729 20269 5732
rect 20303 5729 20315 5763
rect 21542 5760 21548 5772
rect 21503 5732 21548 5760
rect 20257 5723 20315 5729
rect 21542 5720 21548 5732
rect 21600 5720 21606 5772
rect 21637 5763 21695 5769
rect 21637 5729 21649 5763
rect 21683 5760 21695 5763
rect 22646 5760 22652 5772
rect 21683 5732 22652 5760
rect 21683 5729 21695 5732
rect 21637 5723 21695 5729
rect 22646 5720 22652 5732
rect 22704 5720 22710 5772
rect 22922 5760 22928 5772
rect 22883 5732 22928 5760
rect 22922 5720 22928 5732
rect 22980 5720 22986 5772
rect 24026 5760 24032 5772
rect 23032 5732 24032 5760
rect 2700 5664 4752 5692
rect 4801 5695 4859 5701
rect 4801 5661 4813 5695
rect 4847 5692 4859 5695
rect 4982 5692 4988 5704
rect 4847 5664 4988 5692
rect 4847 5661 4859 5664
rect 4801 5655 4859 5661
rect 4982 5652 4988 5664
rect 5040 5692 5046 5704
rect 5442 5692 5448 5704
rect 5040 5664 5448 5692
rect 5040 5652 5046 5664
rect 5442 5652 5448 5664
rect 5500 5652 5506 5704
rect 7285 5695 7343 5701
rect 7285 5661 7297 5695
rect 7331 5692 7343 5695
rect 7742 5692 7748 5704
rect 7331 5664 7748 5692
rect 7331 5661 7343 5664
rect 7285 5655 7343 5661
rect 7742 5652 7748 5664
rect 7800 5652 7806 5704
rect 9674 5692 9680 5704
rect 9587 5664 9680 5692
rect 9674 5652 9680 5664
rect 9732 5692 9738 5704
rect 10226 5692 10232 5704
rect 9732 5664 10232 5692
rect 9732 5652 9738 5664
rect 10226 5652 10232 5664
rect 10284 5652 10290 5704
rect 11517 5695 11575 5701
rect 11517 5661 11529 5695
rect 11563 5692 11575 5695
rect 11698 5692 11704 5704
rect 11563 5664 11704 5692
rect 11563 5661 11575 5664
rect 11517 5655 11575 5661
rect 11698 5652 11704 5664
rect 11756 5652 11762 5704
rect 14185 5695 14243 5701
rect 14185 5661 14197 5695
rect 14231 5692 14243 5695
rect 15565 5695 15623 5701
rect 14231 5664 14780 5692
rect 14231 5661 14243 5664
rect 14185 5655 14243 5661
rect 5166 5584 5172 5636
rect 5224 5624 5230 5636
rect 6273 5627 6331 5633
rect 6273 5624 6285 5627
rect 5224 5596 6285 5624
rect 5224 5584 5230 5596
rect 6273 5593 6285 5596
rect 6319 5624 6331 5627
rect 8110 5624 8116 5636
rect 6319 5596 8116 5624
rect 6319 5593 6331 5596
rect 6273 5587 6331 5593
rect 8110 5584 8116 5596
rect 8168 5624 8174 5636
rect 8297 5627 8355 5633
rect 8297 5624 8309 5627
rect 8168 5596 8309 5624
rect 8168 5584 8174 5596
rect 8297 5593 8309 5596
rect 8343 5624 8355 5627
rect 11054 5624 11060 5636
rect 8343 5596 11060 5624
rect 8343 5593 8355 5596
rect 8297 5587 8355 5593
rect 11054 5584 11060 5596
rect 11112 5584 11118 5636
rect 12526 5584 12532 5636
rect 12584 5624 12590 5636
rect 13081 5627 13139 5633
rect 13081 5624 13093 5627
rect 12584 5596 13093 5624
rect 12584 5584 12590 5596
rect 13081 5593 13093 5596
rect 13127 5593 13139 5627
rect 14090 5624 14096 5636
rect 14051 5596 14096 5624
rect 13081 5587 13139 5593
rect 14090 5584 14096 5596
rect 14148 5584 14154 5636
rect 14752 5633 14780 5664
rect 15565 5661 15577 5695
rect 15611 5661 15623 5695
rect 15565 5655 15623 5661
rect 14737 5627 14795 5633
rect 14737 5593 14749 5627
rect 14783 5624 14795 5627
rect 14918 5624 14924 5636
rect 14783 5596 14924 5624
rect 14783 5593 14795 5596
rect 14737 5587 14795 5593
rect 14918 5584 14924 5596
rect 14976 5624 14982 5636
rect 15580 5624 15608 5655
rect 16574 5652 16580 5704
rect 16632 5692 16638 5704
rect 17405 5695 17463 5701
rect 17405 5692 17417 5695
rect 16632 5664 17417 5692
rect 16632 5652 16638 5664
rect 17405 5661 17417 5664
rect 17451 5692 17463 5695
rect 18046 5692 18052 5704
rect 17451 5664 18052 5692
rect 17451 5661 17463 5664
rect 17405 5655 17463 5661
rect 18046 5652 18052 5664
rect 18104 5652 18110 5704
rect 18509 5695 18567 5701
rect 18509 5661 18521 5695
rect 18555 5692 18567 5695
rect 18555 5664 22508 5692
rect 18555 5661 18567 5664
rect 18509 5655 18567 5661
rect 15930 5624 15936 5636
rect 14976 5596 15516 5624
rect 15580 5596 15936 5624
rect 14976 5584 14982 5596
rect 2314 5516 2320 5568
rect 2372 5556 2378 5568
rect 2409 5559 2467 5565
rect 2409 5556 2421 5559
rect 2372 5528 2421 5556
rect 2372 5516 2378 5528
rect 2409 5525 2421 5528
rect 2455 5525 2467 5559
rect 3510 5556 3516 5568
rect 3471 5528 3516 5556
rect 2409 5519 2467 5525
rect 3510 5516 3516 5528
rect 3568 5516 3574 5568
rect 3786 5556 3792 5568
rect 3747 5528 3792 5556
rect 3786 5516 3792 5528
rect 3844 5556 3850 5568
rect 5626 5556 5632 5568
rect 3844 5528 5632 5556
rect 3844 5516 3850 5528
rect 5626 5516 5632 5528
rect 5684 5516 5690 5568
rect 5718 5516 5724 5568
rect 5776 5556 5782 5568
rect 5905 5559 5963 5565
rect 5905 5556 5917 5559
rect 5776 5528 5917 5556
rect 5776 5516 5782 5528
rect 5905 5525 5917 5528
rect 5951 5525 5963 5559
rect 7006 5556 7012 5568
rect 6967 5528 7012 5556
rect 5905 5519 5963 5525
rect 7006 5516 7012 5528
rect 7064 5516 7070 5568
rect 8757 5559 8815 5565
rect 8757 5525 8769 5559
rect 8803 5556 8815 5559
rect 8846 5556 8852 5568
rect 8803 5528 8852 5556
rect 8803 5525 8815 5528
rect 8757 5519 8815 5525
rect 8846 5516 8852 5528
rect 8904 5516 8910 5568
rect 8938 5516 8944 5568
rect 8996 5556 9002 5568
rect 9953 5559 10011 5565
rect 9953 5556 9965 5559
rect 8996 5528 9965 5556
rect 8996 5516 9002 5528
rect 9953 5525 9965 5528
rect 9999 5525 10011 5559
rect 9953 5519 10011 5525
rect 10410 5516 10416 5568
rect 10468 5556 10474 5568
rect 12345 5559 12403 5565
rect 12345 5556 12357 5559
rect 10468 5528 12357 5556
rect 10468 5516 10474 5528
rect 12345 5525 12357 5528
rect 12391 5525 12403 5559
rect 12802 5556 12808 5568
rect 12763 5528 12808 5556
rect 12345 5519 12403 5525
rect 12802 5516 12808 5528
rect 12860 5516 12866 5568
rect 15102 5556 15108 5568
rect 15063 5528 15108 5556
rect 15102 5516 15108 5528
rect 15160 5516 15166 5568
rect 15488 5556 15516 5596
rect 15930 5584 15936 5596
rect 15988 5624 15994 5636
rect 22370 5624 22376 5636
rect 15988 5596 22376 5624
rect 15988 5584 15994 5596
rect 22370 5584 22376 5596
rect 22428 5584 22434 5636
rect 22480 5624 22508 5664
rect 23032 5624 23060 5732
rect 24026 5720 24032 5732
rect 24084 5720 24090 5772
rect 24136 5769 24164 5800
rect 24854 5788 24860 5800
rect 24912 5788 24918 5840
rect 25314 5788 25320 5840
rect 25372 5828 25378 5840
rect 25501 5831 25559 5837
rect 25501 5828 25513 5831
rect 25372 5800 25513 5828
rect 25372 5788 25378 5800
rect 25501 5797 25513 5800
rect 25547 5797 25559 5831
rect 25501 5791 25559 5797
rect 25590 5788 25596 5840
rect 25648 5828 25654 5840
rect 25869 5831 25927 5837
rect 25869 5828 25881 5831
rect 25648 5800 25881 5828
rect 25648 5788 25654 5800
rect 25869 5797 25881 5800
rect 25915 5797 25927 5831
rect 25869 5791 25927 5797
rect 26329 5831 26387 5837
rect 26329 5797 26341 5831
rect 26375 5828 26387 5831
rect 26418 5828 26424 5840
rect 26375 5800 26424 5828
rect 26375 5797 26387 5800
rect 26329 5791 26387 5797
rect 26418 5788 26424 5800
rect 26476 5828 26482 5840
rect 26605 5831 26663 5837
rect 26605 5828 26617 5831
rect 26476 5800 26617 5828
rect 26476 5788 26482 5800
rect 26605 5797 26617 5800
rect 26651 5797 26663 5831
rect 26605 5791 26663 5797
rect 28629 5831 28687 5837
rect 28629 5797 28641 5831
rect 28675 5828 28687 5831
rect 28675 5800 32168 5828
rect 28675 5797 28687 5800
rect 28629 5791 28687 5797
rect 24121 5763 24179 5769
rect 24121 5729 24133 5763
rect 24167 5729 24179 5763
rect 24394 5760 24400 5772
rect 24355 5732 24400 5760
rect 24121 5723 24179 5729
rect 24394 5720 24400 5732
rect 24452 5760 24458 5772
rect 24670 5760 24676 5772
rect 24452 5732 24676 5760
rect 24452 5720 24458 5732
rect 24670 5720 24676 5732
rect 24728 5720 24734 5772
rect 28537 5763 28595 5769
rect 28537 5729 28549 5763
rect 28583 5729 28595 5763
rect 28537 5723 28595 5729
rect 28905 5763 28963 5769
rect 28905 5729 28917 5763
rect 28951 5760 28963 5763
rect 29086 5760 29092 5772
rect 28951 5732 29092 5760
rect 28951 5729 28963 5732
rect 28905 5723 28963 5729
rect 23198 5652 23204 5704
rect 23256 5692 23262 5704
rect 24857 5695 24915 5701
rect 23256 5664 24532 5692
rect 23256 5652 23262 5664
rect 24213 5627 24271 5633
rect 24213 5624 24225 5627
rect 22480 5596 23060 5624
rect 23124 5596 24225 5624
rect 18509 5559 18567 5565
rect 18509 5556 18521 5559
rect 15488 5528 18521 5556
rect 18509 5525 18521 5528
rect 18555 5525 18567 5559
rect 18509 5519 18567 5525
rect 18690 5516 18696 5568
rect 18748 5556 18754 5568
rect 18785 5559 18843 5565
rect 18785 5556 18797 5559
rect 18748 5528 18797 5556
rect 18748 5516 18754 5528
rect 18785 5525 18797 5528
rect 18831 5556 18843 5559
rect 18969 5559 19027 5565
rect 18969 5556 18981 5559
rect 18831 5528 18981 5556
rect 18831 5525 18843 5528
rect 18785 5519 18843 5525
rect 18969 5525 18981 5528
rect 19015 5525 19027 5559
rect 18969 5519 19027 5525
rect 19245 5559 19303 5565
rect 19245 5525 19257 5559
rect 19291 5556 19303 5559
rect 19334 5556 19340 5568
rect 19291 5528 19340 5556
rect 19291 5525 19303 5528
rect 19245 5519 19303 5525
rect 19334 5516 19340 5528
rect 19392 5556 19398 5568
rect 21361 5559 21419 5565
rect 21361 5556 21373 5559
rect 19392 5528 21373 5556
rect 19392 5516 19398 5528
rect 21361 5525 21373 5528
rect 21407 5556 21419 5559
rect 21726 5556 21732 5568
rect 21407 5528 21732 5556
rect 21407 5525 21419 5528
rect 21361 5519 21419 5525
rect 21726 5516 21732 5528
rect 21784 5516 21790 5568
rect 21821 5559 21879 5565
rect 21821 5525 21833 5559
rect 21867 5556 21879 5559
rect 23124 5556 23152 5596
rect 24213 5593 24225 5596
rect 24259 5624 24271 5627
rect 24394 5624 24400 5636
rect 24259 5596 24400 5624
rect 24259 5593 24271 5596
rect 24213 5587 24271 5593
rect 24394 5584 24400 5596
rect 24452 5584 24458 5636
rect 24504 5624 24532 5664
rect 24857 5661 24869 5695
rect 24903 5692 24915 5695
rect 25038 5692 25044 5704
rect 24903 5664 25044 5692
rect 24903 5661 24915 5664
rect 24857 5655 24915 5661
rect 25038 5652 25044 5664
rect 25096 5692 25102 5704
rect 25133 5695 25191 5701
rect 25133 5692 25145 5695
rect 25096 5664 25145 5692
rect 25096 5652 25102 5664
rect 25133 5661 25145 5664
rect 25179 5661 25191 5695
rect 25133 5655 25191 5661
rect 26694 5652 26700 5704
rect 26752 5701 26758 5704
rect 26752 5695 26810 5701
rect 26752 5661 26764 5695
rect 26798 5661 26810 5695
rect 26752 5655 26810 5661
rect 26752 5652 26758 5655
rect 26970 5652 26976 5704
rect 27028 5692 27034 5704
rect 28552 5692 28580 5723
rect 29086 5720 29092 5732
rect 29144 5720 29150 5772
rect 29454 5760 29460 5772
rect 29415 5732 29460 5760
rect 29454 5720 29460 5732
rect 29512 5720 29518 5772
rect 29546 5720 29552 5772
rect 29604 5760 29610 5772
rect 30006 5760 30012 5772
rect 29604 5732 29649 5760
rect 29967 5732 30012 5760
rect 29604 5720 29610 5732
rect 30006 5720 30012 5732
rect 30064 5720 30070 5772
rect 31018 5760 31024 5772
rect 30979 5732 31024 5760
rect 31018 5720 31024 5732
rect 31076 5720 31082 5772
rect 31294 5720 31300 5772
rect 31352 5760 31358 5772
rect 32140 5769 32168 5800
rect 32950 5788 32956 5840
rect 33008 5828 33014 5840
rect 33045 5831 33103 5837
rect 33045 5828 33057 5831
rect 33008 5800 33057 5828
rect 33008 5788 33014 5800
rect 33045 5797 33057 5800
rect 33091 5797 33103 5831
rect 33045 5791 33103 5797
rect 32125 5763 32183 5769
rect 31352 5732 31616 5760
rect 31352 5720 31358 5732
rect 28626 5692 28632 5704
rect 27028 5664 27073 5692
rect 28539 5664 28632 5692
rect 27028 5652 27034 5664
rect 28626 5652 28632 5664
rect 28684 5692 28690 5704
rect 29822 5692 29828 5704
rect 28684 5664 29828 5692
rect 28684 5652 28690 5664
rect 29822 5652 29828 5664
rect 29880 5652 29886 5704
rect 30024 5692 30052 5720
rect 31478 5692 31484 5704
rect 30024 5664 31484 5692
rect 31478 5652 31484 5664
rect 31536 5652 31542 5704
rect 31588 5692 31616 5732
rect 32125 5729 32137 5763
rect 32171 5760 32183 5763
rect 32490 5760 32496 5772
rect 32171 5732 32496 5760
rect 32171 5729 32183 5732
rect 32125 5723 32183 5729
rect 32490 5720 32496 5732
rect 32548 5720 32554 5772
rect 33244 5769 33272 5868
rect 35250 5856 35256 5908
rect 35308 5896 35314 5908
rect 41322 5896 41328 5908
rect 35308 5868 41328 5896
rect 35308 5856 35314 5868
rect 41322 5856 41328 5868
rect 41380 5856 41386 5908
rect 41598 5896 41604 5908
rect 41559 5868 41604 5896
rect 41598 5856 41604 5868
rect 41656 5896 41662 5908
rect 42061 5899 42119 5905
rect 42061 5896 42073 5899
rect 41656 5868 42073 5896
rect 41656 5856 41662 5868
rect 42061 5865 42073 5868
rect 42107 5865 42119 5899
rect 42061 5859 42119 5865
rect 42242 5856 42248 5908
rect 42300 5896 42306 5908
rect 42613 5899 42671 5905
rect 42613 5896 42625 5899
rect 42300 5868 42625 5896
rect 42300 5856 42306 5868
rect 42613 5865 42625 5868
rect 42659 5865 42671 5899
rect 42978 5896 42984 5908
rect 42939 5868 42984 5896
rect 42613 5859 42671 5865
rect 42978 5856 42984 5868
rect 43036 5856 43042 5908
rect 48222 5896 48228 5908
rect 43272 5868 48228 5896
rect 33873 5831 33931 5837
rect 33873 5797 33885 5831
rect 33919 5828 33931 5831
rect 34146 5828 34152 5840
rect 33919 5800 34152 5828
rect 33919 5797 33931 5800
rect 33873 5791 33931 5797
rect 34146 5788 34152 5800
rect 34204 5788 34210 5840
rect 34333 5831 34391 5837
rect 34333 5797 34345 5831
rect 34379 5828 34391 5831
rect 38378 5828 38384 5840
rect 34379 5800 37872 5828
rect 38339 5800 38384 5828
rect 34379 5797 34391 5800
rect 34333 5791 34391 5797
rect 33229 5763 33287 5769
rect 33229 5729 33241 5763
rect 33275 5760 33287 5763
rect 33594 5760 33600 5772
rect 33275 5732 33600 5760
rect 33275 5729 33287 5732
rect 33229 5723 33287 5729
rect 33594 5720 33600 5732
rect 33652 5720 33658 5772
rect 34882 5760 34888 5772
rect 34843 5732 34888 5760
rect 34882 5720 34888 5732
rect 34940 5720 34946 5772
rect 34974 5720 34980 5772
rect 35032 5760 35038 5772
rect 35158 5760 35164 5772
rect 35032 5732 35077 5760
rect 35119 5732 35164 5760
rect 35032 5720 35038 5732
rect 35158 5720 35164 5732
rect 35216 5720 35222 5772
rect 35342 5760 35348 5772
rect 35303 5732 35348 5760
rect 35342 5720 35348 5732
rect 35400 5720 35406 5772
rect 35434 5720 35440 5772
rect 35492 5760 35498 5772
rect 35621 5763 35679 5769
rect 35621 5760 35633 5763
rect 35492 5732 35633 5760
rect 35492 5720 35498 5732
rect 35621 5729 35633 5732
rect 35667 5729 35679 5763
rect 35621 5723 35679 5729
rect 36633 5763 36691 5769
rect 36633 5729 36645 5763
rect 36679 5760 36691 5763
rect 36998 5760 37004 5772
rect 36679 5732 37004 5760
rect 36679 5729 36691 5732
rect 36633 5723 36691 5729
rect 36998 5720 37004 5732
rect 37056 5720 37062 5772
rect 37274 5720 37280 5772
rect 37332 5760 37338 5772
rect 37461 5763 37519 5769
rect 37461 5760 37473 5763
rect 37332 5732 37473 5760
rect 37332 5720 37338 5732
rect 37461 5729 37473 5732
rect 37507 5729 37519 5763
rect 37734 5760 37740 5772
rect 37695 5732 37740 5760
rect 37461 5723 37519 5729
rect 37734 5720 37740 5732
rect 37792 5720 37798 5772
rect 37844 5760 37872 5800
rect 38378 5788 38384 5800
rect 38436 5788 38442 5840
rect 41874 5828 41880 5840
rect 41623 5800 41880 5828
rect 41623 5760 41651 5800
rect 41874 5788 41880 5800
rect 41932 5788 41938 5840
rect 42797 5831 42855 5837
rect 42797 5797 42809 5831
rect 42843 5828 42855 5831
rect 43272 5828 43300 5868
rect 48222 5856 48228 5868
rect 48280 5856 48286 5908
rect 49142 5896 49148 5908
rect 49103 5868 49148 5896
rect 49142 5856 49148 5868
rect 49200 5856 49206 5908
rect 49970 5896 49976 5908
rect 49931 5868 49976 5896
rect 49970 5856 49976 5868
rect 50028 5856 50034 5908
rect 52178 5896 52184 5908
rect 50080 5868 52184 5896
rect 43438 5828 43444 5840
rect 42843 5800 43300 5828
rect 43399 5800 43444 5828
rect 42843 5797 42855 5800
rect 42797 5791 42855 5797
rect 43438 5788 43444 5800
rect 43496 5788 43502 5840
rect 43993 5831 44051 5837
rect 43993 5797 44005 5831
rect 44039 5828 44051 5831
rect 46290 5828 46296 5840
rect 44039 5800 46296 5828
rect 44039 5797 44051 5800
rect 43993 5791 44051 5797
rect 46290 5788 46296 5800
rect 46348 5788 46354 5840
rect 50080 5828 50108 5868
rect 52178 5856 52184 5868
rect 52236 5856 52242 5908
rect 52270 5856 52276 5908
rect 52328 5896 52334 5908
rect 52328 5868 55628 5896
rect 52328 5856 52334 5868
rect 46584 5800 50108 5828
rect 37844 5732 41651 5760
rect 41690 5720 41696 5772
rect 41748 5760 41754 5772
rect 41785 5763 41843 5769
rect 41785 5760 41797 5763
rect 41748 5732 41797 5760
rect 41748 5720 41754 5732
rect 41785 5729 41797 5732
rect 41831 5729 41843 5763
rect 41966 5760 41972 5772
rect 41927 5732 41972 5760
rect 41785 5723 41843 5729
rect 41966 5720 41972 5732
rect 42024 5720 42030 5772
rect 43625 5763 43683 5769
rect 43625 5729 43637 5763
rect 43671 5760 43683 5763
rect 43898 5760 43904 5772
rect 43671 5732 43904 5760
rect 43671 5729 43683 5732
rect 43625 5723 43683 5729
rect 43898 5720 43904 5732
rect 43956 5720 43962 5772
rect 44082 5720 44088 5772
rect 44140 5760 44146 5772
rect 44269 5763 44327 5769
rect 44269 5760 44281 5763
rect 44140 5732 44281 5760
rect 44140 5720 44146 5732
rect 44269 5729 44281 5732
rect 44315 5729 44327 5763
rect 44269 5723 44327 5729
rect 44358 5720 44364 5772
rect 44416 5760 44422 5772
rect 45002 5760 45008 5772
rect 44416 5732 45008 5760
rect 44416 5720 44422 5732
rect 45002 5720 45008 5732
rect 45060 5720 45066 5772
rect 45094 5720 45100 5772
rect 45152 5760 45158 5772
rect 45833 5763 45891 5769
rect 45833 5760 45845 5763
rect 45152 5732 45845 5760
rect 45152 5720 45158 5732
rect 45833 5729 45845 5732
rect 45879 5729 45891 5763
rect 45833 5723 45891 5729
rect 31588 5664 37228 5692
rect 29362 5624 29368 5636
rect 24504 5596 29368 5624
rect 29362 5584 29368 5596
rect 29420 5584 29426 5636
rect 29454 5584 29460 5636
rect 29512 5624 29518 5636
rect 30098 5624 30104 5636
rect 29512 5596 30104 5624
rect 29512 5584 29518 5596
rect 30098 5584 30104 5596
rect 30156 5624 30162 5636
rect 30929 5627 30987 5633
rect 30929 5624 30941 5627
rect 30156 5596 30941 5624
rect 30156 5584 30162 5596
rect 30929 5593 30941 5596
rect 30975 5624 30987 5627
rect 31202 5624 31208 5636
rect 30975 5596 31208 5624
rect 30975 5593 30987 5596
rect 30929 5587 30987 5593
rect 31202 5584 31208 5596
rect 31260 5584 31266 5636
rect 31297 5627 31355 5633
rect 31297 5593 31309 5627
rect 31343 5624 31355 5627
rect 32309 5627 32367 5633
rect 32309 5624 32321 5627
rect 31343 5596 32321 5624
rect 31343 5593 31355 5596
rect 31297 5587 31355 5593
rect 32309 5593 32321 5596
rect 32355 5593 32367 5627
rect 35158 5624 35164 5636
rect 32309 5587 32367 5593
rect 33520 5596 35164 5624
rect 33520 5568 33548 5596
rect 35158 5584 35164 5596
rect 35216 5624 35222 5636
rect 35986 5624 35992 5636
rect 35216 5596 35992 5624
rect 35216 5584 35222 5596
rect 35986 5584 35992 5596
rect 36044 5584 36050 5636
rect 36170 5584 36176 5636
rect 36228 5624 36234 5636
rect 37093 5627 37151 5633
rect 37093 5624 37105 5627
rect 36228 5596 37105 5624
rect 36228 5584 36234 5596
rect 37093 5593 37105 5596
rect 37139 5593 37151 5627
rect 37200 5624 37228 5664
rect 39022 5652 39028 5704
rect 39080 5692 39086 5704
rect 39298 5692 39304 5704
rect 39080 5664 39304 5692
rect 39080 5652 39086 5664
rect 39298 5652 39304 5664
rect 39356 5652 39362 5704
rect 39574 5692 39580 5704
rect 39535 5664 39580 5692
rect 39574 5652 39580 5664
rect 39632 5652 39638 5704
rect 40218 5652 40224 5704
rect 40276 5692 40282 5704
rect 40681 5695 40739 5701
rect 40681 5692 40693 5695
rect 40276 5664 40693 5692
rect 40276 5652 40282 5664
rect 40681 5661 40693 5664
rect 40727 5692 40739 5695
rect 40862 5692 40868 5704
rect 40727 5664 40868 5692
rect 40727 5661 40739 5664
rect 40681 5655 40739 5661
rect 40862 5652 40868 5664
rect 40920 5652 40926 5704
rect 41138 5652 41144 5704
rect 41196 5692 41202 5704
rect 43714 5692 43720 5704
rect 41196 5664 43720 5692
rect 41196 5652 41202 5664
rect 43714 5652 43720 5664
rect 43772 5652 43778 5704
rect 44450 5652 44456 5704
rect 44508 5692 44514 5704
rect 46584 5692 46612 5800
rect 52822 5788 52828 5840
rect 52880 5828 52886 5840
rect 53837 5831 53895 5837
rect 53837 5828 53849 5831
rect 52880 5800 53849 5828
rect 52880 5788 52886 5800
rect 53837 5797 53849 5800
rect 53883 5797 53895 5831
rect 54754 5828 54760 5840
rect 53837 5791 53895 5797
rect 54588 5800 54760 5828
rect 46658 5720 46664 5772
rect 46716 5760 46722 5772
rect 47121 5763 47179 5769
rect 46716 5732 46761 5760
rect 46716 5720 46722 5732
rect 47121 5729 47133 5763
rect 47167 5760 47179 5763
rect 48038 5760 48044 5772
rect 47167 5732 48044 5760
rect 47167 5729 47179 5732
rect 47121 5723 47179 5729
rect 48038 5720 48044 5732
rect 48096 5720 48102 5772
rect 48222 5720 48228 5772
rect 48280 5760 48286 5772
rect 48961 5763 49019 5769
rect 48961 5760 48973 5763
rect 48280 5732 48973 5760
rect 48280 5720 48286 5732
rect 48961 5729 48973 5732
rect 49007 5760 49019 5763
rect 49513 5763 49571 5769
rect 49513 5760 49525 5763
rect 49007 5732 49525 5760
rect 49007 5729 49019 5732
rect 48961 5723 49019 5729
rect 49513 5729 49525 5732
rect 49559 5760 49571 5763
rect 49694 5760 49700 5772
rect 49559 5732 49700 5760
rect 49559 5729 49571 5732
rect 49513 5723 49571 5729
rect 49694 5720 49700 5732
rect 49752 5720 49758 5772
rect 50246 5760 50252 5772
rect 50207 5732 50252 5760
rect 50246 5720 50252 5732
rect 50304 5760 50310 5772
rect 50430 5760 50436 5772
rect 50304 5732 50436 5760
rect 50304 5720 50310 5732
rect 50430 5720 50436 5732
rect 50488 5720 50494 5772
rect 50890 5760 50896 5772
rect 50851 5732 50896 5760
rect 50890 5720 50896 5732
rect 50948 5720 50954 5772
rect 51810 5720 51816 5772
rect 51868 5760 51874 5772
rect 53009 5763 53067 5769
rect 53009 5760 53021 5763
rect 51868 5732 53021 5760
rect 51868 5720 51874 5732
rect 53009 5729 53021 5732
rect 53055 5729 53067 5763
rect 53374 5760 53380 5772
rect 53287 5732 53380 5760
rect 53009 5723 53067 5729
rect 53374 5720 53380 5732
rect 53432 5760 53438 5772
rect 54588 5769 54616 5800
rect 54754 5788 54760 5800
rect 54812 5828 54818 5840
rect 55033 5831 55091 5837
rect 55033 5828 55045 5831
rect 54812 5800 55045 5828
rect 54812 5788 54818 5800
rect 55033 5797 55045 5800
rect 55079 5828 55091 5831
rect 55122 5828 55128 5840
rect 55079 5800 55128 5828
rect 55079 5797 55091 5800
rect 55033 5791 55091 5797
rect 55122 5788 55128 5800
rect 55180 5788 55186 5840
rect 55600 5769 55628 5868
rect 55858 5856 55864 5908
rect 55916 5896 55922 5908
rect 57057 5899 57115 5905
rect 57057 5896 57069 5899
rect 55916 5868 57069 5896
rect 55916 5856 55922 5868
rect 57057 5865 57069 5868
rect 57103 5896 57115 5899
rect 57790 5896 57796 5908
rect 57103 5868 57796 5896
rect 57103 5865 57115 5868
rect 57057 5859 57115 5865
rect 57790 5856 57796 5868
rect 57848 5856 57854 5908
rect 57974 5856 57980 5908
rect 58032 5896 58038 5908
rect 58342 5896 58348 5908
rect 58032 5868 58348 5896
rect 58032 5856 58038 5868
rect 58342 5856 58348 5868
rect 58400 5856 58406 5908
rect 58710 5856 58716 5908
rect 58768 5896 58774 5908
rect 58805 5899 58863 5905
rect 58805 5896 58817 5899
rect 58768 5868 58817 5896
rect 58768 5856 58774 5868
rect 58805 5865 58817 5868
rect 58851 5865 58863 5899
rect 58805 5859 58863 5865
rect 55766 5788 55772 5840
rect 55824 5828 55830 5840
rect 56597 5831 56655 5837
rect 56597 5828 56609 5831
rect 55824 5800 56609 5828
rect 55824 5788 55830 5800
rect 56597 5797 56609 5800
rect 56643 5828 56655 5831
rect 57330 5828 57336 5840
rect 56643 5800 57336 5828
rect 56643 5797 56655 5800
rect 56597 5791 56655 5797
rect 57330 5788 57336 5800
rect 57388 5788 57394 5840
rect 57606 5788 57612 5840
rect 57664 5828 57670 5840
rect 57664 5800 60136 5828
rect 57664 5788 57670 5800
rect 54205 5763 54263 5769
rect 54205 5760 54217 5763
rect 53432 5732 54217 5760
rect 53432 5720 53438 5732
rect 54205 5729 54217 5732
rect 54251 5729 54263 5763
rect 54205 5723 54263 5729
rect 54573 5763 54631 5769
rect 54573 5729 54585 5763
rect 54619 5729 54631 5763
rect 54573 5723 54631 5729
rect 55585 5763 55643 5769
rect 55585 5729 55597 5763
rect 55631 5760 55643 5763
rect 56502 5760 56508 5772
rect 55631 5732 56508 5760
rect 55631 5729 55643 5732
rect 55585 5723 55643 5729
rect 56502 5720 56508 5732
rect 56560 5720 56566 5772
rect 57701 5763 57759 5769
rect 57701 5729 57713 5763
rect 57747 5760 57759 5763
rect 57790 5760 57796 5772
rect 57747 5732 57796 5760
rect 57747 5729 57759 5732
rect 57701 5723 57759 5729
rect 57790 5720 57796 5732
rect 57848 5720 57854 5772
rect 57977 5763 58035 5769
rect 57977 5729 57989 5763
rect 58023 5760 58035 5763
rect 58066 5760 58072 5772
rect 58023 5732 58072 5760
rect 58023 5729 58035 5732
rect 57977 5723 58035 5729
rect 58066 5720 58072 5732
rect 58124 5720 58130 5772
rect 58250 5720 58256 5772
rect 58308 5760 58314 5772
rect 58894 5760 58900 5772
rect 58308 5732 58900 5760
rect 58308 5720 58314 5732
rect 58894 5720 58900 5732
rect 58952 5760 58958 5772
rect 58989 5763 59047 5769
rect 58989 5760 59001 5763
rect 58952 5732 59001 5760
rect 58952 5720 58958 5732
rect 58989 5729 59001 5732
rect 59035 5729 59047 5763
rect 58989 5723 59047 5729
rect 46750 5692 46756 5704
rect 44508 5664 46612 5692
rect 46663 5664 46756 5692
rect 44508 5652 44514 5664
rect 46750 5652 46756 5664
rect 46808 5692 46814 5704
rect 48133 5695 48191 5701
rect 48133 5692 48145 5695
rect 46808 5664 48145 5692
rect 46808 5652 46814 5664
rect 48133 5661 48145 5664
rect 48179 5661 48191 5695
rect 48133 5655 48191 5661
rect 49142 5652 49148 5704
rect 49200 5692 49206 5704
rect 53469 5695 53527 5701
rect 49200 5664 53420 5692
rect 49200 5652 49206 5664
rect 39114 5624 39120 5636
rect 37200 5596 39120 5624
rect 37093 5587 37151 5593
rect 39114 5584 39120 5596
rect 39172 5584 39178 5636
rect 40770 5584 40776 5636
rect 40828 5624 40834 5636
rect 42797 5627 42855 5633
rect 42797 5624 42809 5627
rect 40828 5596 42809 5624
rect 40828 5584 40834 5596
rect 42797 5593 42809 5596
rect 42843 5593 42855 5627
rect 42797 5587 42855 5593
rect 42886 5584 42892 5636
rect 42944 5624 42950 5636
rect 44637 5627 44695 5633
rect 44637 5624 44649 5627
rect 42944 5596 44649 5624
rect 42944 5584 42950 5596
rect 44637 5593 44649 5596
rect 44683 5624 44695 5627
rect 44726 5624 44732 5636
rect 44683 5596 44732 5624
rect 44683 5593 44695 5596
rect 44637 5587 44695 5593
rect 44726 5584 44732 5596
rect 44784 5584 44790 5636
rect 44818 5584 44824 5636
rect 44876 5624 44882 5636
rect 48682 5624 48688 5636
rect 44876 5596 44921 5624
rect 45296 5596 48688 5624
rect 44876 5584 44882 5596
rect 23934 5556 23940 5568
rect 21867 5528 23152 5556
rect 23895 5528 23940 5556
rect 21867 5525 21879 5528
rect 21821 5519 21879 5525
rect 23934 5516 23940 5528
rect 23992 5516 23998 5568
rect 24026 5516 24032 5568
rect 24084 5556 24090 5568
rect 26602 5556 26608 5568
rect 24084 5528 26608 5556
rect 24084 5516 24090 5528
rect 26602 5516 26608 5528
rect 26660 5516 26666 5568
rect 26786 5516 26792 5568
rect 26844 5556 26850 5568
rect 26881 5559 26939 5565
rect 26881 5556 26893 5559
rect 26844 5528 26893 5556
rect 26844 5516 26850 5528
rect 26881 5525 26893 5528
rect 26927 5525 26939 5559
rect 27798 5556 27804 5568
rect 27759 5528 27804 5556
rect 26881 5519 26939 5525
rect 27798 5516 27804 5528
rect 27856 5516 27862 5568
rect 27982 5516 27988 5568
rect 28040 5556 28046 5568
rect 29270 5556 29276 5568
rect 28040 5528 29276 5556
rect 28040 5516 28046 5528
rect 29270 5516 29276 5528
rect 29328 5516 29334 5568
rect 29546 5516 29552 5568
rect 29604 5556 29610 5568
rect 30282 5556 30288 5568
rect 29604 5528 30288 5556
rect 29604 5516 29610 5528
rect 30282 5516 30288 5528
rect 30340 5556 30346 5568
rect 30469 5559 30527 5565
rect 30469 5556 30481 5559
rect 30340 5528 30481 5556
rect 30340 5516 30346 5528
rect 30469 5525 30481 5528
rect 30515 5525 30527 5559
rect 31110 5556 31116 5568
rect 31071 5528 31116 5556
rect 30469 5519 30527 5525
rect 31110 5516 31116 5528
rect 31168 5516 31174 5568
rect 31846 5556 31852 5568
rect 31807 5528 31852 5556
rect 31846 5516 31852 5528
rect 31904 5516 31910 5568
rect 32582 5516 32588 5568
rect 32640 5556 32646 5568
rect 32677 5559 32735 5565
rect 32677 5556 32689 5559
rect 32640 5528 32689 5556
rect 32640 5516 32646 5528
rect 32677 5525 32689 5528
rect 32723 5525 32735 5559
rect 32677 5519 32735 5525
rect 32766 5516 32772 5568
rect 32824 5556 32830 5568
rect 33413 5559 33471 5565
rect 33413 5556 33425 5559
rect 32824 5528 33425 5556
rect 32824 5516 32830 5528
rect 33413 5525 33425 5528
rect 33459 5556 33471 5559
rect 33502 5556 33508 5568
rect 33459 5528 33508 5556
rect 33459 5525 33471 5528
rect 33413 5519 33471 5525
rect 33502 5516 33508 5528
rect 33560 5516 33566 5568
rect 34241 5559 34299 5565
rect 34241 5525 34253 5559
rect 34287 5556 34299 5559
rect 34514 5556 34520 5568
rect 34287 5528 34520 5556
rect 34287 5525 34299 5528
rect 34241 5519 34299 5525
rect 34514 5516 34520 5528
rect 34572 5556 34578 5568
rect 34974 5556 34980 5568
rect 34572 5528 34980 5556
rect 34572 5516 34578 5528
rect 34974 5516 34980 5528
rect 35032 5516 35038 5568
rect 35250 5516 35256 5568
rect 35308 5556 35314 5568
rect 35710 5556 35716 5568
rect 35308 5528 35716 5556
rect 35308 5516 35314 5528
rect 35710 5516 35716 5528
rect 35768 5516 35774 5568
rect 35894 5516 35900 5568
rect 35952 5556 35958 5568
rect 36081 5559 36139 5565
rect 36081 5556 36093 5559
rect 35952 5528 36093 5556
rect 35952 5516 35958 5528
rect 36081 5525 36093 5528
rect 36127 5556 36139 5559
rect 36354 5556 36360 5568
rect 36127 5528 36360 5556
rect 36127 5525 36139 5528
rect 36081 5519 36139 5525
rect 36354 5516 36360 5528
rect 36412 5556 36418 5568
rect 36449 5559 36507 5565
rect 36449 5556 36461 5559
rect 36412 5528 36461 5556
rect 36412 5516 36418 5528
rect 36449 5525 36461 5528
rect 36495 5525 36507 5559
rect 36722 5556 36728 5568
rect 36683 5528 36728 5556
rect 36449 5519 36507 5525
rect 36722 5516 36728 5528
rect 36780 5516 36786 5568
rect 37918 5556 37924 5568
rect 37879 5528 37924 5556
rect 37918 5516 37924 5528
rect 37976 5516 37982 5568
rect 38378 5516 38384 5568
rect 38436 5556 38442 5568
rect 38746 5556 38752 5568
rect 38436 5528 38752 5556
rect 38436 5516 38442 5528
rect 38746 5516 38752 5528
rect 38804 5516 38810 5568
rect 39209 5559 39267 5565
rect 39209 5525 39221 5559
rect 39255 5556 39267 5559
rect 40586 5556 40592 5568
rect 39255 5528 40592 5556
rect 39255 5525 39267 5528
rect 39209 5519 39267 5525
rect 40586 5516 40592 5528
rect 40644 5516 40650 5568
rect 41325 5559 41383 5565
rect 41325 5525 41337 5559
rect 41371 5556 41383 5559
rect 41782 5556 41788 5568
rect 41371 5528 41788 5556
rect 41371 5525 41383 5528
rect 41325 5519 41383 5525
rect 41782 5516 41788 5528
rect 41840 5516 41846 5568
rect 45296 5565 45324 5596
rect 48682 5584 48688 5596
rect 48740 5584 48746 5636
rect 48777 5627 48835 5633
rect 48777 5593 48789 5627
rect 48823 5624 48835 5627
rect 49326 5624 49332 5636
rect 48823 5596 49332 5624
rect 48823 5593 48835 5596
rect 48777 5587 48835 5593
rect 49326 5584 49332 5596
rect 49384 5584 49390 5636
rect 50246 5584 50252 5636
rect 50304 5624 50310 5636
rect 50982 5624 50988 5636
rect 50304 5596 50988 5624
rect 50304 5584 50310 5596
rect 50982 5584 50988 5596
rect 51040 5624 51046 5636
rect 52273 5627 52331 5633
rect 52273 5624 52285 5627
rect 51040 5596 52285 5624
rect 51040 5584 51046 5596
rect 52273 5593 52285 5596
rect 52319 5593 52331 5627
rect 52273 5587 52331 5593
rect 52825 5627 52883 5633
rect 52825 5593 52837 5627
rect 52871 5624 52883 5627
rect 53282 5624 53288 5636
rect 52871 5596 53288 5624
rect 52871 5593 52883 5596
rect 52825 5587 52883 5593
rect 53282 5584 53288 5596
rect 53340 5584 53346 5636
rect 53392 5624 53420 5664
rect 53469 5661 53481 5695
rect 53515 5692 53527 5695
rect 53834 5692 53840 5704
rect 53515 5664 53840 5692
rect 53515 5661 53527 5664
rect 53469 5655 53527 5661
rect 53834 5652 53840 5664
rect 53892 5652 53898 5704
rect 54938 5652 54944 5704
rect 54996 5692 55002 5704
rect 55953 5695 56011 5701
rect 54996 5664 55904 5692
rect 54996 5652 55002 5664
rect 55582 5624 55588 5636
rect 53392 5596 55588 5624
rect 55582 5584 55588 5596
rect 55640 5584 55646 5636
rect 55766 5633 55772 5636
rect 55750 5627 55772 5633
rect 55750 5593 55762 5627
rect 55750 5587 55772 5593
rect 55766 5584 55772 5587
rect 55824 5584 55830 5636
rect 55876 5624 55904 5664
rect 55953 5661 55965 5695
rect 55999 5692 56011 5695
rect 56134 5692 56140 5704
rect 55999 5664 56140 5692
rect 55999 5661 56011 5664
rect 55953 5655 56011 5661
rect 56134 5652 56140 5664
rect 56192 5652 56198 5704
rect 57146 5692 57152 5704
rect 57107 5664 57152 5692
rect 57146 5652 57152 5664
rect 57204 5652 57210 5704
rect 58158 5692 58164 5704
rect 58071 5664 58164 5692
rect 58158 5652 58164 5664
rect 58216 5692 58222 5704
rect 58437 5695 58495 5701
rect 58437 5692 58449 5695
rect 58216 5664 58449 5692
rect 58216 5652 58222 5664
rect 58437 5661 58449 5664
rect 58483 5661 58495 5695
rect 58437 5655 58495 5661
rect 58176 5624 58204 5652
rect 59630 5624 59636 5636
rect 55876 5596 58204 5624
rect 59188 5596 59636 5624
rect 45281 5559 45339 5565
rect 45281 5525 45293 5559
rect 45327 5525 45339 5559
rect 45281 5519 45339 5525
rect 46106 5516 46112 5568
rect 46164 5556 46170 5568
rect 46201 5559 46259 5565
rect 46201 5556 46213 5559
rect 46164 5528 46213 5556
rect 46164 5516 46170 5528
rect 46201 5525 46213 5528
rect 46247 5525 46259 5559
rect 46201 5519 46259 5525
rect 46658 5516 46664 5568
rect 46716 5556 46722 5568
rect 47489 5559 47547 5565
rect 47489 5556 47501 5559
rect 46716 5528 47501 5556
rect 46716 5516 46722 5528
rect 47489 5525 47501 5528
rect 47535 5556 47547 5559
rect 47762 5556 47768 5568
rect 47535 5528 47768 5556
rect 47535 5525 47547 5528
rect 47489 5519 47547 5525
rect 47762 5516 47768 5528
rect 47820 5516 47826 5568
rect 47857 5559 47915 5565
rect 47857 5525 47869 5559
rect 47903 5556 47915 5559
rect 47946 5556 47952 5568
rect 47903 5528 47952 5556
rect 47903 5525 47915 5528
rect 47857 5519 47915 5525
rect 47946 5516 47952 5528
rect 48004 5516 48010 5568
rect 48406 5516 48412 5568
rect 48464 5556 48470 5568
rect 50154 5556 50160 5568
rect 48464 5528 50160 5556
rect 48464 5516 48470 5528
rect 50154 5516 50160 5528
rect 50212 5516 50218 5568
rect 50338 5556 50344 5568
rect 50299 5528 50344 5556
rect 50338 5516 50344 5528
rect 50396 5516 50402 5568
rect 51353 5559 51411 5565
rect 51353 5525 51365 5559
rect 51399 5556 51411 5559
rect 51442 5556 51448 5568
rect 51399 5528 51448 5556
rect 51399 5525 51411 5528
rect 51353 5519 51411 5525
rect 51442 5516 51448 5528
rect 51500 5556 51506 5568
rect 51721 5559 51779 5565
rect 51721 5556 51733 5559
rect 51500 5528 51733 5556
rect 51500 5516 51506 5528
rect 51721 5525 51733 5528
rect 51767 5525 51779 5559
rect 54662 5556 54668 5568
rect 54623 5528 54668 5556
rect 51721 5519 51779 5525
rect 54662 5516 54668 5528
rect 54720 5516 54726 5568
rect 55490 5556 55496 5568
rect 55451 5528 55496 5556
rect 55490 5516 55496 5528
rect 55548 5516 55554 5568
rect 55861 5559 55919 5565
rect 55861 5525 55873 5559
rect 55907 5556 55919 5559
rect 56042 5556 56048 5568
rect 55907 5528 56048 5556
rect 55907 5525 55919 5528
rect 55861 5519 55919 5525
rect 56042 5516 56048 5528
rect 56100 5516 56106 5568
rect 56226 5556 56232 5568
rect 56187 5528 56232 5556
rect 56226 5516 56232 5528
rect 56284 5516 56290 5568
rect 56594 5516 56600 5568
rect 56652 5556 56658 5568
rect 59188 5565 59216 5596
rect 59630 5584 59636 5596
rect 59688 5584 59694 5636
rect 59173 5559 59231 5565
rect 59173 5556 59185 5559
rect 56652 5528 59185 5556
rect 56652 5516 56658 5528
rect 59173 5525 59185 5528
rect 59219 5525 59231 5559
rect 59173 5519 59231 5525
rect 59262 5516 59268 5568
rect 59320 5556 59326 5568
rect 59541 5559 59599 5565
rect 59541 5556 59553 5559
rect 59320 5528 59553 5556
rect 59320 5516 59326 5528
rect 59541 5525 59553 5528
rect 59587 5525 59599 5559
rect 59541 5519 59599 5525
rect 59722 5516 59728 5568
rect 59780 5556 59786 5568
rect 59909 5559 59967 5565
rect 59909 5556 59921 5559
rect 59780 5528 59921 5556
rect 59780 5516 59786 5528
rect 59909 5525 59921 5528
rect 59955 5525 59967 5559
rect 60108 5556 60136 5800
rect 60185 5763 60243 5769
rect 60185 5729 60197 5763
rect 60231 5760 60243 5763
rect 61286 5760 61292 5772
rect 60231 5732 61292 5760
rect 60231 5729 60243 5732
rect 60185 5723 60243 5729
rect 61286 5720 61292 5732
rect 61344 5720 61350 5772
rect 60458 5692 60464 5704
rect 60419 5664 60464 5692
rect 60458 5652 60464 5664
rect 60516 5652 60522 5704
rect 61746 5556 61752 5568
rect 60108 5528 61752 5556
rect 59909 5519 59967 5525
rect 61746 5516 61752 5528
rect 61804 5516 61810 5568
rect 1104 5466 63480 5488
rect 1104 5414 11378 5466
rect 11430 5414 11442 5466
rect 11494 5414 11506 5466
rect 11558 5414 11570 5466
rect 11622 5414 32170 5466
rect 32222 5414 32234 5466
rect 32286 5414 32298 5466
rect 32350 5414 32362 5466
rect 32414 5414 52962 5466
rect 53014 5414 53026 5466
rect 53078 5414 53090 5466
rect 53142 5414 53154 5466
rect 53206 5414 63480 5466
rect 1104 5392 63480 5414
rect 2317 5355 2375 5361
rect 2317 5321 2329 5355
rect 2363 5352 2375 5355
rect 2682 5352 2688 5364
rect 2363 5324 2688 5352
rect 2363 5321 2375 5324
rect 2317 5315 2375 5321
rect 2682 5312 2688 5324
rect 2740 5312 2746 5364
rect 4062 5312 4068 5364
rect 4120 5352 4126 5364
rect 14090 5352 14096 5364
rect 4120 5324 14096 5352
rect 4120 5312 4126 5324
rect 14090 5312 14096 5324
rect 14148 5312 14154 5364
rect 14461 5355 14519 5361
rect 14461 5321 14473 5355
rect 14507 5352 14519 5355
rect 15010 5352 15016 5364
rect 14507 5324 15016 5352
rect 14507 5321 14519 5324
rect 14461 5315 14519 5321
rect 15010 5312 15016 5324
rect 15068 5312 15074 5364
rect 16298 5312 16304 5364
rect 16356 5352 16362 5364
rect 16393 5355 16451 5361
rect 16393 5352 16405 5355
rect 16356 5324 16405 5352
rect 16356 5312 16362 5324
rect 16393 5321 16405 5324
rect 16439 5321 16451 5355
rect 18049 5355 18107 5361
rect 18049 5352 18061 5355
rect 16393 5315 16451 5321
rect 17420 5324 18061 5352
rect 4982 5284 4988 5296
rect 4943 5256 4988 5284
rect 4982 5244 4988 5256
rect 5040 5244 5046 5296
rect 5166 5244 5172 5296
rect 5224 5284 5230 5296
rect 5261 5287 5319 5293
rect 5261 5284 5273 5287
rect 5224 5256 5273 5284
rect 5224 5244 5230 5256
rect 5261 5253 5273 5256
rect 5307 5253 5319 5287
rect 6178 5284 6184 5296
rect 6139 5256 6184 5284
rect 5261 5247 5319 5253
rect 6178 5244 6184 5256
rect 6236 5244 6242 5296
rect 7742 5244 7748 5296
rect 7800 5284 7806 5296
rect 7837 5287 7895 5293
rect 7837 5284 7849 5287
rect 7800 5256 7849 5284
rect 7800 5244 7806 5256
rect 7837 5253 7849 5256
rect 7883 5253 7895 5287
rect 8294 5284 8300 5296
rect 8207 5256 8300 5284
rect 7837 5247 7895 5253
rect 8294 5244 8300 5256
rect 8352 5284 8358 5296
rect 9490 5284 9496 5296
rect 8352 5256 9496 5284
rect 8352 5244 8358 5256
rect 9490 5244 9496 5256
rect 9548 5244 9554 5296
rect 11882 5284 11888 5296
rect 11843 5256 11888 5284
rect 11882 5244 11888 5256
rect 11940 5244 11946 5296
rect 14829 5287 14887 5293
rect 14829 5253 14841 5287
rect 14875 5284 14887 5287
rect 14875 5256 15700 5284
rect 14875 5253 14887 5256
rect 14829 5247 14887 5253
rect 7193 5219 7251 5225
rect 7193 5185 7205 5219
rect 7239 5216 7251 5219
rect 7926 5216 7932 5228
rect 7239 5188 7932 5216
rect 7239 5185 7251 5188
rect 7193 5179 7251 5185
rect 7926 5176 7932 5188
rect 7984 5176 7990 5228
rect 9398 5216 9404 5228
rect 9359 5188 9404 5216
rect 9398 5176 9404 5188
rect 9456 5176 9462 5228
rect 9766 5176 9772 5228
rect 9824 5216 9830 5228
rect 9824 5188 10456 5216
rect 9824 5176 9830 5188
rect 2314 5108 2320 5160
rect 2372 5148 2378 5160
rect 2961 5151 3019 5157
rect 2961 5148 2973 5151
rect 2372 5120 2973 5148
rect 2372 5108 2378 5120
rect 2961 5117 2973 5120
rect 3007 5117 3019 5151
rect 2961 5111 3019 5117
rect 3237 5151 3295 5157
rect 3237 5117 3249 5151
rect 3283 5148 3295 5151
rect 3510 5148 3516 5160
rect 3283 5120 3516 5148
rect 3283 5117 3295 5120
rect 3237 5111 3295 5117
rect 3510 5108 3516 5120
rect 3568 5148 3574 5160
rect 4062 5148 4068 5160
rect 3568 5120 4068 5148
rect 3568 5108 3574 5120
rect 4062 5108 4068 5120
rect 4120 5108 4126 5160
rect 5626 5148 5632 5160
rect 5587 5120 5632 5148
rect 5626 5108 5632 5120
rect 5684 5108 5690 5160
rect 7006 5148 7012 5160
rect 6967 5120 7012 5148
rect 7006 5108 7012 5120
rect 7064 5108 7070 5160
rect 7561 5151 7619 5157
rect 7561 5117 7573 5151
rect 7607 5148 7619 5151
rect 8018 5148 8024 5160
rect 7607 5120 8024 5148
rect 7607 5117 7619 5120
rect 7561 5111 7619 5117
rect 8018 5108 8024 5120
rect 8076 5108 8082 5160
rect 8481 5151 8539 5157
rect 8481 5117 8493 5151
rect 8527 5148 8539 5151
rect 8846 5148 8852 5160
rect 8527 5120 8852 5148
rect 8527 5117 8539 5120
rect 8481 5111 8539 5117
rect 8846 5108 8852 5120
rect 8904 5108 8910 5160
rect 9306 5148 9312 5160
rect 9219 5120 9312 5148
rect 9306 5108 9312 5120
rect 9364 5108 9370 5160
rect 10318 5148 10324 5160
rect 10244 5120 10324 5148
rect 8294 5080 8300 5092
rect 4448 5052 8300 5080
rect 2590 4972 2596 5024
rect 2648 5012 2654 5024
rect 2685 5015 2743 5021
rect 2685 5012 2697 5015
rect 2648 4984 2697 5012
rect 2648 4972 2654 4984
rect 2685 4981 2697 4984
rect 2731 5012 2743 5015
rect 4448 5012 4476 5052
rect 8294 5040 8300 5052
rect 8352 5040 8358 5092
rect 8570 5080 8576 5092
rect 8531 5052 8576 5080
rect 8570 5040 8576 5052
rect 8628 5040 8634 5092
rect 9324 5080 9352 5108
rect 10244 5080 10272 5120
rect 10318 5108 10324 5120
rect 10376 5108 10382 5160
rect 10428 5157 10456 5188
rect 10502 5176 10508 5228
rect 10560 5216 10566 5228
rect 10873 5219 10931 5225
rect 10873 5216 10885 5219
rect 10560 5188 10885 5216
rect 10560 5176 10566 5188
rect 10873 5185 10885 5188
rect 10919 5185 10931 5219
rect 10873 5179 10931 5185
rect 12342 5176 12348 5228
rect 12400 5216 12406 5228
rect 12437 5219 12495 5225
rect 12437 5216 12449 5219
rect 12400 5188 12449 5216
rect 12400 5176 12406 5188
rect 12437 5185 12449 5188
rect 12483 5185 12495 5219
rect 12437 5179 12495 5185
rect 12713 5219 12771 5225
rect 12713 5185 12725 5219
rect 12759 5216 12771 5219
rect 12802 5216 12808 5228
rect 12759 5188 12808 5216
rect 12759 5185 12771 5188
rect 12713 5179 12771 5185
rect 12802 5176 12808 5188
rect 12860 5216 12866 5228
rect 15672 5225 15700 5256
rect 15838 5244 15844 5296
rect 15896 5284 15902 5296
rect 17420 5293 17448 5324
rect 18049 5321 18061 5324
rect 18095 5352 18107 5355
rect 18138 5352 18144 5364
rect 18095 5324 18144 5352
rect 18095 5321 18107 5324
rect 18049 5315 18107 5321
rect 18138 5312 18144 5324
rect 18196 5352 18202 5364
rect 18877 5355 18935 5361
rect 18877 5352 18889 5355
rect 18196 5324 18889 5352
rect 18196 5312 18202 5324
rect 18877 5321 18889 5324
rect 18923 5321 18935 5355
rect 19058 5352 19064 5364
rect 19019 5324 19064 5352
rect 18877 5315 18935 5321
rect 19058 5312 19064 5324
rect 19116 5312 19122 5364
rect 19150 5312 19156 5364
rect 19208 5352 19214 5364
rect 20806 5352 20812 5364
rect 19208 5324 20812 5352
rect 19208 5312 19214 5324
rect 20806 5312 20812 5324
rect 20864 5352 20870 5364
rect 20864 5324 22140 5352
rect 20864 5312 20870 5324
rect 17405 5287 17463 5293
rect 17405 5284 17417 5287
rect 15896 5256 17417 5284
rect 15896 5244 15902 5256
rect 17405 5253 17417 5256
rect 17451 5253 17463 5287
rect 17405 5247 17463 5253
rect 18598 5244 18604 5296
rect 18656 5284 18662 5296
rect 20254 5284 20260 5296
rect 18656 5256 20260 5284
rect 18656 5244 18662 5256
rect 20254 5244 20260 5256
rect 20312 5244 20318 5296
rect 21910 5284 21916 5296
rect 20364 5256 21916 5284
rect 14921 5219 14979 5225
rect 14921 5216 14933 5219
rect 12860 5188 14933 5216
rect 12860 5176 12866 5188
rect 14921 5185 14933 5188
rect 14967 5185 14979 5219
rect 14921 5179 14979 5185
rect 15657 5219 15715 5225
rect 15657 5185 15669 5219
rect 15703 5216 15715 5219
rect 18785 5219 18843 5225
rect 18785 5216 18797 5219
rect 15703 5188 18797 5216
rect 15703 5185 15715 5188
rect 15657 5179 15715 5185
rect 18785 5185 18797 5188
rect 18831 5185 18843 5219
rect 18785 5179 18843 5185
rect 18877 5219 18935 5225
rect 18877 5185 18889 5219
rect 18923 5216 18935 5219
rect 19334 5216 19340 5228
rect 18923 5188 19340 5216
rect 18923 5185 18935 5188
rect 18877 5179 18935 5185
rect 19334 5176 19340 5188
rect 19392 5216 19398 5228
rect 19429 5219 19487 5225
rect 19429 5216 19441 5219
rect 19392 5188 19441 5216
rect 19392 5176 19398 5188
rect 19429 5185 19441 5188
rect 19475 5185 19487 5219
rect 20364 5216 20392 5256
rect 21910 5244 21916 5256
rect 21968 5244 21974 5296
rect 22112 5284 22140 5324
rect 22186 5312 22192 5364
rect 22244 5352 22250 5364
rect 24029 5355 24087 5361
rect 24029 5352 24041 5355
rect 22244 5324 24041 5352
rect 22244 5312 22250 5324
rect 24029 5321 24041 5324
rect 24075 5321 24087 5355
rect 24210 5352 24216 5364
rect 24171 5324 24216 5352
rect 24029 5315 24087 5321
rect 24210 5312 24216 5324
rect 24268 5312 24274 5364
rect 27246 5352 27252 5364
rect 24504 5324 27252 5352
rect 24504 5284 24532 5324
rect 27246 5312 27252 5324
rect 27304 5312 27310 5364
rect 28166 5312 28172 5364
rect 28224 5352 28230 5364
rect 32217 5355 32275 5361
rect 28224 5324 31340 5352
rect 28224 5312 28230 5324
rect 24670 5284 24676 5296
rect 22112 5256 24532 5284
rect 24631 5256 24676 5284
rect 24670 5244 24676 5256
rect 24728 5244 24734 5296
rect 26786 5244 26792 5296
rect 26844 5284 26850 5296
rect 26881 5287 26939 5293
rect 26881 5284 26893 5287
rect 26844 5256 26893 5284
rect 26844 5244 26850 5256
rect 26881 5253 26893 5256
rect 26927 5253 26939 5287
rect 26881 5247 26939 5253
rect 28721 5287 28779 5293
rect 28721 5253 28733 5287
rect 28767 5284 28779 5287
rect 29086 5284 29092 5296
rect 28767 5256 29092 5284
rect 28767 5253 28779 5256
rect 28721 5247 28779 5253
rect 29086 5244 29092 5256
rect 29144 5284 29150 5296
rect 31205 5287 31263 5293
rect 31205 5284 31217 5287
rect 29144 5256 31217 5284
rect 29144 5244 29150 5256
rect 31205 5253 31217 5256
rect 31251 5253 31263 5287
rect 31312 5284 31340 5324
rect 32217 5321 32229 5355
rect 32263 5352 32275 5355
rect 32490 5352 32496 5364
rect 32263 5324 32496 5352
rect 32263 5321 32275 5324
rect 32217 5315 32275 5321
rect 32490 5312 32496 5324
rect 32548 5312 32554 5364
rect 32858 5312 32864 5364
rect 32916 5352 32922 5364
rect 34425 5355 34483 5361
rect 34425 5352 34437 5355
rect 32916 5324 34437 5352
rect 32916 5312 32922 5324
rect 34425 5321 34437 5324
rect 34471 5321 34483 5355
rect 34425 5315 34483 5321
rect 35342 5312 35348 5364
rect 35400 5352 35406 5364
rect 35621 5355 35679 5361
rect 35621 5352 35633 5355
rect 35400 5324 35633 5352
rect 35400 5312 35406 5324
rect 35621 5321 35633 5324
rect 35667 5321 35679 5355
rect 35986 5352 35992 5364
rect 35947 5324 35992 5352
rect 35621 5315 35679 5321
rect 35986 5312 35992 5324
rect 36044 5312 36050 5364
rect 36446 5312 36452 5364
rect 36504 5352 36510 5364
rect 37734 5352 37740 5364
rect 36504 5324 37740 5352
rect 36504 5312 36510 5324
rect 37734 5312 37740 5324
rect 37792 5312 37798 5364
rect 38010 5312 38016 5364
rect 38068 5352 38074 5364
rect 39393 5355 39451 5361
rect 39393 5352 39405 5355
rect 38068 5324 39405 5352
rect 38068 5312 38074 5324
rect 39393 5321 39405 5324
rect 39439 5321 39451 5355
rect 39574 5352 39580 5364
rect 39535 5324 39580 5352
rect 39393 5315 39451 5321
rect 39574 5312 39580 5324
rect 39632 5312 39638 5364
rect 39758 5312 39764 5364
rect 39816 5352 39822 5364
rect 39945 5355 40003 5361
rect 39945 5352 39957 5355
rect 39816 5324 39957 5352
rect 39816 5312 39822 5324
rect 39945 5321 39957 5324
rect 39991 5321 40003 5355
rect 39945 5315 40003 5321
rect 40862 5312 40868 5364
rect 40920 5352 40926 5364
rect 41417 5355 41475 5361
rect 41417 5352 41429 5355
rect 40920 5324 41429 5352
rect 40920 5312 40926 5324
rect 41417 5321 41429 5324
rect 41463 5321 41475 5355
rect 41782 5352 41788 5364
rect 41743 5324 41788 5352
rect 41417 5315 41475 5321
rect 41782 5312 41788 5324
rect 41840 5312 41846 5364
rect 41966 5312 41972 5364
rect 42024 5352 42030 5364
rect 42705 5355 42763 5361
rect 42705 5352 42717 5355
rect 42024 5324 42717 5352
rect 42024 5312 42030 5324
rect 42705 5321 42717 5324
rect 42751 5321 42763 5355
rect 42705 5315 42763 5321
rect 42886 5312 42892 5364
rect 42944 5352 42950 5364
rect 43073 5355 43131 5361
rect 43073 5352 43085 5355
rect 42944 5324 43085 5352
rect 42944 5312 42950 5324
rect 43073 5321 43085 5324
rect 43119 5321 43131 5355
rect 43073 5315 43131 5321
rect 43346 5312 43352 5364
rect 43404 5352 43410 5364
rect 43533 5355 43591 5361
rect 43533 5352 43545 5355
rect 43404 5324 43545 5352
rect 43404 5312 43410 5324
rect 43533 5321 43545 5324
rect 43579 5352 43591 5355
rect 44269 5355 44327 5361
rect 44269 5352 44281 5355
rect 43579 5324 44281 5352
rect 43579 5321 43591 5324
rect 43533 5315 43591 5321
rect 44269 5321 44281 5324
rect 44315 5352 44327 5355
rect 44450 5352 44456 5364
rect 44315 5324 44456 5352
rect 44315 5321 44327 5324
rect 44269 5315 44327 5321
rect 44450 5312 44456 5324
rect 44508 5312 44514 5364
rect 44726 5312 44732 5364
rect 44784 5352 44790 5364
rect 44913 5355 44971 5361
rect 44913 5352 44925 5355
rect 44784 5324 44925 5352
rect 44784 5312 44790 5324
rect 44913 5321 44925 5324
rect 44959 5321 44971 5355
rect 44913 5315 44971 5321
rect 45002 5312 45008 5364
rect 45060 5352 45066 5364
rect 45833 5355 45891 5361
rect 45833 5352 45845 5355
rect 45060 5324 45845 5352
rect 45060 5312 45066 5324
rect 45833 5321 45845 5324
rect 45879 5321 45891 5355
rect 48866 5352 48872 5364
rect 45833 5315 45891 5321
rect 46216 5324 48872 5352
rect 31662 5284 31668 5296
rect 31312 5256 31668 5284
rect 31205 5247 31263 5253
rect 31662 5244 31668 5256
rect 31720 5244 31726 5296
rect 31938 5244 31944 5296
rect 31996 5284 32002 5296
rect 35250 5284 35256 5296
rect 31996 5256 35256 5284
rect 31996 5244 32002 5256
rect 35250 5244 35256 5256
rect 35308 5244 35314 5296
rect 35437 5287 35495 5293
rect 35437 5253 35449 5287
rect 35483 5284 35495 5287
rect 39022 5284 39028 5296
rect 35483 5256 39028 5284
rect 35483 5253 35495 5256
rect 35437 5247 35495 5253
rect 39022 5244 39028 5256
rect 39080 5244 39086 5296
rect 39114 5244 39120 5296
rect 39172 5284 39178 5296
rect 40770 5284 40776 5296
rect 39172 5256 40776 5284
rect 39172 5244 39178 5256
rect 40770 5244 40776 5256
rect 40828 5244 40834 5296
rect 40954 5244 40960 5296
rect 41012 5284 41018 5296
rect 41984 5284 42012 5312
rect 43898 5284 43904 5296
rect 41012 5256 42012 5284
rect 43859 5256 43904 5284
rect 41012 5244 41018 5256
rect 43898 5244 43904 5256
rect 43956 5244 43962 5296
rect 46106 5284 46112 5296
rect 44468 5256 46112 5284
rect 19429 5179 19487 5185
rect 19536 5188 20392 5216
rect 21269 5219 21327 5225
rect 10413 5151 10471 5157
rect 10413 5117 10425 5151
rect 10459 5117 10471 5151
rect 10413 5111 10471 5117
rect 11609 5151 11667 5157
rect 11609 5117 11621 5151
rect 11655 5148 11667 5151
rect 11698 5148 11704 5160
rect 11655 5120 11704 5148
rect 11655 5117 11667 5120
rect 11609 5111 11667 5117
rect 11698 5108 11704 5120
rect 11756 5148 11762 5160
rect 14550 5148 14556 5160
rect 11756 5120 14556 5148
rect 11756 5108 11762 5120
rect 14550 5108 14556 5120
rect 14608 5108 14614 5160
rect 14642 5108 14648 5160
rect 14700 5148 14706 5160
rect 15562 5148 15568 5160
rect 14700 5120 15568 5148
rect 14700 5108 14706 5120
rect 15562 5108 15568 5120
rect 15620 5108 15626 5160
rect 15930 5148 15936 5160
rect 15891 5120 15936 5148
rect 15930 5108 15936 5120
rect 15988 5108 15994 5160
rect 16022 5108 16028 5160
rect 16080 5148 16086 5160
rect 16761 5151 16819 5157
rect 16761 5148 16773 5151
rect 16080 5120 16773 5148
rect 16080 5108 16086 5120
rect 16761 5117 16773 5120
rect 16807 5117 16819 5151
rect 16761 5111 16819 5117
rect 17770 5108 17776 5160
rect 17828 5148 17834 5160
rect 18325 5151 18383 5157
rect 18325 5148 18337 5151
rect 17828 5120 18337 5148
rect 17828 5108 17834 5120
rect 18325 5117 18337 5120
rect 18371 5117 18383 5151
rect 18325 5111 18383 5117
rect 18506 5108 18512 5160
rect 18564 5148 18570 5160
rect 19536 5148 19564 5188
rect 21269 5185 21281 5219
rect 21315 5216 21327 5219
rect 21542 5216 21548 5228
rect 21315 5188 21548 5216
rect 21315 5185 21327 5188
rect 21269 5179 21327 5185
rect 21542 5176 21548 5188
rect 21600 5176 21606 5228
rect 22278 5176 22284 5228
rect 22336 5216 22342 5228
rect 22830 5216 22836 5228
rect 22336 5188 22836 5216
rect 22336 5176 22342 5188
rect 22830 5176 22836 5188
rect 22888 5176 22894 5228
rect 22922 5176 22928 5228
rect 22980 5216 22986 5228
rect 23109 5219 23167 5225
rect 23109 5216 23121 5219
rect 22980 5188 23121 5216
rect 22980 5176 22986 5188
rect 23109 5185 23121 5188
rect 23155 5216 23167 5219
rect 23155 5188 23704 5216
rect 23155 5185 23167 5188
rect 23109 5179 23167 5185
rect 18564 5120 19564 5148
rect 19613 5151 19671 5157
rect 18564 5108 18570 5120
rect 19613 5117 19625 5151
rect 19659 5148 19671 5151
rect 20346 5148 20352 5160
rect 19659 5120 20352 5148
rect 19659 5117 19671 5120
rect 19613 5111 19671 5117
rect 20346 5108 20352 5120
rect 20404 5108 20410 5160
rect 20714 5108 20720 5160
rect 20772 5148 20778 5160
rect 20901 5151 20959 5157
rect 20901 5148 20913 5151
rect 20772 5120 20913 5148
rect 20772 5108 20778 5120
rect 20901 5117 20913 5120
rect 20947 5117 20959 5151
rect 20901 5111 20959 5117
rect 20990 5108 20996 5160
rect 21048 5148 21054 5160
rect 21453 5151 21511 5157
rect 21453 5148 21465 5151
rect 21048 5120 21465 5148
rect 21048 5108 21054 5120
rect 21453 5117 21465 5120
rect 21499 5148 21511 5151
rect 21913 5151 21971 5157
rect 21913 5148 21925 5151
rect 21499 5120 21925 5148
rect 21499 5117 21511 5120
rect 21453 5111 21511 5117
rect 21913 5117 21925 5120
rect 21959 5148 21971 5151
rect 21959 5120 22416 5148
rect 21959 5117 21971 5120
rect 21913 5111 21971 5117
rect 11149 5083 11207 5089
rect 11149 5080 11161 5083
rect 9324 5052 9904 5080
rect 10244 5052 11161 5080
rect 2731 4984 4476 5012
rect 4525 5015 4583 5021
rect 2731 4981 2743 4984
rect 2685 4975 2743 4981
rect 4525 4981 4537 5015
rect 4571 5012 4583 5015
rect 5350 5012 5356 5024
rect 4571 4984 5356 5012
rect 4571 4981 4583 4984
rect 4525 4975 4583 4981
rect 5350 4972 5356 4984
rect 5408 4972 5414 5024
rect 5810 5012 5816 5024
rect 5771 4984 5816 5012
rect 5810 4972 5816 4984
rect 5868 4972 5874 5024
rect 6641 5015 6699 5021
rect 6641 4981 6653 5015
rect 6687 5012 6699 5015
rect 7834 5012 7840 5024
rect 6687 4984 7840 5012
rect 6687 4981 6699 4984
rect 6641 4975 6699 4981
rect 7834 4972 7840 4984
rect 7892 4972 7898 5024
rect 9876 5021 9904 5052
rect 11149 5049 11161 5052
rect 11195 5080 11207 5083
rect 12066 5080 12072 5092
rect 11195 5052 12072 5080
rect 11195 5049 11207 5052
rect 11149 5043 11207 5049
rect 12066 5040 12072 5052
rect 12124 5040 12130 5092
rect 13630 5040 13636 5092
rect 13688 5080 13694 5092
rect 14093 5083 14151 5089
rect 14093 5080 14105 5083
rect 13688 5052 14105 5080
rect 13688 5040 13694 5052
rect 14093 5049 14105 5052
rect 14139 5080 14151 5083
rect 15948 5080 15976 5108
rect 18230 5080 18236 5092
rect 14139 5052 15976 5080
rect 18143 5052 18236 5080
rect 14139 5049 14151 5052
rect 14093 5043 14151 5049
rect 18230 5040 18236 5052
rect 18288 5040 18294 5092
rect 22186 5080 22192 5092
rect 19352 5052 22192 5080
rect 9861 5015 9919 5021
rect 9861 4981 9873 5015
rect 9907 5012 9919 5015
rect 10042 5012 10048 5024
rect 9907 4984 10048 5012
rect 9907 4981 9919 4984
rect 9861 4975 9919 4981
rect 10042 4972 10048 4984
rect 10100 4972 10106 5024
rect 10226 5012 10232 5024
rect 10139 4984 10232 5012
rect 10226 4972 10232 4984
rect 10284 5012 10290 5024
rect 10962 5012 10968 5024
rect 10284 4984 10968 5012
rect 10284 4972 10290 4984
rect 10962 4972 10968 4984
rect 11020 4972 11026 5024
rect 15746 4972 15752 5024
rect 15804 5012 15810 5024
rect 17773 5015 17831 5021
rect 17773 5012 17785 5015
rect 15804 4984 17785 5012
rect 15804 4972 15810 4984
rect 17773 4981 17785 4984
rect 17819 5012 17831 5015
rect 18248 5012 18276 5040
rect 17819 4984 18276 5012
rect 17819 4981 17831 4984
rect 17773 4975 17831 4981
rect 18322 4972 18328 5024
rect 18380 5012 18386 5024
rect 19352 5012 19380 5052
rect 22186 5040 22192 5052
rect 22244 5040 22250 5092
rect 22388 5080 22416 5120
rect 22462 5108 22468 5160
rect 22520 5148 22526 5160
rect 22520 5120 22565 5148
rect 22520 5108 22526 5120
rect 22646 5108 22652 5160
rect 22704 5148 22710 5160
rect 23676 5157 23704 5188
rect 24118 5176 24124 5228
rect 24176 5216 24182 5228
rect 24489 5219 24547 5225
rect 24176 5188 24348 5216
rect 24176 5176 24182 5188
rect 23385 5151 23443 5157
rect 23385 5148 23397 5151
rect 22704 5120 23397 5148
rect 22704 5108 22710 5120
rect 23385 5117 23397 5120
rect 23431 5117 23443 5151
rect 23385 5111 23443 5117
rect 23661 5151 23719 5157
rect 23661 5117 23673 5151
rect 23707 5148 23719 5151
rect 24210 5148 24216 5160
rect 23707 5120 24216 5148
rect 23707 5117 23719 5120
rect 23661 5111 23719 5117
rect 24210 5108 24216 5120
rect 24268 5108 24274 5160
rect 24320 5148 24348 5188
rect 24489 5185 24501 5219
rect 24535 5216 24547 5219
rect 25038 5216 25044 5228
rect 24535 5188 24900 5216
rect 24999 5188 25044 5216
rect 24535 5185 24547 5188
rect 24489 5179 24547 5185
rect 24765 5151 24823 5157
rect 24765 5148 24777 5151
rect 24320 5120 24777 5148
rect 24765 5117 24777 5120
rect 24811 5117 24823 5151
rect 24872 5148 24900 5188
rect 25038 5176 25044 5188
rect 25096 5176 25102 5228
rect 25222 5176 25228 5228
rect 25280 5216 25286 5228
rect 25280 5188 26188 5216
rect 25280 5176 25286 5188
rect 25958 5148 25964 5160
rect 24872 5120 25964 5148
rect 24765 5111 24823 5117
rect 25958 5108 25964 5120
rect 26016 5108 26022 5160
rect 22388 5052 24808 5080
rect 18380 4984 19380 5012
rect 18380 4972 18386 4984
rect 19518 4972 19524 5024
rect 19576 5012 19582 5024
rect 19797 5015 19855 5021
rect 19797 5012 19809 5015
rect 19576 4984 19809 5012
rect 19576 4972 19582 4984
rect 19797 4981 19809 4984
rect 19843 4981 19855 5015
rect 19797 4975 19855 4981
rect 20257 5015 20315 5021
rect 20257 4981 20269 5015
rect 20303 5012 20315 5015
rect 20346 5012 20352 5024
rect 20303 4984 20352 5012
rect 20303 4981 20315 4984
rect 20257 4975 20315 4981
rect 20346 4972 20352 4984
rect 20404 4972 20410 5024
rect 20809 5015 20867 5021
rect 20809 4981 20821 5015
rect 20855 5012 20867 5015
rect 20898 5012 20904 5024
rect 20855 4984 20904 5012
rect 20855 4981 20867 4984
rect 20809 4975 20867 4981
rect 20898 4972 20904 4984
rect 20956 4972 20962 5024
rect 22278 5012 22284 5024
rect 22239 4984 22284 5012
rect 22278 4972 22284 4984
rect 22336 4972 22342 5024
rect 22554 4972 22560 5024
rect 22612 5012 22618 5024
rect 22649 5015 22707 5021
rect 22649 5012 22661 5015
rect 22612 4984 22661 5012
rect 22612 4972 22618 4984
rect 22649 4981 22661 4984
rect 22695 4981 22707 5015
rect 22649 4975 22707 4981
rect 23845 5015 23903 5021
rect 23845 4981 23857 5015
rect 23891 5012 23903 5015
rect 24029 5015 24087 5021
rect 24029 5012 24041 5015
rect 23891 4984 24041 5012
rect 23891 4981 23903 4984
rect 23845 4975 23903 4981
rect 24029 4981 24041 4984
rect 24075 5012 24087 5015
rect 24489 5015 24547 5021
rect 24489 5012 24501 5015
rect 24075 4984 24501 5012
rect 24075 4981 24087 4984
rect 24029 4975 24087 4981
rect 24489 4981 24501 4984
rect 24535 4981 24547 5015
rect 24780 5012 24808 5052
rect 26050 5012 26056 5024
rect 24780 4984 26056 5012
rect 24489 4975 24547 4981
rect 26050 4972 26056 4984
rect 26108 4972 26114 5024
rect 26160 5012 26188 5188
rect 26234 5176 26240 5228
rect 26292 5216 26298 5228
rect 26421 5219 26479 5225
rect 26421 5216 26433 5219
rect 26292 5188 26433 5216
rect 26292 5176 26298 5188
rect 26421 5185 26433 5188
rect 26467 5216 26479 5219
rect 26970 5216 26976 5228
rect 26467 5188 26976 5216
rect 26467 5185 26479 5188
rect 26421 5179 26479 5185
rect 26970 5176 26976 5188
rect 27028 5176 27034 5228
rect 27249 5219 27307 5225
rect 27249 5185 27261 5219
rect 27295 5216 27307 5219
rect 31846 5216 31852 5228
rect 27295 5188 31852 5216
rect 27295 5185 27307 5188
rect 27249 5179 27307 5185
rect 31846 5176 31852 5188
rect 31904 5176 31910 5228
rect 32122 5176 32128 5228
rect 32180 5216 32186 5228
rect 32180 5188 32720 5216
rect 32180 5176 32186 5188
rect 26694 5108 26700 5160
rect 26752 5148 26758 5160
rect 27801 5151 27859 5157
rect 27801 5148 27813 5151
rect 26752 5120 27813 5148
rect 26752 5108 26758 5120
rect 27801 5117 27813 5120
rect 27847 5148 27859 5151
rect 27890 5148 27896 5160
rect 27847 5120 27896 5148
rect 27847 5117 27859 5120
rect 27801 5111 27859 5117
rect 27890 5108 27896 5120
rect 27948 5108 27954 5160
rect 28074 5148 28080 5160
rect 28035 5120 28080 5148
rect 28074 5108 28080 5120
rect 28132 5108 28138 5160
rect 28258 5148 28264 5160
rect 28171 5120 28264 5148
rect 28258 5108 28264 5120
rect 28316 5108 28322 5160
rect 28350 5108 28356 5160
rect 28408 5148 28414 5160
rect 29273 5151 29331 5157
rect 29273 5148 29285 5151
rect 28408 5120 29285 5148
rect 28408 5108 28414 5120
rect 29273 5117 29285 5120
rect 29319 5117 29331 5151
rect 29822 5148 29828 5160
rect 29735 5120 29828 5148
rect 29273 5111 29331 5117
rect 29822 5108 29828 5120
rect 29880 5108 29886 5160
rect 29914 5108 29920 5160
rect 29972 5148 29978 5160
rect 30098 5148 30104 5160
rect 29972 5120 30017 5148
rect 30059 5120 30104 5148
rect 29972 5108 29978 5120
rect 30098 5108 30104 5120
rect 30156 5108 30162 5160
rect 30282 5148 30288 5160
rect 30243 5120 30288 5148
rect 30282 5108 30288 5120
rect 30340 5108 30346 5160
rect 30653 5151 30711 5157
rect 30653 5117 30665 5151
rect 30699 5148 30711 5151
rect 31386 5148 31392 5160
rect 30699 5120 31392 5148
rect 30699 5117 30711 5120
rect 30653 5111 30711 5117
rect 31386 5108 31392 5120
rect 31444 5108 31450 5160
rect 31573 5151 31631 5157
rect 31573 5117 31585 5151
rect 31619 5148 31631 5151
rect 32582 5148 32588 5160
rect 31619 5120 32588 5148
rect 31619 5117 31631 5120
rect 31573 5111 31631 5117
rect 27154 5040 27160 5092
rect 27212 5080 27218 5092
rect 28276 5080 28304 5108
rect 27212 5052 28304 5080
rect 27212 5040 27218 5052
rect 28994 5040 29000 5092
rect 29052 5080 29058 5092
rect 29840 5080 29868 5108
rect 30190 5080 30196 5092
rect 29052 5052 29097 5080
rect 29840 5052 30196 5080
rect 29052 5040 29058 5052
rect 30190 5040 30196 5052
rect 30248 5040 30254 5092
rect 31588 5080 31616 5111
rect 32582 5108 32588 5120
rect 32640 5108 32646 5160
rect 32692 5157 32720 5188
rect 33502 5176 33508 5228
rect 33560 5216 33566 5228
rect 37918 5216 37924 5228
rect 33560 5188 37924 5216
rect 33560 5176 33566 5188
rect 37918 5176 37924 5188
rect 37976 5216 37982 5228
rect 41138 5216 41144 5228
rect 37976 5188 41144 5216
rect 37976 5176 37982 5188
rect 32677 5151 32735 5157
rect 32677 5117 32689 5151
rect 32723 5148 32735 5151
rect 32953 5151 33011 5157
rect 32953 5148 32965 5151
rect 32723 5120 32965 5148
rect 32723 5117 32735 5120
rect 32677 5111 32735 5117
rect 32953 5117 32965 5120
rect 32999 5117 33011 5151
rect 32953 5111 33011 5117
rect 33226 5108 33232 5160
rect 33284 5148 33290 5160
rect 33689 5151 33747 5157
rect 33689 5148 33701 5151
rect 33284 5120 33701 5148
rect 33284 5108 33290 5120
rect 33689 5117 33701 5120
rect 33735 5148 33747 5151
rect 34238 5148 34244 5160
rect 33735 5120 34244 5148
rect 33735 5117 33747 5120
rect 33689 5111 33747 5117
rect 34238 5108 34244 5120
rect 34296 5108 34302 5160
rect 34425 5151 34483 5157
rect 34425 5117 34437 5151
rect 34471 5148 34483 5151
rect 34701 5151 34759 5157
rect 34701 5148 34713 5151
rect 34471 5120 34713 5148
rect 34471 5117 34483 5120
rect 34425 5111 34483 5117
rect 34701 5117 34713 5120
rect 34747 5148 34759 5151
rect 35069 5151 35127 5157
rect 35069 5148 35081 5151
rect 34747 5120 35081 5148
rect 34747 5117 34759 5120
rect 34701 5111 34759 5117
rect 35069 5117 35081 5120
rect 35115 5148 35127 5151
rect 36078 5148 36084 5160
rect 35115 5120 36084 5148
rect 35115 5117 35127 5120
rect 35069 5111 35127 5117
rect 36078 5108 36084 5120
rect 36136 5108 36142 5160
rect 36170 5108 36176 5160
rect 36228 5148 36234 5160
rect 36354 5148 36360 5160
rect 36228 5120 36273 5148
rect 36315 5120 36360 5148
rect 36228 5108 36234 5120
rect 36354 5108 36360 5120
rect 36412 5108 36418 5160
rect 38010 5148 38016 5160
rect 37971 5120 38016 5148
rect 38010 5108 38016 5120
rect 38068 5108 38074 5160
rect 38378 5148 38384 5160
rect 38339 5120 38384 5148
rect 38378 5108 38384 5120
rect 38436 5108 38442 5160
rect 38749 5151 38807 5157
rect 38749 5117 38761 5151
rect 38795 5148 38807 5151
rect 38795 5120 38884 5148
rect 38795 5117 38807 5120
rect 38749 5111 38807 5117
rect 30944 5052 31616 5080
rect 29730 5012 29736 5024
rect 26160 4984 29736 5012
rect 29730 4972 29736 4984
rect 29788 4972 29794 5024
rect 29914 4972 29920 5024
rect 29972 5012 29978 5024
rect 30944 5012 30972 5052
rect 31662 5040 31668 5092
rect 31720 5080 31726 5092
rect 32493 5083 32551 5089
rect 32493 5080 32505 5083
rect 31720 5052 32505 5080
rect 31720 5040 31726 5052
rect 32493 5049 32505 5052
rect 32539 5049 32551 5083
rect 34514 5080 34520 5092
rect 32493 5043 32551 5049
rect 32600 5052 34520 5080
rect 29972 4984 30972 5012
rect 29972 4972 29978 4984
rect 31018 4972 31024 5024
rect 31076 5012 31082 5024
rect 31205 5015 31263 5021
rect 31076 4984 31121 5012
rect 31076 4972 31082 4984
rect 31205 4981 31217 5015
rect 31251 5012 31263 5015
rect 31757 5015 31815 5021
rect 31757 5012 31769 5015
rect 31251 4984 31769 5012
rect 31251 4981 31263 4984
rect 31205 4975 31263 4981
rect 31757 4981 31769 4984
rect 31803 5012 31815 5015
rect 32600 5012 32628 5052
rect 34514 5040 34520 5052
rect 34572 5040 34578 5092
rect 36096 5080 36124 5108
rect 36538 5080 36544 5092
rect 36096 5052 36544 5080
rect 36538 5040 36544 5052
rect 36596 5040 36602 5092
rect 36725 5083 36783 5089
rect 36725 5049 36737 5083
rect 36771 5080 36783 5083
rect 37550 5080 37556 5092
rect 36771 5052 37556 5080
rect 36771 5049 36783 5052
rect 36725 5043 36783 5049
rect 37550 5040 37556 5052
rect 37608 5040 37614 5092
rect 31803 4984 32628 5012
rect 31803 4981 31815 4984
rect 31757 4975 31815 4981
rect 32674 4972 32680 5024
rect 32732 5012 32738 5024
rect 32769 5015 32827 5021
rect 32769 5012 32781 5015
rect 32732 4984 32781 5012
rect 32732 4972 32738 4984
rect 32769 4981 32781 4984
rect 32815 4981 32827 5015
rect 32769 4975 32827 4981
rect 32953 5015 33011 5021
rect 32953 4981 32965 5015
rect 32999 5012 33011 5015
rect 33229 5015 33287 5021
rect 33229 5012 33241 5015
rect 32999 4984 33241 5012
rect 32999 4981 33011 4984
rect 32953 4975 33011 4981
rect 33229 4981 33241 4984
rect 33275 5012 33287 5015
rect 33318 5012 33324 5024
rect 33275 4984 33324 5012
rect 33275 4981 33287 4984
rect 33229 4975 33287 4981
rect 33318 4972 33324 4984
rect 33376 4972 33382 5024
rect 33594 5012 33600 5024
rect 33507 4984 33600 5012
rect 33594 4972 33600 4984
rect 33652 5012 33658 5024
rect 33873 5015 33931 5021
rect 33873 5012 33885 5015
rect 33652 4984 33885 5012
rect 33652 4972 33658 4984
rect 33873 4981 33885 4984
rect 33919 5012 33931 5015
rect 35437 5015 35495 5021
rect 35437 5012 35449 5015
rect 33919 4984 35449 5012
rect 33919 4981 33931 4984
rect 33873 4975 33931 4981
rect 35437 4981 35449 4984
rect 35483 4981 35495 5015
rect 36998 5012 37004 5024
rect 36959 4984 37004 5012
rect 35437 4975 35495 4981
rect 36998 4972 37004 4984
rect 37056 4972 37062 5024
rect 37366 5012 37372 5024
rect 37327 4984 37372 5012
rect 37366 4972 37372 4984
rect 37424 4972 37430 5024
rect 37458 4972 37464 5024
rect 37516 5012 37522 5024
rect 38856 5012 38884 5120
rect 38930 5108 38936 5160
rect 38988 5148 38994 5160
rect 38988 5120 39033 5148
rect 38988 5108 38994 5120
rect 39298 5108 39304 5160
rect 39356 5148 39362 5160
rect 40494 5148 40500 5160
rect 39356 5120 40500 5148
rect 39356 5108 39362 5120
rect 40494 5108 40500 5120
rect 40552 5108 40558 5160
rect 40604 5157 40632 5188
rect 41138 5176 41144 5188
rect 41196 5176 41202 5228
rect 41417 5219 41475 5225
rect 41417 5185 41429 5219
rect 41463 5216 41475 5219
rect 44082 5216 44088 5228
rect 41463 5188 44088 5216
rect 41463 5185 41475 5188
rect 41417 5179 41475 5185
rect 44082 5176 44088 5188
rect 44140 5176 44146 5228
rect 40589 5151 40647 5157
rect 40589 5117 40601 5151
rect 40635 5117 40647 5151
rect 41966 5148 41972 5160
rect 41927 5120 41972 5148
rect 40589 5111 40647 5117
rect 41966 5108 41972 5120
rect 42024 5108 42030 5160
rect 42429 5151 42487 5157
rect 42429 5117 42441 5151
rect 42475 5148 42487 5151
rect 42886 5148 42892 5160
rect 42475 5120 42892 5148
rect 42475 5117 42487 5120
rect 42429 5111 42487 5117
rect 42886 5108 42892 5120
rect 42944 5108 42950 5160
rect 43349 5151 43407 5157
rect 43349 5117 43361 5151
rect 43395 5148 43407 5151
rect 43622 5148 43628 5160
rect 43395 5120 43628 5148
rect 43395 5117 43407 5120
rect 43349 5111 43407 5117
rect 43622 5108 43628 5120
rect 43680 5108 43686 5160
rect 44468 5157 44496 5256
rect 46106 5244 46112 5256
rect 46164 5244 46170 5296
rect 44818 5176 44824 5228
rect 44876 5216 44882 5228
rect 45557 5219 45615 5225
rect 45557 5216 45569 5219
rect 44876 5188 45569 5216
rect 44876 5176 44882 5188
rect 45557 5185 45569 5188
rect 45603 5216 45615 5219
rect 46216 5216 46244 5324
rect 48866 5312 48872 5324
rect 48924 5312 48930 5364
rect 48961 5355 49019 5361
rect 48961 5321 48973 5355
rect 49007 5352 49019 5355
rect 50246 5352 50252 5364
rect 49007 5324 50252 5352
rect 49007 5321 49019 5324
rect 48961 5315 49019 5321
rect 50246 5312 50252 5324
rect 50304 5312 50310 5364
rect 50430 5312 50436 5364
rect 50488 5352 50494 5364
rect 51261 5355 51319 5361
rect 51261 5352 51273 5355
rect 50488 5324 51273 5352
rect 50488 5312 50494 5324
rect 51261 5321 51273 5324
rect 51307 5321 51319 5355
rect 51261 5315 51319 5321
rect 51810 5312 51816 5364
rect 51868 5352 51874 5364
rect 52365 5355 52423 5361
rect 52365 5352 52377 5355
rect 51868 5324 52377 5352
rect 51868 5312 51874 5324
rect 52365 5321 52377 5324
rect 52411 5321 52423 5355
rect 52365 5315 52423 5321
rect 52564 5324 53512 5352
rect 46290 5244 46296 5296
rect 46348 5284 46354 5296
rect 46348 5256 46393 5284
rect 46348 5244 46354 5256
rect 47118 5244 47124 5296
rect 47176 5284 47182 5296
rect 52564 5284 52592 5324
rect 53374 5284 53380 5296
rect 47176 5256 52592 5284
rect 53335 5256 53380 5284
rect 47176 5244 47182 5256
rect 53374 5244 53380 5256
rect 53432 5244 53438 5296
rect 53484 5284 53512 5324
rect 53834 5312 53840 5364
rect 53892 5352 53898 5364
rect 54297 5355 54355 5361
rect 54297 5352 54309 5355
rect 53892 5324 54309 5352
rect 53892 5312 53898 5324
rect 54297 5321 54309 5324
rect 54343 5321 54355 5355
rect 54297 5315 54355 5321
rect 55214 5312 55220 5364
rect 55272 5352 55278 5364
rect 55766 5352 55772 5364
rect 55272 5324 55772 5352
rect 55272 5312 55278 5324
rect 55766 5312 55772 5324
rect 55824 5312 55830 5364
rect 55953 5355 56011 5361
rect 55953 5321 55965 5355
rect 55999 5352 56011 5355
rect 56042 5352 56048 5364
rect 55999 5324 56048 5352
rect 55999 5321 56011 5324
rect 55953 5315 56011 5321
rect 56042 5312 56048 5324
rect 56100 5312 56106 5364
rect 58894 5352 58900 5364
rect 58855 5324 58900 5352
rect 58894 5312 58900 5324
rect 58952 5312 58958 5364
rect 61286 5312 61292 5364
rect 61344 5352 61350 5364
rect 61473 5355 61531 5361
rect 61473 5352 61485 5355
rect 61344 5324 61485 5352
rect 61344 5312 61350 5324
rect 61473 5321 61485 5324
rect 61519 5321 61531 5355
rect 61473 5315 61531 5321
rect 54018 5284 54024 5296
rect 53484 5256 54024 5284
rect 54018 5244 54024 5256
rect 54076 5244 54082 5296
rect 55600 5256 59400 5284
rect 45603 5188 46244 5216
rect 45603 5185 45615 5188
rect 45557 5179 45615 5185
rect 44453 5151 44511 5157
rect 44453 5148 44465 5151
rect 43732 5120 44465 5148
rect 39022 5040 39028 5092
rect 39080 5080 39086 5092
rect 43732 5080 43760 5120
rect 44453 5117 44465 5120
rect 44499 5117 44511 5151
rect 44453 5111 44511 5117
rect 44542 5108 44548 5160
rect 44600 5148 44606 5160
rect 44729 5151 44787 5157
rect 44729 5148 44741 5151
rect 44600 5120 44741 5148
rect 44600 5108 44606 5120
rect 44729 5117 44741 5120
rect 44775 5148 44787 5151
rect 45002 5148 45008 5160
rect 44775 5120 45008 5148
rect 44775 5117 44787 5120
rect 44729 5111 44787 5117
rect 45002 5108 45008 5120
rect 45060 5108 45066 5160
rect 46308 5148 46336 5244
rect 48130 5176 48136 5228
rect 48188 5216 48194 5228
rect 49145 5219 49203 5225
rect 49145 5216 49157 5219
rect 48188 5188 49157 5216
rect 48188 5176 48194 5188
rect 49145 5185 49157 5188
rect 49191 5185 49203 5219
rect 49145 5179 49203 5185
rect 49510 5176 49516 5228
rect 49568 5216 49574 5228
rect 49605 5219 49663 5225
rect 49605 5216 49617 5219
rect 49568 5188 49617 5216
rect 49568 5176 49574 5188
rect 49605 5185 49617 5188
rect 49651 5185 49663 5219
rect 50525 5219 50583 5225
rect 50525 5216 50537 5219
rect 49605 5179 49663 5185
rect 49712 5188 50537 5216
rect 49712 5160 49740 5188
rect 50525 5185 50537 5188
rect 50571 5185 50583 5219
rect 50525 5179 50583 5185
rect 50614 5176 50620 5228
rect 50672 5216 50678 5228
rect 52730 5216 52736 5228
rect 50672 5188 52736 5216
rect 50672 5176 50678 5188
rect 52730 5176 52736 5188
rect 52788 5176 52794 5228
rect 52932 5188 55444 5216
rect 46477 5151 46535 5157
rect 46477 5148 46489 5151
rect 46308 5120 46489 5148
rect 46477 5117 46489 5120
rect 46523 5117 46535 5151
rect 46477 5111 46535 5117
rect 47213 5151 47271 5157
rect 47213 5117 47225 5151
rect 47259 5117 47271 5151
rect 47213 5111 47271 5117
rect 47489 5151 47547 5157
rect 47489 5117 47501 5151
rect 47535 5148 47547 5151
rect 47854 5148 47860 5160
rect 47535 5120 47860 5148
rect 47535 5117 47547 5120
rect 47489 5111 47547 5117
rect 39080 5052 43760 5080
rect 39080 5040 39086 5052
rect 43806 5040 43812 5092
rect 43864 5080 43870 5092
rect 44637 5083 44695 5089
rect 44637 5080 44649 5083
rect 43864 5052 44649 5080
rect 43864 5040 43870 5052
rect 44637 5049 44649 5052
rect 44683 5049 44695 5083
rect 47228 5080 47256 5111
rect 47854 5108 47860 5120
rect 47912 5148 47918 5160
rect 48225 5151 48283 5157
rect 48225 5148 48237 5151
rect 47912 5120 48237 5148
rect 47912 5108 47918 5120
rect 48225 5117 48237 5120
rect 48271 5117 48283 5151
rect 49326 5148 49332 5160
rect 49287 5120 49332 5148
rect 48225 5111 48283 5117
rect 49326 5108 49332 5120
rect 49384 5108 49390 5160
rect 49694 5148 49700 5160
rect 49655 5120 49700 5148
rect 49694 5108 49700 5120
rect 49752 5108 49758 5160
rect 50890 5148 50896 5160
rect 50851 5120 50896 5148
rect 50890 5108 50896 5120
rect 50948 5108 50954 5160
rect 52638 5148 52644 5160
rect 52599 5120 52644 5148
rect 52638 5108 52644 5120
rect 52696 5108 52702 5160
rect 52822 5108 52828 5160
rect 52880 5148 52886 5160
rect 52932 5157 52960 5188
rect 55416 5160 55444 5188
rect 52917 5151 52975 5157
rect 52917 5148 52929 5151
rect 52880 5120 52929 5148
rect 52880 5108 52886 5120
rect 52917 5117 52929 5120
rect 52963 5117 52975 5151
rect 52917 5111 52975 5117
rect 53377 5151 53435 5157
rect 53377 5117 53389 5151
rect 53423 5148 53435 5151
rect 53929 5151 53987 5157
rect 53929 5148 53941 5151
rect 53423 5120 53941 5148
rect 53423 5117 53435 5120
rect 53377 5111 53435 5117
rect 53929 5117 53941 5120
rect 53975 5148 53987 5151
rect 54662 5148 54668 5160
rect 53975 5120 54668 5148
rect 53975 5117 53987 5120
rect 53929 5111 53987 5117
rect 47946 5080 47952 5092
rect 44637 5043 44695 5049
rect 44744 5052 46704 5080
rect 47228 5052 47952 5080
rect 39206 5012 39212 5024
rect 37516 4984 39212 5012
rect 37516 4972 37522 4984
rect 39206 4972 39212 4984
rect 39264 4972 39270 5024
rect 39393 5015 39451 5021
rect 39393 4981 39405 5015
rect 39439 5012 39451 5015
rect 40218 5012 40224 5024
rect 39439 4984 40224 5012
rect 39439 4981 39451 4984
rect 39393 4975 39451 4981
rect 40218 4972 40224 4984
rect 40276 4972 40282 5024
rect 40862 4972 40868 5024
rect 40920 5012 40926 5024
rect 41601 5015 41659 5021
rect 41601 5012 41613 5015
rect 40920 4984 41613 5012
rect 40920 4972 40926 4984
rect 41601 4981 41613 4984
rect 41647 5012 41659 5015
rect 41966 5012 41972 5024
rect 41647 4984 41972 5012
rect 41647 4981 41659 4984
rect 41601 4975 41659 4981
rect 41966 4972 41972 4984
rect 42024 5012 42030 5024
rect 44744 5012 44772 5052
rect 46566 5012 46572 5024
rect 42024 4984 44772 5012
rect 46527 4984 46572 5012
rect 42024 4972 42030 4984
rect 46566 4972 46572 4984
rect 46624 4972 46630 5024
rect 46676 5012 46704 5052
rect 47946 5040 47952 5052
rect 48004 5040 48010 5092
rect 49344 5080 49372 5108
rect 53392 5080 53420 5111
rect 54662 5108 54668 5120
rect 54720 5108 54726 5160
rect 55125 5151 55183 5157
rect 55125 5117 55137 5151
rect 55171 5148 55183 5151
rect 55214 5148 55220 5160
rect 55171 5120 55220 5148
rect 55171 5117 55183 5120
rect 55125 5111 55183 5117
rect 55214 5108 55220 5120
rect 55272 5108 55278 5160
rect 55398 5148 55404 5160
rect 55311 5120 55404 5148
rect 55398 5108 55404 5120
rect 55456 5108 55462 5160
rect 55490 5108 55496 5160
rect 55548 5148 55554 5160
rect 55600 5157 55628 5256
rect 56410 5176 56416 5228
rect 56468 5216 56474 5228
rect 57974 5216 57980 5228
rect 56468 5188 57652 5216
rect 57935 5188 57980 5216
rect 56468 5176 56474 5188
rect 55585 5151 55643 5157
rect 55585 5148 55597 5151
rect 55548 5120 55597 5148
rect 55548 5108 55554 5120
rect 55585 5117 55597 5120
rect 55631 5117 55643 5151
rect 55585 5111 55643 5117
rect 56781 5151 56839 5157
rect 56781 5117 56793 5151
rect 56827 5148 56839 5151
rect 57146 5148 57152 5160
rect 56827 5120 57152 5148
rect 56827 5117 56839 5120
rect 56781 5111 56839 5117
rect 54570 5080 54576 5092
rect 49344 5052 53420 5080
rect 54531 5052 54576 5080
rect 54570 5040 54576 5052
rect 54628 5040 54634 5092
rect 47857 5015 47915 5021
rect 47857 5012 47869 5015
rect 46676 4984 47869 5012
rect 47857 4981 47869 4984
rect 47903 5012 47915 5015
rect 48038 5012 48044 5024
rect 47903 4984 48044 5012
rect 47903 4981 47915 4984
rect 47857 4975 47915 4981
rect 48038 4972 48044 4984
rect 48096 4972 48102 5024
rect 49510 4972 49516 5024
rect 49568 5012 49574 5024
rect 50157 5015 50215 5021
rect 50157 5012 50169 5015
rect 49568 4984 50169 5012
rect 49568 4972 49574 4984
rect 50157 4981 50169 4984
rect 50203 4981 50215 5015
rect 50157 4975 50215 4981
rect 51534 4972 51540 5024
rect 51592 5012 51598 5024
rect 51905 5015 51963 5021
rect 51905 5012 51917 5015
rect 51592 4984 51917 5012
rect 51592 4972 51598 4984
rect 51905 4981 51917 4984
rect 51951 4981 51963 5015
rect 51905 4975 51963 4981
rect 52546 4972 52552 5024
rect 52604 5012 52610 5024
rect 55600 5012 55628 5111
rect 57146 5108 57152 5120
rect 57204 5148 57210 5160
rect 57624 5157 57652 5188
rect 57974 5176 57980 5188
rect 58032 5176 58038 5228
rect 57333 5151 57391 5157
rect 57333 5148 57345 5151
rect 57204 5120 57345 5148
rect 57204 5108 57210 5120
rect 57333 5117 57345 5120
rect 57379 5117 57391 5151
rect 57333 5111 57391 5117
rect 57425 5151 57483 5157
rect 57425 5117 57437 5151
rect 57471 5117 57483 5151
rect 57425 5111 57483 5117
rect 57609 5151 57667 5157
rect 57609 5117 57621 5151
rect 57655 5148 57667 5151
rect 58345 5151 58403 5157
rect 58345 5148 58357 5151
rect 57655 5120 58357 5148
rect 57655 5117 57667 5120
rect 57609 5111 57667 5117
rect 58345 5117 58357 5120
rect 58391 5148 58403 5151
rect 58618 5148 58624 5160
rect 58391 5120 58624 5148
rect 58391 5117 58403 5120
rect 58345 5111 58403 5117
rect 57440 5080 57468 5111
rect 58618 5108 58624 5120
rect 58676 5108 58682 5160
rect 59078 5148 59084 5160
rect 59039 5120 59084 5148
rect 59078 5108 59084 5120
rect 59136 5108 59142 5160
rect 59262 5148 59268 5160
rect 59223 5120 59268 5148
rect 59262 5108 59268 5120
rect 59320 5108 59326 5160
rect 59372 5148 59400 5256
rect 59722 5148 59728 5160
rect 59372 5120 59728 5148
rect 59722 5108 59728 5120
rect 59780 5108 59786 5160
rect 59814 5108 59820 5160
rect 59872 5148 59878 5160
rect 61010 5148 61016 5160
rect 59872 5120 61016 5148
rect 59872 5108 59878 5120
rect 61010 5108 61016 5120
rect 61068 5108 61074 5160
rect 57072 5052 57468 5080
rect 59740 5080 59768 5108
rect 61194 5080 61200 5092
rect 59740 5052 61200 5080
rect 57072 5024 57100 5052
rect 61194 5040 61200 5052
rect 61252 5040 61258 5092
rect 52604 4984 55628 5012
rect 56321 5015 56379 5021
rect 52604 4972 52610 4984
rect 56321 4981 56333 5015
rect 56367 5012 56379 5015
rect 56502 5012 56508 5024
rect 56367 4984 56508 5012
rect 56367 4981 56379 4984
rect 56321 4975 56379 4981
rect 56502 4972 56508 4984
rect 56560 4972 56566 5024
rect 57054 5012 57060 5024
rect 57015 4984 57060 5012
rect 57054 4972 57060 4984
rect 57112 4972 57118 5024
rect 59998 4972 60004 5024
rect 60056 5012 60062 5024
rect 60277 5015 60335 5021
rect 60277 5012 60289 5015
rect 60056 4984 60289 5012
rect 60056 4972 60062 4984
rect 60277 4981 60289 4984
rect 60323 4981 60335 5015
rect 60277 4975 60335 4981
rect 60458 4972 60464 5024
rect 60516 5012 60522 5024
rect 60737 5015 60795 5021
rect 60737 5012 60749 5015
rect 60516 4984 60749 5012
rect 60516 4972 60522 4984
rect 60737 4981 60749 4984
rect 60783 4981 60795 5015
rect 60737 4975 60795 4981
rect 61010 4972 61016 5024
rect 61068 5012 61074 5024
rect 61105 5015 61163 5021
rect 61105 5012 61117 5015
rect 61068 4984 61117 5012
rect 61068 4972 61074 4984
rect 61105 4981 61117 4984
rect 61151 4981 61163 5015
rect 61105 4975 61163 4981
rect 1104 4922 63480 4944
rect 1104 4870 21774 4922
rect 21826 4870 21838 4922
rect 21890 4870 21902 4922
rect 21954 4870 21966 4922
rect 22018 4870 42566 4922
rect 42618 4870 42630 4922
rect 42682 4870 42694 4922
rect 42746 4870 42758 4922
rect 42810 4870 63480 4922
rect 1104 4848 63480 4870
rect 6457 4811 6515 4817
rect 6457 4808 6469 4811
rect 2608 4780 6469 4808
rect 2498 4700 2504 4752
rect 2556 4740 2562 4752
rect 2608 4749 2636 4780
rect 6457 4777 6469 4780
rect 6503 4777 6515 4811
rect 6457 4771 6515 4777
rect 7653 4811 7711 4817
rect 7653 4777 7665 4811
rect 7699 4808 7711 4811
rect 8297 4811 8355 4817
rect 8297 4808 8309 4811
rect 7699 4780 8309 4808
rect 7699 4777 7711 4780
rect 7653 4771 7711 4777
rect 8297 4777 8309 4780
rect 8343 4808 8355 4811
rect 12158 4808 12164 4820
rect 8343 4780 12164 4808
rect 8343 4777 8355 4780
rect 8297 4771 8355 4777
rect 12158 4768 12164 4780
rect 12216 4768 12222 4820
rect 14918 4808 14924 4820
rect 14879 4780 14924 4808
rect 14918 4768 14924 4780
rect 14976 4768 14982 4820
rect 15562 4768 15568 4820
rect 15620 4808 15626 4820
rect 15933 4811 15991 4817
rect 15933 4808 15945 4811
rect 15620 4780 15945 4808
rect 15620 4768 15626 4780
rect 15933 4777 15945 4780
rect 15979 4808 15991 4811
rect 17218 4808 17224 4820
rect 15979 4780 17224 4808
rect 15979 4777 15991 4780
rect 15933 4771 15991 4777
rect 17218 4768 17224 4780
rect 17276 4768 17282 4820
rect 17770 4768 17776 4820
rect 17828 4808 17834 4820
rect 17865 4811 17923 4817
rect 17865 4808 17877 4811
rect 17828 4780 17877 4808
rect 17828 4768 17834 4780
rect 17865 4777 17877 4780
rect 17911 4777 17923 4811
rect 17865 4771 17923 4777
rect 18046 4768 18052 4820
rect 18104 4808 18110 4820
rect 19429 4811 19487 4817
rect 19429 4808 19441 4811
rect 18104 4780 19441 4808
rect 18104 4768 18110 4780
rect 19429 4777 19441 4780
rect 19475 4777 19487 4811
rect 19429 4771 19487 4777
rect 19613 4811 19671 4817
rect 19613 4777 19625 4811
rect 19659 4808 19671 4811
rect 21542 4808 21548 4820
rect 19659 4780 21548 4808
rect 19659 4777 19671 4780
rect 19613 4771 19671 4777
rect 21542 4768 21548 4780
rect 21600 4768 21606 4820
rect 23934 4808 23940 4820
rect 22112 4780 23940 4808
rect 2593 4743 2651 4749
rect 2593 4740 2605 4743
rect 2556 4712 2605 4740
rect 2556 4700 2562 4712
rect 2593 4709 2605 4712
rect 2639 4709 2651 4743
rect 4062 4740 4068 4752
rect 4023 4712 4068 4740
rect 2593 4703 2651 4709
rect 4062 4700 4068 4712
rect 4120 4700 4126 4752
rect 8481 4743 8539 4749
rect 8481 4740 8493 4743
rect 7024 4712 8493 4740
rect 2777 4675 2835 4681
rect 2777 4641 2789 4675
rect 2823 4672 2835 4675
rect 2866 4672 2872 4684
rect 2823 4644 2872 4672
rect 2823 4641 2835 4644
rect 2777 4635 2835 4641
rect 2866 4632 2872 4644
rect 2924 4632 2930 4684
rect 4522 4672 4528 4684
rect 4483 4644 4528 4672
rect 4522 4632 4528 4644
rect 4580 4632 4586 4684
rect 4709 4675 4767 4681
rect 4709 4641 4721 4675
rect 4755 4641 4767 4675
rect 4709 4635 4767 4641
rect 4893 4675 4951 4681
rect 4893 4641 4905 4675
rect 4939 4672 4951 4675
rect 5166 4672 5172 4684
rect 4939 4644 5172 4672
rect 4939 4641 4951 4644
rect 4893 4635 4951 4641
rect 3145 4607 3203 4613
rect 3145 4573 3157 4607
rect 3191 4604 3203 4607
rect 4724 4604 4752 4635
rect 5166 4632 5172 4644
rect 5224 4672 5230 4684
rect 7024 4681 7052 4712
rect 8481 4709 8493 4712
rect 8527 4740 8539 4743
rect 8754 4740 8760 4752
rect 8527 4712 8760 4740
rect 8527 4709 8539 4712
rect 8481 4703 8539 4709
rect 8754 4700 8760 4712
rect 8812 4700 8818 4752
rect 8846 4700 8852 4752
rect 8904 4740 8910 4752
rect 10781 4743 10839 4749
rect 10781 4740 10793 4743
rect 8904 4712 10793 4740
rect 8904 4700 8910 4712
rect 10781 4709 10793 4712
rect 10827 4709 10839 4743
rect 10781 4703 10839 4709
rect 10980 4712 12020 4740
rect 5353 4675 5411 4681
rect 5353 4672 5365 4675
rect 5224 4644 5365 4672
rect 5224 4632 5230 4644
rect 5353 4641 5365 4644
rect 5399 4641 5411 4675
rect 5353 4635 5411 4641
rect 7009 4675 7067 4681
rect 7009 4641 7021 4675
rect 7055 4641 7067 4675
rect 7009 4635 7067 4641
rect 7377 4675 7435 4681
rect 7377 4641 7389 4675
rect 7423 4672 7435 4675
rect 7653 4675 7711 4681
rect 7653 4672 7665 4675
rect 7423 4644 7665 4672
rect 7423 4641 7435 4644
rect 7377 4635 7435 4641
rect 7653 4641 7665 4644
rect 7699 4641 7711 4675
rect 7653 4635 7711 4641
rect 7834 4632 7840 4684
rect 7892 4672 7898 4684
rect 8389 4675 8447 4681
rect 8389 4672 8401 4675
rect 7892 4644 8401 4672
rect 7892 4632 7898 4644
rect 8389 4641 8401 4644
rect 8435 4672 8447 4675
rect 8662 4672 8668 4684
rect 8435 4644 8668 4672
rect 8435 4641 8447 4644
rect 8389 4635 8447 4641
rect 8662 4632 8668 4644
rect 8720 4632 8726 4684
rect 9674 4672 9680 4684
rect 8772 4644 9680 4672
rect 4798 4604 4804 4616
rect 3191 4576 4804 4604
rect 3191 4573 3203 4576
rect 3145 4567 3203 4573
rect 4798 4564 4804 4576
rect 4856 4564 4862 4616
rect 7101 4607 7159 4613
rect 7101 4573 7113 4607
rect 7147 4573 7159 4607
rect 7282 4604 7288 4616
rect 7195 4576 7288 4604
rect 7101 4567 7159 4573
rect 7116 4536 7144 4567
rect 7282 4564 7288 4576
rect 7340 4604 7346 4616
rect 8772 4604 8800 4644
rect 9674 4632 9680 4644
rect 9732 4632 9738 4684
rect 9766 4632 9772 4684
rect 9824 4672 9830 4684
rect 9861 4675 9919 4681
rect 9861 4672 9873 4675
rect 9824 4644 9873 4672
rect 9824 4632 9830 4644
rect 9861 4641 9873 4644
rect 9907 4641 9919 4675
rect 9861 4635 9919 4641
rect 10045 4675 10103 4681
rect 10045 4641 10057 4675
rect 10091 4672 10103 4675
rect 10134 4672 10140 4684
rect 10091 4644 10140 4672
rect 10091 4641 10103 4644
rect 10045 4635 10103 4641
rect 10134 4632 10140 4644
rect 10192 4632 10198 4684
rect 7340 4576 8800 4604
rect 7340 4564 7346 4576
rect 8846 4564 8852 4616
rect 8904 4564 8910 4616
rect 8941 4607 8999 4613
rect 8941 4573 8953 4607
rect 8987 4604 8999 4607
rect 9493 4607 9551 4613
rect 9493 4604 9505 4607
rect 8987 4576 9505 4604
rect 8987 4573 8999 4576
rect 8941 4567 8999 4573
rect 9493 4573 9505 4576
rect 9539 4604 9551 4607
rect 9582 4604 9588 4616
rect 9539 4576 9588 4604
rect 9539 4573 9551 4576
rect 9493 4567 9551 4573
rect 9582 4564 9588 4576
rect 9640 4604 9646 4616
rect 10413 4607 10471 4613
rect 10413 4604 10425 4607
rect 9640 4576 10425 4604
rect 9640 4564 9646 4576
rect 10413 4573 10425 4576
rect 10459 4604 10471 4607
rect 10980 4604 11008 4712
rect 11609 4675 11667 4681
rect 11609 4641 11621 4675
rect 11655 4672 11667 4675
rect 11698 4672 11704 4684
rect 11655 4644 11704 4672
rect 11655 4641 11667 4644
rect 11609 4635 11667 4641
rect 11698 4632 11704 4644
rect 11756 4632 11762 4684
rect 11793 4675 11851 4681
rect 11793 4641 11805 4675
rect 11839 4672 11851 4675
rect 11882 4672 11888 4684
rect 11839 4644 11888 4672
rect 11839 4641 11851 4644
rect 11793 4635 11851 4641
rect 11882 4632 11888 4644
rect 11940 4632 11946 4684
rect 11992 4672 12020 4712
rect 12066 4700 12072 4752
rect 12124 4740 12130 4752
rect 22112 4740 22140 4780
rect 23934 4768 23940 4780
rect 23992 4768 23998 4820
rect 24029 4811 24087 4817
rect 24029 4777 24041 4811
rect 24075 4808 24087 4811
rect 24210 4808 24216 4820
rect 24075 4780 24216 4808
rect 24075 4777 24087 4780
rect 24029 4771 24087 4777
rect 24210 4768 24216 4780
rect 24268 4768 24274 4820
rect 24394 4808 24400 4820
rect 24355 4780 24400 4808
rect 24394 4768 24400 4780
rect 24452 4768 24458 4820
rect 24854 4808 24860 4820
rect 24815 4780 24860 4808
rect 24854 4768 24860 4780
rect 24912 4768 24918 4820
rect 26050 4768 26056 4820
rect 26108 4808 26114 4820
rect 38841 4811 38899 4817
rect 38841 4808 38853 4811
rect 26108 4780 38853 4808
rect 26108 4768 26114 4780
rect 38841 4777 38853 4780
rect 38887 4777 38899 4811
rect 38841 4771 38899 4777
rect 38933 4811 38991 4817
rect 38933 4777 38945 4811
rect 38979 4808 38991 4811
rect 38979 4780 39712 4808
rect 38979 4777 38991 4780
rect 38933 4771 38991 4777
rect 12124 4712 22140 4740
rect 12124 4700 12130 4712
rect 22186 4700 22192 4752
rect 22244 4740 22250 4752
rect 29822 4740 29828 4752
rect 22244 4712 29828 4740
rect 22244 4700 22250 4712
rect 29822 4700 29828 4712
rect 29880 4700 29886 4752
rect 30466 4740 30472 4752
rect 29932 4712 30472 4740
rect 12805 4675 12863 4681
rect 12805 4672 12817 4675
rect 11992 4644 12817 4672
rect 12805 4641 12817 4644
rect 12851 4641 12863 4675
rect 12805 4635 12863 4641
rect 13265 4675 13323 4681
rect 13265 4641 13277 4675
rect 13311 4641 13323 4675
rect 13265 4635 13323 4641
rect 13725 4675 13783 4681
rect 13725 4641 13737 4675
rect 13771 4672 13783 4675
rect 13906 4672 13912 4684
rect 13771 4644 13912 4672
rect 13771 4641 13783 4644
rect 13725 4635 13783 4641
rect 10459 4576 11008 4604
rect 10459 4573 10471 4576
rect 10413 4567 10471 4573
rect 11054 4564 11060 4616
rect 11112 4604 11118 4616
rect 13280 4604 13308 4635
rect 13906 4632 13912 4644
rect 13964 4672 13970 4684
rect 13964 4644 14228 4672
rect 13964 4632 13970 4644
rect 14001 4607 14059 4613
rect 14001 4604 14013 4607
rect 11112 4576 13216 4604
rect 13280 4576 14013 4604
rect 11112 4564 11118 4576
rect 8864 4536 8892 4564
rect 7116 4508 8892 4536
rect 10210 4539 10268 4545
rect 10210 4505 10222 4539
rect 10256 4536 10268 4539
rect 10778 4536 10784 4548
rect 10256 4508 10784 4536
rect 10256 4505 10268 4508
rect 10210 4499 10268 4505
rect 10778 4496 10784 4508
rect 10836 4496 10842 4548
rect 13078 4536 13084 4548
rect 13039 4508 13084 4536
rect 13078 4496 13084 4508
rect 13136 4496 13142 4548
rect 13188 4536 13216 4576
rect 14001 4573 14013 4576
rect 14047 4604 14059 4607
rect 14090 4604 14096 4616
rect 14047 4576 14096 4604
rect 14047 4573 14059 4576
rect 14001 4567 14059 4573
rect 14090 4564 14096 4576
rect 14148 4564 14154 4616
rect 14200 4604 14228 4644
rect 14734 4632 14740 4684
rect 14792 4672 14798 4684
rect 15289 4675 15347 4681
rect 15289 4672 15301 4675
rect 14792 4644 15301 4672
rect 14792 4632 14798 4644
rect 15289 4641 15301 4644
rect 15335 4672 15347 4675
rect 16574 4672 16580 4684
rect 15335 4644 16344 4672
rect 16535 4644 16580 4672
rect 15335 4641 15347 4644
rect 15289 4635 15347 4641
rect 16206 4604 16212 4616
rect 14200 4576 16212 4604
rect 16206 4564 16212 4576
rect 16264 4564 16270 4616
rect 16316 4604 16344 4644
rect 16574 4632 16580 4644
rect 16632 4632 16638 4684
rect 16666 4632 16672 4684
rect 16724 4672 16730 4684
rect 17037 4675 17095 4681
rect 17037 4672 17049 4675
rect 16724 4644 17049 4672
rect 16724 4632 16730 4644
rect 17037 4641 17049 4644
rect 17083 4641 17095 4675
rect 17037 4635 17095 4641
rect 17144 4644 17632 4672
rect 17144 4604 17172 4644
rect 16316 4576 17172 4604
rect 17402 4564 17408 4616
rect 17460 4604 17466 4616
rect 17604 4604 17632 4644
rect 18138 4632 18144 4684
rect 18196 4672 18202 4684
rect 18233 4675 18291 4681
rect 18233 4672 18245 4675
rect 18196 4644 18245 4672
rect 18196 4632 18202 4644
rect 18233 4641 18245 4644
rect 18279 4672 18291 4675
rect 18417 4675 18475 4681
rect 18417 4672 18429 4675
rect 18279 4644 18429 4672
rect 18279 4641 18291 4644
rect 18233 4635 18291 4641
rect 18417 4641 18429 4644
rect 18463 4641 18475 4675
rect 18598 4672 18604 4684
rect 18559 4644 18604 4672
rect 18417 4635 18475 4641
rect 18598 4632 18604 4644
rect 18656 4632 18662 4684
rect 18693 4675 18751 4681
rect 18693 4641 18705 4675
rect 18739 4672 18751 4675
rect 19334 4672 19340 4684
rect 18739 4644 19340 4672
rect 18739 4641 18751 4644
rect 18693 4635 18751 4641
rect 19334 4632 19340 4644
rect 19392 4672 19398 4684
rect 19978 4672 19984 4684
rect 19392 4644 19984 4672
rect 19392 4632 19398 4644
rect 19978 4632 19984 4644
rect 20036 4632 20042 4684
rect 20898 4672 20904 4684
rect 20859 4644 20904 4672
rect 20898 4632 20904 4644
rect 20956 4632 20962 4684
rect 21174 4672 21180 4684
rect 21135 4644 21180 4672
rect 21174 4632 21180 4644
rect 21232 4632 21238 4684
rect 22373 4675 22431 4681
rect 22373 4641 22385 4675
rect 22419 4672 22431 4675
rect 22465 4675 22523 4681
rect 22465 4672 22477 4675
rect 22419 4644 22477 4672
rect 22419 4641 22431 4644
rect 22373 4635 22431 4641
rect 22465 4641 22477 4644
rect 22511 4641 22523 4675
rect 22465 4635 22523 4641
rect 22649 4675 22707 4681
rect 22649 4641 22661 4675
rect 22695 4672 22707 4675
rect 22922 4672 22928 4684
rect 22695 4644 22928 4672
rect 22695 4641 22707 4644
rect 22649 4635 22707 4641
rect 22922 4632 22928 4644
rect 22980 4632 22986 4684
rect 23842 4672 23848 4684
rect 23803 4644 23848 4672
rect 23842 4632 23848 4644
rect 23900 4632 23906 4684
rect 24486 4632 24492 4684
rect 24544 4672 24550 4684
rect 25130 4672 25136 4684
rect 24544 4644 25136 4672
rect 24544 4632 24550 4644
rect 25130 4632 25136 4644
rect 25188 4632 25194 4684
rect 25314 4672 25320 4684
rect 25275 4644 25320 4672
rect 25314 4632 25320 4644
rect 25372 4672 25378 4684
rect 25869 4675 25927 4681
rect 25869 4672 25881 4675
rect 25372 4644 25881 4672
rect 25372 4632 25378 4644
rect 25869 4641 25881 4644
rect 25915 4672 25927 4675
rect 26881 4675 26939 4681
rect 26881 4672 26893 4675
rect 25915 4644 26893 4672
rect 25915 4641 25927 4644
rect 25869 4635 25927 4641
rect 26881 4641 26893 4644
rect 26927 4641 26939 4675
rect 27154 4672 27160 4684
rect 27115 4644 27160 4672
rect 26881 4635 26939 4641
rect 27154 4632 27160 4644
rect 27212 4632 27218 4684
rect 27430 4672 27436 4684
rect 27391 4644 27436 4672
rect 27430 4632 27436 4644
rect 27488 4632 27494 4684
rect 27985 4675 28043 4681
rect 27985 4641 27997 4675
rect 28031 4641 28043 4675
rect 27985 4635 28043 4641
rect 28445 4675 28503 4681
rect 28445 4641 28457 4675
rect 28491 4672 28503 4675
rect 28626 4672 28632 4684
rect 28491 4644 28632 4672
rect 28491 4641 28503 4644
rect 28445 4635 28503 4641
rect 18322 4604 18328 4616
rect 17460 4576 17505 4604
rect 17604 4576 18328 4604
rect 17460 4564 17466 4576
rect 18322 4564 18328 4576
rect 18380 4564 18386 4616
rect 18966 4564 18972 4616
rect 19024 4604 19030 4616
rect 19153 4607 19211 4613
rect 19153 4604 19165 4607
rect 19024 4576 19165 4604
rect 19024 4564 19030 4576
rect 19153 4573 19165 4576
rect 19199 4573 19211 4607
rect 19153 4567 19211 4573
rect 20714 4564 20720 4616
rect 20772 4604 20778 4616
rect 20993 4607 21051 4613
rect 20993 4604 21005 4607
rect 20772 4576 21005 4604
rect 20772 4564 20778 4576
rect 20993 4573 21005 4576
rect 21039 4573 21051 4607
rect 20993 4567 21051 4573
rect 21266 4564 21272 4616
rect 21324 4604 21330 4616
rect 21361 4607 21419 4613
rect 21361 4604 21373 4607
rect 21324 4576 21373 4604
rect 21324 4564 21330 4576
rect 21361 4573 21373 4576
rect 21407 4573 21419 4607
rect 25774 4604 25780 4616
rect 21361 4567 21419 4573
rect 21468 4576 25780 4604
rect 16666 4536 16672 4548
rect 13188 4508 16672 4536
rect 16666 4496 16672 4508
rect 16724 4496 16730 4548
rect 16761 4539 16819 4545
rect 16761 4505 16773 4539
rect 16807 4536 16819 4539
rect 21468 4536 21496 4576
rect 25774 4564 25780 4576
rect 25832 4564 25838 4616
rect 28000 4604 28028 4635
rect 28626 4632 28632 4644
rect 28684 4672 28690 4684
rect 28902 4672 28908 4684
rect 28684 4644 28908 4672
rect 28684 4632 28690 4644
rect 28902 4632 28908 4644
rect 28960 4632 28966 4684
rect 28994 4632 29000 4684
rect 29052 4672 29058 4684
rect 29365 4675 29423 4681
rect 29365 4672 29377 4675
rect 29052 4644 29377 4672
rect 29052 4632 29058 4644
rect 29365 4641 29377 4644
rect 29411 4672 29423 4675
rect 29454 4672 29460 4684
rect 29411 4644 29460 4672
rect 29411 4641 29423 4644
rect 29365 4635 29423 4641
rect 29454 4632 29460 4644
rect 29512 4632 29518 4684
rect 29932 4681 29960 4712
rect 30466 4700 30472 4712
rect 30524 4700 30530 4752
rect 30650 4700 30656 4752
rect 30708 4740 30714 4752
rect 31573 4743 31631 4749
rect 31573 4740 31585 4743
rect 30708 4712 31585 4740
rect 30708 4700 30714 4712
rect 31573 4709 31585 4712
rect 31619 4709 31631 4743
rect 31754 4740 31760 4752
rect 31715 4712 31760 4740
rect 31573 4703 31631 4709
rect 31754 4700 31760 4712
rect 31812 4700 31818 4752
rect 34149 4743 34207 4749
rect 34149 4709 34161 4743
rect 34195 4740 34207 4743
rect 38654 4740 38660 4752
rect 34195 4712 38660 4740
rect 34195 4709 34207 4712
rect 34149 4703 34207 4709
rect 38654 4700 38660 4712
rect 38712 4700 38718 4752
rect 39209 4743 39267 4749
rect 39209 4709 39221 4743
rect 39255 4740 39267 4743
rect 39574 4740 39580 4752
rect 39255 4712 39580 4740
rect 39255 4709 39267 4712
rect 39209 4703 39267 4709
rect 39574 4700 39580 4712
rect 39632 4700 39638 4752
rect 39684 4740 39712 4780
rect 39758 4768 39764 4820
rect 39816 4808 39822 4820
rect 46566 4808 46572 4820
rect 39816 4780 46572 4808
rect 39816 4768 39822 4780
rect 46566 4768 46572 4780
rect 46624 4768 46630 4820
rect 47210 4768 47216 4820
rect 47268 4808 47274 4820
rect 48130 4808 48136 4820
rect 47268 4780 48136 4808
rect 47268 4768 47274 4780
rect 48130 4768 48136 4780
rect 48188 4808 48194 4820
rect 48685 4811 48743 4817
rect 48685 4808 48697 4811
rect 48188 4780 48697 4808
rect 48188 4768 48194 4780
rect 48685 4777 48697 4780
rect 48731 4777 48743 4811
rect 49786 4808 49792 4820
rect 49747 4780 49792 4808
rect 48685 4771 48743 4777
rect 49786 4768 49792 4780
rect 49844 4768 49850 4820
rect 50062 4768 50068 4820
rect 50120 4808 50126 4820
rect 50890 4808 50896 4820
rect 50120 4780 50896 4808
rect 50120 4768 50126 4780
rect 50890 4768 50896 4780
rect 50948 4768 50954 4820
rect 57054 4808 57060 4820
rect 51368 4780 57060 4808
rect 42521 4743 42579 4749
rect 42521 4740 42533 4743
rect 39684 4712 42533 4740
rect 29917 4675 29975 4681
rect 29917 4641 29929 4675
rect 29963 4641 29975 4675
rect 32766 4672 32772 4684
rect 29917 4635 29975 4641
rect 30116 4644 32772 4672
rect 28813 4607 28871 4613
rect 28813 4604 28825 4607
rect 26068 4576 26740 4604
rect 28000 4576 28825 4604
rect 16807 4508 21496 4536
rect 16807 4505 16819 4508
rect 16761 4499 16819 4505
rect 21542 4496 21548 4548
rect 21600 4536 21606 4548
rect 26068 4536 26096 4576
rect 26513 4539 26571 4545
rect 26513 4536 26525 4539
rect 21600 4508 26096 4536
rect 26160 4508 26525 4536
rect 21600 4496 21606 4508
rect 3510 4468 3516 4480
rect 3471 4440 3516 4468
rect 3510 4428 3516 4440
rect 3568 4428 3574 4480
rect 5350 4428 5356 4480
rect 5408 4468 5414 4480
rect 5813 4471 5871 4477
rect 5813 4468 5825 4471
rect 5408 4440 5825 4468
rect 5408 4428 5414 4440
rect 5813 4437 5825 4440
rect 5859 4468 5871 4471
rect 6273 4471 6331 4477
rect 6273 4468 6285 4471
rect 5859 4440 6285 4468
rect 5859 4437 5871 4440
rect 5813 4431 5871 4437
rect 6273 4437 6285 4440
rect 6319 4468 6331 4471
rect 7834 4468 7840 4480
rect 6319 4440 7840 4468
rect 6319 4437 6331 4440
rect 6273 4431 6331 4437
rect 7834 4428 7840 4440
rect 7892 4428 7898 4480
rect 7929 4471 7987 4477
rect 7929 4437 7941 4471
rect 7975 4468 7987 4471
rect 8018 4468 8024 4480
rect 7975 4440 8024 4468
rect 7975 4437 7987 4440
rect 7929 4431 7987 4437
rect 8018 4428 8024 4440
rect 8076 4428 8082 4480
rect 8662 4428 8668 4480
rect 8720 4468 8726 4480
rect 9490 4468 9496 4480
rect 8720 4440 9496 4468
rect 8720 4428 8726 4440
rect 9490 4428 9496 4440
rect 9548 4428 9554 4480
rect 10321 4471 10379 4477
rect 10321 4437 10333 4471
rect 10367 4468 10379 4471
rect 10686 4468 10692 4480
rect 10367 4440 10692 4468
rect 10367 4437 10379 4440
rect 10321 4431 10379 4437
rect 10686 4428 10692 4440
rect 10744 4428 10750 4480
rect 11238 4468 11244 4480
rect 11199 4440 11244 4468
rect 11238 4428 11244 4440
rect 11296 4428 11302 4480
rect 11885 4471 11943 4477
rect 11885 4437 11897 4471
rect 11931 4468 11943 4471
rect 11974 4468 11980 4480
rect 11931 4440 11980 4468
rect 11931 4437 11943 4440
rect 11885 4431 11943 4437
rect 11974 4428 11980 4440
rect 12032 4428 12038 4480
rect 12526 4468 12532 4480
rect 12487 4440 12532 4468
rect 12526 4428 12532 4440
rect 12584 4428 12590 4480
rect 12710 4428 12716 4480
rect 12768 4468 12774 4480
rect 13354 4468 13360 4480
rect 12768 4440 13360 4468
rect 12768 4428 12774 4440
rect 13354 4428 13360 4440
rect 13412 4428 13418 4480
rect 13630 4428 13636 4480
rect 13688 4468 13694 4480
rect 14645 4471 14703 4477
rect 14645 4468 14657 4471
rect 13688 4440 14657 4468
rect 13688 4428 13694 4440
rect 14645 4437 14657 4440
rect 14691 4468 14703 4471
rect 15194 4468 15200 4480
rect 14691 4440 15200 4468
rect 14691 4437 14703 4440
rect 14645 4431 14703 4437
rect 15194 4428 15200 4440
rect 15252 4428 15258 4480
rect 15470 4428 15476 4480
rect 15528 4468 15534 4480
rect 15528 4440 15573 4468
rect 15528 4428 15534 4440
rect 16114 4428 16120 4480
rect 16172 4468 16178 4480
rect 16301 4471 16359 4477
rect 16301 4468 16313 4471
rect 16172 4440 16313 4468
rect 16172 4428 16178 4440
rect 16301 4437 16313 4440
rect 16347 4468 16359 4471
rect 17494 4468 17500 4480
rect 16347 4440 17500 4468
rect 16347 4437 16359 4440
rect 16301 4431 16359 4437
rect 17494 4428 17500 4440
rect 17552 4428 17558 4480
rect 17954 4428 17960 4480
rect 18012 4468 18018 4480
rect 19613 4471 19671 4477
rect 19613 4468 19625 4471
rect 18012 4440 19625 4468
rect 18012 4428 18018 4440
rect 19613 4437 19625 4440
rect 19659 4437 19671 4471
rect 19794 4468 19800 4480
rect 19755 4440 19800 4468
rect 19613 4431 19671 4437
rect 19794 4428 19800 4440
rect 19852 4428 19858 4480
rect 20254 4468 20260 4480
rect 20215 4440 20260 4468
rect 20254 4428 20260 4440
rect 20312 4468 20318 4480
rect 20530 4468 20536 4480
rect 20312 4440 20536 4468
rect 20312 4428 20318 4440
rect 20530 4428 20536 4440
rect 20588 4428 20594 4480
rect 20714 4468 20720 4480
rect 20675 4440 20720 4468
rect 20714 4428 20720 4440
rect 20772 4428 20778 4480
rect 22186 4468 22192 4480
rect 22147 4440 22192 4468
rect 22186 4428 22192 4440
rect 22244 4468 22250 4480
rect 22373 4471 22431 4477
rect 22373 4468 22385 4471
rect 22244 4440 22385 4468
rect 22244 4428 22250 4440
rect 22373 4437 22385 4440
rect 22419 4437 22431 4471
rect 22373 4431 22431 4437
rect 22646 4428 22652 4480
rect 22704 4468 22710 4480
rect 22741 4471 22799 4477
rect 22741 4468 22753 4471
rect 22704 4440 22753 4468
rect 22704 4428 22710 4440
rect 22741 4437 22753 4440
rect 22787 4437 22799 4471
rect 22741 4431 22799 4437
rect 23014 4428 23020 4480
rect 23072 4468 23078 4480
rect 23293 4471 23351 4477
rect 23293 4468 23305 4471
rect 23072 4440 23305 4468
rect 23072 4428 23078 4440
rect 23293 4437 23305 4440
rect 23339 4437 23351 4471
rect 23658 4468 23664 4480
rect 23619 4440 23664 4468
rect 23293 4431 23351 4437
rect 23658 4428 23664 4440
rect 23716 4428 23722 4480
rect 24486 4428 24492 4480
rect 24544 4468 24550 4480
rect 25501 4471 25559 4477
rect 25501 4468 25513 4471
rect 24544 4440 25513 4468
rect 24544 4428 24550 4440
rect 25501 4437 25513 4440
rect 25547 4437 25559 4471
rect 25501 4431 25559 4437
rect 25774 4428 25780 4480
rect 25832 4468 25838 4480
rect 26160 4468 26188 4508
rect 26513 4505 26525 4508
rect 26559 4536 26571 4539
rect 26602 4536 26608 4548
rect 26559 4508 26608 4536
rect 26559 4505 26571 4508
rect 26513 4499 26571 4505
rect 26602 4496 26608 4508
rect 26660 4496 26666 4548
rect 26712 4536 26740 4576
rect 28813 4573 28825 4576
rect 28859 4604 28871 4607
rect 30116 4604 30144 4644
rect 32766 4632 32772 4644
rect 32824 4632 32830 4684
rect 32953 4675 33011 4681
rect 32953 4641 32965 4675
rect 32999 4641 33011 4675
rect 32953 4635 33011 4641
rect 33689 4675 33747 4681
rect 33689 4641 33701 4675
rect 33735 4672 33747 4675
rect 34422 4672 34428 4684
rect 33735 4644 34428 4672
rect 33735 4641 33747 4644
rect 33689 4635 33747 4641
rect 28859 4576 30144 4604
rect 28859 4573 28871 4576
rect 28813 4567 28871 4573
rect 30190 4564 30196 4616
rect 30248 4604 30254 4616
rect 31389 4607 31447 4613
rect 31389 4604 31401 4607
rect 30248 4576 31401 4604
rect 30248 4564 30254 4576
rect 31389 4573 31401 4576
rect 31435 4573 31447 4607
rect 31389 4567 31447 4573
rect 31573 4607 31631 4613
rect 31573 4573 31585 4607
rect 31619 4604 31631 4607
rect 32968 4604 32996 4635
rect 34422 4632 34428 4644
rect 34480 4672 34486 4684
rect 34609 4675 34667 4681
rect 34609 4672 34621 4675
rect 34480 4644 34621 4672
rect 34480 4632 34486 4644
rect 34609 4641 34621 4644
rect 34655 4641 34667 4675
rect 34609 4635 34667 4641
rect 34793 4675 34851 4681
rect 34793 4641 34805 4675
rect 34839 4641 34851 4675
rect 34974 4672 34980 4684
rect 34935 4644 34980 4672
rect 34793 4635 34851 4641
rect 33502 4604 33508 4616
rect 31619 4576 33508 4604
rect 31619 4573 31631 4576
rect 31573 4567 31631 4573
rect 33502 4564 33508 4576
rect 33560 4564 33566 4616
rect 34514 4564 34520 4616
rect 34572 4604 34578 4616
rect 34808 4604 34836 4635
rect 34974 4632 34980 4644
rect 35032 4632 35038 4684
rect 35253 4675 35311 4681
rect 35253 4641 35265 4675
rect 35299 4641 35311 4675
rect 35434 4672 35440 4684
rect 35395 4644 35440 4672
rect 35253 4635 35311 4641
rect 34572 4576 34836 4604
rect 35268 4604 35296 4635
rect 35434 4632 35440 4644
rect 35492 4632 35498 4684
rect 36446 4672 36452 4684
rect 36407 4644 36452 4672
rect 36446 4632 36452 4644
rect 36504 4632 36510 4684
rect 37918 4672 37924 4684
rect 37879 4644 37924 4672
rect 37918 4632 37924 4644
rect 37976 4632 37982 4684
rect 38749 4675 38807 4681
rect 38749 4641 38761 4675
rect 38795 4672 38807 4675
rect 39022 4672 39028 4684
rect 38795 4644 39028 4672
rect 38795 4641 38807 4644
rect 38749 4635 38807 4641
rect 39022 4632 39028 4644
rect 39080 4632 39086 4684
rect 39850 4672 39856 4684
rect 39811 4644 39856 4672
rect 39850 4632 39856 4644
rect 39908 4632 39914 4684
rect 40218 4672 40224 4684
rect 40179 4644 40224 4672
rect 40218 4632 40224 4644
rect 40276 4632 40282 4684
rect 40310 4632 40316 4684
rect 40368 4672 40374 4684
rect 41892 4681 41920 4712
rect 42521 4709 42533 4712
rect 42567 4709 42579 4743
rect 42521 4703 42579 4709
rect 43165 4743 43223 4749
rect 43165 4709 43177 4743
rect 43211 4740 43223 4743
rect 43806 4740 43812 4752
rect 43211 4712 43812 4740
rect 43211 4709 43223 4712
rect 43165 4703 43223 4709
rect 40405 4675 40463 4681
rect 40405 4672 40417 4675
rect 40368 4644 40417 4672
rect 40368 4632 40374 4644
rect 40405 4641 40417 4644
rect 40451 4672 40463 4675
rect 41233 4675 41291 4681
rect 41233 4672 41245 4675
rect 40451 4644 41245 4672
rect 40451 4641 40463 4644
rect 40405 4635 40463 4641
rect 41233 4641 41245 4644
rect 41279 4641 41291 4675
rect 41233 4635 41291 4641
rect 41693 4675 41751 4681
rect 41693 4641 41705 4675
rect 41739 4641 41751 4675
rect 41693 4635 41751 4641
rect 41877 4675 41935 4681
rect 41877 4641 41889 4675
rect 41923 4641 41935 4675
rect 41877 4635 41935 4641
rect 42061 4675 42119 4681
rect 42061 4641 42073 4675
rect 42107 4672 42119 4675
rect 42150 4672 42156 4684
rect 42107 4644 42156 4672
rect 42107 4641 42119 4644
rect 42061 4635 42119 4641
rect 35802 4604 35808 4616
rect 35268 4576 35808 4604
rect 34572 4564 34578 4576
rect 26712 4508 30144 4536
rect 25832 4440 26188 4468
rect 26329 4471 26387 4477
rect 25832 4428 25838 4440
rect 26329 4437 26341 4471
rect 26375 4468 26387 4471
rect 27890 4468 27896 4480
rect 26375 4440 27896 4468
rect 26375 4437 26387 4440
rect 26329 4431 26387 4437
rect 27890 4428 27896 4440
rect 27948 4428 27954 4480
rect 29638 4468 29644 4480
rect 29599 4440 29644 4468
rect 29638 4428 29644 4440
rect 29696 4428 29702 4480
rect 30116 4477 30144 4508
rect 30282 4496 30288 4548
rect 30340 4536 30346 4548
rect 30340 4508 31156 4536
rect 30340 4496 30346 4508
rect 30101 4471 30159 4477
rect 30101 4437 30113 4471
rect 30147 4437 30159 4471
rect 30101 4431 30159 4437
rect 30466 4428 30472 4480
rect 30524 4468 30530 4480
rect 31128 4477 31156 4508
rect 31846 4496 31852 4548
rect 31904 4536 31910 4548
rect 32306 4536 32312 4548
rect 31904 4508 32312 4536
rect 31904 4496 31910 4508
rect 32306 4496 32312 4508
rect 32364 4496 32370 4548
rect 32401 4539 32459 4545
rect 32401 4505 32413 4539
rect 32447 4536 32459 4539
rect 32490 4536 32496 4548
rect 32447 4508 32496 4536
rect 32447 4505 32459 4508
rect 32401 4499 32459 4505
rect 32490 4496 32496 4508
rect 32548 4496 32554 4548
rect 32861 4539 32919 4545
rect 32861 4505 32873 4539
rect 32907 4536 32919 4539
rect 32950 4536 32956 4548
rect 32907 4508 32956 4536
rect 32907 4505 32919 4508
rect 32861 4499 32919 4505
rect 32950 4496 32956 4508
rect 33008 4496 33014 4548
rect 33134 4536 33140 4548
rect 33095 4508 33140 4536
rect 33134 4496 33140 4508
rect 33192 4496 33198 4548
rect 34808 4536 34836 4576
rect 35802 4564 35808 4576
rect 35860 4604 35866 4616
rect 35897 4607 35955 4613
rect 35897 4604 35909 4607
rect 35860 4576 35909 4604
rect 35860 4564 35866 4576
rect 35897 4573 35909 4576
rect 35943 4573 35955 4607
rect 35897 4567 35955 4573
rect 35986 4564 35992 4616
rect 36044 4604 36050 4616
rect 37001 4607 37059 4613
rect 37001 4604 37013 4607
rect 36044 4576 37013 4604
rect 36044 4564 36050 4576
rect 37001 4573 37013 4576
rect 37047 4604 37059 4607
rect 37182 4604 37188 4616
rect 37047 4576 37188 4604
rect 37047 4573 37059 4576
rect 37001 4567 37059 4573
rect 37182 4564 37188 4576
rect 37240 4564 37246 4616
rect 37550 4564 37556 4616
rect 37608 4604 37614 4616
rect 38933 4607 38991 4613
rect 38933 4604 38945 4607
rect 37608 4576 38945 4604
rect 37608 4564 37614 4576
rect 38764 4548 38792 4576
rect 38933 4573 38945 4576
rect 38979 4604 38991 4607
rect 38979 4576 39068 4604
rect 38979 4573 38991 4576
rect 38933 4567 38991 4573
rect 36265 4539 36323 4545
rect 36265 4536 36277 4539
rect 34808 4508 36277 4536
rect 36265 4505 36277 4508
rect 36311 4505 36323 4539
rect 36265 4499 36323 4505
rect 36633 4539 36691 4545
rect 36633 4505 36645 4539
rect 36679 4536 36691 4539
rect 37918 4536 37924 4548
rect 36679 4508 37924 4536
rect 36679 4505 36691 4508
rect 36633 4499 36691 4505
rect 37918 4496 37924 4508
rect 37976 4496 37982 4548
rect 38105 4539 38163 4545
rect 38105 4505 38117 4539
rect 38151 4536 38163 4539
rect 38562 4536 38568 4548
rect 38151 4508 38568 4536
rect 38151 4505 38163 4508
rect 38105 4499 38163 4505
rect 38562 4496 38568 4508
rect 38620 4496 38626 4548
rect 38746 4496 38752 4548
rect 38804 4496 38810 4548
rect 39040 4545 39068 4576
rect 39574 4564 39580 4616
rect 39632 4604 39638 4616
rect 39945 4607 40003 4613
rect 39945 4604 39957 4607
rect 39632 4576 39957 4604
rect 39632 4564 39638 4576
rect 39945 4573 39957 4576
rect 39991 4604 40003 4607
rect 41049 4607 41107 4613
rect 41049 4604 41061 4607
rect 39991 4576 41061 4604
rect 39991 4573 40003 4576
rect 39945 4567 40003 4573
rect 41049 4573 41061 4576
rect 41095 4573 41107 4607
rect 41708 4604 41736 4635
rect 42150 4632 42156 4644
rect 42208 4632 42214 4684
rect 43180 4672 43208 4703
rect 43806 4700 43812 4712
rect 43864 4700 43870 4752
rect 44082 4700 44088 4752
rect 44140 4740 44146 4752
rect 47118 4740 47124 4752
rect 44140 4712 47124 4740
rect 44140 4700 44146 4712
rect 47118 4700 47124 4712
rect 47176 4700 47182 4752
rect 47486 4740 47492 4752
rect 47399 4712 47492 4740
rect 47486 4700 47492 4712
rect 47544 4740 47550 4752
rect 48958 4740 48964 4752
rect 47544 4712 48964 4740
rect 47544 4700 47550 4712
rect 48958 4700 48964 4712
rect 49016 4740 49022 4752
rect 49602 4740 49608 4752
rect 49016 4712 49608 4740
rect 49016 4700 49022 4712
rect 49602 4700 49608 4712
rect 49660 4700 49666 4752
rect 42352 4644 43208 4672
rect 41966 4604 41972 4616
rect 41708 4576 41972 4604
rect 41049 4567 41107 4573
rect 41966 4564 41972 4576
rect 42024 4564 42030 4616
rect 39025 4539 39083 4545
rect 39025 4505 39037 4539
rect 39071 4505 39083 4539
rect 39025 4499 39083 4505
rect 40034 4496 40040 4548
rect 40092 4536 40098 4548
rect 42352 4536 42380 4644
rect 43622 4632 43628 4684
rect 43680 4672 43686 4684
rect 43993 4675 44051 4681
rect 43993 4672 44005 4675
rect 43680 4644 44005 4672
rect 43680 4632 43686 4644
rect 43993 4641 44005 4644
rect 44039 4672 44051 4675
rect 44729 4675 44787 4681
rect 44729 4672 44741 4675
rect 44039 4644 44741 4672
rect 44039 4641 44051 4644
rect 43993 4635 44051 4641
rect 44729 4641 44741 4644
rect 44775 4641 44787 4675
rect 44729 4635 44787 4641
rect 45741 4675 45799 4681
rect 45741 4641 45753 4675
rect 45787 4641 45799 4675
rect 46106 4672 46112 4684
rect 46067 4644 46112 4672
rect 45741 4635 45799 4641
rect 45646 4604 45652 4616
rect 45607 4576 45652 4604
rect 45646 4564 45652 4576
rect 45704 4564 45710 4616
rect 40092 4508 42380 4536
rect 40092 4496 40098 4508
rect 42426 4496 42432 4548
rect 42484 4536 42490 4548
rect 45756 4536 45784 4635
rect 46106 4632 46112 4644
rect 46164 4632 46170 4684
rect 46290 4672 46296 4684
rect 46251 4644 46296 4672
rect 46290 4632 46296 4644
rect 46348 4632 46354 4684
rect 47305 4675 47363 4681
rect 47305 4641 47317 4675
rect 47351 4641 47363 4675
rect 47305 4635 47363 4641
rect 47397 4675 47455 4681
rect 47397 4641 47409 4675
rect 47443 4672 47455 4675
rect 47578 4672 47584 4684
rect 47443 4644 47584 4672
rect 47443 4641 47455 4644
rect 47397 4635 47455 4641
rect 46124 4604 46152 4632
rect 46937 4607 46995 4613
rect 46937 4604 46949 4607
rect 46124 4576 46949 4604
rect 46937 4573 46949 4576
rect 46983 4573 46995 4607
rect 46937 4567 46995 4573
rect 47320 4536 47348 4635
rect 47578 4632 47584 4644
rect 47636 4632 47642 4684
rect 48130 4632 48136 4684
rect 48188 4672 48194 4684
rect 49694 4672 49700 4684
rect 48188 4644 49700 4672
rect 48188 4632 48194 4644
rect 49694 4632 49700 4644
rect 49752 4632 49758 4684
rect 49804 4672 49832 4768
rect 50157 4743 50215 4749
rect 50157 4709 50169 4743
rect 50203 4740 50215 4743
rect 50338 4740 50344 4752
rect 50203 4712 50344 4740
rect 50203 4709 50215 4712
rect 50157 4703 50215 4709
rect 50338 4700 50344 4712
rect 50396 4740 50402 4752
rect 50985 4743 51043 4749
rect 50985 4740 50997 4743
rect 50396 4712 50997 4740
rect 50396 4700 50402 4712
rect 50985 4709 50997 4712
rect 51031 4709 51043 4743
rect 50985 4703 51043 4709
rect 50249 4675 50307 4681
rect 50249 4672 50261 4675
rect 49804 4644 50261 4672
rect 50249 4641 50261 4644
rect 50295 4641 50307 4675
rect 50249 4635 50307 4641
rect 50709 4675 50767 4681
rect 50709 4641 50721 4675
rect 50755 4672 50767 4675
rect 51368 4672 51396 4780
rect 57054 4768 57060 4780
rect 57112 4768 57118 4820
rect 57330 4808 57336 4820
rect 57291 4780 57336 4808
rect 57330 4768 57336 4780
rect 57388 4768 57394 4820
rect 58066 4808 58072 4820
rect 58027 4780 58072 4808
rect 58066 4768 58072 4780
rect 58124 4768 58130 4820
rect 61562 4808 61568 4820
rect 58176 4780 61568 4808
rect 51534 4740 51540 4752
rect 51495 4712 51540 4740
rect 51534 4700 51540 4712
rect 51592 4700 51598 4752
rect 51810 4700 51816 4752
rect 51868 4740 51874 4752
rect 52270 4740 52276 4752
rect 51868 4712 52276 4740
rect 51868 4700 51874 4712
rect 52270 4700 52276 4712
rect 52328 4700 52334 4752
rect 52362 4700 52368 4752
rect 52420 4740 52426 4752
rect 53650 4740 53656 4752
rect 52420 4712 53656 4740
rect 52420 4700 52426 4712
rect 53650 4700 53656 4712
rect 53708 4740 53714 4752
rect 53929 4743 53987 4749
rect 53929 4740 53941 4743
rect 53708 4712 53941 4740
rect 53708 4700 53714 4712
rect 53929 4709 53941 4712
rect 53975 4709 53987 4743
rect 55398 4740 55404 4752
rect 53929 4703 53987 4709
rect 54404 4712 54800 4740
rect 55359 4712 55404 4740
rect 50755 4644 51396 4672
rect 50755 4641 50767 4644
rect 50709 4635 50767 4641
rect 51994 4632 52000 4684
rect 52052 4672 52058 4684
rect 53101 4675 53159 4681
rect 53101 4672 53113 4675
rect 52052 4644 53113 4672
rect 52052 4632 52058 4644
rect 53101 4641 53113 4644
rect 53147 4672 53159 4675
rect 53190 4672 53196 4684
rect 53147 4644 53196 4672
rect 53147 4641 53159 4644
rect 53101 4635 53159 4641
rect 53190 4632 53196 4644
rect 53248 4632 53254 4684
rect 53285 4675 53343 4681
rect 53285 4641 53297 4675
rect 53331 4672 53343 4675
rect 54404 4672 54432 4712
rect 54772 4684 54800 4712
rect 55398 4700 55404 4712
rect 55456 4700 55462 4752
rect 53331 4644 54432 4672
rect 53331 4641 53343 4644
rect 53285 4635 53343 4641
rect 54478 4632 54484 4684
rect 54536 4672 54542 4684
rect 54573 4675 54631 4681
rect 54573 4672 54585 4675
rect 54536 4644 54585 4672
rect 54536 4632 54542 4644
rect 54573 4641 54585 4644
rect 54619 4641 54631 4675
rect 54573 4635 54631 4641
rect 54754 4632 54760 4684
rect 54812 4672 54818 4684
rect 58176 4672 58204 4780
rect 61562 4768 61568 4780
rect 61620 4768 61626 4820
rect 58253 4743 58311 4749
rect 58253 4709 58265 4743
rect 58299 4740 58311 4743
rect 59814 4740 59820 4752
rect 58299 4712 59820 4740
rect 58299 4709 58311 4712
rect 58253 4703 58311 4709
rect 59814 4700 59820 4712
rect 59872 4700 59878 4752
rect 54812 4644 58204 4672
rect 54812 4632 54818 4644
rect 58342 4632 58348 4684
rect 58400 4672 58406 4684
rect 59078 4672 59084 4684
rect 58400 4644 59084 4672
rect 58400 4632 58406 4644
rect 59078 4632 59084 4644
rect 59136 4672 59142 4684
rect 59909 4675 59967 4681
rect 59909 4672 59921 4675
rect 59136 4644 59921 4672
rect 59136 4632 59142 4644
rect 59909 4641 59921 4644
rect 59955 4641 59967 4675
rect 61010 4672 61016 4684
rect 60971 4644 61016 4672
rect 59909 4635 59967 4641
rect 61010 4632 61016 4644
rect 61068 4632 61074 4684
rect 61194 4672 61200 4684
rect 61155 4644 61200 4672
rect 61194 4632 61200 4644
rect 61252 4632 61258 4684
rect 47854 4604 47860 4616
rect 47815 4576 47860 4604
rect 47854 4564 47860 4576
rect 47912 4564 47918 4616
rect 48866 4564 48872 4616
rect 48924 4604 48930 4616
rect 49973 4607 50031 4613
rect 49973 4604 49985 4607
rect 48924 4576 49985 4604
rect 48924 4564 48930 4576
rect 49973 4573 49985 4576
rect 50019 4604 50031 4607
rect 50614 4604 50620 4616
rect 50019 4576 50620 4604
rect 50019 4573 50031 4576
rect 49973 4567 50031 4573
rect 50614 4564 50620 4576
rect 50672 4564 50678 4616
rect 51905 4607 51963 4613
rect 51905 4573 51917 4607
rect 51951 4604 51963 4607
rect 53653 4607 53711 4613
rect 51951 4576 53604 4604
rect 51951 4573 51963 4576
rect 51905 4567 51963 4573
rect 51166 4536 51172 4548
rect 42484 4508 46704 4536
rect 47320 4508 51172 4536
rect 42484 4496 42490 4508
rect 30653 4471 30711 4477
rect 30653 4468 30665 4471
rect 30524 4440 30665 4468
rect 30524 4428 30530 4440
rect 30653 4437 30665 4440
rect 30699 4437 30711 4471
rect 30653 4431 30711 4437
rect 31113 4471 31171 4477
rect 31113 4437 31125 4471
rect 31159 4468 31171 4471
rect 33318 4468 33324 4480
rect 31159 4440 33324 4468
rect 31159 4437 31171 4440
rect 31113 4431 31171 4437
rect 33318 4428 33324 4440
rect 33376 4428 33382 4480
rect 33962 4468 33968 4480
rect 33923 4440 33968 4468
rect 33962 4428 33968 4440
rect 34020 4468 34026 4480
rect 35434 4468 35440 4480
rect 34020 4440 35440 4468
rect 34020 4428 34026 4440
rect 35434 4428 35440 4440
rect 35492 4468 35498 4480
rect 36446 4468 36452 4480
rect 35492 4440 36452 4468
rect 35492 4428 35498 4440
rect 36446 4428 36452 4440
rect 36504 4468 36510 4480
rect 37366 4468 37372 4480
rect 36504 4440 37372 4468
rect 36504 4428 36510 4440
rect 37366 4428 37372 4440
rect 37424 4428 37430 4480
rect 38841 4471 38899 4477
rect 38841 4437 38853 4471
rect 38887 4468 38899 4471
rect 40773 4471 40831 4477
rect 40773 4468 40785 4471
rect 38887 4440 40785 4468
rect 38887 4437 38899 4440
rect 38841 4431 38899 4437
rect 40773 4437 40785 4440
rect 40819 4468 40831 4471
rect 40862 4468 40868 4480
rect 40819 4440 40868 4468
rect 40819 4437 40831 4440
rect 40773 4431 40831 4437
rect 40862 4428 40868 4440
rect 40920 4428 40926 4480
rect 43622 4468 43628 4480
rect 43583 4440 43628 4468
rect 43622 4428 43628 4440
rect 43680 4428 43686 4480
rect 44174 4468 44180 4480
rect 44135 4440 44180 4468
rect 44174 4428 44180 4440
rect 44232 4428 44238 4480
rect 45189 4471 45247 4477
rect 45189 4437 45201 4471
rect 45235 4468 45247 4471
rect 45554 4468 45560 4480
rect 45235 4440 45560 4468
rect 45235 4437 45247 4440
rect 45189 4431 45247 4437
rect 45554 4428 45560 4440
rect 45612 4428 45618 4480
rect 46676 4477 46704 4508
rect 51166 4496 51172 4508
rect 51224 4496 51230 4548
rect 51442 4536 51448 4548
rect 51276 4508 51448 4536
rect 46661 4471 46719 4477
rect 46661 4437 46673 4471
rect 46707 4468 46719 4471
rect 48130 4468 48136 4480
rect 46707 4440 48136 4468
rect 46707 4437 46719 4440
rect 46661 4431 46719 4437
rect 48130 4428 48136 4440
rect 48188 4428 48194 4480
rect 48409 4471 48467 4477
rect 48409 4437 48421 4471
rect 48455 4468 48467 4471
rect 48682 4468 48688 4480
rect 48455 4440 48688 4468
rect 48455 4437 48467 4440
rect 48409 4431 48467 4437
rect 48682 4428 48688 4440
rect 48740 4428 48746 4480
rect 49142 4468 49148 4480
rect 49103 4440 49148 4468
rect 49142 4428 49148 4440
rect 49200 4428 49206 4480
rect 50982 4428 50988 4480
rect 51040 4468 51046 4480
rect 51276 4468 51304 4508
rect 51442 4496 51448 4508
rect 51500 4536 51506 4548
rect 51702 4539 51760 4545
rect 51702 4536 51714 4539
rect 51500 4508 51714 4536
rect 51500 4496 51506 4508
rect 51702 4505 51714 4508
rect 51748 4536 51760 4539
rect 52362 4536 52368 4548
rect 51748 4508 52368 4536
rect 51748 4505 51760 4508
rect 51702 4499 51760 4505
rect 52362 4496 52368 4508
rect 52420 4496 52426 4548
rect 51040 4440 51304 4468
rect 51353 4471 51411 4477
rect 51040 4428 51046 4440
rect 51353 4437 51365 4471
rect 51399 4468 51411 4471
rect 51534 4468 51540 4480
rect 51399 4440 51540 4468
rect 51399 4437 51411 4440
rect 51353 4431 51411 4437
rect 51534 4428 51540 4440
rect 51592 4428 51598 4480
rect 51813 4471 51871 4477
rect 51813 4437 51825 4471
rect 51859 4468 51871 4471
rect 51902 4468 51908 4480
rect 51859 4440 51908 4468
rect 51859 4437 51871 4440
rect 51813 4431 51871 4437
rect 51902 4428 51908 4440
rect 51960 4428 51966 4480
rect 52178 4428 52184 4480
rect 52236 4468 52242 4480
rect 52549 4471 52607 4477
rect 52549 4468 52561 4471
rect 52236 4440 52561 4468
rect 52236 4428 52242 4440
rect 52549 4437 52561 4440
rect 52595 4437 52607 4471
rect 52549 4431 52607 4437
rect 52730 4428 52736 4480
rect 52788 4468 52794 4480
rect 52917 4471 52975 4477
rect 52917 4468 52929 4471
rect 52788 4440 52929 4468
rect 52788 4428 52794 4440
rect 52917 4437 52929 4440
rect 52963 4437 52975 4471
rect 53576 4468 53604 4576
rect 53653 4573 53665 4607
rect 53699 4604 53711 4607
rect 54018 4604 54024 4616
rect 53699 4576 54024 4604
rect 53699 4573 53711 4576
rect 53653 4567 53711 4573
rect 54018 4564 54024 4576
rect 54076 4564 54082 4616
rect 55769 4607 55827 4613
rect 55769 4573 55781 4607
rect 55815 4573 55827 4607
rect 56042 4604 56048 4616
rect 56003 4576 56048 4604
rect 55769 4567 55827 4573
rect 54294 4536 54300 4548
rect 54255 4508 54300 4536
rect 54294 4496 54300 4508
rect 54352 4496 54358 4548
rect 54662 4496 54668 4548
rect 54720 4536 54726 4548
rect 54757 4539 54815 4545
rect 54757 4536 54769 4539
rect 54720 4508 54769 4536
rect 54720 4496 54726 4508
rect 54757 4505 54769 4508
rect 54803 4505 54815 4539
rect 54757 4499 54815 4505
rect 55122 4468 55128 4480
rect 53576 4440 55128 4468
rect 52917 4431 52975 4437
rect 55122 4428 55128 4440
rect 55180 4428 55186 4480
rect 55784 4468 55812 4567
rect 56042 4564 56048 4576
rect 56100 4564 56106 4616
rect 58805 4607 58863 4613
rect 58805 4573 58817 4607
rect 58851 4604 58863 4607
rect 58894 4604 58900 4616
rect 58851 4576 58900 4604
rect 58851 4573 58863 4576
rect 58805 4567 58863 4573
rect 58894 4564 58900 4576
rect 58952 4564 58958 4616
rect 59262 4604 59268 4616
rect 59223 4576 59268 4604
rect 59262 4564 59268 4576
rect 59320 4564 59326 4616
rect 59354 4564 59360 4616
rect 59412 4604 59418 4616
rect 60185 4607 60243 4613
rect 60185 4604 60197 4607
rect 59412 4576 60197 4604
rect 59412 4564 59418 4576
rect 60185 4573 60197 4576
rect 60231 4573 60243 4607
rect 60185 4567 60243 4573
rect 60737 4607 60795 4613
rect 60737 4573 60749 4607
rect 60783 4604 60795 4607
rect 61746 4604 61752 4616
rect 60783 4576 61752 4604
rect 60783 4573 60795 4576
rect 60737 4567 60795 4573
rect 61746 4564 61752 4576
rect 61804 4564 61810 4616
rect 58912 4536 58940 4564
rect 59446 4536 59452 4548
rect 58912 4508 59452 4536
rect 59446 4496 59452 4508
rect 59504 4496 59510 4548
rect 58434 4468 58440 4480
rect 55784 4440 58440 4468
rect 58434 4428 58440 4440
rect 58492 4428 58498 4480
rect 59538 4468 59544 4480
rect 59499 4440 59544 4468
rect 59538 4428 59544 4440
rect 59596 4428 59602 4480
rect 61470 4468 61476 4480
rect 61431 4440 61476 4468
rect 61470 4428 61476 4440
rect 61528 4428 61534 4480
rect 1104 4378 63480 4400
rect 1104 4326 11378 4378
rect 11430 4326 11442 4378
rect 11494 4326 11506 4378
rect 11558 4326 11570 4378
rect 11622 4326 32170 4378
rect 32222 4326 32234 4378
rect 32286 4326 32298 4378
rect 32350 4326 32362 4378
rect 32414 4326 52962 4378
rect 53014 4326 53026 4378
rect 53078 4326 53090 4378
rect 53142 4326 53154 4378
rect 53206 4326 63480 4378
rect 1104 4304 63480 4326
rect 2498 4264 2504 4276
rect 2459 4236 2504 4264
rect 2498 4224 2504 4236
rect 2556 4224 2562 4276
rect 3602 4264 3608 4276
rect 3563 4236 3608 4264
rect 3602 4224 3608 4236
rect 3660 4224 3666 4276
rect 4522 4224 4528 4276
rect 4580 4264 4586 4276
rect 4709 4267 4767 4273
rect 4709 4264 4721 4267
rect 4580 4236 4721 4264
rect 4580 4224 4586 4236
rect 4709 4233 4721 4236
rect 4755 4233 4767 4267
rect 7282 4264 7288 4276
rect 7243 4236 7288 4264
rect 4709 4227 4767 4233
rect 7282 4224 7288 4236
rect 7340 4224 7346 4276
rect 8754 4264 8760 4276
rect 8715 4236 8760 4264
rect 8754 4224 8760 4236
rect 8812 4224 8818 4276
rect 9582 4224 9588 4276
rect 9640 4264 9646 4276
rect 9953 4267 10011 4273
rect 9953 4264 9965 4267
rect 9640 4236 9965 4264
rect 9640 4224 9646 4236
rect 9953 4233 9965 4236
rect 9999 4233 10011 4267
rect 9953 4227 10011 4233
rect 11698 4224 11704 4276
rect 11756 4264 11762 4276
rect 12250 4264 12256 4276
rect 11756 4236 12256 4264
rect 11756 4224 11762 4236
rect 12250 4224 12256 4236
rect 12308 4224 12314 4276
rect 12434 4224 12440 4276
rect 12492 4264 12498 4276
rect 12575 4267 12633 4273
rect 12575 4264 12587 4267
rect 12492 4236 12587 4264
rect 12492 4224 12498 4236
rect 12575 4233 12587 4236
rect 12621 4233 12633 4267
rect 12710 4264 12716 4276
rect 12671 4236 12716 4264
rect 12575 4227 12633 4233
rect 12710 4224 12716 4236
rect 12768 4224 12774 4276
rect 13906 4264 13912 4276
rect 12912 4236 13124 4264
rect 13867 4236 13912 4264
rect 5166 4196 5172 4208
rect 5127 4168 5172 4196
rect 5166 4156 5172 4168
rect 5224 4156 5230 4208
rect 8481 4199 8539 4205
rect 8481 4165 8493 4199
rect 8527 4196 8539 4199
rect 8846 4196 8852 4208
rect 8527 4168 8852 4196
rect 8527 4165 8539 4168
rect 8481 4159 8539 4165
rect 8846 4156 8852 4168
rect 8904 4156 8910 4208
rect 9490 4156 9496 4208
rect 9548 4196 9554 4208
rect 10410 4196 10416 4208
rect 9548 4168 10416 4196
rect 9548 4156 9554 4168
rect 2133 4131 2191 4137
rect 2133 4097 2145 4131
rect 2179 4128 2191 4131
rect 3694 4128 3700 4140
rect 2179 4100 3700 4128
rect 2179 4097 2191 4100
rect 2133 4091 2191 4097
rect 3694 4088 3700 4100
rect 3752 4088 3758 4140
rect 5813 4131 5871 4137
rect 5813 4097 5825 4131
rect 5859 4128 5871 4131
rect 6641 4131 6699 4137
rect 6641 4128 6653 4131
rect 5859 4100 6653 4128
rect 5859 4097 5871 4100
rect 5813 4091 5871 4097
rect 6641 4097 6653 4100
rect 6687 4128 6699 4131
rect 7006 4128 7012 4140
rect 6687 4100 7012 4128
rect 6687 4097 6699 4100
rect 6641 4091 6699 4097
rect 7006 4088 7012 4100
rect 7064 4088 7070 4140
rect 10060 4137 10088 4168
rect 10410 4156 10416 4168
rect 10468 4156 10474 4208
rect 11425 4199 11483 4205
rect 11425 4165 11437 4199
rect 11471 4165 11483 4199
rect 11882 4196 11888 4208
rect 11843 4168 11888 4196
rect 11425 4159 11483 4165
rect 8113 4131 8171 4137
rect 8113 4097 8125 4131
rect 8159 4128 8171 4131
rect 10045 4131 10103 4137
rect 8159 4100 9996 4128
rect 8159 4097 8171 4100
rect 8113 4091 8171 4097
rect 3050 4020 3056 4072
rect 3108 4060 3114 4072
rect 3510 4069 3516 4072
rect 3476 4063 3516 4069
rect 3476 4060 3488 4063
rect 3108 4032 3488 4060
rect 3108 4020 3114 4032
rect 3476 4029 3488 4032
rect 3568 4060 3574 4072
rect 4062 4060 4068 4072
rect 3568 4032 3624 4060
rect 4023 4032 4068 4060
rect 3476 4023 3516 4029
rect 3510 4020 3516 4023
rect 3568 4020 3574 4032
rect 4062 4020 4068 4032
rect 4120 4020 4126 4072
rect 5350 4060 5356 4072
rect 5311 4032 5356 4060
rect 5350 4020 5356 4032
rect 5408 4020 5414 4072
rect 5721 4063 5779 4069
rect 5721 4029 5733 4063
rect 5767 4060 5779 4063
rect 6273 4063 6331 4069
rect 6273 4060 6285 4063
rect 5767 4032 6285 4060
rect 5767 4029 5779 4032
rect 5721 4023 5779 4029
rect 6273 4029 6285 4032
rect 6319 4060 6331 4063
rect 8018 4060 8024 4072
rect 6319 4032 8024 4060
rect 6319 4029 6331 4032
rect 6273 4023 6331 4029
rect 8018 4020 8024 4032
rect 8076 4020 8082 4072
rect 9858 4069 9864 4072
rect 9217 4063 9275 4069
rect 9217 4029 9229 4063
rect 9263 4060 9275 4063
rect 9824 4063 9864 4069
rect 9824 4060 9836 4063
rect 9263 4032 9836 4060
rect 9263 4029 9275 4032
rect 9217 4023 9275 4029
rect 9824 4029 9836 4032
rect 9824 4023 9864 4029
rect 9858 4020 9864 4023
rect 9916 4020 9922 4072
rect 9968 4060 9996 4100
rect 10045 4097 10057 4131
rect 10091 4097 10103 4131
rect 11054 4128 11060 4140
rect 10045 4091 10103 4097
rect 10244 4100 11060 4128
rect 10244 4060 10272 4100
rect 11054 4088 11060 4100
rect 11112 4088 11118 4140
rect 11440 4128 11468 4159
rect 11882 4156 11888 4168
rect 11940 4156 11946 4208
rect 12912 4196 12940 4236
rect 12268 4168 12940 4196
rect 13096 4196 13124 4236
rect 13906 4224 13912 4236
rect 13964 4224 13970 4276
rect 16209 4267 16267 4273
rect 16209 4233 16221 4267
rect 16255 4264 16267 4267
rect 16574 4264 16580 4276
rect 16255 4236 16580 4264
rect 16255 4233 16267 4236
rect 16209 4227 16267 4233
rect 16574 4224 16580 4236
rect 16632 4224 16638 4276
rect 16666 4224 16672 4276
rect 16724 4264 16730 4276
rect 17313 4267 17371 4273
rect 17313 4264 17325 4267
rect 16724 4236 17325 4264
rect 16724 4224 16730 4236
rect 17313 4233 17325 4236
rect 17359 4233 17371 4267
rect 17313 4227 17371 4233
rect 17494 4224 17500 4276
rect 17552 4264 17558 4276
rect 20806 4264 20812 4276
rect 17552 4236 20812 4264
rect 17552 4224 17558 4236
rect 20806 4224 20812 4236
rect 20864 4224 20870 4276
rect 22097 4267 22155 4273
rect 22097 4233 22109 4267
rect 22143 4264 22155 4267
rect 22186 4264 22192 4276
rect 22143 4236 22192 4264
rect 22143 4233 22155 4236
rect 22097 4227 22155 4233
rect 22186 4224 22192 4236
rect 22244 4264 22250 4276
rect 23566 4264 23572 4276
rect 22244 4236 23572 4264
rect 22244 4224 22250 4236
rect 23566 4224 23572 4236
rect 23624 4224 23630 4276
rect 23842 4264 23848 4276
rect 23803 4236 23848 4264
rect 23842 4224 23848 4236
rect 23900 4224 23906 4276
rect 23934 4224 23940 4276
rect 23992 4264 23998 4276
rect 27430 4264 27436 4276
rect 23992 4236 26280 4264
rect 27391 4236 27436 4264
rect 23992 4224 23998 4236
rect 14826 4196 14832 4208
rect 13096 4168 14504 4196
rect 14787 4168 14832 4196
rect 12268 4128 12296 4168
rect 12897 4131 12955 4137
rect 12897 4128 12909 4131
rect 11440 4100 12296 4128
rect 12360 4100 12909 4128
rect 10778 4060 10784 4072
rect 9968 4032 10272 4060
rect 10336 4032 10784 4060
rect 3237 3995 3295 4001
rect 3237 3961 3249 3995
rect 3283 3992 3295 3995
rect 3326 3992 3332 4004
rect 3283 3964 3332 3992
rect 3283 3961 3295 3964
rect 3237 3955 3295 3961
rect 3326 3952 3332 3964
rect 3384 3952 3390 4004
rect 3602 3952 3608 4004
rect 3660 3992 3666 4004
rect 4341 3995 4399 4001
rect 4341 3992 4353 3995
rect 3660 3964 4353 3992
rect 3660 3952 3666 3964
rect 4341 3961 4353 3964
rect 4387 3961 4399 3995
rect 4341 3955 4399 3961
rect 5626 3952 5632 4004
rect 5684 3992 5690 4004
rect 7377 3995 7435 4001
rect 7377 3992 7389 3995
rect 5684 3964 7389 3992
rect 5684 3952 5690 3964
rect 7377 3961 7389 3964
rect 7423 3961 7435 3995
rect 7377 3955 7435 3961
rect 7745 3995 7803 4001
rect 7745 3961 7757 3995
rect 7791 3992 7803 3995
rect 9490 3992 9496 4004
rect 7791 3964 9496 3992
rect 7791 3961 7803 3964
rect 7745 3955 7803 3961
rect 9490 3952 9496 3964
rect 9548 3952 9554 4004
rect 9585 3995 9643 4001
rect 9585 3961 9597 3995
rect 9631 3992 9643 3995
rect 9677 3995 9735 4001
rect 9677 3992 9689 3995
rect 9631 3964 9689 3992
rect 9631 3961 9643 3964
rect 9585 3955 9643 3961
rect 9677 3961 9689 3964
rect 9723 3992 9735 3995
rect 10336 3992 10364 4032
rect 10778 4020 10784 4032
rect 10836 4020 10842 4072
rect 11238 4060 11244 4072
rect 11151 4032 11244 4060
rect 11238 4020 11244 4032
rect 11296 4060 11302 4072
rect 12360 4060 12388 4100
rect 12897 4097 12909 4100
rect 12943 4097 12955 4131
rect 12897 4091 12955 4097
rect 13354 4088 13360 4140
rect 13412 4128 13418 4140
rect 13449 4131 13507 4137
rect 13449 4128 13461 4131
rect 13412 4100 13461 4128
rect 13412 4088 13418 4100
rect 13449 4097 13461 4100
rect 13495 4128 13507 4131
rect 13722 4128 13728 4140
rect 13495 4100 13728 4128
rect 13495 4097 13507 4100
rect 13449 4091 13507 4097
rect 13722 4088 13728 4100
rect 13780 4088 13786 4140
rect 14476 4072 14504 4168
rect 14826 4156 14832 4168
rect 14884 4156 14890 4208
rect 14918 4156 14924 4208
rect 14976 4196 14982 4208
rect 17402 4196 17408 4208
rect 14976 4168 15056 4196
rect 14976 4156 14982 4168
rect 15028 4137 15056 4168
rect 17052 4168 17408 4196
rect 17052 4137 17080 4168
rect 17402 4156 17408 4168
rect 17460 4196 17466 4208
rect 17681 4199 17739 4205
rect 17681 4196 17693 4199
rect 17460 4168 17693 4196
rect 17460 4156 17466 4168
rect 17681 4165 17693 4168
rect 17727 4165 17739 4199
rect 17681 4159 17739 4165
rect 19242 4156 19248 4208
rect 19300 4196 19306 4208
rect 25590 4196 25596 4208
rect 19300 4168 25596 4196
rect 19300 4156 19306 4168
rect 25590 4156 25596 4168
rect 25648 4156 25654 4208
rect 26145 4199 26203 4205
rect 26145 4196 26157 4199
rect 25700 4168 26157 4196
rect 15013 4131 15071 4137
rect 15013 4097 15025 4131
rect 15059 4097 15071 4131
rect 15013 4091 15071 4097
rect 17037 4131 17095 4137
rect 17037 4097 17049 4131
rect 17083 4097 17095 4131
rect 19429 4131 19487 4137
rect 19429 4128 19441 4131
rect 17037 4091 17095 4097
rect 18800 4100 19441 4128
rect 18800 4072 18828 4100
rect 19429 4097 19441 4100
rect 19475 4097 19487 4131
rect 19429 4091 19487 4097
rect 19981 4131 20039 4137
rect 19981 4097 19993 4131
rect 20027 4128 20039 4131
rect 20898 4128 20904 4140
rect 20027 4100 20904 4128
rect 20027 4097 20039 4100
rect 19981 4091 20039 4097
rect 20898 4088 20904 4100
rect 20956 4088 20962 4140
rect 20993 4131 21051 4137
rect 20993 4097 21005 4131
rect 21039 4128 21051 4131
rect 21082 4128 21088 4140
rect 21039 4100 21088 4128
rect 21039 4097 21051 4100
rect 20993 4091 21051 4097
rect 21082 4088 21088 4100
rect 21140 4088 21146 4140
rect 21174 4088 21180 4140
rect 21232 4128 21238 4140
rect 21361 4131 21419 4137
rect 21361 4128 21373 4131
rect 21232 4100 21373 4128
rect 21232 4088 21238 4100
rect 21361 4097 21373 4100
rect 21407 4128 21419 4131
rect 22002 4128 22008 4140
rect 21407 4100 22008 4128
rect 21407 4097 21419 4100
rect 21361 4091 21419 4097
rect 22002 4088 22008 4100
rect 22060 4088 22066 4140
rect 22094 4088 22100 4140
rect 22152 4128 22158 4140
rect 24213 4131 24271 4137
rect 24213 4128 24225 4131
rect 22152 4100 24225 4128
rect 22152 4088 22158 4100
rect 24213 4097 24225 4100
rect 24259 4097 24271 4131
rect 25314 4128 25320 4140
rect 24213 4091 24271 4097
rect 24504 4100 25320 4128
rect 11296 4032 12388 4060
rect 12776 4063 12834 4069
rect 11296 4020 11302 4032
rect 12776 4029 12788 4063
rect 12822 4060 12834 4063
rect 13170 4060 13176 4072
rect 12822 4032 13176 4060
rect 12822 4029 12834 4032
rect 12776 4023 12834 4029
rect 13170 4020 13176 4032
rect 13228 4020 13234 4072
rect 14182 4020 14188 4072
rect 14240 4060 14246 4072
rect 14366 4060 14372 4072
rect 14240 4032 14372 4060
rect 14240 4020 14246 4032
rect 14366 4020 14372 4032
rect 14424 4020 14430 4072
rect 14458 4020 14464 4072
rect 14516 4060 14522 4072
rect 14921 4063 14979 4069
rect 14921 4060 14933 4063
rect 14516 4032 14933 4060
rect 14516 4020 14522 4032
rect 14921 4029 14933 4032
rect 14967 4029 14979 4063
rect 14921 4023 14979 4029
rect 9723 3964 10364 3992
rect 10413 3995 10471 4001
rect 9723 3961 9735 3964
rect 9677 3955 9735 3961
rect 10413 3961 10425 3995
rect 10459 3992 10471 3995
rect 12437 3995 12495 4001
rect 12437 3992 12449 3995
rect 10459 3964 12449 3992
rect 10459 3961 10471 3964
rect 10413 3955 10471 3961
rect 12437 3961 12449 3964
rect 12483 3992 12495 3995
rect 12526 3992 12532 4004
rect 12483 3964 12532 3992
rect 12483 3961 12495 3964
rect 12437 3955 12495 3961
rect 12526 3952 12532 3964
rect 12584 3952 12590 4004
rect 13630 3992 13636 4004
rect 13004 3964 13636 3992
rect 2866 3924 2872 3936
rect 2827 3896 2872 3924
rect 2866 3884 2872 3896
rect 2924 3884 2930 3936
rect 6546 3884 6552 3936
rect 6604 3924 6610 3936
rect 7098 3924 7104 3936
rect 6604 3896 7104 3924
rect 6604 3884 6610 3896
rect 7098 3884 7104 3896
rect 7156 3884 7162 3936
rect 7466 3884 7472 3936
rect 7524 3924 7530 3936
rect 7561 3927 7619 3933
rect 7561 3924 7573 3927
rect 7524 3896 7573 3924
rect 7524 3884 7530 3896
rect 7561 3893 7573 3896
rect 7607 3893 7619 3927
rect 7561 3887 7619 3893
rect 7653 3927 7711 3933
rect 7653 3893 7665 3927
rect 7699 3924 7711 3927
rect 7834 3924 7840 3936
rect 7699 3896 7840 3924
rect 7699 3893 7711 3896
rect 7653 3887 7711 3893
rect 7834 3884 7840 3896
rect 7892 3884 7898 3936
rect 8018 3884 8024 3936
rect 8076 3924 8082 3936
rect 9766 3924 9772 3936
rect 8076 3896 9772 3924
rect 8076 3884 8082 3896
rect 9766 3884 9772 3896
rect 9824 3884 9830 3936
rect 10686 3924 10692 3936
rect 10647 3896 10692 3924
rect 10686 3884 10692 3896
rect 10744 3884 10750 3936
rect 10778 3884 10784 3936
rect 10836 3924 10842 3936
rect 11149 3927 11207 3933
rect 11149 3924 11161 3927
rect 10836 3896 11161 3924
rect 10836 3884 10842 3896
rect 11149 3893 11161 3896
rect 11195 3924 11207 3927
rect 13004 3924 13032 3964
rect 13630 3952 13636 3964
rect 13688 3952 13694 4004
rect 14936 3992 14964 4023
rect 15194 4020 15200 4072
rect 15252 4060 15258 4072
rect 18782 4060 18788 4072
rect 15252 4032 16712 4060
rect 18743 4032 18788 4060
rect 15252 4020 15258 4032
rect 15473 3995 15531 4001
rect 15473 3992 15485 3995
rect 14936 3964 15485 3992
rect 15473 3961 15485 3964
rect 15519 3992 15531 3995
rect 15654 3992 15660 4004
rect 15519 3964 15660 3992
rect 15519 3961 15531 3964
rect 15473 3955 15531 3961
rect 15654 3952 15660 3964
rect 15712 3952 15718 4004
rect 15930 3952 15936 4004
rect 15988 3992 15994 4004
rect 16684 4001 16712 4032
rect 18782 4020 18788 4032
rect 18840 4020 18846 4072
rect 20530 4060 20536 4072
rect 18892 4032 20392 4060
rect 20491 4032 20536 4060
rect 16301 3995 16359 4001
rect 16301 3992 16313 3995
rect 15988 3964 16313 3992
rect 15988 3952 15994 3964
rect 16301 3961 16313 3964
rect 16347 3961 16359 3995
rect 16301 3955 16359 3961
rect 16669 3995 16727 4001
rect 16669 3961 16681 3995
rect 16715 3992 16727 3995
rect 18230 3992 18236 4004
rect 16715 3964 18236 3992
rect 16715 3961 16727 3964
rect 16669 3955 16727 3961
rect 18230 3952 18236 3964
rect 18288 3952 18294 4004
rect 18509 3995 18567 4001
rect 18509 3961 18521 3995
rect 18555 3992 18567 3995
rect 18601 3995 18659 4001
rect 18601 3992 18613 3995
rect 18555 3964 18613 3992
rect 18555 3961 18567 3964
rect 18509 3955 18567 3961
rect 18601 3961 18613 3964
rect 18647 3992 18659 3995
rect 18892 3992 18920 4032
rect 18647 3964 18920 3992
rect 19153 3995 19211 4001
rect 18647 3961 18659 3964
rect 18601 3955 18659 3961
rect 19153 3961 19165 3995
rect 19199 3992 19211 3995
rect 19889 3995 19947 4001
rect 19889 3992 19901 3995
rect 19199 3964 19901 3992
rect 19199 3961 19211 3964
rect 19153 3955 19211 3961
rect 19889 3961 19901 3964
rect 19935 3992 19947 3995
rect 20162 3992 20168 4004
rect 19935 3964 20168 3992
rect 19935 3961 19947 3964
rect 19889 3955 19947 3961
rect 20162 3952 20168 3964
rect 20220 3952 20226 4004
rect 20364 3992 20392 4032
rect 20530 4020 20536 4032
rect 20588 4020 20594 4072
rect 20622 4020 20628 4072
rect 20680 4060 20686 4072
rect 20809 4063 20867 4069
rect 20809 4060 20821 4063
rect 20680 4032 20821 4060
rect 20680 4020 20686 4032
rect 20809 4029 20821 4032
rect 20855 4029 20867 4063
rect 21100 4060 21128 4088
rect 21637 4063 21695 4069
rect 21637 4060 21649 4063
rect 21100 4032 21649 4060
rect 20809 4023 20867 4029
rect 21637 4029 21649 4032
rect 21683 4060 21695 4063
rect 22373 4063 22431 4069
rect 21683 4032 22324 4060
rect 21683 4029 21695 4032
rect 21637 4023 21695 4029
rect 22186 3992 22192 4004
rect 20364 3964 22192 3992
rect 22186 3952 22192 3964
rect 22244 3952 22250 4004
rect 22296 3992 22324 4032
rect 22373 4029 22385 4063
rect 22419 4060 22431 4063
rect 22646 4060 22652 4072
rect 22419 4032 22652 4060
rect 22419 4029 22431 4032
rect 22373 4023 22431 4029
rect 22646 4020 22652 4032
rect 22704 4020 22710 4072
rect 22741 4063 22799 4069
rect 22741 4029 22753 4063
rect 22787 4060 22799 4063
rect 24302 4060 24308 4072
rect 22787 4032 24308 4060
rect 22787 4029 22799 4032
rect 22741 4023 22799 4029
rect 24302 4020 24308 4032
rect 24360 4020 24366 4072
rect 24504 3992 24532 4100
rect 25314 4088 25320 4100
rect 25372 4088 25378 4140
rect 25406 4088 25412 4140
rect 25464 4128 25470 4140
rect 25700 4128 25728 4168
rect 26145 4165 26157 4168
rect 26191 4165 26203 4199
rect 26252 4196 26280 4236
rect 27430 4224 27436 4236
rect 27488 4224 27494 4276
rect 29454 4264 29460 4276
rect 27540 4236 29460 4264
rect 27540 4196 27568 4236
rect 29454 4224 29460 4236
rect 29512 4264 29518 4276
rect 31018 4264 31024 4276
rect 29512 4236 31024 4264
rect 29512 4224 29518 4236
rect 31018 4224 31024 4236
rect 31076 4224 31082 4276
rect 31113 4267 31171 4273
rect 31113 4233 31125 4267
rect 31159 4264 31171 4267
rect 32030 4264 32036 4276
rect 31159 4236 32036 4264
rect 31159 4233 31171 4236
rect 31113 4227 31171 4233
rect 28813 4199 28871 4205
rect 28813 4196 28825 4199
rect 26252 4168 27568 4196
rect 27632 4168 28825 4196
rect 26145 4159 26203 4165
rect 25464 4100 25728 4128
rect 25464 4088 25470 4100
rect 25774 4088 25780 4140
rect 25832 4128 25838 4140
rect 25869 4131 25927 4137
rect 25869 4128 25881 4131
rect 25832 4100 25881 4128
rect 25832 4088 25838 4100
rect 25869 4097 25881 4100
rect 25915 4097 25927 4131
rect 27632 4128 27660 4168
rect 28813 4165 28825 4168
rect 28859 4165 28871 4199
rect 28813 4159 28871 4165
rect 29362 4156 29368 4208
rect 29420 4196 29426 4208
rect 30282 4196 30288 4208
rect 29420 4168 30288 4196
rect 29420 4156 29426 4168
rect 30282 4156 30288 4168
rect 30340 4156 30346 4208
rect 28997 4131 29055 4137
rect 28997 4128 29009 4131
rect 25869 4091 25927 4097
rect 26252 4100 27660 4128
rect 27724 4100 29009 4128
rect 24670 4060 24676 4072
rect 24583 4032 24676 4060
rect 24670 4020 24676 4032
rect 24728 4020 24734 4072
rect 24762 4020 24768 4072
rect 24820 4060 24826 4072
rect 24857 4063 24915 4069
rect 24857 4060 24869 4063
rect 24820 4032 24869 4060
rect 24820 4020 24826 4032
rect 24857 4029 24869 4032
rect 24903 4060 24915 4063
rect 26252 4060 26280 4100
rect 24903 4032 26280 4060
rect 24903 4029 24915 4032
rect 24857 4023 24915 4029
rect 26326 4020 26332 4072
rect 26384 4060 26390 4072
rect 26789 4063 26847 4069
rect 26384 4032 26429 4060
rect 26384 4020 26390 4032
rect 26789 4029 26801 4063
rect 26835 4060 26847 4063
rect 27246 4060 27252 4072
rect 26835 4032 27252 4060
rect 26835 4029 26847 4032
rect 26789 4023 26847 4029
rect 27246 4020 27252 4032
rect 27304 4020 27310 4072
rect 27614 4020 27620 4072
rect 27672 4060 27678 4072
rect 27724 4069 27752 4100
rect 28997 4097 29009 4100
rect 29043 4097 29055 4131
rect 28997 4091 29055 4097
rect 29638 4088 29644 4140
rect 29696 4128 29702 4140
rect 29733 4131 29791 4137
rect 29733 4128 29745 4131
rect 29696 4100 29745 4128
rect 29696 4088 29702 4100
rect 29733 4097 29745 4100
rect 29779 4128 29791 4131
rect 30193 4131 30251 4137
rect 30193 4128 30205 4131
rect 29779 4100 30205 4128
rect 29779 4097 29791 4100
rect 29733 4091 29791 4097
rect 30193 4097 30205 4100
rect 30239 4128 30251 4131
rect 31128 4128 31156 4227
rect 32030 4224 32036 4236
rect 32088 4224 32094 4276
rect 32401 4267 32459 4273
rect 32401 4233 32413 4267
rect 32447 4264 32459 4267
rect 33962 4264 33968 4276
rect 32447 4236 33968 4264
rect 32447 4233 32459 4236
rect 32401 4227 32459 4233
rect 33962 4224 33968 4236
rect 34020 4224 34026 4276
rect 34238 4264 34244 4276
rect 34199 4236 34244 4264
rect 34238 4224 34244 4236
rect 34296 4224 34302 4276
rect 34514 4224 34520 4276
rect 34572 4264 34578 4276
rect 34609 4267 34667 4273
rect 34609 4264 34621 4267
rect 34572 4236 34621 4264
rect 34572 4224 34578 4236
rect 34609 4233 34621 4236
rect 34655 4233 34667 4267
rect 34609 4227 34667 4233
rect 35802 4224 35808 4276
rect 35860 4264 35866 4276
rect 36262 4264 36268 4276
rect 35860 4236 36268 4264
rect 35860 4224 35866 4236
rect 36262 4224 36268 4236
rect 36320 4264 36326 4276
rect 37093 4267 37151 4273
rect 37093 4264 37105 4267
rect 36320 4236 37105 4264
rect 36320 4224 36326 4236
rect 37093 4233 37105 4236
rect 37139 4233 37151 4267
rect 37093 4227 37151 4233
rect 38841 4267 38899 4273
rect 38841 4233 38853 4267
rect 38887 4264 38899 4267
rect 39022 4264 39028 4276
rect 38887 4236 39028 4264
rect 38887 4233 38899 4236
rect 38841 4227 38899 4233
rect 39022 4224 39028 4236
rect 39080 4224 39086 4276
rect 40310 4264 40316 4276
rect 40271 4236 40316 4264
rect 40310 4224 40316 4236
rect 40368 4224 40374 4276
rect 40402 4224 40408 4276
rect 40460 4264 40466 4276
rect 40589 4267 40647 4273
rect 40589 4264 40601 4267
rect 40460 4236 40601 4264
rect 40460 4224 40466 4236
rect 40589 4233 40601 4236
rect 40635 4233 40647 4267
rect 40589 4227 40647 4233
rect 41966 4224 41972 4276
rect 42024 4264 42030 4276
rect 42024 4236 44128 4264
rect 42024 4224 42030 4236
rect 31294 4156 31300 4208
rect 31352 4196 31358 4208
rect 31481 4199 31539 4205
rect 31481 4196 31493 4199
rect 31352 4168 31493 4196
rect 31352 4156 31358 4168
rect 31481 4165 31493 4168
rect 31527 4196 31539 4199
rect 32585 4199 32643 4205
rect 31527 4168 32352 4196
rect 31527 4165 31539 4168
rect 31481 4159 31539 4165
rect 32214 4128 32220 4140
rect 30239 4100 31156 4128
rect 31772 4100 32220 4128
rect 30239 4097 30251 4100
rect 30193 4091 30251 4097
rect 27709 4063 27767 4069
rect 27709 4060 27721 4063
rect 27672 4032 27721 4060
rect 27672 4020 27678 4032
rect 27709 4029 27721 4032
rect 27755 4029 27767 4063
rect 27890 4060 27896 4072
rect 27851 4032 27896 4060
rect 27709 4023 27767 4029
rect 27890 4020 27896 4032
rect 27948 4020 27954 4072
rect 28166 4020 28172 4072
rect 28224 4060 28230 4072
rect 30006 4060 30012 4072
rect 28224 4032 30012 4060
rect 28224 4020 28230 4032
rect 30006 4020 30012 4032
rect 30064 4020 30070 4072
rect 30101 4063 30159 4069
rect 30101 4029 30113 4063
rect 30147 4060 30159 4063
rect 30285 4063 30343 4069
rect 30285 4060 30297 4063
rect 30147 4032 30297 4060
rect 30147 4029 30159 4032
rect 30101 4023 30159 4029
rect 30285 4029 30297 4032
rect 30331 4060 30343 4063
rect 30466 4060 30472 4072
rect 30331 4032 30472 4060
rect 30331 4029 30343 4032
rect 30285 4023 30343 4029
rect 30466 4020 30472 4032
rect 30524 4020 30530 4072
rect 30742 4060 30748 4072
rect 30703 4032 30748 4060
rect 30742 4020 30748 4032
rect 30800 4020 30806 4072
rect 31386 4020 31392 4072
rect 31444 4060 31450 4072
rect 31598 4063 31656 4069
rect 31598 4060 31610 4063
rect 31444 4032 31610 4060
rect 31444 4020 31450 4032
rect 31598 4029 31610 4032
rect 31644 4060 31656 4063
rect 31772 4060 31800 4100
rect 32214 4088 32220 4100
rect 32272 4088 32278 4140
rect 31644 4032 31800 4060
rect 32324 4060 32352 4168
rect 32585 4165 32597 4199
rect 32631 4196 32643 4199
rect 34422 4196 34428 4208
rect 32631 4168 34428 4196
rect 32631 4165 32643 4168
rect 32585 4159 32643 4165
rect 34422 4156 34428 4168
rect 34480 4196 34486 4208
rect 34885 4199 34943 4205
rect 34885 4196 34897 4199
rect 34480 4168 34897 4196
rect 34480 4156 34486 4168
rect 34885 4165 34897 4168
rect 34931 4196 34943 4199
rect 39758 4196 39764 4208
rect 34931 4168 39764 4196
rect 34931 4165 34943 4168
rect 34885 4159 34943 4165
rect 39758 4156 39764 4168
rect 39816 4156 39822 4208
rect 39850 4156 39856 4208
rect 39908 4196 39914 4208
rect 39945 4199 40003 4205
rect 39945 4196 39957 4199
rect 39908 4168 39957 4196
rect 39908 4156 39914 4168
rect 39945 4165 39957 4168
rect 39991 4196 40003 4199
rect 42245 4199 42303 4205
rect 42245 4196 42257 4199
rect 39991 4168 42257 4196
rect 39991 4165 40003 4168
rect 39945 4159 40003 4165
rect 42245 4165 42257 4168
rect 42291 4196 42303 4199
rect 42426 4196 42432 4208
rect 42291 4168 42432 4196
rect 42291 4165 42303 4168
rect 42245 4159 42303 4165
rect 42426 4156 42432 4168
rect 42484 4156 42490 4208
rect 43622 4196 43628 4208
rect 43535 4168 43628 4196
rect 43622 4156 43628 4168
rect 43680 4196 43686 4208
rect 43993 4199 44051 4205
rect 43993 4196 44005 4199
rect 43680 4168 44005 4196
rect 43680 4156 43686 4168
rect 43993 4165 44005 4168
rect 44039 4165 44051 4199
rect 44100 4196 44128 4236
rect 44174 4224 44180 4276
rect 44232 4264 44238 4276
rect 46750 4264 46756 4276
rect 44232 4236 46756 4264
rect 44232 4224 44238 4236
rect 46750 4224 46756 4236
rect 46808 4224 46814 4276
rect 47026 4224 47032 4276
rect 47084 4264 47090 4276
rect 47305 4267 47363 4273
rect 47305 4264 47317 4267
rect 47084 4236 47317 4264
rect 47084 4224 47090 4236
rect 47305 4233 47317 4236
rect 47351 4264 47363 4267
rect 47857 4267 47915 4273
rect 47857 4264 47869 4267
rect 47351 4236 47869 4264
rect 47351 4233 47363 4236
rect 47305 4227 47363 4233
rect 47857 4233 47869 4236
rect 47903 4233 47915 4267
rect 47857 4227 47915 4233
rect 47946 4224 47952 4276
rect 48004 4264 48010 4276
rect 58345 4267 58403 4273
rect 48004 4236 55444 4264
rect 48004 4224 48010 4236
rect 49142 4196 49148 4208
rect 44100 4168 49148 4196
rect 43993 4159 44051 4165
rect 49142 4156 49148 4168
rect 49200 4196 49206 4208
rect 52546 4196 52552 4208
rect 49200 4168 52552 4196
rect 49200 4156 49206 4168
rect 52546 4156 52552 4168
rect 52604 4156 52610 4208
rect 53009 4199 53067 4205
rect 53009 4165 53021 4199
rect 53055 4196 53067 4199
rect 53282 4196 53288 4208
rect 53055 4168 53288 4196
rect 53055 4165 53067 4168
rect 53009 4159 53067 4165
rect 53282 4156 53288 4168
rect 53340 4196 53346 4208
rect 54478 4196 54484 4208
rect 53340 4168 54484 4196
rect 53340 4156 53346 4168
rect 54478 4156 54484 4168
rect 54536 4156 54542 4208
rect 55030 4156 55036 4208
rect 55088 4196 55094 4208
rect 55088 4168 55352 4196
rect 55088 4156 55094 4168
rect 33229 4131 33287 4137
rect 33229 4128 33241 4131
rect 32692 4100 33241 4128
rect 32582 4060 32588 4072
rect 32324 4032 32588 4060
rect 31644 4029 31656 4032
rect 31598 4023 31656 4029
rect 32582 4020 32588 4032
rect 32640 4020 32646 4072
rect 32692 4069 32720 4100
rect 33229 4097 33241 4100
rect 33275 4128 33287 4131
rect 36078 4128 36084 4140
rect 33275 4100 36084 4128
rect 33275 4097 33287 4100
rect 33229 4091 33287 4097
rect 36078 4088 36084 4100
rect 36136 4088 36142 4140
rect 37182 4088 37188 4140
rect 37240 4128 37246 4140
rect 37461 4131 37519 4137
rect 37461 4128 37473 4131
rect 37240 4100 37473 4128
rect 37240 4088 37246 4100
rect 37461 4097 37473 4100
rect 37507 4097 37519 4131
rect 37461 4091 37519 4097
rect 38289 4131 38347 4137
rect 38289 4097 38301 4131
rect 38335 4128 38347 4131
rect 38657 4131 38715 4137
rect 38657 4128 38669 4131
rect 38335 4100 38669 4128
rect 38335 4097 38347 4100
rect 38289 4091 38347 4097
rect 38657 4097 38669 4100
rect 38703 4128 38715 4131
rect 39574 4128 39580 4140
rect 38703 4100 39252 4128
rect 39535 4100 39580 4128
rect 38703 4097 38715 4100
rect 38657 4091 38715 4097
rect 32677 4063 32735 4069
rect 32677 4029 32689 4063
rect 32723 4029 32735 4063
rect 33502 4060 33508 4072
rect 33463 4032 33508 4060
rect 32677 4023 32735 4029
rect 33502 4020 33508 4032
rect 33560 4020 33566 4072
rect 33689 4063 33747 4069
rect 33689 4029 33701 4063
rect 33735 4060 33747 4063
rect 34238 4060 34244 4072
rect 33735 4032 34244 4060
rect 33735 4029 33747 4032
rect 33689 4023 33747 4029
rect 34238 4020 34244 4032
rect 34296 4020 34302 4072
rect 34514 4020 34520 4072
rect 34572 4060 34578 4072
rect 35345 4063 35403 4069
rect 35345 4060 35357 4063
rect 34572 4032 35357 4060
rect 34572 4020 34578 4032
rect 35345 4029 35357 4032
rect 35391 4029 35403 4063
rect 35986 4060 35992 4072
rect 35947 4032 35992 4060
rect 35345 4023 35403 4029
rect 35986 4020 35992 4032
rect 36044 4020 36050 4072
rect 36262 4060 36268 4072
rect 36223 4032 36268 4060
rect 36262 4020 36268 4032
rect 36320 4020 36326 4072
rect 36446 4020 36452 4072
rect 36504 4060 36510 4072
rect 36541 4063 36599 4069
rect 36541 4060 36553 4063
rect 36504 4032 36553 4060
rect 36504 4020 36510 4032
rect 36541 4029 36553 4032
rect 36587 4029 36599 4063
rect 36541 4023 36599 4029
rect 37645 4063 37703 4069
rect 37645 4029 37657 4063
rect 37691 4060 37703 4063
rect 37918 4060 37924 4072
rect 37691 4032 37924 4060
rect 37691 4029 37703 4032
rect 37645 4023 37703 4029
rect 37918 4020 37924 4032
rect 37976 4060 37982 4072
rect 38304 4060 38332 4091
rect 37976 4032 38332 4060
rect 37976 4020 37982 4032
rect 38930 4020 38936 4072
rect 38988 4060 38994 4072
rect 39117 4063 39175 4069
rect 39117 4060 39129 4063
rect 38988 4032 39129 4060
rect 38988 4020 38994 4032
rect 39117 4029 39129 4032
rect 39163 4029 39175 4063
rect 39224 4060 39252 4100
rect 39574 4088 39580 4100
rect 39632 4088 39638 4140
rect 43640 4128 43668 4156
rect 39684 4100 43668 4128
rect 39684 4060 39712 4100
rect 39224 4032 39712 4060
rect 40773 4063 40831 4069
rect 39117 4023 39175 4029
rect 40773 4029 40785 4063
rect 40819 4060 40831 4063
rect 40954 4060 40960 4072
rect 40819 4032 40960 4060
rect 40819 4029 40831 4032
rect 40773 4023 40831 4029
rect 40954 4020 40960 4032
rect 41012 4020 41018 4072
rect 41233 4063 41291 4069
rect 41233 4029 41245 4063
rect 41279 4060 41291 4063
rect 42058 4060 42064 4072
rect 41279 4032 41644 4060
rect 42019 4032 42064 4060
rect 41279 4029 41291 4032
rect 41233 4023 41291 4029
rect 22296 3964 24532 3992
rect 24688 3992 24716 4020
rect 24688 3964 25084 3992
rect 11195 3896 13032 3924
rect 11195 3893 11207 3896
rect 11149 3887 11207 3893
rect 13446 3884 13452 3936
rect 13504 3924 13510 3936
rect 15102 3924 15108 3936
rect 13504 3896 15108 3924
rect 13504 3884 13510 3896
rect 15102 3884 15108 3896
rect 15160 3924 15166 3936
rect 16482 3924 16488 3936
rect 15160 3896 16488 3924
rect 15160 3884 15166 3896
rect 16482 3884 16488 3896
rect 16540 3884 16546 3936
rect 16574 3884 16580 3936
rect 16632 3924 16638 3936
rect 22370 3924 22376 3936
rect 16632 3896 22376 3924
rect 16632 3884 16638 3896
rect 22370 3884 22376 3896
rect 22428 3884 22434 3936
rect 22646 3884 22652 3936
rect 22704 3924 22710 3936
rect 23017 3927 23075 3933
rect 23017 3924 23029 3927
rect 22704 3896 23029 3924
rect 22704 3884 22710 3896
rect 23017 3893 23029 3896
rect 23063 3893 23075 3927
rect 23382 3924 23388 3936
rect 23343 3896 23388 3924
rect 23017 3887 23075 3893
rect 23382 3884 23388 3896
rect 23440 3884 23446 3936
rect 24946 3924 24952 3936
rect 24907 3896 24952 3924
rect 24946 3884 24952 3896
rect 25004 3884 25010 3936
rect 25056 3924 25084 3964
rect 25130 3952 25136 4004
rect 25188 3992 25194 4004
rect 26510 3992 26516 4004
rect 25188 3964 26516 3992
rect 25188 3952 25194 3964
rect 26510 3952 26516 3964
rect 26568 3952 26574 4004
rect 27798 3992 27804 4004
rect 27759 3964 27804 3992
rect 27798 3952 27804 3964
rect 27856 3952 27862 4004
rect 28350 3992 28356 4004
rect 28311 3964 28356 3992
rect 28350 3952 28356 3964
rect 28408 3952 28414 4004
rect 28813 3995 28871 4001
rect 28460 3964 28764 3992
rect 25501 3927 25559 3933
rect 25501 3924 25513 3927
rect 25056 3896 25513 3924
rect 25501 3893 25513 3896
rect 25547 3893 25559 3927
rect 25501 3887 25559 3893
rect 25590 3884 25596 3936
rect 25648 3924 25654 3936
rect 27154 3924 27160 3936
rect 25648 3896 27160 3924
rect 25648 3884 25654 3896
rect 27154 3884 27160 3896
rect 27212 3924 27218 3936
rect 28460 3924 28488 3964
rect 28626 3924 28632 3936
rect 27212 3896 28488 3924
rect 28587 3896 28632 3924
rect 27212 3884 27218 3896
rect 28626 3884 28632 3896
rect 28684 3884 28690 3936
rect 28736 3924 28764 3964
rect 28813 3961 28825 3995
rect 28859 3992 28871 3995
rect 30190 3992 30196 4004
rect 28859 3964 30196 3992
rect 28859 3961 28871 3964
rect 28813 3955 28871 3961
rect 30190 3952 30196 3964
rect 30248 3952 30254 4004
rect 31938 3952 31944 4004
rect 31996 3992 32002 4004
rect 34974 3992 34980 4004
rect 31996 3964 34980 3992
rect 31996 3952 32002 3964
rect 30650 3924 30656 3936
rect 28736 3896 30656 3924
rect 30650 3884 30656 3896
rect 30708 3884 30714 3936
rect 31478 3884 31484 3936
rect 31536 3924 31542 3936
rect 31757 3927 31815 3933
rect 31757 3924 31769 3927
rect 31536 3896 31769 3924
rect 31536 3884 31542 3896
rect 31757 3893 31769 3896
rect 31803 3924 31815 3927
rect 32401 3927 32459 3933
rect 32401 3924 32413 3927
rect 31803 3896 32413 3924
rect 31803 3893 31815 3896
rect 31757 3887 31815 3893
rect 32401 3893 32413 3896
rect 32447 3893 32459 3927
rect 32766 3924 32772 3936
rect 32727 3896 32772 3924
rect 32401 3887 32459 3893
rect 32766 3884 32772 3896
rect 32824 3884 32830 3936
rect 33888 3933 33916 3964
rect 34974 3952 34980 3964
rect 35032 3952 35038 4004
rect 35253 3995 35311 4001
rect 35253 3961 35265 3995
rect 35299 3992 35311 3995
rect 37734 3992 37740 4004
rect 35299 3964 37740 3992
rect 35299 3961 35311 3964
rect 35253 3955 35311 3961
rect 37734 3952 37740 3964
rect 37792 3952 37798 4004
rect 38746 3952 38752 4004
rect 38804 3992 38810 4004
rect 39025 3995 39083 4001
rect 39025 3992 39037 3995
rect 38804 3964 39037 3992
rect 38804 3952 38810 3964
rect 39025 3961 39037 3964
rect 39071 3961 39083 3995
rect 39025 3955 39083 3961
rect 33873 3927 33931 3933
rect 33873 3893 33885 3927
rect 33919 3893 33931 3927
rect 34992 3924 35020 3952
rect 41616 3936 41644 4032
rect 42058 4020 42064 4032
rect 42116 4060 42122 4072
rect 42613 4063 42671 4069
rect 42613 4060 42625 4063
rect 42116 4032 42625 4060
rect 42116 4020 42122 4032
rect 42613 4029 42625 4032
rect 42659 4029 42671 4063
rect 43640 4060 43668 4100
rect 43717 4131 43775 4137
rect 43717 4097 43729 4131
rect 43763 4128 43775 4131
rect 45646 4128 45652 4140
rect 43763 4100 45652 4128
rect 43763 4097 43775 4100
rect 43717 4091 43775 4097
rect 45646 4088 45652 4100
rect 45704 4088 45710 4140
rect 47305 4131 47363 4137
rect 47305 4128 47317 4131
rect 47182 4100 47317 4128
rect 44729 4063 44787 4069
rect 44729 4060 44741 4063
rect 43640 4032 44741 4060
rect 42613 4023 42671 4029
rect 44729 4029 44741 4032
rect 44775 4029 44787 4063
rect 44729 4023 44787 4029
rect 45005 4063 45063 4069
rect 45005 4029 45017 4063
rect 45051 4029 45063 4063
rect 45005 4023 45063 4029
rect 45189 4063 45247 4069
rect 45189 4029 45201 4063
rect 45235 4060 45247 4063
rect 46201 4063 46259 4069
rect 45235 4032 45269 4060
rect 45235 4029 45247 4032
rect 45189 4023 45247 4029
rect 46201 4029 46213 4063
rect 46247 4060 46259 4063
rect 46934 4060 46940 4072
rect 46247 4032 46940 4060
rect 46247 4029 46259 4032
rect 46201 4023 46259 4029
rect 44174 3992 44180 4004
rect 44135 3964 44180 3992
rect 44174 3952 44180 3964
rect 44232 3952 44238 4004
rect 35986 3924 35992 3936
rect 34992 3896 35992 3924
rect 33873 3887 33931 3893
rect 35986 3884 35992 3896
rect 36044 3884 36050 3936
rect 36170 3884 36176 3936
rect 36228 3924 36234 3936
rect 37829 3927 37887 3933
rect 37829 3924 37841 3927
rect 36228 3896 37841 3924
rect 36228 3884 36234 3896
rect 37829 3893 37841 3896
rect 37875 3893 37887 3927
rect 41598 3924 41604 3936
rect 41559 3896 41604 3924
rect 37829 3887 37887 3893
rect 41598 3884 41604 3896
rect 41656 3884 41662 3936
rect 41969 3927 42027 3933
rect 41969 3893 41981 3927
rect 42015 3924 42027 3927
rect 42150 3924 42156 3936
rect 42015 3896 42156 3924
rect 42015 3893 42027 3896
rect 41969 3887 42027 3893
rect 42150 3884 42156 3896
rect 42208 3884 42214 3936
rect 43349 3927 43407 3933
rect 43349 3893 43361 3927
rect 43395 3924 43407 3927
rect 44726 3924 44732 3936
rect 43395 3896 44732 3924
rect 43395 3893 43407 3896
rect 43349 3887 43407 3893
rect 44726 3884 44732 3896
rect 44784 3884 44790 3936
rect 44818 3884 44824 3936
rect 44876 3924 44882 3936
rect 45020 3924 45048 4023
rect 45094 3952 45100 4004
rect 45152 3992 45158 4004
rect 45204 3992 45232 4023
rect 46934 4020 46940 4032
rect 46992 4020 46998 4072
rect 47026 4020 47032 4072
rect 47084 4060 47090 4072
rect 47182 4069 47210 4100
rect 47305 4097 47317 4100
rect 47351 4097 47363 4131
rect 47305 4091 47363 4097
rect 47946 4088 47952 4140
rect 48004 4128 48010 4140
rect 48041 4131 48099 4137
rect 48041 4128 48053 4131
rect 48004 4100 48053 4128
rect 48004 4088 48010 4100
rect 48041 4097 48053 4100
rect 48087 4097 48099 4131
rect 48041 4091 48099 4097
rect 49234 4088 49240 4140
rect 49292 4128 49298 4140
rect 50614 4128 50620 4140
rect 49292 4100 50620 4128
rect 49292 4088 49298 4100
rect 50614 4088 50620 4100
rect 50672 4088 50678 4140
rect 52178 4128 52184 4140
rect 51736 4100 52184 4128
rect 51736 4072 51764 4100
rect 52178 4088 52184 4100
rect 52236 4088 52242 4140
rect 52273 4131 52331 4137
rect 52273 4097 52285 4131
rect 52319 4128 52331 4131
rect 52822 4128 52828 4140
rect 52319 4100 52828 4128
rect 52319 4097 52331 4100
rect 52273 4091 52331 4097
rect 52822 4088 52828 4100
rect 52880 4088 52886 4140
rect 53208 4100 54064 4128
rect 47167 4063 47225 4069
rect 47084 4032 47129 4060
rect 47084 4020 47090 4032
rect 47167 4029 47179 4063
rect 47213 4029 47225 4063
rect 47489 4063 47547 4069
rect 47489 4060 47501 4063
rect 47167 4023 47225 4029
rect 47320 4032 47501 4060
rect 45465 3995 45523 4001
rect 45465 3992 45477 3995
rect 45152 3964 45477 3992
rect 45152 3952 45158 3964
rect 45465 3961 45477 3964
rect 45511 3961 45523 3995
rect 46290 3992 46296 4004
rect 46251 3964 46296 3992
rect 45465 3955 45523 3961
rect 46290 3952 46296 3964
rect 46348 3952 46354 4004
rect 47044 3992 47072 4020
rect 47320 3992 47348 4032
rect 47489 4029 47501 4032
rect 47535 4060 47547 4063
rect 48406 4060 48412 4072
rect 47535 4032 48412 4060
rect 47535 4029 47547 4032
rect 47489 4023 47547 4029
rect 48406 4020 48412 4032
rect 48464 4020 48470 4072
rect 48498 4020 48504 4072
rect 48556 4060 48562 4072
rect 48593 4063 48651 4069
rect 48593 4060 48605 4063
rect 48556 4032 48605 4060
rect 48556 4020 48562 4032
rect 48593 4029 48605 4032
rect 48639 4029 48651 4063
rect 48593 4023 48651 4029
rect 48682 4020 48688 4072
rect 48740 4060 48746 4072
rect 48869 4063 48927 4069
rect 48869 4060 48881 4063
rect 48740 4032 48881 4060
rect 48740 4020 48746 4032
rect 48869 4029 48881 4032
rect 48915 4029 48927 4063
rect 48869 4023 48927 4029
rect 49053 4063 49111 4069
rect 49053 4029 49065 4063
rect 49099 4060 49111 4063
rect 49145 4063 49203 4069
rect 49145 4060 49157 4063
rect 49099 4032 49157 4060
rect 49099 4029 49111 4032
rect 49053 4023 49111 4029
rect 49145 4029 49157 4032
rect 49191 4029 49203 4063
rect 49145 4023 49203 4029
rect 49786 4020 49792 4072
rect 49844 4060 49850 4072
rect 50065 4063 50123 4069
rect 50065 4060 50077 4063
rect 49844 4032 50077 4060
rect 49844 4020 49850 4032
rect 50065 4029 50077 4032
rect 50111 4060 50123 4063
rect 50709 4063 50767 4069
rect 50709 4060 50721 4063
rect 50111 4032 50721 4060
rect 50111 4029 50123 4032
rect 50065 4023 50123 4029
rect 50709 4029 50721 4032
rect 50755 4029 50767 4063
rect 50709 4023 50767 4029
rect 50893 4063 50951 4069
rect 50893 4029 50905 4063
rect 50939 4060 50951 4063
rect 51718 4060 51724 4072
rect 50939 4032 51488 4060
rect 51679 4032 51724 4060
rect 50939 4029 50951 4032
rect 50893 4023 50951 4029
rect 49697 3995 49755 4001
rect 49697 3992 49709 3995
rect 47044 3964 47348 3992
rect 47412 3964 49709 3992
rect 45925 3927 45983 3933
rect 45925 3924 45937 3927
rect 44876 3896 45937 3924
rect 44876 3884 44882 3896
rect 45925 3893 45937 3896
rect 45971 3924 45983 3927
rect 46014 3924 46020 3936
rect 45971 3896 46020 3924
rect 45971 3893 45983 3896
rect 45925 3887 45983 3893
rect 46014 3884 46020 3896
rect 46072 3884 46078 3936
rect 46198 3884 46204 3936
rect 46256 3924 46262 3936
rect 47412 3924 47440 3964
rect 49697 3961 49709 3964
rect 49743 3992 49755 3995
rect 49881 3995 49939 4001
rect 49881 3992 49893 3995
rect 49743 3964 49893 3992
rect 49743 3961 49755 3964
rect 49697 3955 49755 3961
rect 49881 3961 49893 3964
rect 49927 3961 49939 3995
rect 49881 3955 49939 3961
rect 46256 3896 47440 3924
rect 46256 3884 46262 3896
rect 47486 3884 47492 3936
rect 47544 3924 47550 3936
rect 48314 3924 48320 3936
rect 47544 3896 48320 3924
rect 47544 3884 47550 3896
rect 48314 3884 48320 3896
rect 48372 3884 48378 3936
rect 48866 3884 48872 3936
rect 48924 3924 48930 3936
rect 49329 3927 49387 3933
rect 49329 3924 49341 3927
rect 48924 3896 49341 3924
rect 48924 3884 48930 3896
rect 49329 3893 49341 3896
rect 49375 3893 49387 3927
rect 49329 3887 49387 3893
rect 50062 3884 50068 3936
rect 50120 3924 50126 3936
rect 50157 3927 50215 3933
rect 50157 3924 50169 3927
rect 50120 3896 50169 3924
rect 50120 3884 50126 3896
rect 50157 3893 50169 3896
rect 50203 3893 50215 3927
rect 50157 3887 50215 3893
rect 50246 3884 50252 3936
rect 50304 3924 50310 3936
rect 50893 3927 50951 3933
rect 50893 3924 50905 3927
rect 50304 3896 50905 3924
rect 50304 3884 50310 3896
rect 50893 3893 50905 3896
rect 50939 3893 50951 3927
rect 50893 3887 50951 3893
rect 51074 3884 51080 3936
rect 51132 3924 51138 3936
rect 51460 3924 51488 4032
rect 51718 4020 51724 4032
rect 51776 4020 51782 4072
rect 51810 4020 51816 4072
rect 51868 4060 51874 4072
rect 51868 4032 51913 4060
rect 51868 4020 51874 4032
rect 52546 4020 52552 4072
rect 52604 4060 52610 4072
rect 53208 4060 53236 4100
rect 53374 4060 53380 4072
rect 52604 4032 53236 4060
rect 53335 4032 53380 4060
rect 52604 4020 52610 4032
rect 53374 4020 53380 4032
rect 53432 4020 53438 4072
rect 53469 4063 53527 4069
rect 53469 4029 53481 4063
rect 53515 4060 53527 4063
rect 53558 4060 53564 4072
rect 53515 4032 53564 4060
rect 53515 4029 53527 4032
rect 53469 4023 53527 4029
rect 53558 4020 53564 4032
rect 53616 4020 53622 4072
rect 53650 4020 53656 4072
rect 53708 4060 53714 4072
rect 54036 4060 54064 4100
rect 54110 4088 54116 4140
rect 54168 4128 54174 4140
rect 54205 4131 54263 4137
rect 54205 4128 54217 4131
rect 54168 4100 54217 4128
rect 54168 4088 54174 4100
rect 54205 4097 54217 4100
rect 54251 4128 54263 4131
rect 54754 4128 54760 4140
rect 54251 4100 54760 4128
rect 54251 4097 54263 4100
rect 54205 4091 54263 4097
rect 54754 4088 54760 4100
rect 54812 4088 54818 4140
rect 55214 4128 55220 4140
rect 54864 4100 55220 4128
rect 54864 4069 54892 4100
rect 55214 4088 55220 4100
rect 55272 4088 55278 4140
rect 54849 4063 54907 4069
rect 53708 4032 53753 4060
rect 54036 4032 54800 4060
rect 53708 4020 53714 4032
rect 51537 3995 51595 4001
rect 51537 3961 51549 3995
rect 51583 3992 51595 3995
rect 51994 3992 52000 4004
rect 51583 3964 52000 3992
rect 51583 3961 51595 3964
rect 51537 3955 51595 3961
rect 51994 3952 52000 3964
rect 52052 3992 52058 4004
rect 52641 3995 52699 4001
rect 52641 3992 52653 3995
rect 52052 3964 52653 3992
rect 52052 3952 52058 3964
rect 52641 3961 52653 3964
rect 52687 3992 52699 3995
rect 53926 3992 53932 4004
rect 52687 3964 53932 3992
rect 52687 3961 52699 3964
rect 52641 3955 52699 3961
rect 53926 3952 53932 3964
rect 53984 3952 53990 4004
rect 54662 3992 54668 4004
rect 54623 3964 54668 3992
rect 54662 3952 54668 3964
rect 54720 3952 54726 4004
rect 54772 3992 54800 4032
rect 54849 4029 54861 4063
rect 54895 4029 54907 4063
rect 54849 4023 54907 4029
rect 54941 4063 54999 4069
rect 54941 4029 54953 4063
rect 54987 4060 54999 4063
rect 55122 4060 55128 4072
rect 54987 4032 55128 4060
rect 54987 4029 54999 4032
rect 54941 4023 54999 4029
rect 55122 4020 55128 4032
rect 55180 4020 55186 4072
rect 55324 4060 55352 4168
rect 55416 4137 55444 4236
rect 58345 4233 58357 4267
rect 58391 4264 58403 4267
rect 58713 4267 58771 4273
rect 58713 4264 58725 4267
rect 58391 4236 58725 4264
rect 58391 4233 58403 4236
rect 58345 4227 58403 4233
rect 58713 4233 58725 4236
rect 58759 4264 58771 4267
rect 59262 4264 59268 4276
rect 58759 4236 59268 4264
rect 58759 4233 58771 4236
rect 58713 4227 58771 4233
rect 56134 4156 56140 4208
rect 56192 4196 56198 4208
rect 56192 4168 56548 4196
rect 56192 4156 56198 4168
rect 55401 4131 55459 4137
rect 55401 4097 55413 4131
rect 55447 4097 55459 4131
rect 56520 4128 56548 4168
rect 57425 4131 57483 4137
rect 57425 4128 57437 4131
rect 56520 4100 57437 4128
rect 55401 4091 55459 4097
rect 57425 4097 57437 4100
rect 57471 4128 57483 4131
rect 58360 4128 58388 4227
rect 59262 4224 59268 4236
rect 59320 4264 59326 4276
rect 61105 4267 61163 4273
rect 59320 4236 59768 4264
rect 59320 4224 59326 4236
rect 59740 4196 59768 4236
rect 61105 4233 61117 4267
rect 61151 4264 61163 4267
rect 61194 4264 61200 4276
rect 61151 4236 61200 4264
rect 61151 4233 61163 4236
rect 61105 4227 61163 4233
rect 61194 4224 61200 4236
rect 61252 4224 61258 4276
rect 61473 4199 61531 4205
rect 61473 4196 61485 4199
rect 59740 4168 61485 4196
rect 61473 4165 61485 4168
rect 61519 4165 61531 4199
rect 61473 4159 61531 4165
rect 57471 4100 58388 4128
rect 59081 4131 59139 4137
rect 57471 4097 57483 4100
rect 57425 4091 57483 4097
rect 59081 4097 59093 4131
rect 59127 4128 59139 4131
rect 59538 4128 59544 4140
rect 59127 4100 59544 4128
rect 59127 4097 59139 4100
rect 59081 4091 59139 4097
rect 59538 4088 59544 4100
rect 59596 4088 59602 4140
rect 61010 4088 61016 4140
rect 61068 4128 61074 4140
rect 61068 4100 61608 4128
rect 61068 4088 61074 4100
rect 55677 4063 55735 4069
rect 55677 4060 55689 4063
rect 55324 4032 55689 4060
rect 55677 4029 55689 4032
rect 55723 4060 55735 4063
rect 56413 4063 56471 4069
rect 56413 4060 56425 4063
rect 55723 4032 56425 4060
rect 55723 4029 55735 4032
rect 55677 4023 55735 4029
rect 56413 4029 56425 4032
rect 56459 4029 56471 4063
rect 57517 4063 57575 4069
rect 57517 4060 57529 4063
rect 56413 4023 56471 4029
rect 57072 4032 57529 4060
rect 54772 3964 54984 3992
rect 53282 3924 53288 3936
rect 51132 3896 51177 3924
rect 51460 3896 53288 3924
rect 51132 3884 51138 3896
rect 53282 3884 53288 3896
rect 53340 3884 53346 3936
rect 53374 3884 53380 3936
rect 53432 3924 53438 3936
rect 54846 3924 54852 3936
rect 53432 3896 54852 3924
rect 53432 3884 53438 3896
rect 54846 3884 54852 3896
rect 54904 3884 54910 3936
rect 54956 3924 54984 3964
rect 55030 3952 55036 4004
rect 55088 3992 55094 4004
rect 55088 3964 55133 3992
rect 55088 3952 55094 3964
rect 55214 3952 55220 4004
rect 55272 3992 55278 4004
rect 57072 4001 57100 4032
rect 57517 4029 57529 4032
rect 57563 4029 57575 4063
rect 57517 4023 57575 4029
rect 58066 4020 58072 4072
rect 58124 4060 58130 4072
rect 58434 4060 58440 4072
rect 58124 4032 58440 4060
rect 58124 4020 58130 4032
rect 58434 4020 58440 4032
rect 58492 4060 58498 4072
rect 58805 4063 58863 4069
rect 58805 4060 58817 4063
rect 58492 4032 58817 4060
rect 58492 4020 58498 4032
rect 58805 4029 58817 4032
rect 58851 4029 58863 4063
rect 58805 4023 58863 4029
rect 61289 4063 61347 4069
rect 61289 4029 61301 4063
rect 61335 4060 61347 4063
rect 61470 4060 61476 4072
rect 61335 4032 61476 4060
rect 61335 4029 61347 4032
rect 61289 4023 61347 4029
rect 57057 3995 57115 4001
rect 57057 3992 57069 3995
rect 55272 3964 57069 3992
rect 55272 3952 55278 3964
rect 57057 3961 57069 3964
rect 57103 3961 57115 3995
rect 57057 3955 57115 3961
rect 57606 3952 57612 4004
rect 57664 3992 57670 4004
rect 57977 3995 58035 4001
rect 57977 3992 57989 3995
rect 57664 3964 57989 3992
rect 57664 3952 57670 3964
rect 57977 3961 57989 3964
rect 58023 3961 58035 3995
rect 57977 3955 58035 3961
rect 55582 3924 55588 3936
rect 54956 3896 55588 3924
rect 55582 3884 55588 3896
rect 55640 3884 55646 3936
rect 55674 3884 55680 3936
rect 55732 3924 55738 3936
rect 56042 3924 56048 3936
rect 55732 3896 56048 3924
rect 55732 3884 55738 3896
rect 56042 3884 56048 3896
rect 56100 3884 56106 3936
rect 57330 3884 57336 3936
rect 57388 3924 57394 3936
rect 60185 3927 60243 3933
rect 60185 3924 60197 3927
rect 57388 3896 60197 3924
rect 57388 3884 57394 3896
rect 60185 3893 60197 3896
rect 60231 3924 60243 3927
rect 61304 3924 61332 4023
rect 61470 4020 61476 4032
rect 61528 4020 61534 4072
rect 61580 4060 61608 4100
rect 61746 4088 61752 4140
rect 61804 4128 61810 4140
rect 62209 4131 62267 4137
rect 62209 4128 62221 4131
rect 61804 4100 62221 4128
rect 61804 4088 61810 4100
rect 62209 4097 62221 4100
rect 62255 4097 62267 4131
rect 62209 4091 62267 4097
rect 61841 4063 61899 4069
rect 61841 4060 61853 4063
rect 61580 4032 61853 4060
rect 61841 4029 61853 4032
rect 61887 4029 61899 4063
rect 61841 4023 61899 4029
rect 60231 3896 61332 3924
rect 60231 3893 60243 3896
rect 60185 3887 60243 3893
rect 1104 3834 63480 3856
rect 1104 3782 21774 3834
rect 21826 3782 21838 3834
rect 21890 3782 21902 3834
rect 21954 3782 21966 3834
rect 22018 3782 42566 3834
rect 42618 3782 42630 3834
rect 42682 3782 42694 3834
rect 42746 3782 42758 3834
rect 42810 3782 63480 3834
rect 1104 3760 63480 3782
rect 3326 3680 3332 3732
rect 3384 3720 3390 3732
rect 4157 3723 4215 3729
rect 4157 3720 4169 3723
rect 3384 3692 4169 3720
rect 3384 3680 3390 3692
rect 4157 3689 4169 3692
rect 4203 3689 4215 3723
rect 4157 3683 4215 3689
rect 4798 3680 4804 3732
rect 4856 3720 4862 3732
rect 4893 3723 4951 3729
rect 4893 3720 4905 3723
rect 4856 3692 4905 3720
rect 4856 3680 4862 3692
rect 4893 3689 4905 3692
rect 4939 3689 4951 3723
rect 4893 3683 4951 3689
rect 5718 3680 5724 3732
rect 5776 3720 5782 3732
rect 7466 3720 7472 3732
rect 5776 3692 7472 3720
rect 5776 3680 5782 3692
rect 7466 3680 7472 3692
rect 7524 3720 7530 3732
rect 7834 3720 7840 3732
rect 7524 3692 7840 3720
rect 7524 3680 7530 3692
rect 7834 3680 7840 3692
rect 7892 3680 7898 3732
rect 8570 3680 8576 3732
rect 8628 3720 8634 3732
rect 9401 3723 9459 3729
rect 9401 3720 9413 3723
rect 8628 3692 9413 3720
rect 8628 3680 8634 3692
rect 9401 3689 9413 3692
rect 9447 3720 9459 3723
rect 9582 3720 9588 3732
rect 9447 3692 9588 3720
rect 9447 3689 9459 3692
rect 9401 3683 9459 3689
rect 9582 3680 9588 3692
rect 9640 3680 9646 3732
rect 9858 3680 9864 3732
rect 9916 3720 9922 3732
rect 14090 3720 14096 3732
rect 9916 3692 13952 3720
rect 14051 3692 14096 3720
rect 9916 3680 9922 3692
rect 2222 3612 2228 3664
rect 2280 3652 2286 3664
rect 2280 3624 4108 3652
rect 2280 3612 2286 3624
rect 2685 3587 2743 3593
rect 2685 3553 2697 3587
rect 2731 3584 2743 3587
rect 2866 3584 2872 3596
rect 2731 3556 2872 3584
rect 2731 3553 2743 3556
rect 2685 3547 2743 3553
rect 2866 3544 2872 3556
rect 2924 3584 2930 3596
rect 3418 3584 3424 3596
rect 2924 3556 3424 3584
rect 2924 3544 2930 3556
rect 3418 3544 3424 3556
rect 3476 3544 3482 3596
rect 3513 3587 3571 3593
rect 3513 3553 3525 3587
rect 3559 3584 3571 3587
rect 3786 3584 3792 3596
rect 3559 3556 3792 3584
rect 3559 3553 3571 3556
rect 3513 3547 3571 3553
rect 3786 3544 3792 3556
rect 3844 3544 3850 3596
rect 4080 3593 4108 3624
rect 7926 3612 7932 3664
rect 7984 3652 7990 3664
rect 8665 3655 8723 3661
rect 8665 3652 8677 3655
rect 7984 3624 8677 3652
rect 7984 3612 7990 3624
rect 8665 3621 8677 3624
rect 8711 3621 8723 3655
rect 8665 3615 8723 3621
rect 8938 3612 8944 3664
rect 8996 3652 9002 3664
rect 11977 3655 12035 3661
rect 8996 3624 11652 3652
rect 8996 3612 9002 3624
rect 4065 3587 4123 3593
rect 4065 3553 4077 3587
rect 4111 3584 4123 3587
rect 4525 3587 4583 3593
rect 4525 3584 4537 3587
rect 4111 3556 4537 3584
rect 4111 3553 4123 3556
rect 4065 3547 4123 3553
rect 4525 3553 4537 3556
rect 4571 3553 4583 3587
rect 5902 3584 5908 3596
rect 5863 3556 5908 3584
rect 4525 3547 4583 3553
rect 5902 3544 5908 3556
rect 5960 3544 5966 3596
rect 6273 3587 6331 3593
rect 6273 3553 6285 3587
rect 6319 3584 6331 3587
rect 6638 3584 6644 3596
rect 6319 3556 6644 3584
rect 6319 3553 6331 3556
rect 6273 3547 6331 3553
rect 6638 3544 6644 3556
rect 6696 3544 6702 3596
rect 7561 3587 7619 3593
rect 7561 3553 7573 3587
rect 7607 3584 7619 3587
rect 7742 3584 7748 3596
rect 7607 3556 7748 3584
rect 7607 3553 7619 3556
rect 7561 3547 7619 3553
rect 7742 3544 7748 3556
rect 7800 3544 7806 3596
rect 8021 3587 8079 3593
rect 8021 3553 8033 3587
rect 8067 3584 8079 3587
rect 8294 3584 8300 3596
rect 8067 3556 8300 3584
rect 8067 3553 8079 3556
rect 8021 3547 8079 3553
rect 8294 3544 8300 3556
rect 8352 3544 8358 3596
rect 10134 3584 10140 3596
rect 10095 3556 10140 3584
rect 10134 3544 10140 3556
rect 10192 3544 10198 3596
rect 11057 3587 11115 3593
rect 11057 3553 11069 3587
rect 11103 3553 11115 3587
rect 11624 3584 11652 3624
rect 11977 3621 11989 3655
rect 12023 3652 12035 3655
rect 13924 3652 13952 3692
rect 14090 3680 14096 3692
rect 14148 3680 14154 3732
rect 14737 3723 14795 3729
rect 14737 3689 14749 3723
rect 14783 3720 14795 3723
rect 16574 3720 16580 3732
rect 14783 3692 16580 3720
rect 14783 3689 14795 3692
rect 14737 3683 14795 3689
rect 14752 3652 14780 3683
rect 16574 3680 16580 3692
rect 16632 3680 16638 3732
rect 16684 3692 18000 3720
rect 16684 3652 16712 3692
rect 12023 3624 13124 3652
rect 13924 3624 14780 3652
rect 15580 3624 16712 3652
rect 17221 3655 17279 3661
rect 12023 3621 12035 3624
rect 11977 3615 12035 3621
rect 12820 3596 12848 3624
rect 12250 3584 12256 3596
rect 11624 3556 12256 3584
rect 11057 3547 11115 3553
rect 2593 3519 2651 3525
rect 2593 3485 2605 3519
rect 2639 3516 2651 3519
rect 2774 3516 2780 3528
rect 2639 3488 2780 3516
rect 2639 3485 2651 3488
rect 2593 3479 2651 3485
rect 2774 3476 2780 3488
rect 2832 3476 2838 3528
rect 3145 3519 3203 3525
rect 3145 3485 3157 3519
rect 3191 3516 3203 3519
rect 5813 3519 5871 3525
rect 5813 3516 5825 3519
rect 3191 3488 5825 3516
rect 3191 3485 3203 3488
rect 3145 3479 3203 3485
rect 5813 3485 5825 3488
rect 5859 3516 5871 3519
rect 6178 3516 6184 3528
rect 5859 3488 6184 3516
rect 5859 3485 5871 3488
rect 5813 3479 5871 3485
rect 6178 3476 6184 3488
rect 6236 3476 6242 3528
rect 6365 3519 6423 3525
rect 6365 3485 6377 3519
rect 6411 3485 6423 3519
rect 6365 3479 6423 3485
rect 9125 3519 9183 3525
rect 9125 3485 9137 3519
rect 9171 3516 9183 3519
rect 9306 3516 9312 3528
rect 9171 3488 9312 3516
rect 9171 3485 9183 3488
rect 9125 3479 9183 3485
rect 3881 3451 3939 3457
rect 3881 3417 3893 3451
rect 3927 3448 3939 3451
rect 5718 3448 5724 3460
rect 3927 3420 5724 3448
rect 3927 3417 3939 3420
rect 3881 3411 3939 3417
rect 5718 3408 5724 3420
rect 5776 3408 5782 3460
rect 5350 3380 5356 3392
rect 5311 3352 5356 3380
rect 5350 3340 5356 3352
rect 5408 3340 5414 3392
rect 6380 3380 6408 3479
rect 9306 3476 9312 3488
rect 9364 3516 9370 3528
rect 10229 3519 10287 3525
rect 10229 3516 10241 3519
rect 9364 3488 10241 3516
rect 9364 3476 9370 3488
rect 10229 3485 10241 3488
rect 10275 3485 10287 3519
rect 10229 3479 10287 3485
rect 10781 3519 10839 3525
rect 10781 3485 10793 3519
rect 10827 3485 10839 3519
rect 10781 3479 10839 3485
rect 7006 3408 7012 3460
rect 7064 3448 7070 3460
rect 7377 3451 7435 3457
rect 7377 3448 7389 3451
rect 7064 3420 7389 3448
rect 7064 3408 7070 3420
rect 7377 3417 7389 3420
rect 7423 3417 7435 3451
rect 7377 3411 7435 3417
rect 7650 3408 7656 3460
rect 7708 3448 7714 3460
rect 8297 3451 8355 3457
rect 8297 3448 8309 3451
rect 7708 3420 8309 3448
rect 7708 3408 7714 3420
rect 8297 3417 8309 3420
rect 8343 3448 8355 3451
rect 9030 3448 9036 3460
rect 8343 3420 9036 3448
rect 8343 3417 8355 3420
rect 8297 3411 8355 3417
rect 9030 3408 9036 3420
rect 9088 3408 9094 3460
rect 9398 3408 9404 3460
rect 9456 3448 9462 3460
rect 9674 3448 9680 3460
rect 9456 3420 9680 3448
rect 9456 3408 9462 3420
rect 9674 3408 9680 3420
rect 9732 3448 9738 3460
rect 10796 3448 10824 3479
rect 9732 3420 10824 3448
rect 11072 3448 11100 3547
rect 12250 3544 12256 3556
rect 12308 3584 12314 3596
rect 12618 3584 12624 3596
rect 12308 3556 12624 3584
rect 12308 3544 12314 3556
rect 12618 3544 12624 3556
rect 12676 3544 12682 3596
rect 12802 3584 12808 3596
rect 12715 3556 12808 3584
rect 12802 3544 12808 3556
rect 12860 3544 12866 3596
rect 12894 3544 12900 3596
rect 12952 3584 12958 3596
rect 12989 3587 13047 3593
rect 12989 3584 13001 3587
rect 12952 3556 13001 3584
rect 12952 3544 12958 3556
rect 12989 3553 13001 3556
rect 13035 3553 13047 3587
rect 13096 3584 13124 3624
rect 15580 3584 15608 3624
rect 17221 3621 17233 3655
rect 17267 3652 17279 3655
rect 17678 3652 17684 3664
rect 17267 3624 17684 3652
rect 17267 3621 17279 3624
rect 17221 3615 17279 3621
rect 17678 3612 17684 3624
rect 17736 3612 17742 3664
rect 13096 3556 15608 3584
rect 12989 3547 13047 3553
rect 15654 3544 15660 3596
rect 15712 3584 15718 3596
rect 16206 3584 16212 3596
rect 15712 3556 15757 3584
rect 16167 3556 16212 3584
rect 15712 3544 15718 3556
rect 16206 3544 16212 3556
rect 16264 3544 16270 3596
rect 17402 3584 17408 3596
rect 17363 3556 17408 3584
rect 17402 3544 17408 3556
rect 17460 3544 17466 3596
rect 17773 3587 17831 3593
rect 17773 3553 17785 3587
rect 17819 3584 17831 3587
rect 17862 3584 17868 3596
rect 17819 3556 17868 3584
rect 17819 3553 17831 3556
rect 17773 3547 17831 3553
rect 17862 3544 17868 3556
rect 17920 3544 17926 3596
rect 17972 3584 18000 3692
rect 18046 3680 18052 3732
rect 18104 3720 18110 3732
rect 18141 3723 18199 3729
rect 18141 3720 18153 3723
rect 18104 3692 18153 3720
rect 18104 3680 18110 3692
rect 18141 3689 18153 3692
rect 18187 3720 18199 3723
rect 19518 3720 19524 3732
rect 18187 3692 19524 3720
rect 18187 3689 18199 3692
rect 18141 3683 18199 3689
rect 19518 3680 19524 3692
rect 19576 3680 19582 3732
rect 20438 3720 20444 3732
rect 19628 3692 20444 3720
rect 18230 3612 18236 3664
rect 18288 3652 18294 3664
rect 19628 3652 19656 3692
rect 20438 3680 20444 3692
rect 20496 3680 20502 3732
rect 20806 3680 20812 3732
rect 20864 3720 20870 3732
rect 20864 3692 21864 3720
rect 20864 3680 20870 3692
rect 18288 3624 19656 3652
rect 21836 3652 21864 3692
rect 22370 3680 22376 3732
rect 22428 3720 22434 3732
rect 23014 3720 23020 3732
rect 22428 3692 23020 3720
rect 22428 3680 22434 3692
rect 23014 3680 23020 3692
rect 23072 3680 23078 3732
rect 23106 3680 23112 3732
rect 23164 3720 23170 3732
rect 23201 3723 23259 3729
rect 23201 3720 23213 3723
rect 23164 3692 23213 3720
rect 23164 3680 23170 3692
rect 23201 3689 23213 3692
rect 23247 3689 23259 3723
rect 23201 3683 23259 3689
rect 23842 3680 23848 3732
rect 23900 3720 23906 3732
rect 25038 3720 25044 3732
rect 23900 3692 25044 3720
rect 23900 3680 23906 3692
rect 25038 3680 25044 3692
rect 25096 3680 25102 3732
rect 25501 3723 25559 3729
rect 25501 3689 25513 3723
rect 25547 3720 25559 3723
rect 25590 3720 25596 3732
rect 25547 3692 25596 3720
rect 25547 3689 25559 3692
rect 25501 3683 25559 3689
rect 25590 3680 25596 3692
rect 25648 3680 25654 3732
rect 25961 3723 26019 3729
rect 25961 3689 25973 3723
rect 26007 3720 26019 3723
rect 26326 3720 26332 3732
rect 26007 3692 26332 3720
rect 26007 3689 26019 3692
rect 25961 3683 26019 3689
rect 26326 3680 26332 3692
rect 26384 3680 26390 3732
rect 26418 3680 26424 3732
rect 26476 3720 26482 3732
rect 31846 3720 31852 3732
rect 26476 3692 31852 3720
rect 26476 3680 26482 3692
rect 31846 3680 31852 3692
rect 31904 3680 31910 3732
rect 31941 3723 31999 3729
rect 31941 3689 31953 3723
rect 31987 3720 31999 3723
rect 32030 3720 32036 3732
rect 31987 3692 32036 3720
rect 31987 3689 31999 3692
rect 31941 3683 31999 3689
rect 32030 3680 32036 3692
rect 32088 3720 32094 3732
rect 32401 3723 32459 3729
rect 32401 3720 32413 3723
rect 32088 3692 32413 3720
rect 32088 3680 32094 3692
rect 32401 3689 32413 3692
rect 32447 3689 32459 3723
rect 32401 3683 32459 3689
rect 32766 3680 32772 3732
rect 32824 3720 32830 3732
rect 36541 3723 36599 3729
rect 32824 3692 35296 3720
rect 32824 3680 32830 3692
rect 22557 3655 22615 3661
rect 22557 3652 22569 3655
rect 21836 3624 22569 3652
rect 18288 3612 18294 3624
rect 22557 3621 22569 3624
rect 22603 3652 22615 3655
rect 23658 3652 23664 3664
rect 22603 3624 23664 3652
rect 22603 3621 22615 3624
rect 22557 3615 22615 3621
rect 23658 3612 23664 3624
rect 23716 3612 23722 3664
rect 23750 3612 23756 3664
rect 23808 3652 23814 3664
rect 25222 3652 25228 3664
rect 23808 3624 25228 3652
rect 23808 3612 23814 3624
rect 25222 3612 25228 3624
rect 25280 3612 25286 3664
rect 29086 3652 29092 3664
rect 25332 3624 28304 3652
rect 25332 3596 25360 3624
rect 28276 3596 28304 3624
rect 28552 3624 29092 3652
rect 17972 3556 18552 3584
rect 11238 3516 11244 3528
rect 11151 3488 11244 3516
rect 11238 3476 11244 3488
rect 11296 3516 11302 3528
rect 12069 3519 12127 3525
rect 11296 3488 12020 3516
rect 11296 3476 11302 3488
rect 11606 3448 11612 3460
rect 11072 3420 11612 3448
rect 9732 3408 9738 3420
rect 11606 3408 11612 3420
rect 11664 3408 11670 3460
rect 6822 3380 6828 3392
rect 6380 3352 6828 3380
rect 6822 3340 6828 3352
rect 6880 3340 6886 3392
rect 7190 3380 7196 3392
rect 7151 3352 7196 3380
rect 7190 3340 7196 3352
rect 7248 3340 7254 3392
rect 7282 3340 7288 3392
rect 7340 3380 7346 3392
rect 10870 3380 10876 3392
rect 7340 3352 10876 3380
rect 7340 3340 7346 3352
rect 10870 3340 10876 3352
rect 10928 3340 10934 3392
rect 11992 3380 12020 3488
rect 12069 3485 12081 3519
rect 12115 3485 12127 3519
rect 12069 3479 12127 3485
rect 12084 3448 12112 3479
rect 13446 3476 13452 3528
rect 13504 3516 13510 3528
rect 15010 3516 15016 3528
rect 13504 3488 15016 3516
rect 13504 3476 13510 3488
rect 15010 3476 15016 3488
rect 15068 3476 15074 3528
rect 15473 3519 15531 3525
rect 15473 3485 15485 3519
rect 15519 3516 15531 3519
rect 15930 3516 15936 3528
rect 15519 3488 15936 3516
rect 15519 3485 15531 3488
rect 15473 3479 15531 3485
rect 15930 3476 15936 3488
rect 15988 3476 15994 3528
rect 16393 3519 16451 3525
rect 16393 3485 16405 3519
rect 16439 3516 16451 3519
rect 18322 3516 18328 3528
rect 16439 3488 18328 3516
rect 16439 3485 16451 3488
rect 16393 3479 16451 3485
rect 18322 3476 18328 3488
rect 18380 3516 18386 3528
rect 18417 3519 18475 3525
rect 18417 3516 18429 3519
rect 18380 3488 18429 3516
rect 18380 3476 18386 3488
rect 18417 3485 18429 3488
rect 18463 3485 18475 3519
rect 18524 3516 18552 3556
rect 18690 3544 18696 3596
rect 18748 3584 18754 3596
rect 19245 3587 19303 3593
rect 19245 3584 19257 3587
rect 18748 3556 19257 3584
rect 18748 3544 18754 3556
rect 19245 3553 19257 3556
rect 19291 3553 19303 3587
rect 19245 3547 19303 3553
rect 19981 3587 20039 3593
rect 19981 3553 19993 3587
rect 20027 3584 20039 3587
rect 20625 3587 20683 3593
rect 20625 3584 20637 3587
rect 20027 3556 20637 3584
rect 20027 3553 20039 3556
rect 19981 3547 20039 3553
rect 20625 3553 20637 3556
rect 20671 3584 20683 3587
rect 20990 3584 20996 3596
rect 20671 3556 20996 3584
rect 20671 3553 20683 3556
rect 20625 3547 20683 3553
rect 20990 3544 20996 3556
rect 21048 3544 21054 3596
rect 21177 3587 21235 3593
rect 21177 3553 21189 3587
rect 21223 3584 21235 3587
rect 21266 3584 21272 3596
rect 21223 3556 21272 3584
rect 21223 3553 21235 3556
rect 21177 3547 21235 3553
rect 21266 3544 21272 3556
rect 21324 3544 21330 3596
rect 23566 3544 23572 3596
rect 23624 3584 23630 3596
rect 24213 3587 24271 3593
rect 24213 3584 24225 3587
rect 23624 3556 24225 3584
rect 23624 3544 23630 3556
rect 24213 3553 24225 3556
rect 24259 3584 24271 3587
rect 24854 3584 24860 3596
rect 24259 3556 24860 3584
rect 24259 3553 24271 3556
rect 24213 3547 24271 3553
rect 24854 3544 24860 3556
rect 24912 3544 24918 3596
rect 25314 3584 25320 3596
rect 25275 3556 25320 3584
rect 25314 3544 25320 3556
rect 25372 3544 25378 3596
rect 26510 3584 26516 3596
rect 26471 3556 26516 3584
rect 26510 3544 26516 3556
rect 26568 3544 26574 3596
rect 26786 3544 26792 3596
rect 26844 3584 26850 3596
rect 28074 3584 28080 3596
rect 26844 3556 28080 3584
rect 26844 3544 26850 3556
rect 28074 3544 28080 3556
rect 28132 3544 28138 3596
rect 28258 3584 28264 3596
rect 28171 3556 28264 3584
rect 28258 3544 28264 3556
rect 28316 3544 28322 3596
rect 28552 3593 28580 3624
rect 29086 3612 29092 3624
rect 29144 3652 29150 3664
rect 29365 3655 29423 3661
rect 29365 3652 29377 3655
rect 29144 3624 29377 3652
rect 29144 3612 29150 3624
rect 29365 3621 29377 3624
rect 29411 3621 29423 3655
rect 29365 3615 29423 3621
rect 30466 3612 30472 3664
rect 30524 3652 30530 3664
rect 32493 3655 32551 3661
rect 32493 3652 32505 3655
rect 30524 3624 32505 3652
rect 30524 3612 30530 3624
rect 32493 3621 32505 3624
rect 32539 3652 32551 3655
rect 33502 3652 33508 3664
rect 32539 3624 33508 3652
rect 32539 3621 32551 3624
rect 32493 3615 32551 3621
rect 33502 3612 33508 3624
rect 33560 3612 33566 3664
rect 35069 3655 35127 3661
rect 35069 3652 35081 3655
rect 34256 3624 35081 3652
rect 28537 3587 28595 3593
rect 28537 3553 28549 3587
rect 28583 3553 28595 3587
rect 28537 3547 28595 3553
rect 28721 3587 28779 3593
rect 28721 3553 28733 3587
rect 28767 3584 28779 3587
rect 28902 3584 28908 3596
rect 28767 3556 28908 3584
rect 28767 3553 28779 3556
rect 28721 3547 28779 3553
rect 28902 3544 28908 3556
rect 28960 3544 28966 3596
rect 28997 3587 29055 3593
rect 28997 3553 29009 3587
rect 29043 3584 29055 3587
rect 29733 3587 29791 3593
rect 29733 3584 29745 3587
rect 29043 3556 29745 3584
rect 29043 3553 29055 3556
rect 28997 3547 29055 3553
rect 29733 3553 29745 3556
rect 29779 3584 29791 3587
rect 29914 3584 29920 3596
rect 29779 3556 29920 3584
rect 29779 3553 29791 3556
rect 29733 3547 29791 3553
rect 29914 3544 29920 3556
rect 29972 3544 29978 3596
rect 30193 3587 30251 3593
rect 30193 3553 30205 3587
rect 30239 3584 30251 3587
rect 30282 3584 30288 3596
rect 30239 3556 30288 3584
rect 30239 3553 30251 3556
rect 30193 3547 30251 3553
rect 30282 3544 30288 3556
rect 30340 3544 30346 3596
rect 30558 3584 30564 3596
rect 30519 3556 30564 3584
rect 30558 3544 30564 3556
rect 30616 3544 30622 3596
rect 30650 3544 30656 3596
rect 30708 3584 30714 3596
rect 32309 3587 32367 3593
rect 32309 3584 32321 3587
rect 30708 3556 32321 3584
rect 30708 3544 30714 3556
rect 31956 3528 31984 3556
rect 32309 3553 32321 3556
rect 32355 3553 32367 3587
rect 32309 3547 32367 3553
rect 33962 3544 33968 3596
rect 34020 3584 34026 3596
rect 34256 3593 34284 3624
rect 35069 3621 35081 3624
rect 35115 3621 35127 3655
rect 35268 3652 35296 3692
rect 36541 3689 36553 3723
rect 36587 3720 36599 3723
rect 36722 3720 36728 3732
rect 36587 3692 36728 3720
rect 36587 3689 36599 3692
rect 36541 3683 36599 3689
rect 36722 3680 36728 3692
rect 36780 3680 36786 3732
rect 37734 3680 37740 3732
rect 37792 3720 37798 3732
rect 37921 3723 37979 3729
rect 37921 3720 37933 3723
rect 37792 3692 37933 3720
rect 37792 3680 37798 3692
rect 37921 3689 37933 3692
rect 37967 3689 37979 3723
rect 37921 3683 37979 3689
rect 36262 3652 36268 3664
rect 35268 3624 36268 3652
rect 35069 3615 35127 3621
rect 36262 3612 36268 3624
rect 36320 3652 36326 3664
rect 36817 3655 36875 3661
rect 36817 3652 36829 3655
rect 36320 3624 36829 3652
rect 36320 3612 36326 3624
rect 36817 3621 36829 3624
rect 36863 3621 36875 3655
rect 37936 3652 37964 3683
rect 38010 3680 38016 3732
rect 38068 3720 38074 3732
rect 38838 3720 38844 3732
rect 38068 3692 38844 3720
rect 38068 3680 38074 3692
rect 38838 3680 38844 3692
rect 38896 3680 38902 3732
rect 38930 3680 38936 3732
rect 38988 3720 38994 3732
rect 39853 3723 39911 3729
rect 39853 3720 39865 3723
rect 38988 3692 39865 3720
rect 38988 3680 38994 3692
rect 39853 3689 39865 3692
rect 39899 3689 39911 3723
rect 39853 3683 39911 3689
rect 41230 3680 41236 3732
rect 41288 3720 41294 3732
rect 41966 3720 41972 3732
rect 41288 3692 41972 3720
rect 41288 3680 41294 3692
rect 41966 3680 41972 3692
rect 42024 3680 42030 3732
rect 42245 3723 42303 3729
rect 42245 3689 42257 3723
rect 42291 3689 42303 3723
rect 42245 3683 42303 3689
rect 44361 3723 44419 3729
rect 44361 3689 44373 3723
rect 44407 3720 44419 3723
rect 46198 3720 46204 3732
rect 44407 3692 46204 3720
rect 44407 3689 44419 3692
rect 44361 3683 44419 3689
rect 41414 3652 41420 3664
rect 37936 3624 41420 3652
rect 36817 3615 36875 3621
rect 41414 3612 41420 3624
rect 41472 3612 41478 3664
rect 41598 3652 41604 3664
rect 41511 3624 41604 3652
rect 41598 3612 41604 3624
rect 41656 3652 41662 3664
rect 42260 3652 42288 3683
rect 46198 3680 46204 3692
rect 46256 3680 46262 3732
rect 46290 3680 46296 3732
rect 46348 3720 46354 3732
rect 47581 3723 47639 3729
rect 47581 3720 47593 3723
rect 46348 3692 47593 3720
rect 46348 3680 46354 3692
rect 47581 3689 47593 3692
rect 47627 3689 47639 3723
rect 47581 3683 47639 3689
rect 47949 3723 48007 3729
rect 47949 3689 47961 3723
rect 47995 3720 48007 3723
rect 48038 3720 48044 3732
rect 47995 3692 48044 3720
rect 47995 3689 48007 3692
rect 47949 3683 48007 3689
rect 48038 3680 48044 3692
rect 48096 3680 48102 3732
rect 48777 3723 48835 3729
rect 48777 3689 48789 3723
rect 48823 3720 48835 3723
rect 48958 3720 48964 3732
rect 48823 3692 48964 3720
rect 48823 3689 48835 3692
rect 48777 3683 48835 3689
rect 48958 3680 48964 3692
rect 49016 3680 49022 3732
rect 49050 3680 49056 3732
rect 49108 3720 49114 3732
rect 49145 3723 49203 3729
rect 49145 3720 49157 3723
rect 49108 3692 49157 3720
rect 49108 3680 49114 3692
rect 49145 3689 49157 3692
rect 49191 3689 49203 3723
rect 49878 3720 49884 3732
rect 49839 3692 49884 3720
rect 49145 3683 49203 3689
rect 49878 3680 49884 3692
rect 49936 3680 49942 3732
rect 50062 3680 50068 3732
rect 50120 3720 50126 3732
rect 51813 3723 51871 3729
rect 51813 3720 51825 3723
rect 50120 3692 51825 3720
rect 50120 3680 50126 3692
rect 51813 3689 51825 3692
rect 51859 3720 51871 3723
rect 51859 3692 52316 3720
rect 51859 3689 51871 3692
rect 51813 3683 51871 3689
rect 44818 3652 44824 3664
rect 41656 3624 44824 3652
rect 41656 3612 41662 3624
rect 44818 3612 44824 3624
rect 44876 3612 44882 3664
rect 46934 3612 46940 3664
rect 46992 3652 46998 3664
rect 47210 3652 47216 3664
rect 46992 3624 47216 3652
rect 46992 3612 46998 3624
rect 47210 3612 47216 3624
rect 47268 3612 47274 3664
rect 47394 3612 47400 3664
rect 47452 3652 47458 3664
rect 50798 3652 50804 3664
rect 47452 3624 50804 3652
rect 47452 3612 47458 3624
rect 34241 3587 34299 3593
rect 34241 3584 34253 3587
rect 34020 3556 34253 3584
rect 34020 3544 34026 3556
rect 34241 3553 34253 3556
rect 34287 3553 34299 3587
rect 34241 3547 34299 3553
rect 34422 3544 34428 3596
rect 34480 3584 34486 3596
rect 34609 3587 34667 3593
rect 34609 3584 34621 3587
rect 34480 3556 34621 3584
rect 34480 3544 34486 3556
rect 34609 3553 34621 3556
rect 34655 3553 34667 3587
rect 34609 3547 34667 3553
rect 34698 3544 34704 3596
rect 34756 3584 34762 3596
rect 35713 3587 35771 3593
rect 34756 3556 35112 3584
rect 34756 3544 34762 3556
rect 19610 3516 19616 3528
rect 18524 3488 19472 3516
rect 19523 3488 19616 3516
rect 18417 3479 18475 3485
rect 12342 3448 12348 3460
rect 12084 3420 12348 3448
rect 12342 3408 12348 3420
rect 12400 3448 12406 3460
rect 14090 3448 14096 3460
rect 12400 3420 14096 3448
rect 12400 3408 12406 3420
rect 14090 3408 14096 3420
rect 14148 3408 14154 3460
rect 15028 3448 15056 3476
rect 19444 3448 19472 3488
rect 19610 3476 19616 3488
rect 19668 3516 19674 3528
rect 20070 3516 20076 3528
rect 19668 3488 20076 3516
rect 19668 3476 19674 3488
rect 20070 3476 20076 3488
rect 20128 3476 20134 3528
rect 20901 3519 20959 3525
rect 20901 3485 20913 3519
rect 20947 3516 20959 3519
rect 21358 3516 21364 3528
rect 20947 3488 21364 3516
rect 20947 3485 20959 3488
rect 20901 3479 20959 3485
rect 21358 3476 21364 3488
rect 21416 3476 21422 3528
rect 23382 3516 23388 3528
rect 23343 3488 23388 3516
rect 23382 3476 23388 3488
rect 23440 3476 23446 3528
rect 23750 3476 23756 3528
rect 23808 3516 23814 3528
rect 23937 3519 23995 3525
rect 23937 3516 23949 3519
rect 23808 3488 23949 3516
rect 23808 3476 23814 3488
rect 23937 3485 23949 3488
rect 23983 3485 23995 3519
rect 23937 3479 23995 3485
rect 24397 3519 24455 3525
rect 24397 3485 24409 3519
rect 24443 3516 24455 3519
rect 24578 3516 24584 3528
rect 24443 3488 24584 3516
rect 24443 3485 24455 3488
rect 24397 3479 24455 3485
rect 24578 3476 24584 3488
rect 24636 3476 24642 3528
rect 24762 3476 24768 3528
rect 24820 3516 24826 3528
rect 27614 3516 27620 3528
rect 24820 3488 27620 3516
rect 24820 3476 24826 3488
rect 27614 3476 27620 3488
rect 27672 3476 27678 3528
rect 31573 3519 31631 3525
rect 27724 3488 30972 3516
rect 20254 3448 20260 3460
rect 15028 3420 19380 3448
rect 19444 3420 20260 3448
rect 12894 3380 12900 3392
rect 11992 3352 12900 3380
rect 12894 3340 12900 3352
rect 12952 3340 12958 3392
rect 13262 3380 13268 3392
rect 13223 3352 13268 3380
rect 13262 3340 13268 3352
rect 13320 3340 13326 3392
rect 13814 3380 13820 3392
rect 13775 3352 13820 3380
rect 13814 3340 13820 3352
rect 13872 3340 13878 3392
rect 14366 3340 14372 3392
rect 14424 3380 14430 3392
rect 15930 3380 15936 3392
rect 14424 3352 15936 3380
rect 14424 3340 14430 3352
rect 15930 3340 15936 3352
rect 15988 3340 15994 3392
rect 16114 3340 16120 3392
rect 16172 3380 16178 3392
rect 16669 3383 16727 3389
rect 16669 3380 16681 3383
rect 16172 3352 16681 3380
rect 16172 3340 16178 3352
rect 16669 3349 16681 3352
rect 16715 3349 16727 3383
rect 16669 3343 16727 3349
rect 17129 3383 17187 3389
rect 17129 3349 17141 3383
rect 17175 3380 17187 3383
rect 18598 3380 18604 3392
rect 17175 3352 18604 3380
rect 17175 3349 17187 3352
rect 17129 3343 17187 3349
rect 18598 3340 18604 3352
rect 18656 3340 18662 3392
rect 19153 3383 19211 3389
rect 19153 3349 19165 3383
rect 19199 3380 19211 3383
rect 19242 3380 19248 3392
rect 19199 3352 19248 3380
rect 19199 3349 19211 3352
rect 19153 3343 19211 3349
rect 19242 3340 19248 3352
rect 19300 3340 19306 3392
rect 19352 3380 19380 3420
rect 20254 3408 20260 3420
rect 20312 3408 20318 3460
rect 20349 3451 20407 3457
rect 20349 3417 20361 3451
rect 20395 3448 20407 3451
rect 20438 3448 20444 3460
rect 20395 3420 20444 3448
rect 20395 3417 20407 3420
rect 20349 3411 20407 3417
rect 20438 3408 20444 3420
rect 20496 3408 20502 3460
rect 22462 3408 22468 3460
rect 22520 3448 22526 3460
rect 22520 3420 25176 3448
rect 22520 3408 22526 3420
rect 21818 3380 21824 3392
rect 19352 3352 21824 3380
rect 21818 3340 21824 3352
rect 21876 3340 21882 3392
rect 22738 3340 22744 3392
rect 22796 3380 22802 3392
rect 22833 3383 22891 3389
rect 22833 3380 22845 3383
rect 22796 3352 22845 3380
rect 22796 3340 22802 3352
rect 22833 3349 22845 3352
rect 22879 3380 22891 3383
rect 24486 3380 24492 3392
rect 22879 3352 24492 3380
rect 22879 3349 22891 3352
rect 22833 3343 22891 3349
rect 24486 3340 24492 3352
rect 24544 3340 24550 3392
rect 24578 3340 24584 3392
rect 24636 3380 24642 3392
rect 24673 3383 24731 3389
rect 24673 3380 24685 3383
rect 24636 3352 24685 3380
rect 24636 3340 24642 3352
rect 24673 3349 24685 3352
rect 24719 3380 24731 3383
rect 25041 3383 25099 3389
rect 25041 3380 25053 3383
rect 24719 3352 25053 3380
rect 24719 3349 24731 3352
rect 24673 3343 24731 3349
rect 25041 3349 25053 3352
rect 25087 3349 25099 3383
rect 25148 3380 25176 3420
rect 26510 3408 26516 3460
rect 26568 3448 26574 3460
rect 26697 3451 26755 3457
rect 26697 3448 26709 3451
rect 26568 3420 26709 3448
rect 26568 3408 26574 3420
rect 26697 3417 26709 3420
rect 26743 3417 26755 3451
rect 26697 3411 26755 3417
rect 26786 3408 26792 3460
rect 26844 3448 26850 3460
rect 27724 3448 27752 3488
rect 26844 3420 27752 3448
rect 26844 3408 26850 3420
rect 27890 3408 27896 3460
rect 27948 3448 27954 3460
rect 30009 3451 30067 3457
rect 30009 3448 30021 3451
rect 27948 3420 30021 3448
rect 27948 3408 27954 3420
rect 30009 3417 30021 3420
rect 30055 3417 30067 3451
rect 30009 3411 30067 3417
rect 26142 3380 26148 3392
rect 25148 3352 26148 3380
rect 25041 3343 25099 3349
rect 26142 3340 26148 3352
rect 26200 3340 26206 3392
rect 26326 3380 26332 3392
rect 26239 3352 26332 3380
rect 26326 3340 26332 3352
rect 26384 3380 26390 3392
rect 26970 3380 26976 3392
rect 26384 3352 26976 3380
rect 26384 3340 26390 3352
rect 26970 3340 26976 3352
rect 27028 3340 27034 3392
rect 27157 3383 27215 3389
rect 27157 3349 27169 3383
rect 27203 3380 27215 3383
rect 27246 3380 27252 3392
rect 27203 3352 27252 3380
rect 27203 3349 27215 3352
rect 27157 3343 27215 3349
rect 27246 3340 27252 3352
rect 27304 3340 27310 3392
rect 27430 3380 27436 3392
rect 27391 3352 27436 3380
rect 27430 3340 27436 3352
rect 27488 3340 27494 3392
rect 30944 3380 30972 3488
rect 31573 3485 31585 3519
rect 31619 3516 31631 3519
rect 31754 3516 31760 3528
rect 31619 3488 31760 3516
rect 31619 3485 31631 3488
rect 31573 3479 31631 3485
rect 31754 3476 31760 3488
rect 31812 3476 31818 3528
rect 31938 3476 31944 3528
rect 31996 3476 32002 3528
rect 32125 3519 32183 3525
rect 32125 3485 32137 3519
rect 32171 3516 32183 3519
rect 32674 3516 32680 3528
rect 32171 3488 32680 3516
rect 32171 3485 32183 3488
rect 32125 3479 32183 3485
rect 32674 3476 32680 3488
rect 32732 3476 32738 3528
rect 32861 3519 32919 3525
rect 32861 3485 32873 3519
rect 32907 3485 32919 3519
rect 32861 3479 32919 3485
rect 31018 3408 31024 3460
rect 31076 3448 31082 3460
rect 31113 3451 31171 3457
rect 31113 3448 31125 3451
rect 31076 3420 31125 3448
rect 31076 3408 31082 3420
rect 31113 3417 31125 3420
rect 31159 3448 31171 3451
rect 32876 3448 32904 3479
rect 31159 3420 32904 3448
rect 34057 3451 34115 3457
rect 31159 3417 31171 3420
rect 31113 3411 31171 3417
rect 34057 3417 34069 3451
rect 34103 3448 34115 3451
rect 34330 3448 34336 3460
rect 34103 3420 34336 3448
rect 34103 3417 34115 3420
rect 34057 3411 34115 3417
rect 34330 3408 34336 3420
rect 34388 3408 34394 3460
rect 35084 3448 35112 3556
rect 35713 3553 35725 3587
rect 35759 3584 35771 3587
rect 35894 3584 35900 3596
rect 35759 3556 35900 3584
rect 35759 3553 35771 3556
rect 35713 3547 35771 3553
rect 35894 3544 35900 3556
rect 35952 3544 35958 3596
rect 36354 3544 36360 3596
rect 36412 3584 36418 3596
rect 38470 3584 38476 3596
rect 36412 3556 38476 3584
rect 36412 3544 36418 3556
rect 38470 3544 38476 3556
rect 38528 3584 38534 3596
rect 38657 3587 38715 3593
rect 38657 3584 38669 3587
rect 38528 3556 38669 3584
rect 38528 3544 38534 3556
rect 38657 3553 38669 3556
rect 38703 3553 38715 3587
rect 38657 3547 38715 3553
rect 38746 3544 38752 3596
rect 38804 3584 38810 3596
rect 38841 3587 38899 3593
rect 38841 3584 38853 3587
rect 38804 3556 38853 3584
rect 38804 3544 38810 3556
rect 38841 3553 38853 3556
rect 38887 3553 38899 3587
rect 38841 3547 38899 3553
rect 40310 3544 40316 3596
rect 40368 3584 40374 3596
rect 40678 3584 40684 3596
rect 40368 3556 40684 3584
rect 40368 3544 40374 3556
rect 40678 3544 40684 3556
rect 40736 3544 40742 3596
rect 41049 3587 41107 3593
rect 41049 3553 41061 3587
rect 41095 3584 41107 3587
rect 41616 3584 41644 3612
rect 42058 3584 42064 3596
rect 41095 3556 41644 3584
rect 41971 3556 42064 3584
rect 41095 3553 41107 3556
rect 41049 3547 41107 3553
rect 42058 3544 42064 3556
rect 42116 3584 42122 3596
rect 43070 3584 43076 3596
rect 42116 3556 43076 3584
rect 42116 3544 42122 3556
rect 43070 3544 43076 3556
rect 43128 3544 43134 3596
rect 43714 3584 43720 3596
rect 43675 3556 43720 3584
rect 43714 3544 43720 3556
rect 43772 3544 43778 3596
rect 45186 3584 45192 3596
rect 43916 3556 45192 3584
rect 35345 3519 35403 3525
rect 35345 3485 35357 3519
rect 35391 3516 35403 3519
rect 35621 3519 35679 3525
rect 35621 3516 35633 3519
rect 35391 3488 35633 3516
rect 35391 3485 35403 3488
rect 35345 3479 35403 3485
rect 35621 3485 35633 3488
rect 35667 3485 35679 3519
rect 35621 3479 35679 3485
rect 36173 3519 36231 3525
rect 36173 3485 36185 3519
rect 36219 3485 36231 3519
rect 36173 3479 36231 3485
rect 38565 3519 38623 3525
rect 38565 3485 38577 3519
rect 38611 3516 38623 3519
rect 39206 3516 39212 3528
rect 38611 3488 39212 3516
rect 38611 3485 38623 3488
rect 38565 3479 38623 3485
rect 36188 3448 36216 3479
rect 39206 3476 39212 3488
rect 39264 3476 39270 3528
rect 40586 3516 40592 3528
rect 40547 3488 40592 3516
rect 40586 3476 40592 3488
rect 40644 3476 40650 3528
rect 41141 3519 41199 3525
rect 41141 3485 41153 3519
rect 41187 3516 41199 3519
rect 43625 3519 43683 3525
rect 41187 3488 41552 3516
rect 41187 3485 41199 3488
rect 41141 3479 41199 3485
rect 35084 3420 36216 3448
rect 36630 3408 36636 3460
rect 36688 3448 36694 3460
rect 41524 3448 41552 3488
rect 43625 3485 43637 3519
rect 43671 3516 43683 3519
rect 43916 3516 43944 3556
rect 45186 3544 45192 3556
rect 45244 3544 45250 3596
rect 45554 3584 45560 3596
rect 45515 3556 45560 3584
rect 45554 3544 45560 3556
rect 45612 3584 45618 3596
rect 46198 3584 46204 3596
rect 45612 3556 46204 3584
rect 45612 3544 45618 3556
rect 46198 3544 46204 3556
rect 46256 3544 46262 3596
rect 46750 3544 46756 3596
rect 46808 3584 46814 3596
rect 47489 3587 47547 3593
rect 47489 3584 47501 3587
rect 46808 3556 47501 3584
rect 46808 3544 46814 3556
rect 47489 3553 47501 3556
rect 47535 3584 47547 3587
rect 47765 3587 47823 3593
rect 47765 3584 47777 3587
rect 47535 3556 47777 3584
rect 47535 3553 47547 3556
rect 47489 3547 47547 3553
rect 47765 3553 47777 3556
rect 47811 3553 47823 3587
rect 47765 3547 47823 3553
rect 47854 3544 47860 3596
rect 47912 3584 47918 3596
rect 48866 3584 48872 3596
rect 47912 3556 48872 3584
rect 47912 3544 47918 3556
rect 48866 3544 48872 3556
rect 48924 3544 48930 3596
rect 48976 3593 49004 3624
rect 50798 3612 50804 3624
rect 50856 3612 50862 3664
rect 50908 3624 52040 3652
rect 48961 3587 49019 3593
rect 48961 3553 48973 3587
rect 49007 3553 49019 3587
rect 50062 3584 50068 3596
rect 50023 3556 50068 3584
rect 48961 3547 49019 3553
rect 50062 3544 50068 3556
rect 50120 3544 50126 3596
rect 50908 3593 50936 3624
rect 52012 3596 52040 3624
rect 50893 3587 50951 3593
rect 50893 3553 50905 3587
rect 50939 3553 50951 3587
rect 50893 3547 50951 3553
rect 51074 3544 51080 3596
rect 51132 3584 51138 3596
rect 51718 3584 51724 3596
rect 51132 3556 51724 3584
rect 51132 3544 51138 3556
rect 51718 3544 51724 3556
rect 51776 3544 51782 3596
rect 51994 3584 52000 3596
rect 51955 3556 52000 3584
rect 51994 3544 52000 3556
rect 52052 3544 52058 3596
rect 52089 3587 52147 3593
rect 52089 3553 52101 3587
rect 52135 3584 52147 3587
rect 52178 3584 52184 3596
rect 52135 3556 52184 3584
rect 52135 3553 52147 3556
rect 52089 3547 52147 3553
rect 52178 3544 52184 3556
rect 52236 3544 52242 3596
rect 52288 3593 52316 3692
rect 52362 3680 52368 3732
rect 52420 3720 52426 3732
rect 52420 3692 53604 3720
rect 52420 3680 52426 3692
rect 52733 3655 52791 3661
rect 52733 3621 52745 3655
rect 52779 3652 52791 3655
rect 53576 3652 53604 3692
rect 54018 3680 54024 3732
rect 54076 3720 54082 3732
rect 54205 3723 54263 3729
rect 54205 3720 54217 3723
rect 54076 3692 54217 3720
rect 54076 3680 54082 3692
rect 54205 3689 54217 3692
rect 54251 3689 54263 3723
rect 54757 3723 54815 3729
rect 54757 3720 54769 3723
rect 54205 3683 54263 3689
rect 54312 3692 54769 3720
rect 54312 3652 54340 3692
rect 54757 3689 54769 3692
rect 54803 3689 54815 3723
rect 54757 3683 54815 3689
rect 54846 3680 54852 3732
rect 54904 3720 54910 3732
rect 56226 3720 56232 3732
rect 54904 3692 56088 3720
rect 56187 3692 56232 3720
rect 54904 3680 54910 3692
rect 52779 3624 53512 3652
rect 53576 3624 54340 3652
rect 52779 3621 52791 3624
rect 52733 3615 52791 3621
rect 52273 3587 52331 3593
rect 52273 3553 52285 3587
rect 52319 3553 52331 3587
rect 52273 3547 52331 3553
rect 52362 3544 52368 3596
rect 52420 3584 52426 3596
rect 53374 3584 53380 3596
rect 52420 3556 52592 3584
rect 53335 3556 53380 3584
rect 52420 3544 52426 3556
rect 43671 3488 43944 3516
rect 44085 3519 44143 3525
rect 43671 3485 43683 3488
rect 43625 3479 43683 3485
rect 44085 3485 44097 3519
rect 44131 3516 44143 3519
rect 44634 3516 44640 3528
rect 44131 3488 44640 3516
rect 44131 3485 44143 3488
rect 44085 3479 44143 3485
rect 42705 3451 42763 3457
rect 42705 3448 42717 3451
rect 36688 3420 41460 3448
rect 41524 3420 42717 3448
rect 36688 3408 36694 3420
rect 33042 3380 33048 3392
rect 30944 3352 33048 3380
rect 33042 3340 33048 3352
rect 33100 3340 33106 3392
rect 33226 3380 33232 3392
rect 33187 3352 33232 3380
rect 33226 3340 33232 3352
rect 33284 3340 33290 3392
rect 33502 3380 33508 3392
rect 33463 3352 33508 3380
rect 33502 3340 33508 3352
rect 33560 3340 33566 3392
rect 34514 3340 34520 3392
rect 34572 3380 34578 3392
rect 35345 3383 35403 3389
rect 35345 3380 35357 3383
rect 34572 3352 35357 3380
rect 34572 3340 34578 3352
rect 35345 3349 35357 3352
rect 35391 3380 35403 3383
rect 35437 3383 35495 3389
rect 35437 3380 35449 3383
rect 35391 3352 35449 3380
rect 35391 3349 35403 3352
rect 35345 3343 35403 3349
rect 35437 3349 35449 3352
rect 35483 3380 35495 3383
rect 36446 3380 36452 3392
rect 35483 3352 36452 3380
rect 35483 3349 35495 3352
rect 35437 3343 35495 3349
rect 36446 3340 36452 3352
rect 36504 3380 36510 3392
rect 37185 3383 37243 3389
rect 37185 3380 37197 3383
rect 36504 3352 37197 3380
rect 36504 3340 36510 3352
rect 37185 3349 37197 3352
rect 37231 3349 37243 3383
rect 37185 3343 37243 3349
rect 38470 3340 38476 3392
rect 38528 3380 38534 3392
rect 39482 3380 39488 3392
rect 38528 3352 39488 3380
rect 38528 3340 38534 3352
rect 39482 3340 39488 3352
rect 39540 3340 39546 3392
rect 40126 3380 40132 3392
rect 40087 3352 40132 3380
rect 40126 3340 40132 3352
rect 40184 3340 40190 3392
rect 41432 3380 41460 3420
rect 42705 3417 42717 3420
rect 42751 3448 42763 3451
rect 43640 3448 43668 3479
rect 44634 3476 44640 3488
rect 44692 3476 44698 3528
rect 45281 3519 45339 3525
rect 45281 3485 45293 3519
rect 45327 3485 45339 3519
rect 45281 3479 45339 3485
rect 42751 3420 43668 3448
rect 43882 3451 43940 3457
rect 42751 3417 42763 3420
rect 42705 3411 42763 3417
rect 43882 3417 43894 3451
rect 43928 3448 43940 3451
rect 44818 3448 44824 3460
rect 43928 3420 44824 3448
rect 43928 3417 43940 3420
rect 43882 3411 43940 3417
rect 44818 3408 44824 3420
rect 44876 3408 44882 3460
rect 45094 3448 45100 3460
rect 45055 3420 45100 3448
rect 45094 3408 45100 3420
rect 45152 3408 45158 3460
rect 42794 3380 42800 3392
rect 41432 3352 42800 3380
rect 42794 3340 42800 3352
rect 42852 3340 42858 3392
rect 42978 3380 42984 3392
rect 42939 3352 42984 3380
rect 42978 3340 42984 3352
rect 43036 3340 43042 3392
rect 43990 3380 43996 3392
rect 43951 3352 43996 3380
rect 43990 3340 43996 3352
rect 44048 3340 44054 3392
rect 44266 3340 44272 3392
rect 44324 3380 44330 3392
rect 45296 3380 45324 3479
rect 45462 3476 45468 3528
rect 45520 3516 45526 3528
rect 52564 3516 52592 3556
rect 53374 3544 53380 3556
rect 53432 3544 53438 3596
rect 53484 3584 53512 3624
rect 54662 3612 54668 3664
rect 54720 3652 54726 3664
rect 54720 3624 55628 3652
rect 54720 3612 54726 3624
rect 53742 3584 53748 3596
rect 53484 3556 53748 3584
rect 53742 3544 53748 3556
rect 53800 3544 53806 3596
rect 54570 3544 54576 3596
rect 54628 3584 54634 3596
rect 54938 3584 54944 3596
rect 54628 3556 54944 3584
rect 54628 3544 54634 3556
rect 54938 3544 54944 3556
rect 54996 3544 55002 3596
rect 55030 3544 55036 3596
rect 55088 3584 55094 3596
rect 55217 3587 55275 3593
rect 55088 3556 55133 3584
rect 55088 3544 55094 3556
rect 55217 3553 55229 3587
rect 55263 3584 55275 3587
rect 55306 3584 55312 3596
rect 55263 3556 55312 3584
rect 55263 3553 55275 3556
rect 55217 3547 55275 3553
rect 55306 3544 55312 3556
rect 55364 3544 55370 3596
rect 55600 3584 55628 3624
rect 55674 3612 55680 3664
rect 55732 3652 55738 3664
rect 56060 3652 56088 3692
rect 56226 3680 56232 3692
rect 56284 3680 56290 3732
rect 56781 3723 56839 3729
rect 56781 3720 56793 3723
rect 56336 3692 56793 3720
rect 56336 3652 56364 3692
rect 56781 3689 56793 3692
rect 56827 3720 56839 3723
rect 57885 3723 57943 3729
rect 57885 3720 57897 3723
rect 56827 3692 57897 3720
rect 56827 3689 56839 3692
rect 56781 3683 56839 3689
rect 57885 3689 57897 3692
rect 57931 3689 57943 3723
rect 57885 3683 57943 3689
rect 58069 3723 58127 3729
rect 58069 3689 58081 3723
rect 58115 3720 58127 3723
rect 59906 3720 59912 3732
rect 58115 3692 59912 3720
rect 58115 3689 58127 3692
rect 58069 3683 58127 3689
rect 59906 3680 59912 3692
rect 59964 3680 59970 3732
rect 57330 3652 57336 3664
rect 55732 3624 55777 3652
rect 56060 3624 56364 3652
rect 56428 3624 57336 3652
rect 55732 3612 55738 3624
rect 56428 3584 56456 3624
rect 57330 3612 57336 3624
rect 57388 3612 57394 3664
rect 59265 3655 59323 3661
rect 59265 3621 59277 3655
rect 59311 3652 59323 3655
rect 60458 3652 60464 3664
rect 59311 3624 60464 3652
rect 59311 3621 59323 3624
rect 59265 3615 59323 3621
rect 60458 3612 60464 3624
rect 60516 3612 60522 3664
rect 55600 3556 56456 3584
rect 56502 3544 56508 3596
rect 56560 3584 56566 3596
rect 56689 3587 56747 3593
rect 56560 3556 56605 3584
rect 56560 3544 56566 3556
rect 56689 3553 56701 3587
rect 56735 3584 56747 3587
rect 57238 3584 57244 3596
rect 56735 3556 57244 3584
rect 56735 3553 56747 3556
rect 56689 3547 56747 3553
rect 57238 3544 57244 3556
rect 57296 3544 57302 3596
rect 57885 3587 57943 3593
rect 57885 3553 57897 3587
rect 57931 3584 57943 3587
rect 58342 3584 58348 3596
rect 57931 3556 58348 3584
rect 57931 3553 57943 3556
rect 57885 3547 57943 3553
rect 58342 3544 58348 3556
rect 58400 3544 58406 3596
rect 58526 3584 58532 3596
rect 58487 3556 58532 3584
rect 58526 3544 58532 3556
rect 58584 3544 58590 3596
rect 58710 3544 58716 3596
rect 58768 3584 58774 3596
rect 58805 3587 58863 3593
rect 58805 3584 58817 3587
rect 58768 3556 58817 3584
rect 58768 3544 58774 3556
rect 58805 3553 58817 3556
rect 58851 3553 58863 3587
rect 58805 3547 58863 3553
rect 59446 3544 59452 3596
rect 59504 3584 59510 3596
rect 59541 3587 59599 3593
rect 59541 3584 59553 3587
rect 59504 3556 59553 3584
rect 59504 3544 59510 3556
rect 59541 3553 59553 3556
rect 59587 3553 59599 3587
rect 59541 3547 59599 3553
rect 59630 3544 59636 3596
rect 59688 3584 59694 3596
rect 59909 3587 59967 3593
rect 59909 3584 59921 3587
rect 59688 3556 59921 3584
rect 59688 3544 59694 3556
rect 59909 3553 59921 3556
rect 59955 3584 59967 3587
rect 60185 3587 60243 3593
rect 60185 3584 60197 3587
rect 59955 3556 60197 3584
rect 59955 3553 59967 3556
rect 59909 3547 59967 3553
rect 60185 3553 60197 3556
rect 60231 3553 60243 3587
rect 60185 3547 60243 3553
rect 60274 3544 60280 3596
rect 60332 3584 60338 3596
rect 60369 3587 60427 3593
rect 60369 3584 60381 3587
rect 60332 3556 60381 3584
rect 60332 3544 60338 3556
rect 60369 3553 60381 3556
rect 60415 3553 60427 3587
rect 60369 3547 60427 3553
rect 57054 3516 57060 3528
rect 45520 3488 52500 3516
rect 52564 3488 57060 3516
rect 45520 3476 45526 3488
rect 46382 3408 46388 3460
rect 46440 3448 46446 3460
rect 46661 3451 46719 3457
rect 46661 3448 46673 3451
rect 46440 3420 46673 3448
rect 46440 3408 46446 3420
rect 46661 3417 46673 3420
rect 46707 3417 46719 3451
rect 46661 3411 46719 3417
rect 44324 3352 45324 3380
rect 46676 3380 46704 3411
rect 46842 3408 46848 3460
rect 46900 3448 46906 3460
rect 50246 3448 50252 3460
rect 46900 3420 50252 3448
rect 46900 3408 46906 3420
rect 50246 3408 50252 3420
rect 50304 3408 50310 3460
rect 50614 3408 50620 3460
rect 50672 3448 50678 3460
rect 50801 3451 50859 3457
rect 50801 3448 50813 3451
rect 50672 3420 50813 3448
rect 50672 3408 50678 3420
rect 50801 3417 50813 3420
rect 50847 3417 50859 3451
rect 50801 3411 50859 3417
rect 51166 3408 51172 3460
rect 51224 3448 51230 3460
rect 52086 3448 52092 3460
rect 51224 3420 52092 3448
rect 51224 3408 51230 3420
rect 52086 3408 52092 3420
rect 52144 3408 52150 3460
rect 52472 3448 52500 3488
rect 57054 3476 57060 3488
rect 57112 3476 57118 3528
rect 57974 3476 57980 3528
rect 58032 3516 58038 3528
rect 58621 3519 58679 3525
rect 58621 3516 58633 3519
rect 58032 3488 58633 3516
rect 58032 3476 58038 3488
rect 58621 3485 58633 3488
rect 58667 3516 58679 3519
rect 59354 3516 59360 3528
rect 58667 3488 59360 3516
rect 58667 3485 58679 3488
rect 58621 3479 58679 3485
rect 59354 3476 59360 3488
rect 59412 3476 59418 3528
rect 59814 3476 59820 3528
rect 59872 3516 59878 3528
rect 62298 3516 62304 3528
rect 59872 3488 62304 3516
rect 59872 3476 59878 3488
rect 62298 3476 62304 3488
rect 62356 3476 62362 3528
rect 53834 3448 53840 3460
rect 52472 3420 53840 3448
rect 53834 3408 53840 3420
rect 53892 3408 53898 3460
rect 53926 3408 53932 3460
rect 53984 3448 53990 3460
rect 61286 3448 61292 3460
rect 53984 3420 61292 3448
rect 53984 3408 53990 3420
rect 61286 3408 61292 3420
rect 61344 3408 61350 3460
rect 47302 3380 47308 3392
rect 46676 3352 47308 3380
rect 44324 3340 44330 3352
rect 47302 3340 47308 3352
rect 47360 3340 47366 3392
rect 47489 3383 47547 3389
rect 47489 3349 47501 3383
rect 47535 3380 47547 3383
rect 48409 3383 48467 3389
rect 48409 3380 48421 3383
rect 47535 3352 48421 3380
rect 47535 3349 47547 3352
rect 47489 3343 47547 3349
rect 48409 3349 48421 3352
rect 48455 3380 48467 3383
rect 48682 3380 48688 3392
rect 48455 3352 48688 3380
rect 48455 3349 48467 3352
rect 48409 3343 48467 3349
rect 48682 3340 48688 3352
rect 48740 3340 48746 3392
rect 49326 3340 49332 3392
rect 49384 3380 49390 3392
rect 49513 3383 49571 3389
rect 49513 3380 49525 3383
rect 49384 3352 49525 3380
rect 49384 3340 49390 3352
rect 49513 3349 49525 3352
rect 49559 3349 49571 3383
rect 51534 3380 51540 3392
rect 51495 3352 51540 3380
rect 49513 3343 49571 3349
rect 51534 3340 51540 3352
rect 51592 3340 51598 3392
rect 51810 3340 51816 3392
rect 51868 3380 51874 3392
rect 52454 3380 52460 3392
rect 51868 3352 52460 3380
rect 51868 3340 51874 3352
rect 52454 3340 52460 3352
rect 52512 3340 52518 3392
rect 52638 3340 52644 3392
rect 52696 3380 52702 3392
rect 53009 3383 53067 3389
rect 53009 3380 53021 3383
rect 52696 3352 53021 3380
rect 52696 3340 52702 3352
rect 53009 3349 53021 3352
rect 53055 3349 53067 3383
rect 53009 3343 53067 3349
rect 53282 3340 53288 3392
rect 53340 3380 53346 3392
rect 58526 3380 58532 3392
rect 53340 3352 58532 3380
rect 53340 3340 53346 3352
rect 58526 3340 58532 3352
rect 58584 3340 58590 3392
rect 59814 3340 59820 3392
rect 59872 3380 59878 3392
rect 60461 3383 60519 3389
rect 60461 3380 60473 3383
rect 59872 3352 60473 3380
rect 59872 3340 59878 3352
rect 60461 3349 60473 3352
rect 60507 3349 60519 3383
rect 60461 3343 60519 3349
rect 60550 3340 60556 3392
rect 60608 3380 60614 3392
rect 61105 3383 61163 3389
rect 61105 3380 61117 3383
rect 60608 3352 61117 3380
rect 60608 3340 60614 3352
rect 61105 3349 61117 3352
rect 61151 3349 61163 3383
rect 61105 3343 61163 3349
rect 61565 3383 61623 3389
rect 61565 3349 61577 3383
rect 61611 3380 61623 3383
rect 62206 3380 62212 3392
rect 61611 3352 62212 3380
rect 61611 3349 61623 3352
rect 61565 3343 61623 3349
rect 62206 3340 62212 3352
rect 62264 3340 62270 3392
rect 1104 3290 63480 3312
rect 1104 3238 11378 3290
rect 11430 3238 11442 3290
rect 11494 3238 11506 3290
rect 11558 3238 11570 3290
rect 11622 3238 32170 3290
rect 32222 3238 32234 3290
rect 32286 3238 32298 3290
rect 32350 3238 32362 3290
rect 32414 3238 52962 3290
rect 53014 3238 53026 3290
rect 53078 3238 53090 3290
rect 53142 3238 53154 3290
rect 53206 3238 63480 3290
rect 1104 3216 63480 3238
rect 2685 3179 2743 3185
rect 2685 3145 2697 3179
rect 2731 3176 2743 3179
rect 2774 3176 2780 3188
rect 2731 3148 2780 3176
rect 2731 3145 2743 3148
rect 2685 3139 2743 3145
rect 2774 3136 2780 3148
rect 2832 3136 2838 3188
rect 2866 3136 2872 3188
rect 2924 3176 2930 3188
rect 2961 3179 3019 3185
rect 2961 3176 2973 3179
rect 2924 3148 2973 3176
rect 2924 3136 2930 3148
rect 2961 3145 2973 3148
rect 3007 3145 3019 3179
rect 2961 3139 3019 3145
rect 3878 3136 3884 3188
rect 3936 3176 3942 3188
rect 5077 3179 5135 3185
rect 5077 3176 5089 3179
rect 3936 3148 5089 3176
rect 3936 3136 3942 3148
rect 5077 3145 5089 3148
rect 5123 3145 5135 3179
rect 5902 3176 5908 3188
rect 5863 3148 5908 3176
rect 5077 3139 5135 3145
rect 5902 3136 5908 3148
rect 5960 3136 5966 3188
rect 6365 3179 6423 3185
rect 6365 3145 6377 3179
rect 6411 3176 6423 3179
rect 6638 3176 6644 3188
rect 6411 3148 6644 3176
rect 6411 3145 6423 3148
rect 6365 3139 6423 3145
rect 6638 3136 6644 3148
rect 6696 3136 6702 3188
rect 7742 3136 7748 3188
rect 7800 3176 7806 3188
rect 8297 3179 8355 3185
rect 8297 3176 8309 3179
rect 7800 3148 8309 3176
rect 7800 3136 7806 3148
rect 8297 3145 8309 3148
rect 8343 3176 8355 3179
rect 10229 3179 10287 3185
rect 10229 3176 10241 3179
rect 8343 3148 10241 3176
rect 8343 3145 8355 3148
rect 8297 3139 8355 3145
rect 10229 3145 10241 3148
rect 10275 3145 10287 3179
rect 10229 3139 10287 3145
rect 10873 3179 10931 3185
rect 10873 3145 10885 3179
rect 10919 3176 10931 3179
rect 11238 3176 11244 3188
rect 10919 3148 11244 3176
rect 10919 3145 10931 3148
rect 10873 3139 10931 3145
rect 11238 3136 11244 3148
rect 11296 3136 11302 3188
rect 11609 3179 11667 3185
rect 11609 3145 11621 3179
rect 11655 3176 11667 3179
rect 11885 3179 11943 3185
rect 11885 3176 11897 3179
rect 11655 3148 11897 3176
rect 11655 3145 11667 3148
rect 11609 3139 11667 3145
rect 11885 3145 11897 3148
rect 11931 3176 11943 3179
rect 12526 3176 12532 3188
rect 11931 3148 12532 3176
rect 11931 3145 11943 3148
rect 11885 3139 11943 3145
rect 12526 3136 12532 3148
rect 12584 3136 12590 3188
rect 14458 3176 14464 3188
rect 14419 3148 14464 3176
rect 14458 3136 14464 3148
rect 14516 3136 14522 3188
rect 15654 3136 15660 3188
rect 15712 3176 15718 3188
rect 16761 3179 16819 3185
rect 16761 3176 16773 3179
rect 15712 3148 16773 3176
rect 15712 3136 15718 3148
rect 16761 3145 16773 3148
rect 16807 3145 16819 3179
rect 17770 3176 17776 3188
rect 17731 3148 17776 3176
rect 16761 3139 16819 3145
rect 3602 3068 3608 3120
rect 3660 3108 3666 3120
rect 3660 3080 3740 3108
rect 3660 3068 3666 3080
rect 3712 3049 3740 3080
rect 6822 3068 6828 3120
rect 6880 3108 6886 3120
rect 13262 3108 13268 3120
rect 6880 3080 13268 3108
rect 6880 3068 6886 3080
rect 13262 3068 13268 3080
rect 13320 3068 13326 3120
rect 13814 3108 13820 3120
rect 13556 3080 13820 3108
rect 3697 3043 3755 3049
rect 3697 3009 3709 3043
rect 3743 3009 3755 3043
rect 3973 3043 4031 3049
rect 3973 3040 3985 3043
rect 3697 3003 3755 3009
rect 3804 3012 3985 3040
rect 2314 2972 2320 2984
rect 2275 2944 2320 2972
rect 2314 2932 2320 2944
rect 2372 2932 2378 2984
rect 3605 2975 3663 2981
rect 3605 2941 3617 2975
rect 3651 2972 3663 2975
rect 3804 2972 3832 3012
rect 3973 3009 3985 3012
rect 4019 3040 4031 3043
rect 5350 3040 5356 3052
rect 4019 3012 5356 3040
rect 4019 3009 4031 3012
rect 3973 3003 4031 3009
rect 5350 3000 5356 3012
rect 5408 3000 5414 3052
rect 7190 3000 7196 3052
rect 7248 3040 7254 3052
rect 7377 3043 7435 3049
rect 7377 3040 7389 3043
rect 7248 3012 7389 3040
rect 7248 3000 7254 3012
rect 7377 3009 7389 3012
rect 7423 3040 7435 3043
rect 7742 3040 7748 3052
rect 7423 3012 7748 3040
rect 7423 3009 7435 3012
rect 7377 3003 7435 3009
rect 7742 3000 7748 3012
rect 7800 3000 7806 3052
rect 7926 3040 7932 3052
rect 7887 3012 7932 3040
rect 7926 3000 7932 3012
rect 7984 3000 7990 3052
rect 8386 3000 8392 3052
rect 8444 3040 8450 3052
rect 8665 3043 8723 3049
rect 8665 3040 8677 3043
rect 8444 3012 8677 3040
rect 8444 3000 8450 3012
rect 8665 3009 8677 3012
rect 8711 3009 8723 3043
rect 8665 3003 8723 3009
rect 9306 3000 9312 3052
rect 9364 3040 9370 3052
rect 9493 3043 9551 3049
rect 9493 3040 9505 3043
rect 9364 3012 9505 3040
rect 9364 3000 9370 3012
rect 9493 3009 9505 3012
rect 9539 3009 9551 3043
rect 9493 3003 9551 3009
rect 9582 3000 9588 3052
rect 9640 3040 9646 3052
rect 9953 3043 10011 3049
rect 9953 3040 9965 3043
rect 9640 3012 9965 3040
rect 9640 3000 9646 3012
rect 9953 3009 9965 3012
rect 9999 3009 10011 3043
rect 10410 3040 10416 3052
rect 9953 3003 10011 3009
rect 10060 3012 10416 3040
rect 3651 2944 3832 2972
rect 3651 2941 3663 2944
rect 3605 2935 3663 2941
rect 5902 2932 5908 2984
rect 5960 2972 5966 2984
rect 7469 2975 7527 2981
rect 7469 2972 7481 2975
rect 5960 2944 7481 2972
rect 5960 2932 5966 2944
rect 7469 2941 7481 2944
rect 7515 2972 7527 2975
rect 7650 2972 7656 2984
rect 7515 2944 7656 2972
rect 7515 2941 7527 2944
rect 7469 2935 7527 2941
rect 7650 2932 7656 2944
rect 7708 2932 7714 2984
rect 7834 2972 7840 2984
rect 7795 2944 7840 2972
rect 7834 2932 7840 2944
rect 7892 2932 7898 2984
rect 9030 2932 9036 2984
rect 9088 2972 9094 2984
rect 9415 2975 9473 2981
rect 9415 2972 9427 2975
rect 9088 2944 9427 2972
rect 9088 2932 9094 2944
rect 9415 2941 9427 2944
rect 9461 2941 9473 2975
rect 9415 2935 9473 2941
rect 9766 2932 9772 2984
rect 9824 2972 9830 2984
rect 9861 2975 9919 2981
rect 9861 2972 9873 2975
rect 9824 2944 9873 2972
rect 9824 2932 9830 2944
rect 9861 2941 9873 2944
rect 9907 2972 9919 2975
rect 10060 2972 10088 3012
rect 10410 3000 10416 3012
rect 10468 3000 10474 3052
rect 11517 3043 11575 3049
rect 11517 3009 11529 3043
rect 11563 3040 11575 3043
rect 12342 3040 12348 3052
rect 11563 3012 12348 3040
rect 11563 3009 11575 3012
rect 11517 3003 11575 3009
rect 12342 3000 12348 3012
rect 12400 3000 12406 3052
rect 12713 3043 12771 3049
rect 12713 3009 12725 3043
rect 12759 3040 12771 3043
rect 12802 3040 12808 3052
rect 12759 3012 12808 3040
rect 12759 3009 12771 3012
rect 12713 3003 12771 3009
rect 12802 3000 12808 3012
rect 12860 3000 12866 3052
rect 13556 3040 13584 3080
rect 13814 3068 13820 3080
rect 13872 3068 13878 3120
rect 16206 3068 16212 3120
rect 16264 3108 16270 3120
rect 16393 3111 16451 3117
rect 16393 3108 16405 3111
rect 16264 3080 16405 3108
rect 16264 3068 16270 3080
rect 16393 3077 16405 3080
rect 16439 3077 16451 3111
rect 16776 3108 16804 3139
rect 17770 3136 17776 3148
rect 17828 3136 17834 3188
rect 18046 3176 18052 3188
rect 18007 3148 18052 3176
rect 18046 3136 18052 3148
rect 18104 3136 18110 3188
rect 18138 3136 18144 3188
rect 18196 3176 18202 3188
rect 21266 3176 21272 3188
rect 18196 3148 20852 3176
rect 21227 3148 21272 3176
rect 18196 3136 18202 3148
rect 18690 3108 18696 3120
rect 16776 3080 18696 3108
rect 16393 3071 16451 3077
rect 18690 3068 18696 3080
rect 18748 3068 18754 3120
rect 18966 3068 18972 3120
rect 19024 3108 19030 3120
rect 19024 3080 20576 3108
rect 19024 3068 19030 3080
rect 13722 3040 13728 3052
rect 13280 3012 13584 3040
rect 13683 3012 13728 3040
rect 9907 2944 10088 2972
rect 10229 2975 10287 2981
rect 9907 2941 9919 2944
rect 9861 2935 9919 2941
rect 10229 2941 10241 2975
rect 10275 2972 10287 2975
rect 11146 2972 11152 2984
rect 10275 2944 11008 2972
rect 11107 2944 11152 2972
rect 10275 2941 10287 2944
rect 10229 2935 10287 2941
rect 4706 2864 4712 2916
rect 4764 2904 4770 2916
rect 6825 2907 6883 2913
rect 6825 2904 6837 2907
rect 4764 2876 6837 2904
rect 4764 2864 4770 2876
rect 6825 2873 6837 2876
rect 6871 2873 6883 2907
rect 6825 2867 6883 2873
rect 8110 2864 8116 2916
rect 8168 2904 8174 2916
rect 8849 2907 8907 2913
rect 8849 2904 8861 2907
rect 8168 2876 8861 2904
rect 8168 2864 8174 2876
rect 8849 2873 8861 2876
rect 8895 2873 8907 2907
rect 8849 2867 8907 2873
rect 9582 2864 9588 2916
rect 9640 2904 9646 2916
rect 10980 2913 11008 2944
rect 11146 2932 11152 2944
rect 11204 2932 11210 2984
rect 12250 2972 12256 2984
rect 12211 2944 12256 2972
rect 12250 2932 12256 2944
rect 12308 2932 12314 2984
rect 13280 2981 13308 3012
rect 13722 3000 13728 3012
rect 13780 3040 13786 3052
rect 14001 3043 14059 3049
rect 14001 3040 14013 3043
rect 13780 3012 14013 3040
rect 13780 3000 13786 3012
rect 14001 3009 14013 3012
rect 14047 3009 14059 3043
rect 14001 3003 14059 3009
rect 14829 3043 14887 3049
rect 14829 3009 14841 3043
rect 14875 3040 14887 3043
rect 15657 3043 15715 3049
rect 15657 3040 15669 3043
rect 14875 3012 15669 3040
rect 14875 3009 14887 3012
rect 14829 3003 14887 3009
rect 15657 3009 15669 3012
rect 15703 3040 15715 3043
rect 18785 3043 18843 3049
rect 18785 3040 18797 3043
rect 15703 3012 18797 3040
rect 15703 3009 15715 3012
rect 15657 3003 15715 3009
rect 18785 3009 18797 3012
rect 18831 3009 18843 3043
rect 18785 3003 18843 3009
rect 19058 3000 19064 3052
rect 19116 3040 19122 3052
rect 20346 3040 20352 3052
rect 19116 3012 20352 3040
rect 19116 3000 19122 3012
rect 20346 3000 20352 3012
rect 20404 3000 20410 3052
rect 13265 2975 13323 2981
rect 13265 2941 13277 2975
rect 13311 2941 13323 2975
rect 13265 2935 13323 2941
rect 13541 2975 13599 2981
rect 13541 2941 13553 2975
rect 13587 2941 13599 2975
rect 13541 2935 13599 2941
rect 10965 2907 11023 2913
rect 9640 2876 10916 2904
rect 9640 2864 9646 2876
rect 1949 2839 2007 2845
rect 1949 2805 1961 2839
rect 1995 2836 2007 2839
rect 2130 2836 2136 2848
rect 1995 2808 2136 2836
rect 1995 2805 2007 2808
rect 1949 2799 2007 2805
rect 2130 2796 2136 2808
rect 2188 2796 2194 2848
rect 8294 2796 8300 2848
rect 8352 2836 8358 2848
rect 10318 2836 10324 2848
rect 8352 2808 10324 2836
rect 8352 2796 8358 2808
rect 10318 2796 10324 2808
rect 10376 2796 10382 2848
rect 10888 2836 10916 2876
rect 10965 2873 10977 2907
rect 11011 2904 11023 2907
rect 11609 2907 11667 2913
rect 11609 2904 11621 2907
rect 11011 2876 11621 2904
rect 11011 2873 11023 2876
rect 10965 2867 11023 2873
rect 11609 2873 11621 2876
rect 11655 2873 11667 2907
rect 13446 2904 13452 2916
rect 11609 2867 11667 2873
rect 12084 2876 13452 2904
rect 12084 2836 12112 2876
rect 13446 2864 13452 2876
rect 13504 2864 13510 2916
rect 13556 2904 13584 2935
rect 15010 2932 15016 2984
rect 15068 2972 15074 2984
rect 15565 2975 15623 2981
rect 15565 2972 15577 2975
rect 15068 2944 15577 2972
rect 15068 2932 15074 2944
rect 15565 2941 15577 2944
rect 15611 2941 15623 2975
rect 15930 2972 15936 2984
rect 15891 2944 15936 2972
rect 15565 2935 15623 2941
rect 15930 2932 15936 2944
rect 15988 2932 15994 2984
rect 16114 2972 16120 2984
rect 16075 2944 16120 2972
rect 16114 2932 16120 2944
rect 16172 2932 16178 2984
rect 16390 2932 16396 2984
rect 16448 2972 16454 2984
rect 18046 2972 18052 2984
rect 16448 2944 18052 2972
rect 16448 2932 16454 2944
rect 18046 2932 18052 2944
rect 18104 2932 18110 2984
rect 18322 2972 18328 2984
rect 18283 2944 18328 2972
rect 18322 2932 18328 2944
rect 18380 2932 18386 2984
rect 19889 2975 19947 2981
rect 19889 2941 19901 2975
rect 19935 2941 19947 2975
rect 20070 2972 20076 2984
rect 20031 2944 20076 2972
rect 19889 2935 19947 2941
rect 14090 2904 14096 2916
rect 13556 2876 14096 2904
rect 14090 2864 14096 2876
rect 14148 2864 14154 2916
rect 14921 2907 14979 2913
rect 14921 2873 14933 2907
rect 14967 2904 14979 2907
rect 15194 2904 15200 2916
rect 14967 2876 15200 2904
rect 14967 2873 14979 2876
rect 14921 2867 14979 2873
rect 15194 2864 15200 2876
rect 15252 2864 15258 2916
rect 15378 2864 15384 2916
rect 15436 2904 15442 2916
rect 16132 2904 16160 2932
rect 17402 2904 17408 2916
rect 15436 2876 16160 2904
rect 16316 2876 17408 2904
rect 15436 2864 15442 2876
rect 10888 2808 12112 2836
rect 14550 2796 14556 2848
rect 14608 2836 14614 2848
rect 16316 2836 16344 2876
rect 17402 2864 17408 2876
rect 17460 2864 17466 2916
rect 17678 2864 17684 2916
rect 17736 2904 17742 2916
rect 17862 2904 17868 2916
rect 17736 2876 17868 2904
rect 17736 2864 17742 2876
rect 17862 2864 17868 2876
rect 17920 2904 17926 2916
rect 18233 2907 18291 2913
rect 18233 2904 18245 2907
rect 17920 2876 18245 2904
rect 17920 2864 17926 2876
rect 18233 2873 18245 2876
rect 18279 2904 18291 2907
rect 19061 2907 19119 2913
rect 19061 2904 19073 2907
rect 18279 2876 19073 2904
rect 18279 2873 18291 2876
rect 18233 2867 18291 2873
rect 19061 2873 19073 2876
rect 19107 2873 19119 2907
rect 19904 2904 19932 2935
rect 20070 2932 20076 2944
rect 20128 2932 20134 2984
rect 20162 2932 20168 2984
rect 20220 2972 20226 2984
rect 20548 2972 20576 3080
rect 20625 3043 20683 3049
rect 20625 3009 20637 3043
rect 20671 3040 20683 3043
rect 20714 3040 20720 3052
rect 20671 3012 20720 3040
rect 20671 3009 20683 3012
rect 20625 3003 20683 3009
rect 20714 3000 20720 3012
rect 20772 3000 20778 3052
rect 20824 3040 20852 3148
rect 21266 3136 21272 3148
rect 21324 3136 21330 3188
rect 21453 3179 21511 3185
rect 21453 3145 21465 3179
rect 21499 3176 21511 3179
rect 22646 3176 22652 3188
rect 21499 3148 22652 3176
rect 21499 3145 21511 3148
rect 21453 3139 21511 3145
rect 22646 3136 22652 3148
rect 22704 3136 22710 3188
rect 23474 3136 23480 3188
rect 23532 3176 23538 3188
rect 25314 3176 25320 3188
rect 23532 3148 23796 3176
rect 25275 3148 25320 3176
rect 23532 3136 23538 3148
rect 21542 3068 21548 3120
rect 21600 3108 21606 3120
rect 21637 3111 21695 3117
rect 21637 3108 21649 3111
rect 21600 3080 21649 3108
rect 21600 3068 21606 3080
rect 21637 3077 21649 3080
rect 21683 3077 21695 3111
rect 21637 3071 21695 3077
rect 21818 3068 21824 3120
rect 21876 3108 21882 3120
rect 21876 3080 22508 3108
rect 21876 3068 21882 3080
rect 22094 3040 22100 3052
rect 20824 3012 22100 3040
rect 22094 3000 22100 3012
rect 22152 3000 22158 3052
rect 22281 3043 22339 3049
rect 22281 3009 22293 3043
rect 22327 3040 22339 3043
rect 22370 3040 22376 3052
rect 22327 3012 22376 3040
rect 22327 3009 22339 3012
rect 22281 3003 22339 3009
rect 22370 3000 22376 3012
rect 22428 3000 22434 3052
rect 22480 3040 22508 3080
rect 23106 3040 23112 3052
rect 22480 3012 23112 3040
rect 21453 2975 21511 2981
rect 21453 2972 21465 2975
rect 20220 2944 20265 2972
rect 20548 2944 21465 2972
rect 20220 2932 20226 2944
rect 21453 2941 21465 2944
rect 21499 2941 21511 2975
rect 21453 2935 21511 2941
rect 22189 2975 22247 2981
rect 22189 2941 22201 2975
rect 22235 2972 22247 2975
rect 22480 2972 22508 3012
rect 23106 3000 23112 3012
rect 23164 3000 23170 3052
rect 23477 3043 23535 3049
rect 23477 3009 23489 3043
rect 23523 3040 23535 3043
rect 23566 3040 23572 3052
rect 23523 3012 23572 3040
rect 23523 3009 23535 3012
rect 23477 3003 23535 3009
rect 23566 3000 23572 3012
rect 23624 3000 23630 3052
rect 23768 3049 23796 3148
rect 25314 3136 25320 3148
rect 25372 3136 25378 3188
rect 27430 3176 27436 3188
rect 25516 3148 27436 3176
rect 24486 3068 24492 3120
rect 24544 3108 24550 3120
rect 25516 3108 25544 3148
rect 27430 3136 27436 3148
rect 27488 3136 27494 3188
rect 28166 3176 28172 3188
rect 27724 3148 28172 3176
rect 24544 3080 25544 3108
rect 25593 3111 25651 3117
rect 24544 3068 24550 3080
rect 25593 3077 25605 3111
rect 25639 3108 25651 3111
rect 27724 3108 27752 3148
rect 28166 3136 28172 3148
rect 28224 3136 28230 3188
rect 28258 3136 28264 3188
rect 28316 3176 28322 3188
rect 28353 3179 28411 3185
rect 28353 3176 28365 3179
rect 28316 3148 28365 3176
rect 28316 3136 28322 3148
rect 28353 3145 28365 3148
rect 28399 3145 28411 3179
rect 28353 3139 28411 3145
rect 28718 3136 28724 3188
rect 28776 3176 28782 3188
rect 32030 3176 32036 3188
rect 28776 3148 32036 3176
rect 28776 3136 28782 3148
rect 32030 3136 32036 3148
rect 32088 3136 32094 3188
rect 32217 3179 32275 3185
rect 32217 3145 32229 3179
rect 32263 3176 32275 3179
rect 32674 3176 32680 3188
rect 32263 3148 32680 3176
rect 32263 3145 32275 3148
rect 32217 3139 32275 3145
rect 32674 3136 32680 3148
rect 32732 3176 32738 3188
rect 34514 3176 34520 3188
rect 32732 3148 34520 3176
rect 32732 3136 32738 3148
rect 34514 3136 34520 3148
rect 34572 3136 34578 3188
rect 34698 3176 34704 3188
rect 34659 3148 34704 3176
rect 34698 3136 34704 3148
rect 34756 3136 34762 3188
rect 35621 3179 35679 3185
rect 35621 3145 35633 3179
rect 35667 3176 35679 3179
rect 38010 3176 38016 3188
rect 35667 3148 38016 3176
rect 35667 3145 35679 3148
rect 35621 3139 35679 3145
rect 38010 3136 38016 3148
rect 38068 3136 38074 3188
rect 38105 3179 38163 3185
rect 38105 3145 38117 3179
rect 38151 3176 38163 3179
rect 41230 3176 41236 3188
rect 38151 3148 41236 3176
rect 38151 3145 38163 3148
rect 38105 3139 38163 3145
rect 41230 3136 41236 3148
rect 41288 3136 41294 3188
rect 42058 3136 42064 3188
rect 42116 3176 42122 3188
rect 42705 3179 42763 3185
rect 42116 3148 42161 3176
rect 42116 3136 42122 3148
rect 42705 3145 42717 3179
rect 42751 3176 42763 3179
rect 43438 3176 43444 3188
rect 42751 3148 43444 3176
rect 42751 3145 42763 3148
rect 42705 3139 42763 3145
rect 43438 3136 43444 3148
rect 43496 3136 43502 3188
rect 43622 3136 43628 3188
rect 43680 3176 43686 3188
rect 43990 3176 43996 3188
rect 43680 3148 43996 3176
rect 43680 3136 43686 3148
rect 43990 3136 43996 3148
rect 44048 3176 44054 3188
rect 45465 3179 45523 3185
rect 45465 3176 45477 3179
rect 44048 3148 45477 3176
rect 44048 3136 44054 3148
rect 45465 3145 45477 3148
rect 45511 3145 45523 3179
rect 45465 3139 45523 3145
rect 46106 3136 46112 3188
rect 46164 3176 46170 3188
rect 48590 3176 48596 3188
rect 46164 3148 48596 3176
rect 46164 3136 46170 3148
rect 48590 3136 48596 3148
rect 48648 3176 48654 3188
rect 48777 3179 48835 3185
rect 48777 3176 48789 3179
rect 48648 3148 48789 3176
rect 48648 3136 48654 3148
rect 48777 3145 48789 3148
rect 48823 3145 48835 3179
rect 48777 3139 48835 3145
rect 49237 3179 49295 3185
rect 49237 3145 49249 3179
rect 49283 3176 49295 3179
rect 50062 3176 50068 3188
rect 49283 3148 50068 3176
rect 49283 3145 49295 3148
rect 49237 3139 49295 3145
rect 50062 3136 50068 3148
rect 50120 3136 50126 3188
rect 51537 3179 51595 3185
rect 51537 3145 51549 3179
rect 51583 3176 51595 3179
rect 52362 3176 52368 3188
rect 51583 3148 52368 3176
rect 51583 3145 51595 3148
rect 51537 3139 51595 3145
rect 52362 3136 52368 3148
rect 52420 3136 52426 3188
rect 52549 3179 52607 3185
rect 52549 3145 52561 3179
rect 52595 3176 52607 3179
rect 52638 3176 52644 3188
rect 52595 3148 52644 3176
rect 52595 3145 52607 3148
rect 52549 3139 52607 3145
rect 52638 3136 52644 3148
rect 52696 3136 52702 3188
rect 53834 3176 53840 3188
rect 53795 3148 53840 3176
rect 53834 3136 53840 3148
rect 53892 3136 53898 3188
rect 54662 3136 54668 3188
rect 54720 3176 54726 3188
rect 55122 3176 55128 3188
rect 54720 3148 55128 3176
rect 54720 3136 54726 3148
rect 55122 3136 55128 3148
rect 55180 3176 55186 3188
rect 55953 3179 56011 3185
rect 55953 3176 55965 3179
rect 55180 3148 55965 3176
rect 55180 3136 55186 3148
rect 55953 3145 55965 3148
rect 55999 3145 56011 3179
rect 56318 3176 56324 3188
rect 56279 3148 56324 3176
rect 55953 3139 56011 3145
rect 56318 3136 56324 3148
rect 56376 3136 56382 3188
rect 56502 3136 56508 3188
rect 56560 3176 56566 3188
rect 56689 3179 56747 3185
rect 56689 3176 56701 3179
rect 56560 3148 56701 3176
rect 56560 3136 56566 3148
rect 56689 3145 56701 3148
rect 56735 3145 56747 3179
rect 56689 3139 56747 3145
rect 57149 3179 57207 3185
rect 57149 3145 57161 3179
rect 57195 3176 57207 3179
rect 57238 3176 57244 3188
rect 57195 3148 57244 3176
rect 57195 3145 57207 3148
rect 57149 3139 57207 3145
rect 57238 3136 57244 3148
rect 57296 3136 57302 3188
rect 57606 3176 57612 3188
rect 57567 3148 57612 3176
rect 57606 3136 57612 3148
rect 57664 3136 57670 3188
rect 57974 3136 57980 3188
rect 58032 3176 58038 3188
rect 58618 3176 58624 3188
rect 58032 3148 58077 3176
rect 58579 3148 58624 3176
rect 58032 3136 58038 3148
rect 58618 3136 58624 3148
rect 58676 3136 58682 3188
rect 58897 3179 58955 3185
rect 58897 3145 58909 3179
rect 58943 3176 58955 3179
rect 59538 3176 59544 3188
rect 58943 3148 59544 3176
rect 58943 3145 58955 3148
rect 58897 3139 58955 3145
rect 59538 3136 59544 3148
rect 59596 3136 59602 3188
rect 60550 3136 60556 3188
rect 60608 3176 60614 3188
rect 61105 3179 61163 3185
rect 61105 3176 61117 3179
rect 60608 3148 61117 3176
rect 60608 3136 60614 3148
rect 61105 3145 61117 3148
rect 61151 3145 61163 3179
rect 61286 3176 61292 3188
rect 61247 3148 61292 3176
rect 61105 3139 61163 3145
rect 61286 3136 61292 3148
rect 61344 3136 61350 3188
rect 62298 3176 62304 3188
rect 62259 3148 62304 3176
rect 62298 3136 62304 3148
rect 62356 3136 62362 3188
rect 25639 3080 27752 3108
rect 25639 3077 25651 3080
rect 25593 3071 25651 3077
rect 27798 3068 27804 3120
rect 27856 3108 27862 3120
rect 27856 3080 29776 3108
rect 27856 3068 27862 3080
rect 23753 3043 23811 3049
rect 23753 3009 23765 3043
rect 23799 3009 23811 3043
rect 23753 3003 23811 3009
rect 25222 3000 25228 3052
rect 25280 3040 25286 3052
rect 25685 3043 25743 3049
rect 25685 3040 25697 3043
rect 25280 3012 25697 3040
rect 25280 3000 25286 3012
rect 25685 3009 25697 3012
rect 25731 3009 25743 3043
rect 25685 3003 25743 3009
rect 26513 3043 26571 3049
rect 26513 3009 26525 3043
rect 26559 3040 26571 3043
rect 27341 3043 27399 3049
rect 27341 3040 27353 3043
rect 26559 3012 27353 3040
rect 26559 3009 26571 3012
rect 26513 3003 26571 3009
rect 27341 3009 27353 3012
rect 27387 3040 27399 3043
rect 28350 3040 28356 3052
rect 27387 3012 28356 3040
rect 27387 3009 27399 3012
rect 27341 3003 27399 3009
rect 28350 3000 28356 3012
rect 28408 3000 28414 3052
rect 28442 3000 28448 3052
rect 28500 3040 28506 3052
rect 29748 3049 29776 3080
rect 30742 3068 30748 3120
rect 30800 3108 30806 3120
rect 31481 3111 31539 3117
rect 31481 3108 31493 3111
rect 30800 3080 31493 3108
rect 30800 3068 30806 3080
rect 31481 3077 31493 3080
rect 31527 3077 31539 3111
rect 31481 3071 31539 3077
rect 31846 3068 31852 3120
rect 31904 3108 31910 3120
rect 32122 3108 32128 3120
rect 31904 3080 32128 3108
rect 31904 3068 31910 3080
rect 32122 3068 32128 3080
rect 32180 3068 32186 3120
rect 33318 3068 33324 3120
rect 33376 3108 33382 3120
rect 35069 3111 35127 3117
rect 35069 3108 35081 3111
rect 33376 3080 35081 3108
rect 33376 3068 33382 3080
rect 35069 3077 35081 3080
rect 35115 3108 35127 3111
rect 37458 3108 37464 3120
rect 35115 3080 37464 3108
rect 35115 3077 35127 3080
rect 35069 3071 35127 3077
rect 37458 3068 37464 3080
rect 37516 3068 37522 3120
rect 37829 3111 37887 3117
rect 37829 3077 37841 3111
rect 37875 3108 37887 3111
rect 39758 3108 39764 3120
rect 37875 3080 39764 3108
rect 37875 3077 37887 3080
rect 37829 3071 37887 3077
rect 39758 3068 39764 3080
rect 39816 3068 39822 3120
rect 39942 3108 39948 3120
rect 39903 3080 39948 3108
rect 39942 3068 39948 3080
rect 40000 3068 40006 3120
rect 40310 3108 40316 3120
rect 40271 3080 40316 3108
rect 40310 3068 40316 3080
rect 40368 3068 40374 3120
rect 41966 3068 41972 3120
rect 42024 3108 42030 3120
rect 42797 3111 42855 3117
rect 42797 3108 42809 3111
rect 42024 3080 42809 3108
rect 42024 3068 42030 3080
rect 42797 3077 42809 3080
rect 42843 3077 42855 3111
rect 42797 3071 42855 3077
rect 29733 3043 29791 3049
rect 28500 3012 29592 3040
rect 28500 3000 28506 3012
rect 22235 2944 22508 2972
rect 22235 2941 22247 2944
rect 22189 2935 22247 2941
rect 22554 2932 22560 2984
rect 22612 2972 22618 2984
rect 22738 2972 22744 2984
rect 22612 2944 22657 2972
rect 22699 2944 22744 2972
rect 22612 2932 22618 2944
rect 22738 2932 22744 2944
rect 22796 2932 22802 2984
rect 24578 2972 24584 2984
rect 23032 2944 24584 2972
rect 20438 2904 20444 2916
rect 19904 2876 20444 2904
rect 19061 2867 19119 2873
rect 20438 2864 20444 2876
rect 20496 2904 20502 2916
rect 22830 2904 22836 2916
rect 20496 2876 22836 2904
rect 20496 2864 20502 2876
rect 22830 2864 22836 2876
rect 22888 2864 22894 2916
rect 14608 2808 16344 2836
rect 14608 2796 14614 2808
rect 18690 2796 18696 2848
rect 18748 2836 18754 2848
rect 19429 2839 19487 2845
rect 19429 2836 19441 2839
rect 18748 2808 19441 2836
rect 18748 2796 18754 2808
rect 19429 2805 19441 2808
rect 19475 2805 19487 2839
rect 19429 2799 19487 2805
rect 20714 2796 20720 2848
rect 20772 2836 20778 2848
rect 22186 2836 22192 2848
rect 20772 2808 22192 2836
rect 20772 2796 20778 2808
rect 22186 2796 22192 2808
rect 22244 2796 22250 2848
rect 22554 2796 22560 2848
rect 22612 2836 22618 2848
rect 23032 2845 23060 2944
rect 24578 2932 24584 2944
rect 24636 2932 24642 2984
rect 24719 2975 24777 2981
rect 24719 2941 24731 2975
rect 24765 2972 24777 2975
rect 24854 2972 24860 2984
rect 24765 2944 24860 2972
rect 24765 2941 24777 2944
rect 24719 2935 24777 2941
rect 24854 2932 24860 2944
rect 24912 2932 24918 2984
rect 26970 2932 26976 2984
rect 27028 2972 27034 2984
rect 27249 2975 27307 2981
rect 27249 2972 27261 2975
rect 27028 2944 27261 2972
rect 27028 2932 27034 2944
rect 27249 2941 27261 2944
rect 27295 2941 27307 2975
rect 27249 2935 27307 2941
rect 27617 2975 27675 2981
rect 27617 2941 27629 2975
rect 27663 2941 27675 2975
rect 27617 2935 27675 2941
rect 23845 2907 23903 2913
rect 23845 2873 23857 2907
rect 23891 2904 23903 2907
rect 24302 2904 24308 2916
rect 23891 2876 24308 2904
rect 23891 2873 23903 2876
rect 23845 2867 23903 2873
rect 24302 2864 24308 2876
rect 24360 2904 24366 2916
rect 26053 2907 26111 2913
rect 26053 2904 26065 2907
rect 24360 2876 26065 2904
rect 24360 2864 24366 2876
rect 26053 2873 26065 2876
rect 26099 2873 26111 2907
rect 26602 2904 26608 2916
rect 26563 2876 26608 2904
rect 26053 2867 26111 2873
rect 26602 2864 26608 2876
rect 26660 2864 26666 2916
rect 27632 2904 27660 2935
rect 27706 2932 27712 2984
rect 27764 2972 27770 2984
rect 29270 2972 29276 2984
rect 27764 2944 27809 2972
rect 29231 2944 29276 2972
rect 27764 2932 27770 2944
rect 29270 2932 29276 2944
rect 29328 2932 29334 2984
rect 29454 2972 29460 2984
rect 29415 2944 29460 2972
rect 29454 2932 29460 2944
rect 29512 2932 29518 2984
rect 29564 2972 29592 3012
rect 29733 3009 29745 3043
rect 29779 3009 29791 3043
rect 29733 3003 29791 3009
rect 30190 3000 30196 3052
rect 30248 3040 30254 3052
rect 30837 3043 30895 3049
rect 30837 3040 30849 3043
rect 30248 3012 30849 3040
rect 30248 3000 30254 3012
rect 30837 3009 30849 3012
rect 30883 3040 30895 3043
rect 32490 3040 32496 3052
rect 30883 3012 32496 3040
rect 30883 3009 30895 3012
rect 30837 3003 30895 3009
rect 32490 3000 32496 3012
rect 32548 3000 32554 3052
rect 32585 3043 32643 3049
rect 32585 3009 32597 3043
rect 32631 3040 32643 3043
rect 33962 3040 33968 3052
rect 32631 3012 33548 3040
rect 33923 3012 33968 3040
rect 32631 3009 32643 3012
rect 32585 3003 32643 3009
rect 33520 2984 33548 3012
rect 33962 3000 33968 3012
rect 34020 3000 34026 3052
rect 34057 3043 34115 3049
rect 34057 3009 34069 3043
rect 34103 3040 34115 3043
rect 34333 3043 34391 3049
rect 34333 3040 34345 3043
rect 34103 3012 34345 3040
rect 34103 3009 34115 3012
rect 34057 3003 34115 3009
rect 34333 3009 34345 3012
rect 34379 3040 34391 3043
rect 35621 3043 35679 3049
rect 35621 3040 35633 3043
rect 34379 3012 35633 3040
rect 34379 3009 34391 3012
rect 34333 3003 34391 3009
rect 35621 3009 35633 3012
rect 35667 3009 35679 3043
rect 35621 3003 35679 3009
rect 36081 3043 36139 3049
rect 36081 3009 36093 3043
rect 36127 3040 36139 3043
rect 36722 3040 36728 3052
rect 36127 3012 36728 3040
rect 36127 3009 36139 3012
rect 36081 3003 36139 3009
rect 36722 3000 36728 3012
rect 36780 3000 36786 3052
rect 36906 3000 36912 3052
rect 36964 3040 36970 3052
rect 39577 3043 39635 3049
rect 36964 3012 39160 3040
rect 36964 3000 36970 3012
rect 30285 2975 30343 2981
rect 30285 2972 30297 2975
rect 29564 2944 30297 2972
rect 30285 2941 30297 2944
rect 30331 2941 30343 2975
rect 31018 2972 31024 2984
rect 30979 2944 31024 2972
rect 30285 2935 30343 2941
rect 31018 2932 31024 2944
rect 31076 2972 31082 2984
rect 31202 2972 31208 2984
rect 31076 2944 31208 2972
rect 31076 2932 31082 2944
rect 31202 2932 31208 2944
rect 31260 2932 31266 2984
rect 31478 2972 31484 2984
rect 31439 2944 31484 2972
rect 31478 2932 31484 2944
rect 31536 2932 31542 2984
rect 33226 2972 33232 2984
rect 31956 2944 33232 2972
rect 28813 2907 28871 2913
rect 28813 2904 28825 2907
rect 27632 2876 28825 2904
rect 23017 2839 23075 2845
rect 23017 2836 23029 2839
rect 22612 2808 23029 2836
rect 22612 2796 22618 2808
rect 23017 2805 23029 2808
rect 23063 2805 23075 2839
rect 23017 2799 23075 2805
rect 23382 2796 23388 2848
rect 23440 2836 23446 2848
rect 25593 2839 25651 2845
rect 25593 2836 25605 2839
rect 23440 2808 25605 2836
rect 23440 2796 23446 2808
rect 25593 2805 25605 2808
rect 25639 2805 25651 2839
rect 25593 2799 25651 2805
rect 26510 2796 26516 2848
rect 26568 2836 26574 2848
rect 27632 2836 27660 2876
rect 28813 2873 28825 2876
rect 28859 2904 28871 2907
rect 30469 2907 30527 2913
rect 30469 2904 30481 2907
rect 28859 2876 30481 2904
rect 28859 2873 28871 2876
rect 28813 2867 28871 2873
rect 30469 2873 30481 2876
rect 30515 2904 30527 2907
rect 30558 2904 30564 2916
rect 30515 2876 30564 2904
rect 30515 2873 30527 2876
rect 30469 2867 30527 2873
rect 30558 2864 30564 2876
rect 30616 2904 30622 2916
rect 31956 2904 31984 2944
rect 33226 2932 33232 2944
rect 33284 2972 33290 2984
rect 33321 2975 33379 2981
rect 33321 2972 33333 2975
rect 33284 2944 33333 2972
rect 33284 2932 33290 2944
rect 33321 2941 33333 2944
rect 33367 2941 33379 2975
rect 33502 2972 33508 2984
rect 33415 2944 33508 2972
rect 33321 2935 33379 2941
rect 33502 2932 33508 2944
rect 33560 2932 33566 2984
rect 34790 2932 34796 2984
rect 34848 2972 34854 2984
rect 34885 2975 34943 2981
rect 34885 2972 34897 2975
rect 34848 2944 34897 2972
rect 34848 2932 34854 2944
rect 34885 2941 34897 2944
rect 34931 2972 34943 2975
rect 36262 2972 36268 2984
rect 34931 2944 36124 2972
rect 36223 2944 36268 2972
rect 34931 2941 34943 2944
rect 34885 2935 34943 2941
rect 32674 2904 32680 2916
rect 30616 2876 31984 2904
rect 32048 2876 32680 2904
rect 30616 2864 30622 2876
rect 26568 2808 27660 2836
rect 26568 2796 26574 2808
rect 29454 2796 29460 2848
rect 29512 2836 29518 2848
rect 30101 2839 30159 2845
rect 30101 2836 30113 2839
rect 29512 2808 30113 2836
rect 29512 2796 29518 2808
rect 30101 2805 30113 2808
rect 30147 2805 30159 2839
rect 30101 2799 30159 2805
rect 30285 2839 30343 2845
rect 30285 2805 30297 2839
rect 30331 2836 30343 2839
rect 32048 2836 32076 2876
rect 32674 2864 32680 2876
rect 32732 2864 32738 2916
rect 33410 2904 33416 2916
rect 33323 2876 33416 2904
rect 33410 2864 33416 2876
rect 33468 2864 33474 2916
rect 33520 2904 33548 2932
rect 36096 2904 36124 2944
rect 36262 2932 36268 2944
rect 36320 2932 36326 2984
rect 36354 2932 36360 2984
rect 36412 2972 36418 2984
rect 36412 2944 36457 2972
rect 36412 2932 36418 2944
rect 36538 2932 36544 2984
rect 36596 2972 36602 2984
rect 36817 2975 36875 2981
rect 36817 2972 36829 2975
rect 36596 2944 36829 2972
rect 36596 2932 36602 2944
rect 36817 2941 36829 2944
rect 36863 2941 36875 2975
rect 36817 2935 36875 2941
rect 37734 2932 37740 2984
rect 37792 2972 37798 2984
rect 37921 2975 37979 2981
rect 37921 2972 37933 2975
rect 37792 2944 37933 2972
rect 37792 2932 37798 2944
rect 37921 2941 37933 2944
rect 37967 2941 37979 2975
rect 37921 2935 37979 2941
rect 38010 2932 38016 2984
rect 38068 2972 38074 2984
rect 38838 2972 38844 2984
rect 38068 2944 38844 2972
rect 38068 2932 38074 2944
rect 38838 2932 38844 2944
rect 38896 2932 38902 2984
rect 36170 2904 36176 2916
rect 33520 2876 35848 2904
rect 36096 2876 36176 2904
rect 32950 2836 32956 2848
rect 30331 2808 32076 2836
rect 32911 2808 32956 2836
rect 30331 2805 30343 2808
rect 30285 2799 30343 2805
rect 32950 2796 32956 2808
rect 33008 2796 33014 2848
rect 33428 2836 33456 2864
rect 35820 2845 35848 2876
rect 36170 2864 36176 2876
rect 36228 2864 36234 2916
rect 36449 2907 36507 2913
rect 36449 2873 36461 2907
rect 36495 2873 36507 2907
rect 38470 2904 38476 2916
rect 38431 2876 38476 2904
rect 36449 2867 36507 2873
rect 34057 2839 34115 2845
rect 34057 2836 34069 2839
rect 33428 2808 34069 2836
rect 34057 2805 34069 2808
rect 34103 2805 34115 2839
rect 34057 2799 34115 2805
rect 35805 2839 35863 2845
rect 35805 2805 35817 2839
rect 35851 2836 35863 2839
rect 35894 2836 35900 2848
rect 35851 2808 35900 2836
rect 35851 2805 35863 2808
rect 35805 2799 35863 2805
rect 35894 2796 35900 2808
rect 35952 2796 35958 2848
rect 36464 2836 36492 2867
rect 38470 2864 38476 2876
rect 38528 2904 38534 2916
rect 39025 2907 39083 2913
rect 39025 2904 39037 2907
rect 38528 2876 39037 2904
rect 38528 2864 38534 2876
rect 39025 2873 39037 2876
rect 39071 2873 39083 2907
rect 39132 2904 39160 3012
rect 39577 3009 39589 3043
rect 39623 3040 39635 3043
rect 40034 3040 40040 3052
rect 39623 3012 40040 3040
rect 39623 3009 39635 3012
rect 39577 3003 39635 3009
rect 40034 3000 40040 3012
rect 40092 3000 40098 3052
rect 40126 3000 40132 3052
rect 40184 3040 40190 3052
rect 40770 3040 40776 3052
rect 40184 3012 40776 3040
rect 40184 3000 40190 3012
rect 40770 3000 40776 3012
rect 40828 3000 40834 3052
rect 42705 3043 42763 3049
rect 42705 3040 42717 3043
rect 40880 3012 42717 3040
rect 39209 2975 39267 2981
rect 39209 2941 39221 2975
rect 39255 2972 39267 2975
rect 39298 2972 39304 2984
rect 39255 2944 39304 2972
rect 39255 2941 39267 2944
rect 39209 2935 39267 2941
rect 39298 2932 39304 2944
rect 39356 2972 39362 2984
rect 39942 2972 39948 2984
rect 39356 2944 39948 2972
rect 39356 2932 39362 2944
rect 39942 2932 39948 2944
rect 40000 2932 40006 2984
rect 40494 2972 40500 2984
rect 40455 2944 40500 2972
rect 40494 2932 40500 2944
rect 40552 2932 40558 2984
rect 40880 2972 40908 3012
rect 42705 3009 42717 3012
rect 42751 3009 42763 3043
rect 42812 3040 42840 3071
rect 42886 3068 42892 3120
rect 42944 3108 42950 3120
rect 42944 3080 44772 3108
rect 42944 3068 42950 3080
rect 44744 3040 44772 3080
rect 45002 3068 45008 3120
rect 45060 3108 45066 3120
rect 46290 3108 46296 3120
rect 45060 3080 46296 3108
rect 45060 3068 45066 3080
rect 46290 3068 46296 3080
rect 46348 3068 46354 3120
rect 47026 3068 47032 3120
rect 47084 3108 47090 3120
rect 47581 3111 47639 3117
rect 47581 3108 47593 3111
rect 47084 3080 47593 3108
rect 47084 3068 47090 3080
rect 47581 3077 47593 3080
rect 47627 3108 47639 3111
rect 49050 3108 49056 3120
rect 47627 3080 49056 3108
rect 47627 3077 47639 3080
rect 47581 3071 47639 3077
rect 49050 3068 49056 3080
rect 49108 3068 49114 3120
rect 52178 3068 52184 3120
rect 52236 3108 52242 3120
rect 52733 3111 52791 3117
rect 52733 3108 52745 3111
rect 52236 3080 52745 3108
rect 52236 3068 52242 3080
rect 52733 3077 52745 3080
rect 52779 3077 52791 3111
rect 52733 3071 52791 3077
rect 53466 3068 53472 3120
rect 53524 3108 53530 3120
rect 56134 3108 56140 3120
rect 53524 3080 56140 3108
rect 53524 3068 53530 3080
rect 56134 3068 56140 3080
rect 56192 3068 56198 3120
rect 50430 3040 50436 3052
rect 42812 3012 44680 3040
rect 44744 3012 50436 3040
rect 42705 3003 42763 3009
rect 42978 2972 42984 2984
rect 40604 2944 40908 2972
rect 41800 2944 42984 2972
rect 40604 2904 40632 2944
rect 39132 2876 40632 2904
rect 39025 2867 39083 2873
rect 37093 2839 37151 2845
rect 37093 2836 37105 2839
rect 36464 2808 37105 2836
rect 37093 2805 37105 2808
rect 37139 2836 37151 2839
rect 37274 2836 37280 2848
rect 37139 2808 37280 2836
rect 37139 2805 37151 2808
rect 37093 2799 37151 2805
rect 37274 2796 37280 2808
rect 37332 2796 37338 2848
rect 38746 2796 38752 2848
rect 38804 2836 38810 2848
rect 38841 2839 38899 2845
rect 38841 2836 38853 2839
rect 38804 2808 38853 2836
rect 38804 2796 38810 2808
rect 38841 2805 38853 2808
rect 38887 2805 38899 2839
rect 38841 2799 38899 2805
rect 40310 2796 40316 2848
rect 40368 2836 40374 2848
rect 41800 2836 41828 2944
rect 42978 2932 42984 2944
rect 43036 2932 43042 2984
rect 44652 2981 44680 3012
rect 50430 3000 50436 3012
rect 50488 3000 50494 3052
rect 50801 3043 50859 3049
rect 50801 3009 50813 3043
rect 50847 3040 50859 3043
rect 51166 3040 51172 3052
rect 50847 3012 51172 3040
rect 50847 3009 50859 3012
rect 50801 3003 50859 3009
rect 51166 3000 51172 3012
rect 51224 3000 51230 3052
rect 51718 3000 51724 3052
rect 51776 3040 51782 3052
rect 52641 3043 52699 3049
rect 52641 3040 52653 3043
rect 51776 3012 52653 3040
rect 51776 3000 51782 3012
rect 52641 3009 52653 3012
rect 52687 3040 52699 3043
rect 53285 3043 53343 3049
rect 53285 3040 53297 3043
rect 52687 3012 53297 3040
rect 52687 3009 52699 3012
rect 52641 3003 52699 3009
rect 53285 3009 53297 3012
rect 53331 3009 53343 3043
rect 54386 3040 54392 3052
rect 53285 3003 53343 3009
rect 53392 3012 54392 3040
rect 44637 2975 44695 2981
rect 44637 2941 44649 2975
rect 44683 2941 44695 2975
rect 44637 2935 44695 2941
rect 44726 2932 44732 2984
rect 44784 2972 44790 2984
rect 45002 2972 45008 2984
rect 44784 2944 44829 2972
rect 44963 2944 45008 2972
rect 44784 2932 44790 2944
rect 45002 2932 45008 2944
rect 45060 2932 45066 2984
rect 45186 2972 45192 2984
rect 45099 2944 45192 2972
rect 45186 2932 45192 2944
rect 45244 2972 45250 2984
rect 45244 2944 45968 2972
rect 45244 2932 45250 2944
rect 42521 2907 42579 2913
rect 42521 2873 42533 2907
rect 42567 2904 42579 2907
rect 42886 2904 42892 2916
rect 42567 2876 42892 2904
rect 42567 2873 42579 2876
rect 42521 2867 42579 2873
rect 42886 2864 42892 2876
rect 42944 2864 42950 2916
rect 43990 2904 43996 2916
rect 43951 2876 43996 2904
rect 43990 2864 43996 2876
rect 44048 2864 44054 2916
rect 45370 2864 45376 2916
rect 45428 2904 45434 2916
rect 45833 2907 45891 2913
rect 45833 2904 45845 2907
rect 45428 2876 45845 2904
rect 45428 2864 45434 2876
rect 45833 2873 45845 2876
rect 45879 2873 45891 2907
rect 45833 2867 45891 2873
rect 43070 2836 43076 2848
rect 40368 2808 41828 2836
rect 43031 2808 43076 2836
rect 40368 2796 40374 2808
rect 43070 2796 43076 2808
rect 43128 2796 43134 2848
rect 43714 2796 43720 2848
rect 43772 2836 43778 2848
rect 43809 2839 43867 2845
rect 43809 2836 43821 2839
rect 43772 2808 43821 2836
rect 43772 2796 43778 2808
rect 43809 2805 43821 2808
rect 43855 2836 43867 2839
rect 45554 2836 45560 2848
rect 43855 2808 45560 2836
rect 43855 2805 43867 2808
rect 43809 2799 43867 2805
rect 45554 2796 45560 2808
rect 45612 2796 45618 2848
rect 45940 2836 45968 2944
rect 46106 2932 46112 2984
rect 46164 2972 46170 2984
rect 46201 2975 46259 2981
rect 46201 2972 46213 2975
rect 46164 2944 46213 2972
rect 46164 2932 46170 2944
rect 46201 2941 46213 2944
rect 46247 2941 46259 2975
rect 46201 2935 46259 2941
rect 46290 2932 46296 2984
rect 46348 2972 46354 2984
rect 47026 2972 47032 2984
rect 46348 2944 46393 2972
rect 46987 2944 47032 2972
rect 46348 2932 46354 2944
rect 47026 2932 47032 2944
rect 47084 2932 47090 2984
rect 47121 2975 47179 2981
rect 47121 2941 47133 2975
rect 47167 2972 47179 2975
rect 47949 2975 48007 2981
rect 47949 2972 47961 2975
rect 47167 2944 47961 2972
rect 47167 2941 47179 2944
rect 47121 2935 47179 2941
rect 47949 2941 47961 2944
rect 47995 2972 48007 2975
rect 48222 2972 48228 2984
rect 47995 2944 48228 2972
rect 47995 2941 48007 2944
rect 47949 2935 48007 2941
rect 46014 2864 46020 2916
rect 46072 2904 46078 2916
rect 47136 2904 47164 2935
rect 48222 2932 48228 2944
rect 48280 2932 48286 2984
rect 49326 2972 49332 2984
rect 49287 2944 49332 2972
rect 49326 2932 49332 2944
rect 49384 2932 49390 2984
rect 49878 2972 49884 2984
rect 49839 2944 49884 2972
rect 49878 2932 49884 2944
rect 49936 2932 49942 2984
rect 50341 2975 50399 2981
rect 50341 2941 50353 2975
rect 50387 2941 50399 2975
rect 50341 2935 50399 2941
rect 46072 2876 47164 2904
rect 46072 2864 46078 2876
rect 48130 2864 48136 2916
rect 48188 2904 48194 2916
rect 50356 2904 50384 2935
rect 50522 2932 50528 2984
rect 50580 2972 50586 2984
rect 50709 2975 50767 2981
rect 50709 2972 50721 2975
rect 50580 2944 50721 2972
rect 50580 2932 50586 2944
rect 50709 2941 50721 2944
rect 50755 2972 50767 2975
rect 51534 2972 51540 2984
rect 50755 2944 51540 2972
rect 50755 2941 50767 2944
rect 50709 2935 50767 2941
rect 51534 2932 51540 2944
rect 51592 2932 51598 2984
rect 52181 2975 52239 2981
rect 52181 2941 52193 2975
rect 52227 2972 52239 2975
rect 52420 2975 52478 2981
rect 52420 2972 52432 2975
rect 52227 2944 52432 2972
rect 52227 2941 52239 2944
rect 52181 2935 52239 2941
rect 52420 2941 52432 2944
rect 52466 2972 52478 2975
rect 53392 2972 53420 3012
rect 54386 3000 54392 3012
rect 54444 3000 54450 3052
rect 54573 3043 54631 3049
rect 54573 3009 54585 3043
rect 54619 3040 54631 3043
rect 55030 3040 55036 3052
rect 54619 3012 55036 3040
rect 54619 3009 54631 3012
rect 54573 3003 54631 3009
rect 55030 3000 55036 3012
rect 55088 3040 55094 3052
rect 55585 3043 55643 3049
rect 55585 3040 55597 3043
rect 55088 3012 55597 3040
rect 55088 3000 55094 3012
rect 55585 3009 55597 3012
rect 55631 3009 55643 3043
rect 57624 3040 57652 3136
rect 57882 3068 57888 3120
rect 57940 3108 57946 3120
rect 60826 3108 60832 3120
rect 57940 3080 60832 3108
rect 57940 3068 57946 3080
rect 60826 3068 60832 3080
rect 60884 3068 60890 3120
rect 60994 3111 61052 3117
rect 60994 3077 61006 3111
rect 61040 3108 61052 3111
rect 62206 3108 62212 3120
rect 61040 3080 62212 3108
rect 61040 3077 61052 3080
rect 60994 3071 61052 3077
rect 62206 3068 62212 3080
rect 62264 3068 62270 3120
rect 59357 3043 59415 3049
rect 59357 3040 59369 3043
rect 57624 3012 59369 3040
rect 55585 3003 55643 3009
rect 59357 3009 59369 3012
rect 59403 3009 59415 3043
rect 59357 3003 59415 3009
rect 61194 3000 61200 3052
rect 61252 3040 61258 3052
rect 61252 3012 61294 3040
rect 61252 3000 61258 3012
rect 54110 2972 54116 2984
rect 52466 2944 53420 2972
rect 54071 2944 54116 2972
rect 52466 2941 52478 2944
rect 52420 2935 52478 2941
rect 54110 2932 54116 2944
rect 54168 2932 54174 2984
rect 54849 2975 54907 2981
rect 54849 2972 54861 2975
rect 54220 2944 54861 2972
rect 51074 2904 51080 2916
rect 48188 2876 48544 2904
rect 50356 2876 51080 2904
rect 48188 2864 48194 2876
rect 46934 2836 46940 2848
rect 45940 2808 46940 2836
rect 46934 2796 46940 2808
rect 46992 2796 46998 2848
rect 48314 2796 48320 2848
rect 48372 2836 48378 2848
rect 48409 2839 48467 2845
rect 48409 2836 48421 2839
rect 48372 2808 48421 2836
rect 48372 2796 48378 2808
rect 48409 2805 48421 2808
rect 48455 2805 48467 2839
rect 48516 2836 48544 2876
rect 51074 2864 51080 2876
rect 51132 2904 51138 2916
rect 51169 2907 51227 2913
rect 51169 2904 51181 2907
rect 51132 2876 51181 2904
rect 51132 2864 51138 2876
rect 51169 2873 51181 2876
rect 51215 2904 51227 2907
rect 51994 2904 52000 2916
rect 51215 2876 52000 2904
rect 51215 2873 51227 2876
rect 51169 2867 51227 2873
rect 51994 2864 52000 2876
rect 52052 2864 52058 2916
rect 52270 2904 52276 2916
rect 52231 2876 52276 2904
rect 52270 2864 52276 2876
rect 52328 2864 52334 2916
rect 53558 2864 53564 2916
rect 53616 2904 53622 2916
rect 54021 2907 54079 2913
rect 54021 2904 54033 2907
rect 53616 2876 54033 2904
rect 53616 2864 53622 2876
rect 54021 2873 54033 2876
rect 54067 2904 54079 2907
rect 54220 2904 54248 2944
rect 54849 2941 54861 2944
rect 54895 2941 54907 2975
rect 55306 2972 55312 2984
rect 55267 2944 55312 2972
rect 54849 2935 54907 2941
rect 55306 2932 55312 2944
rect 55364 2932 55370 2984
rect 56137 2975 56195 2981
rect 56137 2941 56149 2975
rect 56183 2972 56195 2975
rect 56226 2972 56232 2984
rect 56183 2944 56232 2972
rect 56183 2941 56195 2944
rect 56137 2935 56195 2941
rect 56226 2932 56232 2944
rect 56284 2932 56290 2984
rect 59449 2975 59507 2981
rect 59449 2941 59461 2975
rect 59495 2941 59507 2975
rect 59814 2972 59820 2984
rect 59775 2944 59820 2972
rect 59449 2935 59507 2941
rect 55122 2904 55128 2916
rect 54067 2876 54248 2904
rect 54772 2876 55128 2904
rect 54067 2873 54079 2876
rect 54021 2867 54079 2873
rect 51810 2836 51816 2848
rect 48516 2808 51816 2836
rect 48409 2799 48467 2805
rect 51810 2796 51816 2808
rect 51868 2796 51874 2848
rect 53742 2836 53748 2848
rect 53703 2808 53748 2836
rect 53742 2796 53748 2808
rect 53800 2836 53806 2848
rect 54772 2836 54800 2876
rect 55122 2864 55128 2876
rect 55180 2864 55186 2916
rect 55582 2864 55588 2916
rect 55640 2904 55646 2916
rect 58253 2907 58311 2913
rect 58253 2904 58265 2907
rect 55640 2876 58265 2904
rect 55640 2864 55646 2876
rect 58253 2873 58265 2876
rect 58299 2904 58311 2907
rect 59464 2904 59492 2935
rect 59814 2932 59820 2944
rect 59872 2932 59878 2984
rect 59998 2972 60004 2984
rect 59959 2944 60004 2972
rect 59998 2932 60004 2944
rect 60056 2932 60062 2984
rect 64138 2972 64144 2984
rect 60108 2944 64144 2972
rect 58299 2876 59492 2904
rect 58299 2873 58311 2876
rect 58253 2867 58311 2873
rect 53800 2808 54800 2836
rect 53800 2796 53806 2808
rect 59446 2796 59452 2848
rect 59504 2836 59510 2848
rect 60108 2836 60136 2944
rect 64138 2932 64144 2944
rect 64196 2932 64202 2984
rect 60274 2904 60280 2916
rect 60235 2876 60280 2904
rect 60274 2864 60280 2876
rect 60332 2864 60338 2916
rect 60737 2907 60795 2913
rect 60737 2873 60749 2907
rect 60783 2904 60795 2907
rect 60829 2907 60887 2913
rect 60829 2904 60841 2907
rect 60783 2876 60841 2904
rect 60783 2873 60795 2876
rect 60737 2867 60795 2873
rect 60829 2873 60841 2876
rect 60875 2904 60887 2907
rect 63218 2904 63224 2916
rect 60875 2876 63224 2904
rect 60875 2873 60887 2876
rect 60829 2867 60887 2873
rect 63218 2864 63224 2876
rect 63276 2864 63282 2916
rect 59504 2808 60136 2836
rect 59504 2796 59510 2808
rect 61194 2796 61200 2848
rect 61252 2836 61258 2848
rect 61841 2839 61899 2845
rect 61841 2836 61853 2839
rect 61252 2808 61853 2836
rect 61252 2796 61258 2808
rect 61841 2805 61853 2808
rect 61887 2805 61899 2839
rect 61841 2799 61899 2805
rect 1104 2746 63480 2768
rect 1104 2694 21774 2746
rect 21826 2694 21838 2746
rect 21890 2694 21902 2746
rect 21954 2694 21966 2746
rect 22018 2694 42566 2746
rect 42618 2694 42630 2746
rect 42682 2694 42694 2746
rect 42746 2694 42758 2746
rect 42810 2694 63480 2746
rect 1104 2672 63480 2694
rect 3050 2632 3056 2644
rect 3011 2604 3056 2632
rect 3050 2592 3056 2604
rect 3108 2592 3114 2644
rect 5718 2632 5724 2644
rect 5679 2604 5724 2632
rect 5718 2592 5724 2604
rect 5776 2592 5782 2644
rect 6178 2592 6184 2644
rect 6236 2632 6242 2644
rect 6273 2635 6331 2641
rect 6273 2632 6285 2635
rect 6236 2604 6285 2632
rect 6236 2592 6242 2604
rect 6273 2601 6285 2604
rect 6319 2601 6331 2635
rect 6273 2595 6331 2601
rect 9030 2592 9036 2644
rect 9088 2632 9094 2644
rect 9493 2635 9551 2641
rect 9493 2632 9505 2635
rect 9088 2604 9505 2632
rect 9088 2592 9094 2604
rect 9493 2601 9505 2604
rect 9539 2632 9551 2635
rect 9582 2632 9588 2644
rect 9539 2604 9588 2632
rect 9539 2601 9551 2604
rect 9493 2595 9551 2601
rect 9582 2592 9588 2604
rect 9640 2592 9646 2644
rect 10410 2592 10416 2644
rect 10468 2632 10474 2644
rect 10689 2635 10747 2641
rect 10689 2632 10701 2635
rect 10468 2604 10701 2632
rect 10468 2592 10474 2604
rect 10689 2601 10701 2604
rect 10735 2632 10747 2635
rect 10781 2635 10839 2641
rect 10781 2632 10793 2635
rect 10735 2604 10793 2632
rect 10735 2601 10747 2604
rect 10689 2595 10747 2601
rect 10781 2601 10793 2604
rect 10827 2632 10839 2635
rect 12161 2635 12219 2641
rect 12161 2632 12173 2635
rect 10827 2604 12173 2632
rect 10827 2601 10839 2604
rect 10781 2595 10839 2601
rect 12161 2601 12173 2604
rect 12207 2601 12219 2635
rect 12342 2632 12348 2644
rect 12303 2604 12348 2632
rect 12161 2595 12219 2601
rect 12342 2592 12348 2604
rect 12400 2592 12406 2644
rect 12894 2632 12900 2644
rect 12855 2604 12900 2632
rect 12894 2592 12900 2604
rect 12952 2592 12958 2644
rect 13354 2592 13360 2644
rect 13412 2632 13418 2644
rect 13449 2635 13507 2641
rect 13449 2632 13461 2635
rect 13412 2604 13461 2632
rect 13412 2592 13418 2604
rect 13449 2601 13461 2604
rect 13495 2632 13507 2635
rect 14737 2635 14795 2641
rect 14737 2632 14749 2635
rect 13495 2604 14749 2632
rect 13495 2601 13507 2604
rect 13449 2595 13507 2601
rect 8849 2567 8907 2573
rect 8849 2533 8861 2567
rect 8895 2564 8907 2567
rect 9217 2567 9275 2573
rect 9217 2564 9229 2567
rect 8895 2536 9229 2564
rect 8895 2533 8907 2536
rect 8849 2527 8907 2533
rect 9217 2533 9229 2536
rect 9263 2564 9275 2567
rect 9398 2564 9404 2576
rect 9263 2536 9404 2564
rect 9263 2533 9275 2536
rect 9217 2527 9275 2533
rect 9398 2524 9404 2536
rect 9456 2524 9462 2576
rect 10137 2567 10195 2573
rect 10137 2533 10149 2567
rect 10183 2564 10195 2567
rect 10183 2536 11284 2564
rect 10183 2533 10195 2536
rect 10137 2527 10195 2533
rect 2958 2496 2964 2508
rect 2919 2468 2964 2496
rect 2958 2456 2964 2468
rect 3016 2496 3022 2508
rect 3421 2499 3479 2505
rect 3421 2496 3433 2499
rect 3016 2468 3433 2496
rect 3016 2456 3022 2468
rect 3421 2465 3433 2468
rect 3467 2465 3479 2499
rect 3421 2459 3479 2465
rect 3881 2499 3939 2505
rect 3881 2465 3893 2499
rect 3927 2496 3939 2499
rect 4617 2499 4675 2505
rect 4617 2496 4629 2499
rect 3927 2468 4629 2496
rect 3927 2465 3939 2468
rect 3881 2459 3939 2465
rect 4617 2465 4629 2468
rect 4663 2496 4675 2499
rect 4706 2496 4712 2508
rect 4663 2468 4712 2496
rect 4663 2465 4675 2468
rect 4617 2459 4675 2465
rect 4706 2456 4712 2468
rect 4764 2456 4770 2508
rect 6733 2499 6791 2505
rect 6733 2465 6745 2499
rect 6779 2496 6791 2499
rect 7469 2499 7527 2505
rect 7469 2496 7481 2499
rect 6779 2468 7481 2496
rect 6779 2465 6791 2468
rect 6733 2459 6791 2465
rect 7469 2465 7481 2468
rect 7515 2496 7527 2499
rect 8110 2496 8116 2508
rect 7515 2468 8116 2496
rect 7515 2465 7527 2468
rect 7469 2459 7527 2465
rect 8110 2456 8116 2468
rect 8168 2456 8174 2508
rect 11256 2505 11284 2536
rect 10689 2499 10747 2505
rect 10689 2465 10701 2499
rect 10735 2496 10747 2499
rect 10965 2499 11023 2505
rect 10965 2496 10977 2499
rect 10735 2468 10977 2496
rect 10735 2465 10747 2468
rect 10689 2459 10747 2465
rect 10965 2465 10977 2468
rect 11011 2465 11023 2499
rect 10965 2459 11023 2465
rect 11149 2499 11207 2505
rect 11149 2465 11161 2499
rect 11195 2465 11207 2499
rect 11149 2459 11207 2465
rect 11241 2499 11299 2505
rect 11241 2465 11253 2499
rect 11287 2496 11299 2499
rect 11974 2496 11980 2508
rect 11287 2468 11980 2496
rect 11287 2465 11299 2468
rect 11241 2459 11299 2465
rect 2314 2388 2320 2440
rect 2372 2428 2378 2440
rect 2501 2431 2559 2437
rect 2501 2428 2513 2431
rect 2372 2400 2513 2428
rect 2372 2388 2378 2400
rect 2501 2397 2513 2400
rect 2547 2428 2559 2431
rect 2869 2431 2927 2437
rect 2869 2428 2881 2431
rect 2547 2400 2881 2428
rect 2547 2397 2559 2400
rect 2501 2391 2559 2397
rect 2869 2397 2881 2400
rect 2915 2428 2927 2431
rect 3602 2428 3608 2440
rect 2915 2400 3608 2428
rect 2915 2397 2927 2400
rect 2869 2391 2927 2397
rect 3602 2388 3608 2400
rect 3660 2428 3666 2440
rect 4341 2431 4399 2437
rect 4341 2428 4353 2431
rect 3660 2400 4353 2428
rect 3660 2388 3666 2400
rect 4341 2397 4353 2400
rect 4387 2428 4399 2431
rect 7193 2431 7251 2437
rect 7193 2428 7205 2431
rect 4387 2400 7205 2428
rect 4387 2397 4399 2400
rect 4341 2391 4399 2397
rect 7193 2397 7205 2400
rect 7239 2397 7251 2431
rect 7193 2391 7251 2397
rect 10505 2431 10563 2437
rect 10505 2397 10517 2431
rect 10551 2428 10563 2431
rect 11164 2428 11192 2459
rect 11974 2456 11980 2468
rect 12032 2456 12038 2508
rect 14016 2505 14044 2604
rect 14737 2601 14749 2604
rect 14783 2601 14795 2635
rect 15194 2632 15200 2644
rect 15155 2604 15200 2632
rect 14737 2595 14795 2601
rect 15194 2592 15200 2604
rect 15252 2592 15258 2644
rect 16390 2632 16396 2644
rect 15396 2604 16396 2632
rect 15396 2564 15424 2604
rect 16390 2592 16396 2604
rect 16448 2592 16454 2644
rect 17773 2635 17831 2641
rect 17773 2601 17785 2635
rect 17819 2632 17831 2635
rect 19334 2632 19340 2644
rect 17819 2604 19340 2632
rect 17819 2601 17831 2604
rect 17773 2595 17831 2601
rect 19334 2592 19340 2604
rect 19392 2592 19398 2644
rect 19610 2632 19616 2644
rect 19571 2604 19616 2632
rect 19610 2592 19616 2604
rect 19668 2592 19674 2644
rect 20272 2604 24256 2632
rect 14292 2536 15424 2564
rect 17129 2567 17187 2573
rect 14001 2499 14059 2505
rect 14001 2465 14013 2499
rect 14047 2465 14059 2499
rect 14001 2459 14059 2465
rect 13078 2428 13084 2440
rect 10551 2400 13084 2428
rect 10551 2397 10563 2400
rect 10505 2391 10563 2397
rect 13078 2388 13084 2400
rect 13136 2388 13142 2440
rect 14292 2428 14320 2536
rect 17129 2533 17141 2567
rect 17175 2564 17187 2567
rect 17862 2564 17868 2576
rect 17175 2536 17868 2564
rect 17175 2533 17187 2536
rect 17129 2527 17187 2533
rect 17862 2524 17868 2536
rect 17920 2524 17926 2576
rect 18877 2567 18935 2573
rect 18064 2536 18552 2564
rect 14369 2499 14427 2505
rect 14369 2465 14381 2499
rect 14415 2465 14427 2499
rect 14369 2459 14427 2465
rect 13740 2400 14320 2428
rect 14384 2428 14412 2459
rect 14458 2456 14464 2508
rect 14516 2496 14522 2508
rect 14516 2468 14561 2496
rect 14516 2456 14522 2468
rect 15286 2456 15292 2508
rect 15344 2496 15350 2508
rect 15473 2499 15531 2505
rect 15473 2496 15485 2499
rect 15344 2468 15485 2496
rect 15344 2456 15350 2468
rect 15473 2465 15485 2468
rect 15519 2465 15531 2499
rect 15746 2496 15752 2508
rect 15707 2468 15752 2496
rect 15473 2459 15531 2465
rect 15746 2456 15752 2468
rect 15804 2456 15810 2508
rect 17586 2456 17592 2508
rect 17644 2496 17650 2508
rect 18064 2496 18092 2536
rect 18524 2505 18552 2536
rect 18877 2533 18889 2567
rect 18923 2564 18935 2567
rect 19794 2564 19800 2576
rect 18923 2536 19800 2564
rect 18923 2533 18935 2536
rect 18877 2527 18935 2533
rect 19794 2524 19800 2536
rect 19852 2524 19858 2576
rect 20272 2573 20300 2604
rect 20257 2567 20315 2573
rect 20257 2533 20269 2567
rect 20303 2533 20315 2567
rect 20257 2527 20315 2533
rect 23014 2524 23020 2576
rect 23072 2564 23078 2576
rect 23109 2567 23167 2573
rect 23109 2564 23121 2567
rect 23072 2536 23121 2564
rect 23072 2524 23078 2536
rect 23109 2533 23121 2536
rect 23155 2533 23167 2567
rect 23474 2564 23480 2576
rect 23435 2536 23480 2564
rect 23109 2527 23167 2533
rect 23474 2524 23480 2536
rect 23532 2524 23538 2576
rect 24228 2573 24256 2604
rect 24854 2592 24860 2644
rect 24912 2632 24918 2644
rect 25133 2635 25191 2641
rect 25133 2632 25145 2635
rect 24912 2604 25145 2632
rect 24912 2592 24918 2604
rect 25133 2601 25145 2604
rect 25179 2632 25191 2635
rect 26418 2632 26424 2644
rect 25179 2604 26424 2632
rect 25179 2601 25191 2604
rect 25133 2595 25191 2601
rect 26418 2592 26424 2604
rect 26476 2592 26482 2644
rect 26602 2632 26608 2644
rect 26563 2604 26608 2632
rect 26602 2592 26608 2604
rect 26660 2592 26666 2644
rect 26694 2592 26700 2644
rect 26752 2632 26758 2644
rect 28261 2635 28319 2641
rect 28261 2632 28273 2635
rect 26752 2604 28273 2632
rect 26752 2592 26758 2604
rect 28261 2601 28273 2604
rect 28307 2601 28319 2635
rect 28261 2595 28319 2601
rect 28994 2592 29000 2644
rect 29052 2632 29058 2644
rect 29181 2635 29239 2641
rect 29181 2632 29193 2635
rect 29052 2604 29193 2632
rect 29052 2592 29058 2604
rect 29181 2601 29193 2604
rect 29227 2601 29239 2635
rect 29181 2595 29239 2601
rect 31938 2592 31944 2644
rect 31996 2632 32002 2644
rect 32309 2635 32367 2641
rect 32309 2632 32321 2635
rect 31996 2604 32321 2632
rect 31996 2592 32002 2604
rect 32309 2601 32321 2604
rect 32355 2601 32367 2635
rect 32309 2595 32367 2601
rect 32674 2592 32680 2644
rect 32732 2632 32738 2644
rect 34790 2632 34796 2644
rect 32732 2604 34796 2632
rect 32732 2592 32738 2604
rect 34790 2592 34796 2604
rect 34848 2632 34854 2644
rect 34885 2635 34943 2641
rect 34885 2632 34897 2635
rect 34848 2604 34897 2632
rect 34848 2592 34854 2604
rect 34885 2601 34897 2604
rect 34931 2601 34943 2635
rect 34885 2595 34943 2601
rect 35894 2592 35900 2644
rect 35952 2632 35958 2644
rect 36081 2635 36139 2641
rect 36081 2632 36093 2635
rect 35952 2604 36093 2632
rect 35952 2592 35958 2604
rect 36081 2601 36093 2604
rect 36127 2601 36139 2635
rect 36081 2595 36139 2601
rect 38565 2635 38623 2641
rect 38565 2601 38577 2635
rect 38611 2632 38623 2635
rect 39022 2632 39028 2644
rect 38611 2604 39028 2632
rect 38611 2601 38623 2604
rect 38565 2595 38623 2601
rect 39022 2592 39028 2604
rect 39080 2632 39086 2644
rect 39301 2635 39359 2641
rect 39301 2632 39313 2635
rect 39080 2604 39313 2632
rect 39080 2592 39086 2604
rect 24213 2567 24271 2573
rect 24213 2533 24225 2567
rect 24259 2564 24271 2567
rect 25409 2567 25467 2573
rect 25409 2564 25421 2567
rect 24259 2536 25421 2564
rect 24259 2533 24271 2536
rect 24213 2527 24271 2533
rect 25409 2533 25421 2536
rect 25455 2533 25467 2567
rect 25409 2527 25467 2533
rect 17644 2468 18092 2496
rect 18141 2499 18199 2505
rect 17644 2456 17650 2468
rect 18141 2465 18153 2499
rect 18187 2496 18199 2499
rect 18325 2499 18383 2505
rect 18325 2496 18337 2499
rect 18187 2468 18337 2496
rect 18187 2465 18199 2468
rect 18141 2459 18199 2465
rect 18325 2465 18337 2468
rect 18371 2465 18383 2499
rect 18325 2459 18383 2465
rect 18509 2499 18567 2505
rect 18509 2465 18521 2499
rect 18555 2496 18567 2499
rect 19153 2499 19211 2505
rect 19153 2496 19165 2499
rect 18555 2468 19165 2496
rect 18555 2465 18567 2468
rect 18509 2459 18567 2465
rect 19153 2465 19165 2468
rect 19199 2465 19211 2499
rect 19153 2459 19211 2465
rect 19705 2499 19763 2505
rect 19705 2465 19717 2499
rect 19751 2465 19763 2499
rect 19705 2459 19763 2465
rect 19889 2499 19947 2505
rect 19889 2465 19901 2499
rect 19935 2496 19947 2499
rect 19978 2496 19984 2508
rect 19935 2468 19984 2496
rect 19935 2465 19947 2468
rect 19889 2459 19947 2465
rect 14645 2431 14703 2437
rect 14645 2428 14657 2431
rect 14384 2400 14657 2428
rect 2130 2292 2136 2304
rect 2091 2264 2136 2292
rect 2130 2252 2136 2264
rect 2188 2252 2194 2304
rect 7834 2252 7840 2304
rect 7892 2292 7898 2304
rect 11425 2295 11483 2301
rect 11425 2292 11437 2295
rect 7892 2264 11437 2292
rect 7892 2252 7898 2264
rect 11425 2261 11437 2264
rect 11471 2261 11483 2295
rect 11425 2255 11483 2261
rect 12161 2295 12219 2301
rect 12161 2261 12173 2295
rect 12207 2292 12219 2295
rect 13740 2292 13768 2400
rect 14645 2397 14657 2400
rect 14691 2397 14703 2431
rect 14645 2391 14703 2397
rect 14737 2431 14795 2437
rect 14737 2397 14749 2431
rect 14783 2428 14795 2431
rect 18340 2428 18368 2459
rect 19242 2428 19248 2440
rect 14783 2400 17816 2428
rect 18340 2400 19248 2428
rect 14783 2397 14795 2400
rect 14737 2391 14795 2397
rect 13817 2363 13875 2369
rect 13817 2329 13829 2363
rect 13863 2360 13875 2363
rect 15378 2360 15384 2372
rect 13863 2332 15384 2360
rect 13863 2329 13875 2332
rect 13817 2323 13875 2329
rect 15378 2320 15384 2332
rect 15436 2320 15442 2372
rect 12207 2264 13768 2292
rect 14645 2295 14703 2301
rect 12207 2261 12219 2264
rect 12161 2255 12219 2261
rect 14645 2261 14657 2295
rect 14691 2292 14703 2295
rect 14921 2295 14979 2301
rect 14921 2292 14933 2295
rect 14691 2264 14933 2292
rect 14691 2261 14703 2264
rect 14645 2255 14703 2261
rect 14921 2261 14933 2264
rect 14967 2292 14979 2295
rect 17678 2292 17684 2304
rect 14967 2264 17684 2292
rect 14967 2261 14979 2264
rect 14921 2255 14979 2261
rect 17678 2252 17684 2264
rect 17736 2252 17742 2304
rect 17788 2292 17816 2400
rect 19242 2388 19248 2400
rect 19300 2428 19306 2440
rect 19720 2428 19748 2459
rect 19978 2456 19984 2468
rect 20036 2496 20042 2508
rect 20533 2499 20591 2505
rect 20533 2496 20545 2499
rect 20036 2468 20545 2496
rect 20036 2456 20042 2468
rect 20533 2465 20545 2468
rect 20579 2465 20591 2499
rect 20533 2459 20591 2465
rect 20993 2499 21051 2505
rect 20993 2465 21005 2499
rect 21039 2496 21051 2499
rect 21542 2496 21548 2508
rect 21039 2468 21548 2496
rect 21039 2465 21051 2468
rect 20993 2459 21051 2465
rect 21542 2456 21548 2468
rect 21600 2496 21606 2508
rect 21729 2499 21787 2505
rect 21729 2496 21741 2499
rect 21600 2468 21741 2496
rect 21600 2456 21606 2468
rect 21729 2465 21741 2468
rect 21775 2465 21787 2499
rect 21729 2459 21787 2465
rect 24302 2456 24308 2508
rect 24360 2496 24366 2508
rect 24360 2468 24405 2496
rect 24360 2456 24366 2468
rect 25038 2456 25044 2508
rect 25096 2496 25102 2508
rect 25593 2499 25651 2505
rect 25593 2496 25605 2499
rect 25096 2468 25605 2496
rect 25096 2456 25102 2468
rect 25593 2465 25605 2468
rect 25639 2496 25651 2499
rect 26145 2499 26203 2505
rect 26145 2496 26157 2499
rect 25639 2468 26157 2496
rect 25639 2465 25651 2468
rect 25593 2459 25651 2465
rect 26145 2465 26157 2468
rect 26191 2465 26203 2499
rect 26620 2496 26648 2592
rect 28074 2524 28080 2576
rect 28132 2564 28138 2576
rect 28813 2567 28871 2573
rect 28813 2564 28825 2567
rect 28132 2536 28825 2564
rect 28132 2524 28138 2536
rect 28813 2533 28825 2536
rect 28859 2533 28871 2567
rect 36998 2564 37004 2576
rect 28813 2527 28871 2533
rect 36004 2536 37004 2564
rect 27157 2499 27215 2505
rect 27157 2496 27169 2499
rect 26620 2468 27169 2496
rect 26145 2459 26203 2465
rect 27157 2465 27169 2468
rect 27203 2465 27215 2499
rect 27157 2459 27215 2465
rect 30101 2499 30159 2505
rect 30101 2465 30113 2499
rect 30147 2496 30159 2499
rect 30742 2496 30748 2508
rect 30147 2468 30748 2496
rect 30147 2465 30159 2468
rect 30101 2459 30159 2465
rect 30742 2456 30748 2468
rect 30800 2456 30806 2508
rect 31110 2496 31116 2508
rect 31071 2468 31116 2496
rect 31110 2456 31116 2468
rect 31168 2496 31174 2508
rect 31941 2499 31999 2505
rect 31941 2496 31953 2499
rect 31168 2468 31953 2496
rect 31168 2456 31174 2468
rect 31941 2465 31953 2468
rect 31987 2465 31999 2499
rect 31941 2459 31999 2465
rect 32585 2499 32643 2505
rect 32585 2465 32597 2499
rect 32631 2496 32643 2499
rect 33686 2496 33692 2508
rect 32631 2468 33692 2496
rect 32631 2465 32643 2468
rect 32585 2459 32643 2465
rect 33686 2456 33692 2468
rect 33744 2456 33750 2508
rect 36004 2505 36032 2536
rect 36998 2524 37004 2536
rect 37056 2524 37062 2576
rect 35897 2499 35955 2505
rect 35897 2465 35909 2499
rect 35943 2496 35955 2499
rect 35989 2499 36047 2505
rect 35989 2496 36001 2499
rect 35943 2468 36001 2496
rect 35943 2465 35955 2468
rect 35897 2459 35955 2465
rect 35989 2465 36001 2468
rect 36035 2465 36047 2499
rect 35989 2459 36047 2465
rect 36078 2456 36084 2508
rect 36136 2496 36142 2508
rect 36630 2496 36636 2508
rect 36136 2468 36636 2496
rect 36136 2456 36142 2468
rect 36630 2456 36636 2468
rect 36688 2456 36694 2508
rect 36817 2499 36875 2505
rect 36817 2465 36829 2499
rect 36863 2496 36875 2499
rect 37274 2496 37280 2508
rect 36863 2468 37280 2496
rect 36863 2465 36875 2468
rect 36817 2459 36875 2465
rect 37274 2456 37280 2468
rect 37332 2456 37338 2508
rect 38381 2499 38439 2505
rect 38381 2465 38393 2499
rect 38427 2465 38439 2499
rect 39132 2496 39160 2604
rect 39301 2601 39313 2604
rect 39347 2601 39359 2635
rect 40770 2632 40776 2644
rect 40731 2604 40776 2632
rect 39301 2595 39359 2601
rect 40770 2592 40776 2604
rect 40828 2592 40834 2644
rect 41414 2592 41420 2644
rect 41472 2632 41478 2644
rect 43809 2635 43867 2641
rect 41472 2604 43760 2632
rect 41472 2592 41478 2604
rect 39206 2524 39212 2576
rect 39264 2564 39270 2576
rect 39669 2567 39727 2573
rect 39669 2564 39681 2567
rect 39264 2536 39681 2564
rect 39264 2524 39270 2536
rect 39669 2533 39681 2536
rect 39715 2533 39727 2567
rect 39669 2527 39727 2533
rect 40221 2567 40279 2573
rect 40221 2533 40233 2567
rect 40267 2564 40279 2567
rect 40586 2564 40592 2576
rect 40267 2536 40592 2564
rect 40267 2533 40279 2536
rect 40221 2527 40279 2533
rect 40586 2524 40592 2536
rect 40644 2524 40650 2576
rect 41046 2524 41052 2576
rect 41104 2564 41110 2576
rect 41104 2536 42196 2564
rect 41104 2524 41110 2536
rect 39485 2499 39543 2505
rect 39485 2496 39497 2499
rect 39132 2468 39497 2496
rect 38381 2459 38439 2465
rect 39485 2465 39497 2468
rect 39531 2465 39543 2499
rect 39758 2496 39764 2508
rect 39671 2468 39764 2496
rect 39485 2459 39543 2465
rect 21450 2428 21456 2440
rect 19300 2400 19748 2428
rect 21411 2400 21456 2428
rect 19300 2388 19306 2400
rect 21450 2388 21456 2400
rect 21508 2388 21514 2440
rect 22370 2388 22376 2440
rect 22428 2428 22434 2440
rect 24765 2431 24823 2437
rect 24765 2428 24777 2431
rect 22428 2400 24777 2428
rect 22428 2388 22434 2400
rect 24765 2397 24777 2400
rect 24811 2397 24823 2431
rect 26881 2431 26939 2437
rect 26881 2428 26893 2431
rect 24765 2391 24823 2397
rect 24872 2400 26893 2428
rect 18046 2320 18052 2372
rect 18104 2360 18110 2372
rect 18874 2360 18880 2372
rect 18104 2332 18880 2360
rect 18104 2320 18110 2332
rect 18874 2320 18880 2332
rect 18932 2320 18938 2372
rect 24118 2320 24124 2372
rect 24176 2360 24182 2372
rect 24872 2360 24900 2400
rect 26881 2397 26893 2400
rect 26927 2397 26939 2431
rect 26881 2391 26939 2397
rect 30469 2431 30527 2437
rect 30469 2397 30481 2431
rect 30515 2428 30527 2431
rect 31202 2428 31208 2440
rect 30515 2400 31208 2428
rect 30515 2397 30527 2400
rect 30469 2391 30527 2397
rect 31202 2388 31208 2400
rect 31260 2428 31266 2440
rect 31389 2431 31447 2437
rect 31389 2428 31401 2431
rect 31260 2400 31401 2428
rect 31260 2388 31266 2400
rect 31389 2397 31401 2400
rect 31435 2397 31447 2431
rect 32861 2431 32919 2437
rect 32861 2428 32873 2431
rect 31389 2391 31447 2397
rect 32508 2400 32873 2428
rect 24176 2332 24900 2360
rect 25777 2363 25835 2369
rect 24176 2320 24182 2332
rect 25777 2329 25789 2363
rect 25823 2360 25835 2363
rect 25866 2360 25872 2372
rect 25823 2332 25872 2360
rect 25823 2329 25835 2332
rect 25777 2323 25835 2329
rect 25866 2320 25872 2332
rect 25924 2320 25930 2372
rect 30837 2363 30895 2369
rect 30837 2329 30849 2363
rect 30883 2360 30895 2363
rect 32508 2360 32536 2400
rect 32861 2397 32873 2400
rect 32907 2428 32919 2431
rect 32950 2428 32956 2440
rect 32907 2400 32956 2428
rect 32907 2397 32919 2400
rect 32861 2391 32919 2397
rect 32950 2388 32956 2400
rect 33008 2388 33014 2440
rect 36648 2428 36676 2456
rect 37369 2431 37427 2437
rect 37369 2428 37381 2431
rect 36648 2400 37381 2428
rect 37369 2397 37381 2400
rect 37415 2397 37427 2431
rect 38396 2428 38424 2459
rect 39758 2456 39764 2468
rect 39816 2496 39822 2508
rect 40402 2496 40408 2508
rect 39816 2468 40408 2496
rect 39816 2456 39822 2468
rect 40402 2456 40408 2468
rect 40460 2456 40466 2508
rect 41785 2499 41843 2505
rect 41785 2465 41797 2499
rect 41831 2496 41843 2499
rect 41831 2468 41865 2496
rect 41831 2465 41843 2468
rect 41785 2459 41843 2465
rect 38654 2428 38660 2440
rect 38396 2400 38660 2428
rect 37369 2391 37427 2397
rect 38654 2388 38660 2400
rect 38712 2428 38718 2440
rect 39022 2428 39028 2440
rect 38712 2400 39028 2428
rect 38712 2388 38718 2400
rect 39022 2388 39028 2400
rect 39080 2388 39086 2440
rect 41693 2431 41751 2437
rect 41693 2397 41705 2431
rect 41739 2428 41751 2431
rect 41800 2428 41828 2459
rect 41966 2428 41972 2440
rect 41739 2400 41972 2428
rect 41739 2397 41751 2400
rect 41693 2391 41751 2397
rect 41966 2388 41972 2400
rect 42024 2388 42030 2440
rect 42168 2437 42196 2536
rect 42153 2431 42211 2437
rect 42153 2397 42165 2431
rect 42199 2428 42211 2431
rect 42797 2431 42855 2437
rect 42797 2428 42809 2431
rect 42199 2400 42809 2428
rect 42199 2397 42211 2400
rect 42153 2391 42211 2397
rect 42797 2397 42809 2400
rect 42843 2397 42855 2431
rect 42797 2391 42855 2397
rect 30883 2332 32536 2360
rect 42061 2363 42119 2369
rect 30883 2329 30895 2332
rect 30837 2323 30895 2329
rect 42061 2329 42073 2363
rect 42107 2360 42119 2363
rect 43070 2360 43076 2372
rect 42107 2332 43076 2360
rect 42107 2329 42119 2332
rect 42061 2323 42119 2329
rect 43070 2320 43076 2332
rect 43128 2360 43134 2372
rect 43165 2363 43223 2369
rect 43165 2360 43177 2363
rect 43128 2332 43177 2360
rect 43128 2320 43134 2332
rect 43165 2329 43177 2332
rect 43211 2329 43223 2363
rect 43165 2323 43223 2329
rect 22738 2292 22744 2304
rect 17788 2264 22744 2292
rect 22738 2252 22744 2264
rect 22796 2252 22802 2304
rect 22830 2252 22836 2304
rect 22888 2292 22894 2304
rect 23845 2295 23903 2301
rect 23845 2292 23857 2295
rect 22888 2264 23857 2292
rect 22888 2252 22894 2264
rect 23845 2261 23857 2264
rect 23891 2292 23903 2295
rect 24029 2295 24087 2301
rect 24029 2292 24041 2295
rect 23891 2264 24041 2292
rect 23891 2261 23903 2264
rect 23845 2255 23903 2261
rect 24029 2261 24041 2264
rect 24075 2292 24087 2295
rect 24762 2292 24768 2304
rect 24075 2264 24768 2292
rect 24075 2261 24087 2264
rect 24029 2255 24087 2261
rect 24762 2252 24768 2264
rect 24820 2252 24826 2304
rect 32582 2252 32588 2304
rect 32640 2292 32646 2304
rect 33965 2295 34023 2301
rect 33965 2292 33977 2295
rect 32640 2264 33977 2292
rect 32640 2252 32646 2264
rect 33965 2261 33977 2264
rect 34011 2292 34023 2295
rect 34422 2292 34428 2304
rect 34011 2264 34428 2292
rect 34011 2261 34023 2264
rect 33965 2255 34023 2261
rect 34422 2252 34428 2264
rect 34480 2292 34486 2304
rect 34517 2295 34575 2301
rect 34517 2292 34529 2295
rect 34480 2264 34529 2292
rect 34480 2252 34486 2264
rect 34517 2261 34529 2264
rect 34563 2261 34575 2295
rect 34517 2255 34575 2261
rect 37274 2252 37280 2304
rect 37332 2292 37338 2304
rect 37829 2295 37887 2301
rect 37829 2292 37841 2295
rect 37332 2264 37841 2292
rect 37332 2252 37338 2264
rect 37829 2261 37841 2264
rect 37875 2292 37887 2295
rect 38470 2292 38476 2304
rect 37875 2264 38476 2292
rect 37875 2261 37887 2264
rect 37829 2255 37887 2261
rect 38470 2252 38476 2264
rect 38528 2252 38534 2304
rect 41950 2295 42008 2301
rect 41950 2261 41962 2295
rect 41996 2292 42008 2295
rect 42150 2292 42156 2304
rect 41996 2264 42156 2292
rect 41996 2261 42008 2264
rect 41950 2255 42008 2261
rect 42150 2252 42156 2264
rect 42208 2252 42214 2304
rect 42426 2292 42432 2304
rect 42387 2264 42432 2292
rect 42426 2252 42432 2264
rect 42484 2252 42490 2304
rect 43732 2292 43760 2604
rect 43809 2601 43821 2635
rect 43855 2632 43867 2635
rect 43990 2632 43996 2644
rect 43855 2604 43996 2632
rect 43855 2601 43867 2604
rect 43809 2595 43867 2601
rect 43990 2592 43996 2604
rect 44048 2592 44054 2644
rect 46198 2632 46204 2644
rect 46159 2604 46204 2632
rect 46198 2592 46204 2604
rect 46256 2592 46262 2644
rect 46934 2592 46940 2644
rect 46992 2632 46998 2644
rect 47029 2635 47087 2641
rect 47029 2632 47041 2635
rect 46992 2604 47041 2632
rect 46992 2592 46998 2604
rect 47029 2601 47041 2604
rect 47075 2632 47087 2635
rect 48130 2632 48136 2644
rect 47075 2604 48136 2632
rect 47075 2601 47087 2604
rect 47029 2595 47087 2601
rect 48130 2592 48136 2604
rect 48188 2592 48194 2644
rect 49878 2632 49884 2644
rect 49839 2604 49884 2632
rect 49878 2592 49884 2604
rect 49936 2592 49942 2644
rect 51902 2632 51908 2644
rect 51863 2604 51908 2632
rect 51902 2592 51908 2604
rect 51960 2592 51966 2644
rect 51994 2592 52000 2644
rect 52052 2632 52058 2644
rect 53837 2635 53895 2641
rect 53837 2632 53849 2635
rect 52052 2604 53849 2632
rect 52052 2592 52058 2604
rect 53837 2601 53849 2604
rect 53883 2601 53895 2635
rect 54662 2632 54668 2644
rect 54623 2604 54668 2632
rect 53837 2595 53895 2601
rect 54662 2592 54668 2604
rect 54720 2592 54726 2644
rect 54938 2632 54944 2644
rect 54899 2604 54944 2632
rect 54938 2592 54944 2604
rect 54996 2592 55002 2644
rect 55677 2635 55735 2641
rect 55677 2601 55689 2635
rect 55723 2632 55735 2635
rect 57238 2632 57244 2644
rect 55723 2604 57244 2632
rect 55723 2601 55735 2604
rect 55677 2595 55735 2601
rect 57238 2592 57244 2604
rect 57296 2592 57302 2644
rect 58526 2632 58532 2644
rect 58487 2604 58532 2632
rect 58526 2592 58532 2604
rect 58584 2592 58590 2644
rect 62206 2632 62212 2644
rect 62167 2604 62212 2632
rect 62206 2592 62212 2604
rect 62264 2592 62270 2644
rect 44008 2496 44036 2592
rect 45925 2567 45983 2573
rect 45925 2533 45937 2567
rect 45971 2564 45983 2567
rect 47578 2564 47584 2576
rect 45971 2536 47584 2564
rect 45971 2533 45983 2536
rect 45925 2527 45983 2533
rect 47578 2524 47584 2536
rect 47636 2524 47642 2576
rect 48777 2567 48835 2573
rect 48777 2533 48789 2567
rect 48823 2564 48835 2567
rect 49786 2564 49792 2576
rect 48823 2536 49792 2564
rect 48823 2533 48835 2536
rect 48777 2527 48835 2533
rect 49786 2524 49792 2536
rect 49844 2524 49850 2576
rect 50065 2567 50123 2573
rect 50065 2533 50077 2567
rect 50111 2564 50123 2567
rect 50522 2564 50528 2576
rect 50111 2536 50528 2564
rect 50111 2533 50123 2536
rect 50065 2527 50123 2533
rect 50522 2524 50528 2536
rect 50580 2524 50586 2576
rect 50801 2567 50859 2573
rect 50801 2533 50813 2567
rect 50847 2564 50859 2567
rect 51258 2564 51264 2576
rect 50847 2536 51264 2564
rect 50847 2533 50859 2536
rect 50801 2527 50859 2533
rect 51258 2524 51264 2536
rect 51316 2524 51322 2576
rect 52365 2567 52423 2573
rect 52365 2533 52377 2567
rect 52411 2564 52423 2567
rect 53193 2567 53251 2573
rect 53193 2564 53205 2567
rect 52411 2536 53205 2564
rect 52411 2533 52423 2536
rect 52365 2527 52423 2533
rect 53193 2533 53205 2536
rect 53239 2564 53251 2567
rect 53466 2564 53472 2576
rect 53239 2536 53472 2564
rect 53239 2533 53251 2536
rect 53193 2527 53251 2533
rect 53466 2524 53472 2536
rect 53524 2524 53530 2576
rect 58989 2567 59047 2573
rect 58989 2533 59001 2567
rect 59035 2564 59047 2567
rect 59446 2564 59452 2576
rect 59035 2536 59452 2564
rect 59035 2533 59047 2536
rect 58989 2527 59047 2533
rect 59446 2524 59452 2536
rect 59504 2524 59510 2576
rect 44545 2499 44603 2505
rect 44545 2496 44557 2499
rect 44008 2468 44557 2496
rect 44545 2465 44557 2468
rect 44591 2465 44603 2499
rect 46845 2499 46903 2505
rect 46845 2496 46857 2499
rect 44545 2459 44603 2465
rect 46584 2468 46857 2496
rect 44266 2428 44272 2440
rect 44227 2400 44272 2428
rect 44266 2388 44272 2400
rect 44324 2388 44330 2440
rect 46584 2301 46612 2468
rect 46845 2465 46857 2468
rect 46891 2465 46903 2499
rect 46845 2459 46903 2465
rect 47949 2499 48007 2505
rect 47949 2465 47961 2499
rect 47995 2496 48007 2499
rect 48041 2499 48099 2505
rect 48041 2496 48053 2499
rect 47995 2468 48053 2496
rect 47995 2465 48007 2468
rect 47949 2459 48007 2465
rect 48041 2465 48053 2468
rect 48087 2496 48099 2499
rect 49050 2496 49056 2508
rect 48087 2468 49056 2496
rect 48087 2465 48099 2468
rect 48041 2459 48099 2465
rect 49050 2456 49056 2468
rect 49108 2456 49114 2508
rect 50893 2499 50951 2505
rect 50893 2465 50905 2499
rect 50939 2496 50951 2499
rect 51074 2496 51080 2508
rect 50939 2468 51080 2496
rect 50939 2465 50951 2468
rect 50893 2459 50951 2465
rect 51074 2456 51080 2468
rect 51132 2456 51138 2508
rect 53340 2499 53398 2505
rect 53340 2465 53352 2499
rect 53386 2496 53398 2499
rect 53742 2496 53748 2508
rect 53386 2468 53748 2496
rect 53386 2465 53398 2468
rect 53340 2459 53398 2465
rect 53742 2456 53748 2468
rect 53800 2456 53806 2508
rect 59596 2499 59654 2505
rect 59596 2465 59608 2499
rect 59642 2496 59654 2499
rect 60829 2499 60887 2505
rect 60829 2496 60841 2499
rect 59642 2468 60841 2496
rect 59642 2465 59654 2468
rect 59596 2459 59654 2465
rect 60829 2465 60841 2468
rect 60875 2465 60887 2499
rect 60829 2459 60887 2465
rect 61105 2499 61163 2505
rect 61105 2465 61117 2499
rect 61151 2496 61163 2499
rect 61470 2496 61476 2508
rect 61151 2468 61476 2496
rect 61151 2465 61163 2468
rect 61105 2459 61163 2465
rect 48314 2388 48320 2440
rect 48372 2428 48378 2440
rect 48409 2431 48467 2437
rect 48409 2428 48421 2431
rect 48372 2400 48421 2428
rect 48372 2388 48378 2400
rect 48409 2397 48421 2400
rect 48455 2397 48467 2431
rect 48409 2391 48467 2397
rect 49326 2388 49332 2440
rect 49384 2428 49390 2440
rect 50433 2431 50491 2437
rect 50433 2428 50445 2431
rect 49384 2400 50445 2428
rect 49384 2388 49390 2400
rect 50433 2397 50445 2400
rect 50479 2397 50491 2431
rect 50433 2391 50491 2397
rect 47302 2320 47308 2372
rect 47360 2360 47366 2372
rect 47360 2332 48360 2360
rect 47360 2320 47366 2332
rect 48222 2301 48228 2304
rect 46569 2295 46627 2301
rect 46569 2292 46581 2295
rect 43732 2264 46581 2292
rect 46569 2261 46581 2264
rect 46615 2261 46627 2295
rect 46569 2255 46627 2261
rect 47581 2295 47639 2301
rect 47581 2261 47593 2295
rect 47627 2292 47639 2295
rect 48206 2295 48228 2301
rect 48206 2292 48218 2295
rect 47627 2264 48218 2292
rect 47627 2261 47639 2264
rect 47581 2255 47639 2261
rect 48206 2261 48218 2264
rect 48206 2255 48228 2261
rect 48222 2252 48228 2255
rect 48280 2252 48286 2304
rect 48332 2301 48360 2332
rect 49878 2320 49884 2372
rect 49936 2360 49942 2372
rect 50341 2363 50399 2369
rect 50341 2360 50353 2363
rect 49936 2332 50353 2360
rect 49936 2320 49942 2332
rect 50341 2329 50353 2332
rect 50387 2329 50399 2363
rect 50448 2360 50476 2391
rect 50798 2388 50804 2440
rect 50856 2428 50862 2440
rect 53561 2431 53619 2437
rect 53561 2428 53573 2431
rect 50856 2400 53573 2428
rect 50856 2388 50862 2400
rect 53561 2397 53573 2400
rect 53607 2428 53619 2431
rect 54205 2431 54263 2437
rect 54205 2428 54217 2431
rect 53607 2400 54217 2428
rect 53607 2397 53619 2400
rect 53561 2391 53619 2397
rect 54205 2397 54217 2400
rect 54251 2397 54263 2431
rect 54205 2391 54263 2397
rect 56781 2431 56839 2437
rect 56781 2397 56793 2431
rect 56827 2428 56839 2431
rect 57977 2431 58035 2437
rect 57977 2428 57989 2431
rect 56827 2400 57989 2428
rect 56827 2397 56839 2400
rect 56781 2391 56839 2397
rect 57977 2397 57989 2400
rect 58023 2428 58035 2431
rect 58066 2428 58072 2440
rect 58023 2400 58072 2428
rect 58023 2397 58035 2400
rect 57977 2391 58035 2397
rect 58066 2388 58072 2400
rect 58124 2388 58130 2440
rect 58802 2388 58808 2440
rect 58860 2428 58866 2440
rect 59817 2431 59875 2437
rect 59817 2428 59829 2431
rect 58860 2400 59829 2428
rect 58860 2388 58866 2400
rect 59817 2397 59829 2400
rect 59863 2428 59875 2431
rect 60461 2431 60519 2437
rect 60461 2428 60473 2431
rect 59863 2400 60473 2428
rect 59863 2397 59875 2400
rect 59817 2391 59875 2397
rect 60461 2397 60473 2400
rect 60507 2397 60519 2431
rect 60844 2428 60872 2459
rect 61470 2456 61476 2468
rect 61528 2456 61534 2508
rect 62117 2499 62175 2505
rect 62117 2465 62129 2499
rect 62163 2496 62175 2499
rect 62390 2496 62396 2508
rect 62163 2468 62396 2496
rect 62163 2465 62175 2468
rect 62117 2459 62175 2465
rect 62390 2456 62396 2468
rect 62448 2456 62454 2508
rect 61197 2431 61255 2437
rect 61197 2428 61209 2431
rect 60844 2400 61209 2428
rect 60461 2391 60519 2397
rect 61197 2397 61209 2400
rect 61243 2397 61255 2431
rect 61197 2391 61255 2397
rect 51077 2363 51135 2369
rect 51077 2360 51089 2363
rect 50448 2332 51089 2360
rect 50341 2323 50399 2329
rect 51077 2329 51089 2332
rect 51123 2329 51135 2363
rect 51077 2323 51135 2329
rect 53101 2363 53159 2369
rect 53101 2329 53113 2363
rect 53147 2360 53159 2363
rect 59357 2363 59415 2369
rect 53147 2332 53512 2360
rect 53147 2329 53159 2332
rect 53101 2323 53159 2329
rect 53484 2304 53512 2332
rect 59357 2329 59369 2363
rect 59403 2360 59415 2363
rect 59403 2332 59768 2360
rect 59403 2329 59415 2332
rect 59357 2323 59415 2329
rect 59740 2304 59768 2332
rect 48317 2295 48375 2301
rect 48317 2261 48329 2295
rect 48363 2292 48375 2295
rect 49053 2295 49111 2301
rect 49053 2292 49065 2295
rect 48363 2264 49065 2292
rect 48363 2261 48375 2264
rect 48317 2255 48375 2261
rect 49053 2261 49065 2264
rect 49099 2261 49111 2295
rect 49053 2255 49111 2261
rect 49513 2295 49571 2301
rect 49513 2261 49525 2295
rect 49559 2292 49571 2295
rect 50203 2295 50261 2301
rect 50203 2292 50215 2295
rect 49559 2264 50215 2292
rect 49559 2261 49571 2264
rect 49513 2255 49571 2261
rect 50203 2261 50215 2264
rect 50249 2292 50261 2295
rect 50893 2295 50951 2301
rect 50893 2292 50905 2295
rect 50249 2264 50905 2292
rect 50249 2261 50261 2264
rect 50203 2255 50261 2261
rect 50893 2261 50905 2264
rect 50939 2261 50951 2295
rect 51534 2292 51540 2304
rect 51495 2264 51540 2292
rect 50893 2255 50951 2261
rect 51534 2252 51540 2264
rect 51592 2252 51598 2304
rect 53466 2292 53472 2304
rect 53427 2264 53472 2292
rect 53466 2252 53472 2264
rect 53524 2252 53530 2304
rect 55950 2292 55956 2304
rect 55911 2264 55956 2292
rect 55950 2252 55956 2264
rect 56008 2292 56014 2304
rect 56321 2295 56379 2301
rect 56321 2292 56333 2295
rect 56008 2264 56333 2292
rect 56008 2252 56014 2264
rect 56321 2261 56333 2264
rect 56367 2261 56379 2295
rect 59722 2292 59728 2304
rect 59683 2264 59728 2292
rect 56321 2255 56379 2261
rect 59722 2252 59728 2264
rect 59780 2252 59786 2304
rect 59906 2292 59912 2304
rect 59867 2264 59912 2292
rect 59906 2252 59912 2264
rect 59964 2252 59970 2304
rect 61470 2252 61476 2304
rect 61528 2292 61534 2304
rect 61565 2295 61623 2301
rect 61565 2292 61577 2295
rect 61528 2264 61577 2292
rect 61528 2252 61534 2264
rect 61565 2261 61577 2264
rect 61611 2261 61623 2295
rect 61565 2255 61623 2261
rect 62390 2252 62396 2304
rect 62448 2292 62454 2304
rect 62577 2295 62635 2301
rect 62577 2292 62589 2295
rect 62448 2264 62589 2292
rect 62448 2252 62454 2264
rect 62577 2261 62589 2264
rect 62623 2261 62635 2295
rect 62577 2255 62635 2261
rect 1104 2202 63480 2224
rect 1104 2150 11378 2202
rect 11430 2150 11442 2202
rect 11494 2150 11506 2202
rect 11558 2150 11570 2202
rect 11622 2150 32170 2202
rect 32222 2150 32234 2202
rect 32286 2150 32298 2202
rect 32350 2150 32362 2202
rect 32414 2150 52962 2202
rect 53014 2150 53026 2202
rect 53078 2150 53090 2202
rect 53142 2150 53154 2202
rect 53206 2150 63480 2202
rect 1104 2128 63480 2150
rect 2130 2048 2136 2100
rect 2188 2088 2194 2100
rect 9585 2091 9643 2097
rect 9585 2088 9597 2091
rect 2188 2060 9597 2088
rect 2188 2048 2194 2060
rect 9585 2057 9597 2060
rect 9631 2057 9643 2091
rect 9585 2051 9643 2057
rect 15194 2048 15200 2100
rect 15252 2088 15258 2100
rect 15746 2088 15752 2100
rect 15252 2060 15752 2088
rect 15252 2048 15258 2060
rect 15746 2048 15752 2060
rect 15804 2048 15810 2100
rect 42150 2048 42156 2100
rect 42208 2088 42214 2100
rect 42702 2088 42708 2100
rect 42208 2060 42708 2088
rect 42208 2048 42214 2060
rect 42702 2048 42708 2060
rect 42760 2048 42766 2100
rect 48222 2048 48228 2100
rect 48280 2088 48286 2100
rect 49970 2088 49976 2100
rect 48280 2060 49976 2088
rect 48280 2048 48286 2060
rect 49970 2048 49976 2060
rect 50028 2048 50034 2100
rect 51534 2048 51540 2100
rect 51592 2088 51598 2100
rect 59906 2088 59912 2100
rect 51592 2060 59912 2088
rect 51592 2048 51598 2060
rect 59906 2048 59912 2060
rect 59964 2048 59970 2100
rect 9214 1980 9220 2032
rect 9272 2020 9278 2032
rect 19978 2020 19984 2032
rect 9272 1992 19984 2020
rect 9272 1980 9278 1992
rect 19978 1980 19984 1992
rect 20036 1980 20042 2032
rect 42426 1980 42432 2032
rect 42484 2020 42490 2032
rect 49326 2020 49332 2032
rect 42484 1992 49332 2020
rect 42484 1980 42490 1992
rect 49326 1980 49332 1992
rect 49384 1980 49390 2032
rect 9585 1955 9643 1961
rect 9585 1921 9597 1955
rect 9631 1952 9643 1955
rect 15286 1952 15292 1964
rect 9631 1924 15292 1952
rect 9631 1921 9643 1924
rect 9585 1915 9643 1921
rect 15286 1912 15292 1924
rect 15344 1912 15350 1964
rect 40494 1912 40500 1964
rect 40552 1952 40558 1964
rect 44266 1952 44272 1964
rect 40552 1924 44272 1952
rect 40552 1912 40558 1924
rect 44266 1912 44272 1924
rect 44324 1952 44330 1964
rect 55950 1952 55956 1964
rect 44324 1924 55956 1952
rect 44324 1912 44330 1924
rect 55950 1912 55956 1924
rect 56008 1912 56014 1964
rect 15304 1816 15332 1912
rect 16298 1844 16304 1896
rect 16356 1884 16362 1896
rect 17586 1884 17592 1896
rect 16356 1856 17592 1884
rect 16356 1844 16362 1856
rect 17586 1844 17592 1856
rect 17644 1844 17650 1896
rect 21450 1816 21456 1828
rect 15304 1788 21456 1816
rect 21450 1776 21456 1788
rect 21508 1776 21514 1828
rect 1210 1368 1216 1420
rect 1268 1408 1274 1420
rect 7282 1408 7288 1420
rect 1268 1380 7288 1408
rect 1268 1368 1274 1380
rect 7282 1368 7288 1380
rect 7340 1368 7346 1420
rect 32214 1368 32220 1420
rect 32272 1408 32278 1420
rect 36906 1408 36912 1420
rect 32272 1380 36912 1408
rect 32272 1368 32278 1380
rect 36906 1368 36912 1380
rect 36964 1368 36970 1420
rect 4062 1300 4068 1352
rect 4120 1340 4126 1352
rect 24946 1340 24952 1352
rect 4120 1312 24952 1340
rect 4120 1300 4126 1312
rect 24946 1300 24952 1312
rect 25004 1300 25010 1352
rect 30466 1300 30472 1352
rect 30524 1340 30530 1352
rect 32766 1340 32772 1352
rect 30524 1312 32772 1340
rect 30524 1300 30530 1312
rect 32766 1300 32772 1312
rect 32824 1300 32830 1352
<< via1 >>
rect 11378 17382 11430 17434
rect 11442 17382 11494 17434
rect 11506 17382 11558 17434
rect 11570 17382 11622 17434
rect 32170 17382 32222 17434
rect 32234 17382 32286 17434
rect 32298 17382 32350 17434
rect 32362 17382 32414 17434
rect 52962 17382 53014 17434
rect 53026 17382 53078 17434
rect 53090 17382 53142 17434
rect 53154 17382 53206 17434
rect 14648 17280 14700 17332
rect 19156 17212 19208 17264
rect 12256 17144 12308 17196
rect 15752 17144 15804 17196
rect 22744 17212 22796 17264
rect 24400 17280 24452 17332
rect 28356 17280 28408 17332
rect 28908 17280 28960 17332
rect 42064 17280 42116 17332
rect 45928 17280 45980 17332
rect 48136 17280 48188 17332
rect 53840 17280 53892 17332
rect 33784 17255 33836 17264
rect 33784 17221 33793 17255
rect 33793 17221 33827 17255
rect 33827 17221 33836 17255
rect 33784 17212 33836 17221
rect 49976 17255 50028 17264
rect 49976 17221 49985 17255
rect 49985 17221 50019 17255
rect 50019 17221 50028 17255
rect 49976 17212 50028 17221
rect 13912 17076 13964 17128
rect 18512 17076 18564 17128
rect 18328 17051 18380 17060
rect 18328 17017 18337 17051
rect 18337 17017 18371 17051
rect 18371 17017 18380 17051
rect 18328 17008 18380 17017
rect 19248 17008 19300 17060
rect 22744 17119 22796 17128
rect 22744 17085 22753 17119
rect 22753 17085 22787 17119
rect 22787 17085 22796 17119
rect 22744 17076 22796 17085
rect 23112 17076 23164 17128
rect 27528 17144 27580 17196
rect 23572 17008 23624 17060
rect 20444 16940 20496 16992
rect 20720 16983 20772 16992
rect 20720 16949 20729 16983
rect 20729 16949 20763 16983
rect 20763 16949 20772 16983
rect 20720 16940 20772 16949
rect 28356 17076 28408 17128
rect 28724 17076 28776 17128
rect 30564 17119 30616 17128
rect 30564 17085 30573 17119
rect 30573 17085 30607 17119
rect 30607 17085 30616 17119
rect 30564 17076 30616 17085
rect 30748 17076 30800 17128
rect 34244 17144 34296 17196
rect 34152 17119 34204 17128
rect 34152 17085 34161 17119
rect 34161 17085 34195 17119
rect 34195 17085 34204 17119
rect 34152 17076 34204 17085
rect 34336 17119 34388 17128
rect 34336 17085 34345 17119
rect 34345 17085 34379 17119
rect 34379 17085 34388 17119
rect 34336 17076 34388 17085
rect 39488 17119 39540 17128
rect 39488 17085 39497 17119
rect 39497 17085 39531 17119
rect 39531 17085 39540 17119
rect 39488 17076 39540 17085
rect 39028 17051 39080 17060
rect 39028 17017 39037 17051
rect 39037 17017 39071 17051
rect 39071 17017 39080 17051
rect 39028 17008 39080 17017
rect 29368 16983 29420 16992
rect 29368 16949 29377 16983
rect 29377 16949 29411 16983
rect 29411 16949 29420 16983
rect 29368 16940 29420 16949
rect 39212 16940 39264 16992
rect 39856 17119 39908 17128
rect 39856 17085 39865 17119
rect 39865 17085 39899 17119
rect 39899 17085 39908 17119
rect 39856 17076 39908 17085
rect 40224 17076 40276 17128
rect 43628 17076 43680 17128
rect 46940 17076 46992 17128
rect 47124 17119 47176 17128
rect 47124 17085 47133 17119
rect 47133 17085 47167 17119
rect 47167 17085 47176 17119
rect 47124 17076 47176 17085
rect 49884 17076 49936 17128
rect 50344 17119 50396 17128
rect 50344 17085 50353 17119
rect 50353 17085 50387 17119
rect 50387 17085 50396 17119
rect 50344 17076 50396 17085
rect 48780 17008 48832 17060
rect 43076 16983 43128 16992
rect 43076 16949 43085 16983
rect 43085 16949 43119 16983
rect 43119 16949 43128 16983
rect 43076 16940 43128 16949
rect 52828 17008 52880 17060
rect 53932 17076 53984 17128
rect 53472 16940 53524 16992
rect 21774 16838 21826 16890
rect 21838 16838 21890 16890
rect 21902 16838 21954 16890
rect 21966 16838 22018 16890
rect 42566 16838 42618 16890
rect 42630 16838 42682 16890
rect 42694 16838 42746 16890
rect 42758 16838 42810 16890
rect 12624 16779 12676 16788
rect 12624 16745 12633 16779
rect 12633 16745 12667 16779
rect 12667 16745 12676 16779
rect 12624 16736 12676 16745
rect 16672 16736 16724 16788
rect 17132 16779 17184 16788
rect 17132 16745 17141 16779
rect 17141 16745 17175 16779
rect 17175 16745 17184 16779
rect 17132 16736 17184 16745
rect 19248 16736 19300 16788
rect 22468 16779 22520 16788
rect 22468 16745 22477 16779
rect 22477 16745 22511 16779
rect 22511 16745 22520 16779
rect 22468 16736 22520 16745
rect 24492 16736 24544 16788
rect 34244 16736 34296 16788
rect 40132 16736 40184 16788
rect 48780 16779 48832 16788
rect 48780 16745 48789 16779
rect 48789 16745 48823 16779
rect 48823 16745 48832 16779
rect 48780 16736 48832 16745
rect 49884 16736 49936 16788
rect 53932 16736 53984 16788
rect 8116 16600 8168 16652
rect 7932 16532 7984 16584
rect 9496 16600 9548 16652
rect 12256 16600 12308 16652
rect 13912 16600 13964 16652
rect 18052 16643 18104 16652
rect 18052 16609 18061 16643
rect 18061 16609 18095 16643
rect 18095 16609 18104 16643
rect 18052 16600 18104 16609
rect 22100 16600 22152 16652
rect 11244 16532 11296 16584
rect 15752 16575 15804 16584
rect 15752 16541 15761 16575
rect 15761 16541 15795 16575
rect 15795 16541 15804 16575
rect 15752 16532 15804 16541
rect 16028 16575 16080 16584
rect 16028 16541 16037 16575
rect 16037 16541 16071 16575
rect 16071 16541 16080 16575
rect 16028 16532 16080 16541
rect 18512 16575 18564 16584
rect 18512 16541 18521 16575
rect 18521 16541 18555 16575
rect 18555 16541 18564 16575
rect 18512 16532 18564 16541
rect 19984 16532 20036 16584
rect 20720 16532 20772 16584
rect 21456 16532 21508 16584
rect 25044 16600 25096 16652
rect 30288 16643 30340 16652
rect 30288 16609 30297 16643
rect 30297 16609 30331 16643
rect 30331 16609 30340 16643
rect 30288 16600 30340 16609
rect 30656 16643 30708 16652
rect 30656 16609 30665 16643
rect 30665 16609 30699 16643
rect 30699 16609 30708 16643
rect 30656 16600 30708 16609
rect 33324 16600 33376 16652
rect 34152 16600 34204 16652
rect 47308 16600 47360 16652
rect 47952 16668 48004 16720
rect 23848 16575 23900 16584
rect 23848 16541 23857 16575
rect 23857 16541 23891 16575
rect 23891 16541 23900 16575
rect 23848 16532 23900 16541
rect 27620 16575 27672 16584
rect 27620 16541 27629 16575
rect 27629 16541 27663 16575
rect 27663 16541 27672 16575
rect 27620 16532 27672 16541
rect 30748 16575 30800 16584
rect 30748 16541 30757 16575
rect 30757 16541 30791 16575
rect 30791 16541 30800 16575
rect 30748 16532 30800 16541
rect 31944 16532 31996 16584
rect 32588 16532 32640 16584
rect 34612 16575 34664 16584
rect 34612 16541 34621 16575
rect 34621 16541 34655 16575
rect 34655 16541 34664 16575
rect 34612 16532 34664 16541
rect 35072 16532 35124 16584
rect 8208 16464 8260 16516
rect 4804 16396 4856 16448
rect 9036 16439 9088 16448
rect 9036 16405 9045 16439
rect 9045 16405 9079 16439
rect 9079 16405 9088 16439
rect 9036 16396 9088 16405
rect 9496 16439 9548 16448
rect 9496 16405 9505 16439
rect 9505 16405 9539 16439
rect 9539 16405 9548 16439
rect 9496 16396 9548 16405
rect 10876 16439 10928 16448
rect 10876 16405 10885 16439
rect 10885 16405 10919 16439
rect 10919 16405 10928 16439
rect 10876 16396 10928 16405
rect 26332 16464 26384 16516
rect 30104 16507 30156 16516
rect 11980 16396 12032 16448
rect 14280 16439 14332 16448
rect 14280 16405 14289 16439
rect 14289 16405 14323 16439
rect 14323 16405 14332 16439
rect 14280 16396 14332 16405
rect 20352 16439 20404 16448
rect 20352 16405 20361 16439
rect 20361 16405 20395 16439
rect 20395 16405 20404 16439
rect 20352 16396 20404 16405
rect 22560 16396 22612 16448
rect 22744 16396 22796 16448
rect 25412 16396 25464 16448
rect 26148 16396 26200 16448
rect 30104 16473 30113 16507
rect 30113 16473 30147 16507
rect 30147 16473 30156 16507
rect 30104 16464 30156 16473
rect 28724 16439 28776 16448
rect 28724 16405 28733 16439
rect 28733 16405 28767 16439
rect 28767 16405 28776 16439
rect 28724 16396 28776 16405
rect 29552 16439 29604 16448
rect 29552 16405 29561 16439
rect 29561 16405 29595 16439
rect 29595 16405 29604 16439
rect 29552 16396 29604 16405
rect 31116 16439 31168 16448
rect 31116 16405 31125 16439
rect 31125 16405 31159 16439
rect 31159 16405 31168 16439
rect 31116 16396 31168 16405
rect 32496 16396 32548 16448
rect 32864 16396 32916 16448
rect 33692 16396 33744 16448
rect 37372 16439 37424 16448
rect 37372 16405 37381 16439
rect 37381 16405 37415 16439
rect 37415 16405 37424 16439
rect 37372 16396 37424 16405
rect 38108 16532 38160 16584
rect 38200 16532 38252 16584
rect 39488 16532 39540 16584
rect 40224 16575 40276 16584
rect 38476 16396 38528 16448
rect 40224 16541 40233 16575
rect 40233 16541 40267 16575
rect 40267 16541 40276 16575
rect 40224 16532 40276 16541
rect 40960 16532 41012 16584
rect 47032 16532 47084 16584
rect 48228 16532 48280 16584
rect 49424 16532 49476 16584
rect 41604 16464 41656 16516
rect 43076 16464 43128 16516
rect 47216 16464 47268 16516
rect 53380 16600 53432 16652
rect 52092 16575 52144 16584
rect 39856 16396 39908 16448
rect 40684 16396 40736 16448
rect 42156 16439 42208 16448
rect 42156 16405 42165 16439
rect 42165 16405 42199 16439
rect 42199 16405 42208 16439
rect 42156 16396 42208 16405
rect 46940 16439 46992 16448
rect 46940 16405 46949 16439
rect 46949 16405 46983 16439
rect 46983 16405 46992 16439
rect 46940 16396 46992 16405
rect 47400 16396 47452 16448
rect 48320 16439 48372 16448
rect 48320 16405 48329 16439
rect 48329 16405 48363 16439
rect 48363 16405 48372 16439
rect 48320 16396 48372 16405
rect 50620 16464 50672 16516
rect 52092 16541 52101 16575
rect 52101 16541 52135 16575
rect 52135 16541 52144 16575
rect 52092 16532 52144 16541
rect 49700 16396 49752 16448
rect 50344 16396 50396 16448
rect 51816 16396 51868 16448
rect 53288 16396 53340 16448
rect 53748 16439 53800 16448
rect 53748 16405 53757 16439
rect 53757 16405 53791 16439
rect 53791 16405 53800 16439
rect 53748 16396 53800 16405
rect 11378 16294 11430 16346
rect 11442 16294 11494 16346
rect 11506 16294 11558 16346
rect 11570 16294 11622 16346
rect 32170 16294 32222 16346
rect 32234 16294 32286 16346
rect 32298 16294 32350 16346
rect 32362 16294 32414 16346
rect 52962 16294 53014 16346
rect 53026 16294 53078 16346
rect 53090 16294 53142 16346
rect 53154 16294 53206 16346
rect 8116 16192 8168 16244
rect 10692 16192 10744 16244
rect 11244 16235 11296 16244
rect 11244 16201 11253 16235
rect 11253 16201 11287 16235
rect 11287 16201 11296 16235
rect 11244 16192 11296 16201
rect 12256 16235 12308 16244
rect 12256 16201 12265 16235
rect 12265 16201 12299 16235
rect 12299 16201 12308 16235
rect 12256 16192 12308 16201
rect 14648 16235 14700 16244
rect 14648 16201 14657 16235
rect 14657 16201 14691 16235
rect 14691 16201 14700 16235
rect 14648 16192 14700 16201
rect 16028 16192 16080 16244
rect 18052 16192 18104 16244
rect 19984 16235 20036 16244
rect 19984 16201 19993 16235
rect 19993 16201 20027 16235
rect 20027 16201 20036 16235
rect 19984 16192 20036 16201
rect 20536 16192 20588 16244
rect 20996 16192 21048 16244
rect 49700 16235 49752 16244
rect 940 15852 992 15904
rect 3608 15852 3660 15904
rect 7288 15852 7340 15904
rect 9036 16056 9088 16108
rect 19800 16124 19852 16176
rect 21088 16124 21140 16176
rect 22376 16124 22428 16176
rect 22560 16124 22612 16176
rect 25412 16167 25464 16176
rect 25412 16133 25421 16167
rect 25421 16133 25455 16167
rect 25455 16133 25464 16167
rect 25412 16124 25464 16133
rect 27620 16124 27672 16176
rect 10876 16031 10928 16040
rect 10876 15997 10885 16031
rect 10885 15997 10919 16031
rect 10919 15997 10928 16031
rect 10876 15988 10928 15997
rect 12256 15988 12308 16040
rect 14648 16056 14700 16108
rect 16764 16056 16816 16108
rect 17040 16056 17092 16108
rect 18052 16056 18104 16108
rect 11152 15920 11204 15972
rect 13360 15963 13412 15972
rect 13360 15929 13369 15963
rect 13369 15929 13403 15963
rect 13403 15929 13412 15963
rect 13360 15920 13412 15929
rect 7932 15852 7984 15904
rect 13268 15852 13320 15904
rect 14280 16031 14332 16040
rect 14280 15997 14289 16031
rect 14289 15997 14323 16031
rect 14323 15997 14332 16031
rect 14280 15988 14332 15997
rect 16396 15988 16448 16040
rect 17132 15988 17184 16040
rect 19156 15988 19208 16040
rect 20352 16031 20404 16040
rect 20352 15997 20361 16031
rect 20361 15997 20395 16031
rect 20395 15997 20404 16031
rect 20352 15988 20404 15997
rect 23664 16031 23716 16040
rect 23664 15997 23673 16031
rect 23673 15997 23707 16031
rect 23707 15997 23716 16031
rect 23664 15988 23716 15997
rect 23848 16056 23900 16108
rect 25044 16099 25096 16108
rect 25044 16065 25053 16099
rect 25053 16065 25087 16099
rect 25087 16065 25096 16099
rect 25044 16056 25096 16065
rect 26148 16056 26200 16108
rect 15568 15852 15620 15904
rect 15752 15895 15804 15904
rect 15752 15861 15761 15895
rect 15761 15861 15795 15895
rect 15795 15861 15804 15895
rect 15752 15852 15804 15861
rect 22100 15963 22152 15972
rect 22100 15929 22109 15963
rect 22109 15929 22143 15963
rect 22143 15929 22152 15963
rect 22100 15920 22152 15929
rect 22560 15920 22612 15972
rect 23572 15920 23624 15972
rect 24124 15988 24176 16040
rect 26976 15988 27028 16040
rect 27068 15988 27120 16040
rect 29276 16124 29328 16176
rect 30288 16124 30340 16176
rect 30748 16124 30800 16176
rect 32680 16124 32732 16176
rect 33692 16167 33744 16176
rect 28356 16099 28408 16108
rect 28356 16065 28365 16099
rect 28365 16065 28399 16099
rect 28399 16065 28408 16099
rect 28356 16056 28408 16065
rect 33324 16099 33376 16108
rect 28264 15988 28316 16040
rect 29368 15988 29420 16040
rect 29552 16031 29604 16040
rect 29552 15997 29561 16031
rect 29561 15997 29595 16031
rect 29595 15997 29604 16031
rect 29552 15988 29604 15997
rect 20444 15852 20496 15904
rect 23664 15852 23716 15904
rect 27712 15852 27764 15904
rect 28540 15852 28592 15904
rect 29368 15852 29420 15904
rect 30656 15852 30708 15904
rect 32864 16031 32916 16040
rect 32864 15997 32873 16031
rect 32873 15997 32907 16031
rect 32907 15997 32916 16031
rect 32864 15988 32916 15997
rect 33324 16065 33333 16099
rect 33333 16065 33367 16099
rect 33367 16065 33376 16099
rect 33324 16056 33376 16065
rect 33692 16133 33701 16167
rect 33701 16133 33735 16167
rect 33735 16133 33744 16167
rect 33692 16124 33744 16133
rect 35716 16124 35768 16176
rect 40132 16124 40184 16176
rect 43444 16167 43496 16176
rect 43444 16133 43453 16167
rect 43453 16133 43487 16167
rect 43487 16133 43496 16167
rect 43444 16124 43496 16133
rect 43996 16124 44048 16176
rect 47032 16124 47084 16176
rect 47308 16124 47360 16176
rect 34336 15988 34388 16040
rect 37372 16031 37424 16040
rect 37372 15997 37381 16031
rect 37381 15997 37415 16031
rect 37415 15997 37424 16031
rect 37372 15988 37424 15997
rect 32312 15920 32364 15972
rect 33692 15920 33744 15972
rect 38936 15988 38988 16040
rect 41604 16056 41656 16108
rect 39212 16031 39264 16040
rect 39212 15997 39221 16031
rect 39221 15997 39255 16031
rect 39255 15997 39264 16031
rect 39212 15988 39264 15997
rect 42156 16031 42208 16040
rect 38660 15920 38712 15972
rect 42156 15997 42165 16031
rect 42165 15997 42199 16031
rect 42199 15997 42208 16031
rect 42156 15988 42208 15997
rect 46204 16031 46256 16040
rect 46204 15997 46213 16031
rect 46213 15997 46247 16031
rect 46247 15997 46256 16031
rect 46756 16031 46808 16040
rect 46204 15988 46256 15997
rect 46756 15997 46765 16031
rect 46765 15997 46799 16031
rect 46799 15997 46808 16031
rect 46756 15988 46808 15997
rect 47400 15988 47452 16040
rect 48320 16056 48372 16108
rect 49700 16201 49709 16235
rect 49709 16201 49743 16235
rect 49743 16201 49752 16235
rect 49700 16192 49752 16201
rect 52092 16192 52144 16244
rect 53932 16192 53984 16244
rect 51632 16124 51684 16176
rect 51448 15988 51500 16040
rect 51540 16031 51592 16040
rect 51540 15997 51549 16031
rect 51549 15997 51583 16031
rect 51583 15997 51592 16031
rect 51540 15988 51592 15997
rect 52460 15988 52512 16040
rect 53748 16056 53800 16108
rect 31944 15895 31996 15904
rect 31944 15861 31953 15895
rect 31953 15861 31987 15895
rect 31987 15861 31996 15895
rect 31944 15852 31996 15861
rect 32588 15852 32640 15904
rect 32772 15852 32824 15904
rect 34612 15895 34664 15904
rect 34612 15861 34621 15895
rect 34621 15861 34655 15895
rect 34655 15861 34664 15895
rect 34612 15852 34664 15861
rect 35072 15895 35124 15904
rect 35072 15861 35081 15895
rect 35081 15861 35115 15895
rect 35115 15861 35124 15895
rect 35072 15852 35124 15861
rect 35624 15852 35676 15904
rect 35900 15852 35952 15904
rect 37924 15852 37976 15904
rect 38108 15895 38160 15904
rect 38108 15861 38117 15895
rect 38117 15861 38151 15895
rect 38151 15861 38160 15895
rect 38108 15852 38160 15861
rect 40776 15852 40828 15904
rect 41052 15895 41104 15904
rect 41052 15861 41061 15895
rect 41061 15861 41095 15895
rect 41095 15861 41104 15895
rect 41052 15852 41104 15861
rect 41604 15895 41656 15904
rect 41604 15861 41613 15895
rect 41613 15861 41647 15895
rect 41647 15861 41656 15895
rect 41604 15852 41656 15861
rect 47952 15852 48004 15904
rect 49424 15852 49476 15904
rect 50620 15852 50672 15904
rect 50988 15852 51040 15904
rect 51080 15852 51132 15904
rect 52644 15852 52696 15904
rect 57152 15988 57204 16040
rect 53380 15852 53432 15904
rect 56968 15852 57020 15904
rect 21774 15750 21826 15802
rect 21838 15750 21890 15802
rect 21902 15750 21954 15802
rect 21966 15750 22018 15802
rect 42566 15750 42618 15802
rect 42630 15750 42682 15802
rect 42694 15750 42746 15802
rect 42758 15750 42810 15802
rect 6736 15648 6788 15700
rect 7840 15648 7892 15700
rect 10876 15648 10928 15700
rect 8208 15623 8260 15632
rect 8208 15589 8217 15623
rect 8217 15589 8251 15623
rect 8251 15589 8260 15623
rect 8208 15580 8260 15589
rect 9036 15580 9088 15632
rect 8300 15555 8352 15564
rect 8300 15521 8309 15555
rect 8309 15521 8343 15555
rect 8343 15521 8352 15555
rect 8300 15512 8352 15521
rect 5356 15487 5408 15496
rect 5356 15453 5365 15487
rect 5365 15453 5399 15487
rect 5399 15453 5408 15487
rect 5356 15444 5408 15453
rect 5632 15487 5684 15496
rect 5632 15453 5641 15487
rect 5641 15453 5675 15487
rect 5675 15453 5684 15487
rect 5632 15444 5684 15453
rect 7288 15444 7340 15496
rect 12164 15512 12216 15564
rect 14280 15648 14332 15700
rect 19156 15691 19208 15700
rect 19156 15657 19165 15691
rect 19165 15657 19199 15691
rect 19199 15657 19208 15691
rect 19156 15648 19208 15657
rect 13360 15580 13412 15632
rect 11244 15487 11296 15496
rect 11244 15453 11253 15487
rect 11253 15453 11287 15487
rect 11287 15453 11296 15487
rect 11244 15444 11296 15453
rect 14004 15512 14056 15564
rect 15200 15512 15252 15564
rect 14096 15444 14148 15496
rect 15752 15444 15804 15496
rect 18328 15580 18380 15632
rect 18512 15580 18564 15632
rect 19340 15512 19392 15564
rect 19524 15555 19576 15564
rect 19524 15521 19533 15555
rect 19533 15521 19567 15555
rect 19567 15521 19576 15555
rect 19524 15512 19576 15521
rect 23572 15648 23624 15700
rect 19800 15555 19852 15564
rect 19800 15521 19809 15555
rect 19809 15521 19843 15555
rect 19843 15521 19852 15555
rect 21088 15580 21140 15632
rect 21456 15623 21508 15632
rect 21456 15589 21465 15623
rect 21465 15589 21499 15623
rect 21499 15589 21508 15623
rect 21456 15580 21508 15589
rect 23112 15580 23164 15632
rect 26976 15648 27028 15700
rect 30288 15648 30340 15700
rect 31116 15691 31168 15700
rect 31116 15657 31125 15691
rect 31125 15657 31159 15691
rect 31159 15657 31168 15691
rect 31116 15648 31168 15657
rect 31944 15691 31996 15700
rect 31944 15657 31953 15691
rect 31953 15657 31987 15691
rect 31987 15657 31996 15691
rect 31944 15648 31996 15657
rect 32772 15648 32824 15700
rect 33692 15691 33744 15700
rect 33692 15657 33701 15691
rect 33701 15657 33735 15691
rect 33735 15657 33744 15691
rect 33692 15648 33744 15657
rect 26056 15623 26108 15632
rect 26056 15589 26065 15623
rect 26065 15589 26099 15623
rect 26099 15589 26108 15623
rect 26056 15580 26108 15589
rect 27160 15623 27212 15632
rect 27160 15589 27169 15623
rect 27169 15589 27203 15623
rect 27203 15589 27212 15623
rect 27160 15580 27212 15589
rect 27528 15580 27580 15632
rect 27620 15580 27672 15632
rect 28172 15580 28224 15632
rect 28540 15623 28592 15632
rect 28540 15589 28549 15623
rect 28549 15589 28583 15623
rect 28583 15589 28592 15623
rect 28540 15580 28592 15589
rect 19800 15512 19852 15521
rect 20444 15512 20496 15564
rect 32312 15623 32364 15632
rect 32312 15589 32321 15623
rect 32321 15589 32355 15623
rect 32355 15589 32364 15623
rect 32312 15580 32364 15589
rect 33784 15580 33836 15632
rect 36176 15648 36228 15700
rect 40040 15648 40092 15700
rect 40224 15648 40276 15700
rect 41604 15648 41656 15700
rect 47216 15691 47268 15700
rect 47216 15657 47225 15691
rect 47225 15657 47259 15691
rect 47259 15657 47268 15691
rect 47216 15648 47268 15657
rect 35072 15580 35124 15632
rect 24124 15512 24176 15564
rect 24676 15512 24728 15564
rect 27068 15555 27120 15564
rect 7196 15376 7248 15428
rect 7472 15376 7524 15428
rect 10876 15376 10928 15428
rect 7656 15351 7708 15360
rect 7656 15317 7665 15351
rect 7665 15317 7699 15351
rect 7699 15317 7708 15351
rect 7656 15308 7708 15317
rect 8944 15308 8996 15360
rect 9496 15308 9548 15360
rect 10508 15308 10560 15360
rect 11980 15308 12032 15360
rect 13820 15376 13872 15428
rect 16120 15376 16172 15428
rect 16396 15376 16448 15428
rect 16856 15376 16908 15428
rect 13268 15351 13320 15360
rect 13268 15317 13277 15351
rect 13277 15317 13311 15351
rect 13311 15317 13320 15351
rect 13268 15308 13320 15317
rect 13912 15351 13964 15360
rect 13912 15317 13921 15351
rect 13921 15317 13955 15351
rect 13955 15317 13964 15351
rect 13912 15308 13964 15317
rect 16764 15308 16816 15360
rect 17868 15308 17920 15360
rect 18144 15376 18196 15428
rect 19800 15308 19852 15360
rect 21640 15487 21692 15496
rect 21640 15453 21649 15487
rect 21649 15453 21683 15487
rect 21683 15453 21692 15487
rect 21640 15444 21692 15453
rect 22008 15487 22060 15496
rect 22008 15453 22017 15487
rect 22017 15453 22051 15487
rect 22051 15453 22060 15487
rect 22008 15444 22060 15453
rect 23296 15351 23348 15360
rect 23296 15317 23305 15351
rect 23305 15317 23339 15351
rect 23339 15317 23348 15351
rect 23296 15308 23348 15317
rect 23664 15351 23716 15360
rect 23664 15317 23673 15351
rect 23673 15317 23707 15351
rect 23707 15317 23716 15351
rect 23664 15308 23716 15317
rect 25044 15308 25096 15360
rect 25964 15308 26016 15360
rect 27068 15521 27077 15555
rect 27077 15521 27111 15555
rect 27111 15521 27120 15555
rect 27068 15512 27120 15521
rect 28080 15512 28132 15564
rect 28908 15512 28960 15564
rect 29184 15555 29236 15564
rect 29184 15521 29193 15555
rect 29193 15521 29227 15555
rect 29227 15521 29236 15555
rect 29184 15512 29236 15521
rect 29368 15555 29420 15564
rect 29368 15521 29377 15555
rect 29377 15521 29411 15555
rect 29411 15521 29420 15555
rect 29368 15512 29420 15521
rect 31300 15512 31352 15564
rect 31760 15512 31812 15564
rect 34796 15512 34848 15564
rect 36544 15555 36596 15564
rect 27436 15444 27488 15496
rect 29276 15444 29328 15496
rect 32036 15444 32088 15496
rect 36544 15521 36553 15555
rect 36553 15521 36587 15555
rect 36587 15521 36596 15555
rect 36544 15512 36596 15521
rect 43444 15580 43496 15632
rect 48780 15648 48832 15700
rect 49976 15691 50028 15700
rect 48320 15580 48372 15632
rect 49976 15657 49985 15691
rect 49985 15657 50019 15691
rect 50019 15657 50028 15691
rect 49976 15648 50028 15657
rect 52460 15691 52512 15700
rect 52460 15657 52469 15691
rect 52469 15657 52503 15691
rect 52503 15657 52512 15691
rect 52460 15648 52512 15657
rect 54024 15691 54076 15700
rect 54024 15657 54033 15691
rect 54033 15657 54067 15691
rect 54067 15657 54076 15691
rect 54024 15648 54076 15657
rect 50712 15580 50764 15632
rect 52644 15623 52696 15632
rect 52644 15589 52653 15623
rect 52653 15589 52687 15623
rect 52687 15589 52696 15623
rect 52644 15580 52696 15589
rect 42248 15555 42300 15564
rect 30748 15376 30800 15428
rect 35716 15444 35768 15496
rect 38476 15444 38528 15496
rect 40132 15444 40184 15496
rect 42248 15521 42257 15555
rect 42257 15521 42291 15555
rect 42291 15521 42300 15555
rect 42248 15512 42300 15521
rect 46204 15555 46256 15564
rect 46204 15521 46213 15555
rect 46213 15521 46247 15555
rect 46247 15521 46256 15555
rect 46204 15512 46256 15521
rect 47584 15555 47636 15564
rect 47584 15521 47593 15555
rect 47593 15521 47627 15555
rect 47627 15521 47636 15555
rect 47584 15512 47636 15521
rect 49608 15512 49660 15564
rect 51632 15555 51684 15564
rect 32588 15351 32640 15360
rect 32588 15317 32597 15351
rect 32597 15317 32631 15351
rect 32631 15317 32640 15351
rect 32588 15308 32640 15317
rect 32864 15308 32916 15360
rect 34336 15308 34388 15360
rect 35164 15351 35216 15360
rect 35164 15317 35173 15351
rect 35173 15317 35207 15351
rect 35207 15317 35216 15351
rect 35164 15308 35216 15317
rect 36176 15351 36228 15360
rect 36176 15317 36185 15351
rect 36185 15317 36219 15351
rect 36219 15317 36228 15351
rect 36176 15308 36228 15317
rect 37188 15351 37240 15360
rect 37188 15317 37197 15351
rect 37197 15317 37231 15351
rect 37231 15317 37240 15351
rect 37188 15308 37240 15317
rect 37464 15351 37516 15360
rect 37464 15317 37473 15351
rect 37473 15317 37507 15351
rect 37507 15317 37516 15351
rect 37464 15308 37516 15317
rect 38016 15308 38068 15360
rect 39856 15376 39908 15428
rect 42340 15444 42392 15496
rect 50252 15444 50304 15496
rect 41696 15419 41748 15428
rect 41696 15385 41705 15419
rect 41705 15385 41739 15419
rect 41739 15385 41748 15419
rect 41696 15376 41748 15385
rect 48780 15376 48832 15428
rect 51632 15521 51641 15555
rect 51641 15521 51675 15555
rect 51675 15521 51684 15555
rect 51632 15512 51684 15521
rect 53288 15512 53340 15564
rect 53472 15555 53524 15564
rect 53472 15521 53481 15555
rect 53481 15521 53515 15555
rect 53515 15521 53524 15555
rect 53472 15512 53524 15521
rect 51724 15487 51776 15496
rect 51724 15453 51733 15487
rect 51733 15453 51767 15487
rect 51767 15453 51776 15487
rect 51724 15444 51776 15453
rect 51356 15376 51408 15428
rect 61660 15648 61712 15700
rect 57704 15580 57756 15632
rect 56876 15555 56928 15564
rect 56876 15521 56885 15555
rect 56885 15521 56919 15555
rect 56919 15521 56928 15555
rect 56876 15512 56928 15521
rect 56968 15512 57020 15564
rect 55864 15444 55916 15496
rect 56784 15444 56836 15496
rect 58164 15444 58216 15496
rect 58900 15376 58952 15428
rect 59728 15376 59780 15428
rect 38936 15308 38988 15360
rect 40500 15351 40552 15360
rect 40500 15317 40509 15351
rect 40509 15317 40543 15351
rect 40543 15317 40552 15351
rect 40500 15308 40552 15317
rect 42892 15351 42944 15360
rect 42892 15317 42901 15351
rect 42901 15317 42935 15351
rect 42935 15317 42944 15351
rect 42892 15308 42944 15317
rect 43076 15308 43128 15360
rect 43904 15351 43956 15360
rect 43904 15317 43913 15351
rect 43913 15317 43947 15351
rect 43947 15317 43956 15351
rect 43904 15308 43956 15317
rect 47308 15351 47360 15360
rect 47308 15317 47317 15351
rect 47317 15317 47351 15351
rect 47351 15317 47360 15351
rect 47308 15308 47360 15317
rect 49148 15308 49200 15360
rect 49424 15351 49476 15360
rect 49424 15317 49433 15351
rect 49433 15317 49467 15351
rect 49467 15317 49476 15351
rect 49424 15308 49476 15317
rect 50344 15351 50396 15360
rect 50344 15317 50353 15351
rect 50353 15317 50387 15351
rect 50387 15317 50396 15351
rect 50344 15308 50396 15317
rect 52276 15308 52328 15360
rect 55680 15351 55732 15360
rect 55680 15317 55689 15351
rect 55689 15317 55723 15351
rect 55723 15317 55732 15351
rect 55680 15308 55732 15317
rect 57980 15308 58032 15360
rect 11378 15206 11430 15258
rect 11442 15206 11494 15258
rect 11506 15206 11558 15258
rect 11570 15206 11622 15258
rect 32170 15206 32222 15258
rect 32234 15206 32286 15258
rect 32298 15206 32350 15258
rect 32362 15206 32414 15258
rect 52962 15206 53014 15258
rect 53026 15206 53078 15258
rect 53090 15206 53142 15258
rect 53154 15206 53206 15258
rect 5356 15104 5408 15156
rect 5632 15104 5684 15156
rect 6276 15104 6328 15156
rect 7196 15147 7248 15156
rect 7196 15113 7205 15147
rect 7205 15113 7239 15147
rect 7239 15113 7248 15147
rect 7196 15104 7248 15113
rect 2872 15036 2924 15088
rect 8760 15036 8812 15088
rect 4068 14968 4120 15020
rect 5356 14943 5408 14952
rect 5356 14909 5365 14943
rect 5365 14909 5399 14943
rect 5399 14909 5408 14943
rect 5356 14900 5408 14909
rect 5540 14900 5592 14952
rect 5908 14875 5960 14884
rect 5908 14841 5917 14875
rect 5917 14841 5951 14875
rect 5951 14841 5960 14875
rect 5908 14832 5960 14841
rect 5448 14764 5500 14816
rect 7104 14764 7156 14816
rect 7748 14968 7800 15020
rect 7288 14943 7340 14952
rect 7288 14909 7297 14943
rect 7297 14909 7331 14943
rect 7331 14909 7340 14943
rect 7288 14900 7340 14909
rect 7656 14900 7708 14952
rect 8024 14900 8076 14952
rect 14096 15079 14148 15088
rect 14096 15045 14105 15079
rect 14105 15045 14139 15079
rect 14139 15045 14148 15079
rect 14096 15036 14148 15045
rect 15568 15079 15620 15088
rect 15568 15045 15577 15079
rect 15577 15045 15611 15079
rect 15611 15045 15620 15079
rect 15568 15036 15620 15045
rect 17040 15036 17092 15088
rect 10416 14943 10468 14952
rect 10416 14909 10425 14943
rect 10425 14909 10459 14943
rect 10459 14909 10468 14943
rect 10416 14900 10468 14909
rect 10508 14900 10560 14952
rect 8300 14832 8352 14884
rect 11152 14900 11204 14952
rect 11520 14832 11572 14884
rect 12164 14832 12216 14884
rect 12624 14900 12676 14952
rect 13268 14943 13320 14952
rect 13268 14909 13277 14943
rect 13277 14909 13311 14943
rect 13311 14909 13320 14943
rect 13268 14900 13320 14909
rect 13452 14900 13504 14952
rect 14188 14968 14240 15020
rect 15200 15011 15252 15020
rect 15200 14977 15209 15011
rect 15209 14977 15243 15011
rect 15243 14977 15252 15011
rect 15200 14968 15252 14977
rect 14280 14943 14332 14952
rect 14280 14909 14289 14943
rect 14289 14909 14323 14943
rect 14323 14909 14332 14943
rect 14280 14900 14332 14909
rect 16028 14900 16080 14952
rect 18144 15036 18196 15088
rect 20812 15036 20864 15088
rect 20996 15079 21048 15088
rect 20996 15045 21005 15079
rect 21005 15045 21039 15079
rect 21039 15045 21048 15079
rect 20996 15036 21048 15045
rect 21088 15036 21140 15088
rect 22008 15036 22060 15088
rect 22468 15104 22520 15156
rect 28264 15147 28316 15156
rect 23112 15079 23164 15088
rect 23112 15045 23121 15079
rect 23121 15045 23155 15079
rect 23155 15045 23164 15079
rect 23112 15036 23164 15045
rect 23296 15036 23348 15088
rect 27068 15079 27120 15088
rect 27068 15045 27077 15079
rect 27077 15045 27111 15079
rect 27111 15045 27120 15079
rect 27068 15036 27120 15045
rect 27436 15036 27488 15088
rect 28264 15113 28273 15147
rect 28273 15113 28307 15147
rect 28307 15113 28316 15147
rect 28264 15104 28316 15113
rect 29000 15147 29052 15156
rect 29000 15113 29009 15147
rect 29009 15113 29043 15147
rect 29043 15113 29052 15147
rect 29000 15104 29052 15113
rect 29276 15147 29328 15156
rect 29276 15113 29285 15147
rect 29285 15113 29319 15147
rect 29319 15113 29328 15147
rect 29276 15104 29328 15113
rect 29552 15104 29604 15156
rect 30104 15104 30156 15156
rect 31300 15147 31352 15156
rect 31300 15113 31309 15147
rect 31309 15113 31343 15147
rect 31343 15113 31352 15147
rect 31300 15104 31352 15113
rect 31760 15147 31812 15156
rect 31760 15113 31769 15147
rect 31769 15113 31803 15147
rect 31803 15113 31812 15147
rect 32036 15147 32088 15156
rect 31760 15104 31812 15113
rect 32036 15113 32045 15147
rect 32045 15113 32079 15147
rect 32079 15113 32088 15147
rect 32864 15147 32916 15156
rect 32036 15104 32088 15113
rect 32864 15113 32873 15147
rect 32873 15113 32907 15147
rect 32907 15113 32916 15147
rect 32864 15104 32916 15113
rect 32404 15036 32456 15088
rect 32680 15036 32732 15088
rect 20352 14968 20404 15020
rect 20536 15011 20588 15020
rect 20536 14977 20545 15011
rect 20545 14977 20579 15011
rect 20579 14977 20588 15011
rect 22376 15011 22428 15020
rect 20536 14968 20588 14977
rect 22376 14977 22385 15011
rect 22385 14977 22419 15011
rect 22419 14977 22428 15011
rect 22376 14968 22428 14977
rect 22560 14968 22612 15020
rect 25044 15011 25096 15020
rect 25044 14977 25053 15011
rect 25053 14977 25087 15011
rect 25087 14977 25096 15011
rect 25044 14968 25096 14977
rect 25228 14968 25280 15020
rect 17868 14900 17920 14952
rect 18328 14943 18380 14952
rect 18328 14909 18337 14943
rect 18337 14909 18371 14943
rect 18371 14909 18380 14943
rect 18328 14900 18380 14909
rect 19984 14900 20036 14952
rect 20444 14943 20496 14952
rect 18880 14832 18932 14884
rect 20444 14909 20453 14943
rect 20453 14909 20487 14943
rect 20487 14909 20496 14943
rect 20444 14900 20496 14909
rect 21916 14943 21968 14952
rect 21916 14909 21925 14943
rect 21925 14909 21959 14943
rect 21959 14909 21968 14943
rect 21916 14900 21968 14909
rect 23112 14900 23164 14952
rect 23664 14943 23716 14952
rect 23664 14909 23673 14943
rect 23673 14909 23707 14943
rect 23707 14909 23716 14943
rect 23664 14900 23716 14909
rect 23940 14943 23992 14952
rect 23940 14909 23949 14943
rect 23949 14909 23983 14943
rect 23983 14909 23992 14943
rect 23940 14900 23992 14909
rect 20996 14832 21048 14884
rect 23848 14875 23900 14884
rect 23848 14841 23857 14875
rect 23857 14841 23891 14875
rect 23891 14841 23900 14875
rect 23848 14832 23900 14841
rect 24676 14875 24728 14884
rect 24676 14841 24685 14875
rect 24685 14841 24719 14875
rect 24719 14841 24728 14875
rect 24676 14832 24728 14841
rect 25136 14832 25188 14884
rect 26056 14900 26108 14952
rect 27344 14900 27396 14952
rect 27804 14943 27856 14952
rect 27804 14909 27810 14943
rect 27810 14909 27856 14943
rect 27804 14900 27856 14909
rect 28172 14968 28224 15020
rect 29184 14968 29236 15020
rect 30380 14968 30432 15020
rect 34244 15104 34296 15156
rect 38660 15104 38712 15156
rect 39212 15104 39264 15156
rect 39856 15147 39908 15156
rect 39856 15113 39865 15147
rect 39865 15113 39899 15147
rect 39899 15113 39908 15147
rect 39856 15104 39908 15113
rect 35348 15036 35400 15088
rect 35716 15079 35768 15088
rect 35716 15045 35725 15079
rect 35725 15045 35759 15079
rect 35759 15045 35768 15079
rect 35716 15036 35768 15045
rect 36084 15036 36136 15088
rect 41788 15104 41840 15156
rect 42064 15104 42116 15156
rect 42432 15104 42484 15156
rect 47124 15104 47176 15156
rect 51356 15147 51408 15156
rect 51356 15113 51365 15147
rect 51365 15113 51399 15147
rect 51399 15113 51408 15147
rect 51356 15104 51408 15113
rect 51724 15104 51776 15156
rect 53288 15104 53340 15156
rect 56876 15147 56928 15156
rect 56876 15113 56885 15147
rect 56885 15113 56919 15147
rect 56919 15113 56928 15147
rect 56876 15104 56928 15113
rect 58900 15147 58952 15156
rect 58900 15113 58909 15147
rect 58909 15113 58943 15147
rect 58943 15113 58952 15147
rect 58900 15104 58952 15113
rect 43076 15036 43128 15088
rect 47308 15036 47360 15088
rect 49148 15036 49200 15088
rect 50988 15036 51040 15088
rect 53472 15036 53524 15088
rect 29552 14943 29604 14952
rect 29552 14909 29561 14943
rect 29561 14909 29595 14943
rect 29595 14909 29604 14943
rect 29552 14900 29604 14909
rect 29828 14900 29880 14952
rect 32680 14900 32732 14952
rect 33692 14968 33744 15020
rect 36452 14968 36504 15020
rect 36544 14968 36596 15020
rect 38660 14968 38712 15020
rect 26424 14875 26476 14884
rect 26424 14841 26433 14875
rect 26433 14841 26467 14875
rect 26467 14841 26476 14875
rect 26424 14832 26476 14841
rect 27896 14832 27948 14884
rect 30104 14832 30156 14884
rect 11244 14764 11296 14816
rect 12900 14764 12952 14816
rect 16028 14807 16080 14816
rect 16028 14773 16037 14807
rect 16037 14773 16071 14807
rect 16071 14773 16080 14807
rect 16028 14764 16080 14773
rect 16856 14764 16908 14816
rect 17868 14807 17920 14816
rect 17868 14773 17877 14807
rect 17877 14773 17911 14807
rect 17911 14773 17920 14807
rect 17868 14764 17920 14773
rect 19524 14807 19576 14816
rect 19524 14773 19533 14807
rect 19533 14773 19567 14807
rect 19567 14773 19576 14807
rect 19524 14764 19576 14773
rect 20168 14764 20220 14816
rect 22376 14764 22428 14816
rect 33784 14943 33836 14952
rect 33784 14909 33793 14943
rect 33793 14909 33827 14943
rect 33827 14909 33836 14943
rect 33784 14900 33836 14909
rect 30288 14764 30340 14816
rect 34152 14832 34204 14884
rect 34336 14764 34388 14816
rect 35164 14900 35216 14952
rect 35440 14943 35492 14952
rect 35440 14909 35449 14943
rect 35449 14909 35483 14943
rect 35483 14909 35492 14943
rect 35440 14900 35492 14909
rect 35624 14832 35676 14884
rect 37832 14900 37884 14952
rect 37924 14900 37976 14952
rect 41052 14968 41104 15020
rect 42064 14968 42116 15020
rect 43444 14968 43496 15020
rect 43628 15011 43680 15020
rect 43628 14977 43637 15011
rect 43637 14977 43671 15011
rect 43671 14977 43680 15011
rect 43628 14968 43680 14977
rect 51632 14968 51684 15020
rect 52368 15011 52420 15020
rect 52368 14977 52377 15011
rect 52377 14977 52411 15011
rect 52411 14977 52420 15011
rect 52368 14968 52420 14977
rect 53748 14968 53800 15020
rect 37188 14832 37240 14884
rect 36452 14764 36504 14816
rect 38384 14832 38436 14884
rect 37740 14807 37792 14816
rect 37740 14773 37749 14807
rect 37749 14773 37783 14807
rect 37783 14773 37792 14807
rect 37740 14764 37792 14773
rect 40132 14832 40184 14884
rect 41604 14900 41656 14952
rect 41880 14943 41932 14952
rect 41880 14909 41889 14943
rect 41889 14909 41923 14943
rect 41923 14909 41932 14943
rect 41880 14900 41932 14909
rect 42340 14900 42392 14952
rect 42892 14943 42944 14952
rect 42892 14909 42901 14943
rect 42901 14909 42935 14943
rect 42935 14909 42944 14943
rect 42892 14900 42944 14909
rect 43076 14943 43128 14952
rect 43076 14909 43085 14943
rect 43085 14909 43119 14943
rect 43119 14909 43128 14943
rect 43076 14900 43128 14909
rect 43168 14943 43220 14952
rect 43168 14909 43177 14943
rect 43177 14909 43211 14943
rect 43211 14909 43220 14943
rect 43168 14900 43220 14909
rect 43904 14900 43956 14952
rect 48136 14943 48188 14952
rect 41144 14832 41196 14884
rect 41236 14832 41288 14884
rect 46204 14832 46256 14884
rect 46848 14832 46900 14884
rect 40592 14764 40644 14816
rect 40684 14807 40736 14816
rect 40684 14773 40693 14807
rect 40693 14773 40727 14807
rect 40727 14773 40736 14807
rect 40684 14764 40736 14773
rect 41788 14764 41840 14816
rect 45192 14764 45244 14816
rect 48136 14909 48145 14943
rect 48145 14909 48179 14943
rect 48179 14909 48188 14943
rect 48136 14900 48188 14909
rect 48228 14900 48280 14952
rect 48780 14900 48832 14952
rect 49792 14943 49844 14952
rect 49792 14909 49801 14943
rect 49801 14909 49835 14943
rect 49835 14909 49844 14943
rect 49792 14900 49844 14909
rect 50344 14900 50396 14952
rect 52276 14900 52328 14952
rect 52828 14900 52880 14952
rect 53840 14900 53892 14952
rect 48964 14764 49016 14816
rect 52736 14832 52788 14884
rect 63592 14968 63644 15020
rect 55680 14943 55732 14952
rect 55680 14909 55689 14943
rect 55689 14909 55723 14943
rect 55723 14909 55732 14943
rect 55680 14900 55732 14909
rect 55864 14943 55916 14952
rect 55864 14909 55873 14943
rect 55873 14909 55907 14943
rect 55907 14909 55916 14943
rect 55864 14900 55916 14909
rect 56232 14900 56284 14952
rect 57244 14900 57296 14952
rect 57980 14900 58032 14952
rect 58716 14900 58768 14952
rect 56416 14875 56468 14884
rect 56416 14841 56425 14875
rect 56425 14841 56459 14875
rect 56459 14841 56468 14875
rect 56416 14832 56468 14841
rect 55496 14764 55548 14816
rect 21774 14662 21826 14714
rect 21838 14662 21890 14714
rect 21902 14662 21954 14714
rect 21966 14662 22018 14714
rect 42566 14662 42618 14714
rect 42630 14662 42682 14714
rect 42694 14662 42746 14714
rect 42758 14662 42810 14714
rect 4896 14560 4948 14612
rect 10784 14560 10836 14612
rect 18880 14603 18932 14612
rect 7472 14492 7524 14544
rect 7932 14492 7984 14544
rect 6000 14467 6052 14476
rect 6000 14433 6009 14467
rect 6009 14433 6043 14467
rect 6043 14433 6052 14467
rect 6000 14424 6052 14433
rect 7840 14467 7892 14476
rect 7840 14433 7849 14467
rect 7849 14433 7883 14467
rect 7883 14433 7892 14467
rect 7840 14424 7892 14433
rect 8116 14424 8168 14476
rect 14096 14492 14148 14544
rect 18880 14569 18889 14603
rect 18889 14569 18923 14603
rect 18923 14569 18932 14603
rect 18880 14560 18932 14569
rect 20536 14603 20588 14612
rect 20536 14569 20545 14603
rect 20545 14569 20579 14603
rect 20579 14569 20588 14603
rect 20536 14560 20588 14569
rect 20720 14492 20772 14544
rect 21640 14492 21692 14544
rect 23848 14535 23900 14544
rect 23848 14501 23857 14535
rect 23857 14501 23891 14535
rect 23891 14501 23900 14535
rect 23848 14492 23900 14501
rect 26424 14492 26476 14544
rect 28264 14492 28316 14544
rect 29368 14535 29420 14544
rect 29368 14501 29377 14535
rect 29377 14501 29411 14535
rect 29411 14501 29420 14535
rect 29368 14492 29420 14501
rect 9680 14467 9732 14476
rect 9680 14433 9689 14467
rect 9689 14433 9723 14467
rect 9723 14433 9732 14467
rect 9680 14424 9732 14433
rect 9864 14467 9916 14476
rect 9864 14433 9873 14467
rect 9873 14433 9907 14467
rect 9907 14433 9916 14467
rect 9864 14424 9916 14433
rect 10416 14424 10468 14476
rect 13452 14467 13504 14476
rect 13452 14433 13461 14467
rect 13461 14433 13495 14467
rect 13495 14433 13504 14467
rect 13452 14424 13504 14433
rect 14280 14424 14332 14476
rect 15936 14424 15988 14476
rect 16028 14424 16080 14476
rect 8944 14356 8996 14408
rect 10324 14356 10376 14408
rect 11520 14399 11572 14408
rect 11520 14365 11529 14399
rect 11529 14365 11563 14399
rect 11563 14365 11572 14399
rect 11520 14356 11572 14365
rect 12440 14356 12492 14408
rect 16856 14399 16908 14408
rect 16856 14365 16865 14399
rect 16865 14365 16899 14399
rect 16899 14365 16908 14399
rect 16856 14356 16908 14365
rect 17132 14399 17184 14408
rect 17132 14365 17141 14399
rect 17141 14365 17175 14399
rect 17175 14365 17184 14399
rect 17132 14356 17184 14365
rect 19892 14424 19944 14476
rect 24860 14467 24912 14476
rect 24860 14433 24869 14467
rect 24869 14433 24903 14467
rect 24903 14433 24912 14467
rect 24860 14424 24912 14433
rect 25136 14467 25188 14476
rect 25136 14433 25145 14467
rect 25145 14433 25179 14467
rect 25179 14433 25188 14467
rect 25136 14424 25188 14433
rect 25780 14424 25832 14476
rect 27160 14467 27212 14476
rect 27160 14433 27169 14467
rect 27169 14433 27203 14467
rect 27203 14433 27212 14467
rect 27160 14424 27212 14433
rect 29552 14424 29604 14476
rect 30196 14467 30248 14476
rect 30196 14433 30205 14467
rect 30205 14433 30239 14467
rect 30239 14433 30248 14467
rect 30196 14424 30248 14433
rect 30380 14560 30432 14612
rect 32312 14560 32364 14612
rect 32496 14560 32548 14612
rect 34152 14603 34204 14612
rect 31760 14492 31812 14544
rect 34152 14569 34161 14603
rect 34161 14569 34195 14603
rect 34195 14569 34204 14603
rect 34152 14560 34204 14569
rect 34336 14560 34388 14612
rect 34704 14560 34756 14612
rect 37188 14560 37240 14612
rect 40316 14560 40368 14612
rect 42248 14560 42300 14612
rect 32496 14424 32548 14476
rect 33324 14424 33376 14476
rect 34152 14424 34204 14476
rect 21548 14356 21600 14408
rect 21640 14356 21692 14408
rect 22560 14356 22612 14408
rect 25044 14399 25096 14408
rect 25044 14365 25053 14399
rect 25053 14365 25087 14399
rect 25087 14365 25096 14399
rect 25044 14356 25096 14365
rect 27528 14356 27580 14408
rect 27988 14356 28040 14408
rect 28172 14356 28224 14408
rect 28356 14356 28408 14408
rect 30104 14356 30156 14408
rect 5356 14288 5408 14340
rect 11152 14288 11204 14340
rect 5724 14220 5776 14272
rect 6276 14263 6328 14272
rect 6276 14229 6285 14263
rect 6285 14229 6319 14263
rect 6319 14229 6328 14263
rect 6276 14220 6328 14229
rect 7104 14220 7156 14272
rect 9496 14220 9548 14272
rect 16396 14288 16448 14340
rect 29276 14288 29328 14340
rect 31208 14356 31260 14408
rect 32772 14399 32824 14408
rect 32772 14365 32781 14399
rect 32781 14365 32815 14399
rect 32815 14365 32824 14399
rect 32772 14356 32824 14365
rect 33048 14399 33100 14408
rect 33048 14365 33057 14399
rect 33057 14365 33091 14399
rect 33091 14365 33100 14399
rect 33048 14356 33100 14365
rect 35348 14492 35400 14544
rect 36360 14492 36412 14544
rect 39028 14492 39080 14544
rect 39856 14492 39908 14544
rect 36268 14424 36320 14476
rect 37924 14467 37976 14476
rect 37924 14433 37933 14467
rect 37933 14433 37967 14467
rect 37967 14433 37976 14467
rect 37924 14424 37976 14433
rect 38200 14467 38252 14476
rect 38200 14433 38209 14467
rect 38209 14433 38243 14467
rect 38243 14433 38252 14467
rect 38200 14424 38252 14433
rect 38384 14424 38436 14476
rect 36084 14356 36136 14408
rect 14004 14220 14056 14272
rect 14740 14263 14792 14272
rect 14740 14229 14749 14263
rect 14749 14229 14783 14263
rect 14783 14229 14792 14263
rect 14740 14220 14792 14229
rect 14832 14220 14884 14272
rect 15936 14263 15988 14272
rect 15936 14229 15945 14263
rect 15945 14229 15979 14263
rect 15979 14229 15988 14263
rect 15936 14220 15988 14229
rect 16580 14220 16632 14272
rect 16764 14263 16816 14272
rect 16764 14229 16773 14263
rect 16773 14229 16807 14263
rect 16807 14229 16816 14263
rect 16764 14220 16816 14229
rect 18328 14220 18380 14272
rect 19984 14220 20036 14272
rect 20720 14220 20772 14272
rect 21364 14220 21416 14272
rect 23388 14263 23440 14272
rect 23388 14229 23397 14263
rect 23397 14229 23431 14263
rect 23431 14229 23440 14263
rect 23388 14220 23440 14229
rect 23572 14220 23624 14272
rect 23940 14220 23992 14272
rect 25780 14220 25832 14272
rect 26240 14263 26292 14272
rect 26240 14229 26249 14263
rect 26249 14229 26283 14263
rect 26283 14229 26292 14263
rect 26240 14220 26292 14229
rect 26792 14263 26844 14272
rect 26792 14229 26801 14263
rect 26801 14229 26835 14263
rect 26835 14229 26844 14263
rect 26792 14220 26844 14229
rect 27344 14220 27396 14272
rect 28816 14263 28868 14272
rect 28816 14229 28825 14263
rect 28825 14229 28859 14263
rect 28859 14229 28868 14263
rect 28816 14220 28868 14229
rect 28908 14220 28960 14272
rect 34796 14331 34848 14340
rect 30380 14263 30432 14272
rect 30380 14229 30404 14263
rect 30404 14229 30432 14263
rect 30380 14220 30432 14229
rect 30472 14263 30524 14272
rect 30472 14229 30481 14263
rect 30481 14229 30515 14263
rect 30515 14229 30524 14263
rect 31944 14263 31996 14272
rect 30472 14220 30524 14229
rect 31944 14229 31953 14263
rect 31953 14229 31987 14263
rect 31987 14229 31996 14263
rect 31944 14220 31996 14229
rect 34796 14297 34805 14331
rect 34805 14297 34839 14331
rect 34839 14297 34848 14331
rect 34796 14288 34848 14297
rect 39028 14288 39080 14340
rect 40040 14424 40092 14476
rect 40776 14492 40828 14544
rect 41604 14492 41656 14544
rect 41696 14492 41748 14544
rect 39304 14399 39356 14408
rect 39304 14365 39313 14399
rect 39313 14365 39347 14399
rect 39347 14365 39356 14399
rect 39304 14356 39356 14365
rect 39488 14399 39540 14408
rect 39488 14365 39497 14399
rect 39497 14365 39531 14399
rect 39531 14365 39540 14399
rect 39488 14356 39540 14365
rect 40592 14424 40644 14476
rect 42064 14492 42116 14544
rect 42156 14492 42208 14544
rect 40408 14356 40460 14408
rect 41972 14424 42024 14476
rect 47492 14560 47544 14612
rect 52736 14560 52788 14612
rect 52828 14560 52880 14612
rect 55772 14560 55824 14612
rect 57704 14560 57756 14612
rect 43444 14424 43496 14476
rect 47400 14424 47452 14476
rect 48228 14424 48280 14476
rect 48964 14467 49016 14476
rect 48964 14433 48973 14467
rect 48973 14433 49007 14467
rect 49007 14433 49016 14467
rect 48964 14424 49016 14433
rect 49148 14492 49200 14544
rect 52276 14492 52328 14544
rect 52368 14492 52420 14544
rect 52644 14467 52696 14476
rect 52644 14433 52653 14467
rect 52653 14433 52687 14467
rect 52687 14433 52696 14467
rect 52644 14424 52696 14433
rect 56784 14492 56836 14544
rect 55864 14424 55916 14476
rect 56416 14424 56468 14476
rect 41236 14288 41288 14340
rect 42984 14356 43036 14408
rect 45836 14399 45888 14408
rect 45836 14365 45845 14399
rect 45845 14365 45879 14399
rect 45879 14365 45888 14399
rect 45836 14356 45888 14365
rect 46756 14356 46808 14408
rect 47768 14356 47820 14408
rect 41788 14288 41840 14340
rect 42892 14288 42944 14340
rect 43628 14288 43680 14340
rect 47400 14288 47452 14340
rect 48044 14288 48096 14340
rect 50528 14356 50580 14408
rect 50620 14356 50672 14408
rect 51356 14356 51408 14408
rect 53380 14356 53432 14408
rect 53748 14356 53800 14408
rect 55220 14356 55272 14408
rect 55496 14356 55548 14408
rect 56968 14356 57020 14408
rect 32956 14220 33008 14272
rect 34888 14220 34940 14272
rect 35716 14263 35768 14272
rect 35716 14229 35725 14263
rect 35725 14229 35759 14263
rect 35759 14229 35768 14263
rect 35716 14220 35768 14229
rect 36268 14263 36320 14272
rect 36268 14229 36277 14263
rect 36277 14229 36311 14263
rect 36311 14229 36320 14263
rect 36268 14220 36320 14229
rect 36728 14263 36780 14272
rect 36728 14229 36737 14263
rect 36737 14229 36771 14263
rect 36771 14229 36780 14263
rect 36728 14220 36780 14229
rect 37004 14263 37056 14272
rect 37004 14229 37013 14263
rect 37013 14229 37047 14263
rect 37047 14229 37056 14263
rect 37004 14220 37056 14229
rect 38108 14220 38160 14272
rect 41420 14263 41472 14272
rect 41420 14229 41429 14263
rect 41429 14229 41463 14263
rect 41463 14229 41472 14263
rect 41420 14220 41472 14229
rect 43536 14263 43588 14272
rect 43536 14229 43545 14263
rect 43545 14229 43579 14263
rect 43579 14229 43588 14263
rect 43536 14220 43588 14229
rect 43812 14220 43864 14272
rect 48320 14220 48372 14272
rect 49148 14263 49200 14272
rect 49148 14229 49157 14263
rect 49157 14229 49191 14263
rect 49191 14229 49200 14263
rect 49148 14220 49200 14229
rect 49608 14220 49660 14272
rect 57244 14356 57296 14408
rect 50620 14220 50672 14272
rect 52828 14263 52880 14272
rect 52828 14229 52837 14263
rect 52837 14229 52871 14263
rect 52871 14229 52880 14263
rect 52828 14220 52880 14229
rect 53840 14220 53892 14272
rect 54576 14220 54628 14272
rect 55588 14220 55640 14272
rect 56784 14220 56836 14272
rect 56968 14220 57020 14272
rect 11378 14118 11430 14170
rect 11442 14118 11494 14170
rect 11506 14118 11558 14170
rect 11570 14118 11622 14170
rect 32170 14118 32222 14170
rect 32234 14118 32286 14170
rect 32298 14118 32350 14170
rect 32362 14118 32414 14170
rect 52962 14118 53014 14170
rect 53026 14118 53078 14170
rect 53090 14118 53142 14170
rect 53154 14118 53206 14170
rect 4896 14059 4948 14068
rect 4896 14025 4905 14059
rect 4905 14025 4939 14059
rect 4939 14025 4948 14059
rect 4896 14016 4948 14025
rect 6000 14016 6052 14068
rect 7472 14059 7524 14068
rect 7472 14025 7481 14059
rect 7481 14025 7515 14059
rect 7515 14025 7524 14059
rect 7472 14016 7524 14025
rect 8024 14059 8076 14068
rect 8024 14025 8033 14059
rect 8033 14025 8067 14059
rect 8067 14025 8076 14059
rect 8024 14016 8076 14025
rect 8116 14016 8168 14068
rect 8944 14059 8996 14068
rect 8944 14025 8953 14059
rect 8953 14025 8987 14059
rect 8987 14025 8996 14059
rect 8944 14016 8996 14025
rect 10784 14059 10836 14068
rect 10784 14025 10793 14059
rect 10793 14025 10827 14059
rect 10827 14025 10836 14059
rect 10784 14016 10836 14025
rect 11244 14059 11296 14068
rect 11244 14025 11253 14059
rect 11253 14025 11287 14059
rect 11287 14025 11296 14059
rect 11244 14016 11296 14025
rect 14372 14016 14424 14068
rect 14740 14016 14792 14068
rect 15292 14016 15344 14068
rect 16396 14059 16448 14068
rect 16396 14025 16405 14059
rect 16405 14025 16439 14059
rect 16439 14025 16448 14059
rect 16396 14016 16448 14025
rect 3148 13948 3200 14000
rect 4896 13880 4948 13932
rect 4160 13855 4212 13864
rect 4160 13821 4169 13855
rect 4169 13821 4203 13855
rect 4203 13821 4212 13855
rect 4528 13855 4580 13864
rect 4160 13812 4212 13821
rect 4528 13821 4537 13855
rect 4537 13821 4571 13855
rect 4571 13821 4580 13855
rect 4528 13812 4580 13821
rect 5632 13880 5684 13932
rect 8760 13880 8812 13932
rect 9956 13880 10008 13932
rect 4712 13744 4764 13796
rect 6920 13812 6972 13864
rect 7748 13855 7800 13864
rect 7748 13821 7757 13855
rect 7757 13821 7791 13855
rect 7791 13821 7800 13855
rect 7748 13812 7800 13821
rect 8024 13812 8076 13864
rect 9496 13812 9548 13864
rect 11244 13880 11296 13932
rect 9588 13744 9640 13796
rect 11152 13812 11204 13864
rect 11704 13744 11756 13796
rect 12440 13812 12492 13864
rect 13268 13880 13320 13932
rect 14280 13948 14332 14000
rect 13452 13880 13504 13932
rect 13912 13880 13964 13932
rect 14188 13880 14240 13932
rect 14924 13948 14976 14000
rect 14740 13923 14792 13932
rect 14740 13889 14749 13923
rect 14749 13889 14783 13923
rect 14783 13889 14792 13923
rect 14740 13880 14792 13889
rect 13820 13812 13872 13864
rect 17684 13948 17736 14000
rect 15936 13880 15988 13932
rect 17040 13880 17092 13932
rect 17132 13880 17184 13932
rect 21088 14016 21140 14068
rect 21180 14016 21232 14068
rect 22376 14016 22428 14068
rect 22560 14059 22612 14068
rect 22560 14025 22569 14059
rect 22569 14025 22603 14059
rect 22603 14025 22612 14059
rect 22560 14016 22612 14025
rect 24124 14016 24176 14068
rect 26056 14016 26108 14068
rect 18696 13948 18748 14000
rect 21824 13948 21876 14000
rect 22100 13948 22152 14000
rect 24492 13948 24544 14000
rect 25228 13948 25280 14000
rect 23296 13923 23348 13932
rect 23296 13889 23305 13923
rect 23305 13889 23339 13923
rect 23339 13889 23348 13923
rect 23296 13880 23348 13889
rect 24860 13923 24912 13932
rect 24860 13889 24869 13923
rect 24869 13889 24903 13923
rect 24903 13889 24912 13923
rect 24860 13880 24912 13889
rect 5724 13676 5776 13728
rect 9312 13676 9364 13728
rect 9956 13676 10008 13728
rect 10600 13676 10652 13728
rect 13636 13744 13688 13796
rect 14740 13744 14792 13796
rect 15568 13812 15620 13864
rect 16212 13855 16264 13864
rect 16212 13821 16221 13855
rect 16221 13821 16255 13855
rect 16255 13821 16264 13855
rect 16212 13812 16264 13821
rect 16764 13812 16816 13864
rect 18236 13812 18288 13864
rect 18604 13812 18656 13864
rect 18696 13855 18748 13864
rect 18696 13821 18705 13855
rect 18705 13821 18739 13855
rect 18739 13821 18748 13855
rect 18696 13812 18748 13821
rect 19892 13855 19944 13864
rect 19892 13821 19901 13855
rect 19901 13821 19935 13855
rect 19935 13821 19944 13855
rect 19892 13812 19944 13821
rect 20720 13855 20772 13864
rect 20720 13821 20729 13855
rect 20729 13821 20763 13855
rect 20763 13821 20772 13855
rect 20720 13812 20772 13821
rect 20996 13812 21048 13864
rect 20444 13744 20496 13796
rect 21640 13812 21692 13864
rect 21824 13812 21876 13864
rect 22100 13855 22152 13864
rect 22100 13821 22109 13855
rect 22109 13821 22143 13855
rect 22143 13821 22152 13855
rect 22100 13812 22152 13821
rect 23480 13812 23532 13864
rect 26240 13923 26292 13932
rect 26240 13889 26249 13923
rect 26249 13889 26283 13923
rect 26283 13889 26292 13923
rect 26240 13880 26292 13889
rect 22192 13744 22244 13796
rect 22928 13787 22980 13796
rect 22928 13753 22937 13787
rect 22937 13753 22971 13787
rect 22971 13753 22980 13787
rect 22928 13744 22980 13753
rect 23020 13744 23072 13796
rect 25136 13744 25188 13796
rect 27988 14016 28040 14068
rect 28080 14059 28132 14068
rect 28080 14025 28089 14059
rect 28089 14025 28123 14059
rect 28123 14025 28132 14059
rect 28080 14016 28132 14025
rect 28264 14016 28316 14068
rect 30380 14016 30432 14068
rect 33048 14016 33100 14068
rect 35716 14016 35768 14068
rect 36084 14016 36136 14068
rect 36360 14059 36412 14068
rect 36360 14025 36369 14059
rect 36369 14025 36403 14059
rect 36403 14025 36412 14059
rect 36360 14016 36412 14025
rect 38200 14016 38252 14068
rect 27436 13948 27488 14000
rect 28816 13948 28868 14000
rect 35348 13948 35400 14000
rect 35440 13948 35492 14000
rect 37924 13948 37976 14000
rect 38292 13991 38344 14000
rect 38292 13957 38301 13991
rect 38301 13957 38335 13991
rect 38335 13957 38344 13991
rect 38292 13948 38344 13957
rect 41788 14016 41840 14068
rect 42064 14016 42116 14068
rect 42524 14016 42576 14068
rect 43168 14016 43220 14068
rect 43536 14016 43588 14068
rect 43996 14059 44048 14068
rect 43996 14025 44005 14059
rect 44005 14025 44039 14059
rect 44039 14025 44048 14059
rect 43996 14016 44048 14025
rect 45836 14059 45888 14068
rect 45836 14025 45845 14059
rect 45845 14025 45879 14059
rect 45879 14025 45888 14059
rect 45836 14016 45888 14025
rect 47492 14059 47544 14068
rect 27344 13880 27396 13932
rect 28172 13880 28224 13932
rect 28908 13880 28960 13932
rect 26240 13744 26292 13796
rect 27528 13812 27580 13864
rect 28540 13812 28592 13864
rect 29828 13880 29880 13932
rect 30196 13880 30248 13932
rect 31944 13880 31996 13932
rect 35716 13880 35768 13932
rect 37464 13923 37516 13932
rect 37464 13889 37473 13923
rect 37473 13889 37507 13923
rect 37507 13889 37516 13923
rect 37464 13880 37516 13889
rect 29736 13812 29788 13864
rect 30104 13812 30156 13864
rect 33048 13855 33100 13864
rect 31208 13787 31260 13796
rect 31208 13753 31217 13787
rect 31217 13753 31251 13787
rect 31251 13753 31260 13787
rect 31208 13744 31260 13753
rect 32128 13787 32180 13796
rect 32128 13753 32137 13787
rect 32137 13753 32171 13787
rect 32171 13753 32180 13787
rect 33048 13821 33057 13855
rect 33057 13821 33091 13855
rect 33091 13821 33100 13855
rect 33048 13812 33100 13821
rect 33140 13812 33192 13864
rect 33876 13855 33928 13864
rect 33876 13821 33885 13855
rect 33885 13821 33919 13855
rect 33919 13821 33928 13855
rect 33876 13812 33928 13821
rect 34152 13812 34204 13864
rect 32128 13744 32180 13753
rect 34888 13787 34940 13796
rect 17408 13676 17460 13728
rect 17868 13719 17920 13728
rect 17868 13685 17877 13719
rect 17877 13685 17911 13719
rect 17911 13685 17920 13719
rect 17868 13676 17920 13685
rect 19524 13676 19576 13728
rect 22744 13676 22796 13728
rect 29828 13676 29880 13728
rect 30012 13676 30064 13728
rect 33508 13676 33560 13728
rect 33968 13676 34020 13728
rect 34888 13753 34897 13787
rect 34897 13753 34931 13787
rect 34931 13753 34940 13787
rect 34888 13744 34940 13753
rect 35348 13812 35400 13864
rect 38108 13812 38160 13864
rect 39028 13855 39080 13864
rect 39028 13821 39034 13855
rect 39034 13821 39080 13855
rect 39028 13812 39080 13821
rect 39304 13880 39356 13932
rect 40040 13923 40092 13932
rect 40040 13889 40049 13923
rect 40049 13889 40083 13923
rect 40083 13889 40092 13923
rect 40040 13880 40092 13889
rect 40500 13923 40552 13932
rect 40500 13889 40509 13923
rect 40509 13889 40543 13923
rect 40543 13889 40552 13923
rect 40500 13880 40552 13889
rect 41236 13948 41288 14000
rect 43812 13991 43864 14000
rect 43812 13957 43821 13991
rect 43821 13957 43855 13991
rect 43855 13957 43864 13991
rect 43812 13948 43864 13957
rect 40592 13855 40644 13864
rect 40592 13821 40601 13855
rect 40601 13821 40635 13855
rect 40635 13821 40644 13855
rect 40592 13812 40644 13821
rect 40684 13812 40736 13864
rect 41972 13855 42024 13864
rect 41972 13821 41981 13855
rect 41981 13821 42015 13855
rect 42015 13821 42024 13855
rect 41972 13812 42024 13821
rect 42156 13855 42208 13864
rect 42156 13821 42162 13855
rect 42162 13821 42208 13855
rect 42156 13812 42208 13821
rect 42524 13880 42576 13932
rect 43536 13855 43588 13864
rect 35256 13787 35308 13796
rect 35256 13753 35265 13787
rect 35265 13753 35299 13787
rect 35299 13753 35308 13787
rect 38844 13787 38896 13796
rect 35256 13744 35308 13753
rect 38844 13753 38853 13787
rect 38853 13753 38887 13787
rect 38887 13753 38896 13787
rect 38844 13744 38896 13753
rect 41420 13744 41472 13796
rect 43536 13821 43545 13855
rect 43545 13821 43579 13855
rect 43579 13821 43588 13855
rect 43536 13812 43588 13821
rect 43628 13812 43680 13864
rect 43904 13923 43956 13932
rect 43904 13889 43913 13923
rect 43913 13889 43947 13923
rect 43947 13889 43956 13923
rect 43904 13880 43956 13889
rect 47492 14025 47501 14059
rect 47501 14025 47535 14059
rect 47535 14025 47544 14059
rect 47492 14016 47544 14025
rect 48320 14059 48372 14068
rect 48320 14025 48329 14059
rect 48329 14025 48363 14059
rect 48363 14025 48372 14059
rect 48320 14016 48372 14025
rect 48964 14016 49016 14068
rect 49148 14016 49200 14068
rect 46848 13948 46900 14000
rect 51448 14016 51500 14068
rect 52276 14016 52328 14068
rect 55680 14016 55732 14068
rect 55772 14016 55824 14068
rect 56416 14016 56468 14068
rect 53288 13948 53340 14000
rect 53748 13948 53800 14000
rect 55128 13991 55180 14000
rect 48228 13923 48280 13932
rect 48228 13889 48234 13923
rect 48234 13889 48280 13923
rect 48228 13880 48280 13889
rect 48412 13923 48464 13932
rect 48412 13889 48421 13923
rect 48421 13889 48455 13923
rect 48455 13889 48464 13923
rect 48412 13880 48464 13889
rect 43904 13744 43956 13796
rect 45652 13744 45704 13796
rect 46112 13787 46164 13796
rect 46112 13753 46121 13787
rect 46121 13753 46155 13787
rect 46155 13753 46164 13787
rect 46112 13744 46164 13753
rect 46756 13855 46808 13864
rect 46756 13821 46765 13855
rect 46765 13821 46799 13855
rect 46799 13821 46808 13855
rect 46756 13812 46808 13821
rect 46848 13812 46900 13864
rect 50252 13855 50304 13864
rect 50252 13821 50261 13855
rect 50261 13821 50295 13855
rect 50295 13821 50304 13855
rect 50252 13812 50304 13821
rect 52460 13880 52512 13932
rect 55128 13957 55137 13991
rect 55137 13957 55171 13991
rect 55171 13957 55180 13991
rect 55128 13948 55180 13957
rect 55588 13948 55640 14000
rect 58440 13948 58492 14000
rect 58900 14016 58952 14068
rect 50528 13812 50580 13864
rect 52092 13812 52144 13864
rect 52184 13812 52236 13864
rect 52644 13855 52696 13864
rect 52644 13821 52653 13855
rect 52653 13821 52687 13855
rect 52687 13821 52696 13855
rect 52644 13812 52696 13821
rect 52736 13812 52788 13864
rect 55220 13812 55272 13864
rect 55496 13855 55548 13864
rect 55496 13821 55505 13855
rect 55505 13821 55539 13855
rect 55539 13821 55548 13855
rect 55496 13812 55548 13821
rect 55864 13812 55916 13864
rect 56968 13812 57020 13864
rect 47308 13744 47360 13796
rect 35348 13676 35400 13728
rect 35532 13676 35584 13728
rect 39212 13676 39264 13728
rect 39304 13676 39356 13728
rect 43444 13676 43496 13728
rect 45100 13676 45152 13728
rect 45560 13719 45612 13728
rect 45560 13685 45569 13719
rect 45569 13685 45603 13719
rect 45603 13685 45612 13719
rect 45560 13676 45612 13685
rect 46204 13676 46256 13728
rect 52368 13744 52420 13796
rect 58164 13855 58216 13864
rect 58164 13821 58173 13855
rect 58173 13821 58207 13855
rect 58207 13821 58216 13855
rect 58164 13812 58216 13821
rect 57888 13744 57940 13796
rect 50988 13676 51040 13728
rect 51080 13676 51132 13728
rect 52092 13676 52144 13728
rect 21774 13574 21826 13626
rect 21838 13574 21890 13626
rect 21902 13574 21954 13626
rect 21966 13574 22018 13626
rect 42566 13574 42618 13626
rect 42630 13574 42682 13626
rect 42694 13574 42746 13626
rect 42758 13574 42810 13626
rect 4528 13472 4580 13524
rect 5448 13472 5500 13524
rect 5540 13404 5592 13456
rect 4988 13379 5040 13388
rect 4988 13345 4997 13379
rect 4997 13345 5031 13379
rect 5031 13345 5040 13379
rect 7748 13515 7800 13524
rect 7748 13481 7757 13515
rect 7757 13481 7791 13515
rect 7791 13481 7800 13515
rect 7748 13472 7800 13481
rect 8116 13472 8168 13524
rect 13728 13472 13780 13524
rect 10600 13447 10652 13456
rect 4988 13336 5040 13345
rect 7012 13336 7064 13388
rect 6552 13268 6604 13320
rect 6920 13200 6972 13252
rect 7288 13379 7340 13388
rect 7288 13345 7297 13379
rect 7297 13345 7331 13379
rect 7331 13345 7340 13379
rect 7288 13336 7340 13345
rect 9772 13379 9824 13388
rect 9772 13345 9781 13379
rect 9781 13345 9815 13379
rect 9815 13345 9824 13379
rect 9772 13336 9824 13345
rect 10600 13413 10609 13447
rect 10609 13413 10643 13447
rect 10643 13413 10652 13447
rect 10600 13404 10652 13413
rect 11704 13447 11756 13456
rect 11704 13413 11713 13447
rect 11713 13413 11747 13447
rect 11747 13413 11756 13447
rect 11704 13404 11756 13413
rect 14740 13472 14792 13524
rect 14924 13472 14976 13524
rect 16856 13472 16908 13524
rect 18236 13472 18288 13524
rect 20996 13472 21048 13524
rect 25044 13472 25096 13524
rect 13912 13404 13964 13456
rect 11980 13336 12032 13388
rect 7380 13311 7432 13320
rect 7380 13277 7389 13311
rect 7389 13277 7423 13311
rect 7423 13277 7432 13311
rect 7380 13268 7432 13277
rect 9588 13268 9640 13320
rect 9680 13311 9732 13320
rect 9680 13277 9699 13311
rect 9699 13277 9732 13311
rect 9680 13268 9732 13277
rect 10692 13268 10744 13320
rect 12624 13379 12676 13388
rect 12624 13345 12633 13379
rect 12633 13345 12667 13379
rect 12667 13345 12676 13379
rect 13084 13379 13136 13388
rect 12624 13336 12676 13345
rect 13084 13345 13093 13379
rect 13093 13345 13127 13379
rect 13127 13345 13136 13379
rect 13084 13336 13136 13345
rect 14096 13336 14148 13388
rect 14648 13336 14700 13388
rect 14924 13336 14976 13388
rect 16028 13336 16080 13388
rect 16580 13379 16632 13388
rect 16580 13345 16589 13379
rect 16589 13345 16623 13379
rect 16623 13345 16632 13379
rect 17592 13404 17644 13456
rect 17868 13404 17920 13456
rect 19616 13404 19668 13456
rect 20812 13404 20864 13456
rect 17408 13379 17460 13388
rect 16580 13336 16632 13345
rect 17408 13345 17417 13379
rect 17417 13345 17451 13379
rect 17451 13345 17460 13379
rect 17408 13336 17460 13345
rect 17684 13336 17736 13388
rect 22100 13404 22152 13456
rect 21548 13336 21600 13388
rect 21824 13379 21876 13388
rect 21824 13345 21833 13379
rect 21833 13345 21867 13379
rect 21867 13345 21876 13379
rect 21824 13336 21876 13345
rect 21916 13336 21968 13388
rect 23388 13336 23440 13388
rect 14188 13268 14240 13320
rect 14832 13268 14884 13320
rect 15568 13268 15620 13320
rect 17316 13311 17368 13320
rect 2412 13175 2464 13184
rect 2412 13141 2421 13175
rect 2421 13141 2455 13175
rect 2455 13141 2464 13175
rect 2412 13132 2464 13141
rect 3884 13175 3936 13184
rect 3884 13141 3893 13175
rect 3893 13141 3927 13175
rect 3927 13141 3936 13175
rect 3884 13132 3936 13141
rect 4712 13175 4764 13184
rect 4712 13141 4721 13175
rect 4721 13141 4755 13175
rect 4755 13141 4764 13175
rect 4712 13132 4764 13141
rect 5172 13132 5224 13184
rect 8024 13132 8076 13184
rect 8484 13175 8536 13184
rect 8484 13141 8493 13175
rect 8493 13141 8527 13175
rect 8527 13141 8536 13175
rect 8484 13132 8536 13141
rect 9404 13175 9456 13184
rect 9404 13141 9413 13175
rect 9413 13141 9447 13175
rect 9447 13141 9456 13175
rect 9404 13132 9456 13141
rect 10508 13200 10560 13252
rect 10232 13132 10284 13184
rect 11152 13175 11204 13184
rect 11152 13141 11161 13175
rect 11161 13141 11195 13175
rect 11195 13141 11204 13175
rect 11152 13132 11204 13141
rect 12624 13200 12676 13252
rect 12716 13200 12768 13252
rect 17316 13277 17325 13311
rect 17325 13277 17359 13311
rect 17359 13277 17368 13311
rect 17316 13268 17368 13277
rect 19524 13311 19576 13320
rect 19524 13277 19533 13311
rect 19533 13277 19567 13311
rect 19567 13277 19576 13311
rect 19524 13268 19576 13277
rect 12072 13132 12124 13184
rect 17040 13132 17092 13184
rect 18604 13175 18656 13184
rect 18604 13141 18613 13175
rect 18613 13141 18647 13175
rect 18647 13141 18656 13175
rect 18604 13132 18656 13141
rect 20904 13200 20956 13252
rect 23296 13268 23348 13320
rect 24216 13311 24268 13320
rect 24216 13277 24225 13311
rect 24225 13277 24259 13311
rect 24259 13277 24268 13311
rect 26056 13336 26108 13388
rect 26240 13515 26292 13524
rect 26240 13481 26249 13515
rect 26249 13481 26283 13515
rect 26283 13481 26292 13515
rect 26240 13472 26292 13481
rect 27712 13472 27764 13524
rect 28172 13515 28224 13524
rect 28172 13481 28181 13515
rect 28181 13481 28215 13515
rect 28215 13481 28224 13515
rect 28172 13472 28224 13481
rect 28540 13515 28592 13524
rect 28540 13481 28549 13515
rect 28549 13481 28583 13515
rect 28583 13481 28592 13515
rect 28540 13472 28592 13481
rect 28816 13472 28868 13524
rect 29276 13515 29328 13524
rect 29276 13481 29285 13515
rect 29285 13481 29319 13515
rect 29319 13481 29328 13515
rect 29276 13472 29328 13481
rect 29736 13515 29788 13524
rect 29736 13481 29745 13515
rect 29745 13481 29779 13515
rect 29779 13481 29788 13515
rect 29736 13472 29788 13481
rect 30472 13515 30524 13524
rect 30472 13481 30481 13515
rect 30481 13481 30515 13515
rect 30515 13481 30524 13515
rect 30472 13472 30524 13481
rect 31208 13472 31260 13524
rect 35532 13472 35584 13524
rect 41052 13472 41104 13524
rect 41144 13472 41196 13524
rect 41696 13472 41748 13524
rect 42984 13472 43036 13524
rect 43536 13472 43588 13524
rect 28724 13379 28776 13388
rect 28724 13345 28733 13379
rect 28733 13345 28767 13379
rect 28767 13345 28776 13379
rect 28724 13336 28776 13345
rect 29828 13379 29880 13388
rect 24216 13268 24268 13277
rect 28172 13268 28224 13320
rect 29092 13268 29144 13320
rect 29828 13345 29837 13379
rect 29837 13345 29871 13379
rect 29871 13345 29880 13379
rect 29828 13336 29880 13345
rect 30932 13379 30984 13388
rect 30932 13345 30941 13379
rect 30941 13345 30975 13379
rect 30975 13345 30984 13379
rect 33048 13404 33100 13456
rect 30932 13336 30984 13345
rect 31668 13268 31720 13320
rect 32496 13336 32548 13388
rect 33508 13379 33560 13388
rect 33508 13345 33517 13379
rect 33517 13345 33551 13379
rect 33551 13345 33560 13379
rect 33508 13336 33560 13345
rect 34244 13379 34296 13388
rect 22560 13200 22612 13252
rect 22836 13200 22888 13252
rect 23664 13200 23716 13252
rect 27160 13200 27212 13252
rect 29184 13200 29236 13252
rect 32680 13268 32732 13320
rect 33232 13268 33284 13320
rect 34244 13345 34253 13379
rect 34253 13345 34287 13379
rect 34287 13345 34296 13379
rect 34244 13336 34296 13345
rect 35440 13404 35492 13456
rect 38200 13404 38252 13456
rect 39304 13404 39356 13456
rect 39488 13404 39540 13456
rect 40132 13447 40184 13456
rect 40132 13413 40141 13447
rect 40141 13413 40175 13447
rect 40175 13413 40184 13447
rect 40132 13404 40184 13413
rect 34612 13379 34664 13388
rect 34612 13345 34621 13379
rect 34621 13345 34655 13379
rect 34655 13345 34664 13379
rect 34612 13336 34664 13345
rect 35900 13336 35952 13388
rect 38108 13379 38160 13388
rect 38108 13345 38117 13379
rect 38117 13345 38151 13379
rect 38151 13345 38160 13379
rect 38108 13336 38160 13345
rect 38292 13336 38344 13388
rect 39396 13379 39448 13388
rect 39396 13345 39405 13379
rect 39405 13345 39439 13379
rect 39439 13345 39448 13379
rect 39396 13336 39448 13345
rect 39672 13379 39724 13388
rect 39672 13345 39681 13379
rect 39681 13345 39715 13379
rect 39715 13345 39724 13379
rect 39672 13336 39724 13345
rect 34152 13268 34204 13320
rect 36360 13311 36412 13320
rect 33048 13200 33100 13252
rect 34336 13200 34388 13252
rect 36360 13277 36369 13311
rect 36369 13277 36403 13311
rect 36403 13277 36412 13311
rect 36360 13268 36412 13277
rect 36820 13268 36872 13320
rect 37924 13268 37976 13320
rect 39948 13268 40000 13320
rect 36636 13200 36688 13252
rect 40408 13379 40460 13388
rect 40408 13345 40417 13379
rect 40417 13345 40451 13379
rect 40451 13345 40460 13379
rect 40408 13336 40460 13345
rect 40684 13336 40736 13388
rect 41052 13336 41104 13388
rect 43352 13379 43404 13388
rect 43352 13345 43361 13379
rect 43361 13345 43395 13379
rect 43395 13345 43404 13379
rect 43352 13336 43404 13345
rect 43536 13336 43588 13388
rect 44548 13379 44600 13388
rect 44548 13345 44557 13379
rect 44557 13345 44591 13379
rect 44591 13345 44600 13379
rect 44548 13336 44600 13345
rect 45652 13404 45704 13456
rect 45836 13404 45888 13456
rect 47308 13447 47360 13456
rect 47308 13413 47317 13447
rect 47317 13413 47351 13447
rect 47351 13413 47360 13447
rect 47308 13404 47360 13413
rect 48320 13472 48372 13524
rect 48228 13404 48280 13456
rect 49792 13472 49844 13524
rect 50252 13515 50304 13524
rect 50252 13481 50261 13515
rect 50261 13481 50295 13515
rect 50295 13481 50304 13515
rect 50252 13472 50304 13481
rect 50988 13472 51040 13524
rect 55128 13472 55180 13524
rect 57152 13515 57204 13524
rect 57152 13481 57161 13515
rect 57161 13481 57195 13515
rect 57195 13481 57204 13515
rect 57152 13472 57204 13481
rect 56784 13404 56836 13456
rect 57796 13404 57848 13456
rect 58440 13447 58492 13456
rect 58440 13413 58449 13447
rect 58449 13413 58483 13447
rect 58483 13413 58492 13447
rect 58440 13404 58492 13413
rect 46848 13379 46900 13388
rect 46848 13345 46857 13379
rect 46857 13345 46891 13379
rect 46891 13345 46900 13379
rect 46848 13336 46900 13345
rect 46940 13336 46992 13388
rect 48964 13379 49016 13388
rect 48964 13345 48973 13379
rect 48973 13345 49007 13379
rect 49007 13345 49016 13379
rect 48964 13336 49016 13345
rect 51080 13379 51132 13388
rect 51080 13345 51089 13379
rect 51089 13345 51123 13379
rect 51123 13345 51132 13379
rect 51080 13336 51132 13345
rect 52368 13379 52420 13388
rect 41144 13243 41196 13252
rect 41144 13209 41168 13243
rect 41168 13209 41196 13243
rect 41144 13200 41196 13209
rect 41420 13268 41472 13320
rect 41972 13268 42024 13320
rect 46204 13268 46256 13320
rect 46572 13268 46624 13320
rect 47032 13268 47084 13320
rect 48412 13268 48464 13320
rect 48688 13268 48740 13320
rect 49424 13268 49476 13320
rect 52368 13345 52377 13379
rect 52377 13345 52411 13379
rect 52411 13345 52420 13379
rect 52368 13336 52420 13345
rect 52092 13268 52144 13320
rect 55680 13336 55732 13388
rect 58256 13379 58308 13388
rect 58256 13345 58265 13379
rect 58265 13345 58299 13379
rect 58299 13345 58308 13379
rect 58256 13336 58308 13345
rect 59176 13336 59228 13388
rect 55588 13268 55640 13320
rect 56048 13311 56100 13320
rect 56048 13277 56057 13311
rect 56057 13277 56091 13311
rect 56091 13277 56100 13311
rect 56048 13268 56100 13277
rect 53472 13243 53524 13252
rect 24216 13132 24268 13184
rect 24860 13175 24912 13184
rect 24860 13141 24869 13175
rect 24869 13141 24903 13175
rect 24903 13141 24912 13175
rect 24860 13132 24912 13141
rect 26332 13132 26384 13184
rect 27436 13175 27488 13184
rect 27436 13141 27445 13175
rect 27445 13141 27479 13175
rect 27479 13141 27488 13175
rect 27436 13132 27488 13141
rect 28264 13132 28316 13184
rect 29736 13132 29788 13184
rect 30012 13175 30064 13184
rect 30012 13141 30021 13175
rect 30021 13141 30055 13175
rect 30055 13141 30064 13175
rect 30012 13132 30064 13141
rect 32036 13132 32088 13184
rect 32588 13175 32640 13184
rect 32588 13141 32597 13175
rect 32597 13141 32631 13175
rect 32631 13141 32640 13175
rect 32588 13132 32640 13141
rect 33416 13132 33468 13184
rect 34060 13132 34112 13184
rect 34888 13132 34940 13184
rect 34980 13132 35032 13184
rect 35256 13132 35308 13184
rect 36176 13175 36228 13184
rect 36176 13141 36200 13175
rect 36200 13141 36228 13175
rect 36176 13132 36228 13141
rect 36452 13132 36504 13184
rect 36820 13132 36872 13184
rect 39212 13175 39264 13184
rect 39212 13141 39221 13175
rect 39221 13141 39255 13175
rect 39255 13141 39264 13175
rect 39212 13132 39264 13141
rect 40592 13132 40644 13184
rect 41236 13175 41288 13184
rect 41236 13141 41245 13175
rect 41245 13141 41279 13175
rect 41279 13141 41288 13175
rect 41236 13132 41288 13141
rect 41788 13132 41840 13184
rect 41972 13175 42024 13184
rect 41972 13141 41981 13175
rect 41981 13141 42015 13175
rect 42015 13141 42024 13175
rect 41972 13132 42024 13141
rect 43076 13175 43128 13184
rect 43076 13141 43085 13175
rect 43085 13141 43119 13175
rect 43119 13141 43128 13175
rect 43076 13132 43128 13141
rect 43720 13132 43772 13184
rect 45192 13175 45244 13184
rect 45192 13141 45201 13175
rect 45201 13141 45235 13175
rect 45235 13141 45244 13175
rect 45192 13132 45244 13141
rect 47216 13132 47268 13184
rect 48044 13175 48096 13184
rect 48044 13141 48053 13175
rect 48053 13141 48087 13175
rect 48087 13141 48096 13175
rect 48044 13132 48096 13141
rect 48136 13175 48188 13184
rect 48136 13141 48145 13175
rect 48145 13141 48179 13175
rect 48179 13141 48188 13175
rect 48688 13175 48740 13184
rect 48136 13132 48188 13141
rect 48688 13141 48697 13175
rect 48697 13141 48731 13175
rect 48731 13141 48740 13175
rect 48688 13132 48740 13141
rect 48780 13132 48832 13184
rect 49240 13175 49292 13184
rect 49240 13141 49249 13175
rect 49249 13141 49283 13175
rect 49283 13141 49292 13175
rect 49240 13132 49292 13141
rect 51724 13132 51776 13184
rect 51908 13132 51960 13184
rect 52552 13175 52604 13184
rect 52552 13141 52561 13175
rect 52561 13141 52595 13175
rect 52595 13141 52604 13175
rect 52552 13132 52604 13141
rect 53472 13209 53481 13243
rect 53481 13209 53515 13243
rect 53515 13209 53524 13243
rect 53472 13200 53524 13209
rect 54208 13200 54260 13252
rect 57336 13200 57388 13252
rect 58716 13175 58768 13184
rect 58716 13141 58725 13175
rect 58725 13141 58759 13175
rect 58759 13141 58768 13175
rect 58716 13132 58768 13141
rect 59268 13175 59320 13184
rect 59268 13141 59277 13175
rect 59277 13141 59311 13175
rect 59311 13141 59320 13175
rect 59268 13132 59320 13141
rect 11378 13030 11430 13082
rect 11442 13030 11494 13082
rect 11506 13030 11558 13082
rect 11570 13030 11622 13082
rect 32170 13030 32222 13082
rect 32234 13030 32286 13082
rect 32298 13030 32350 13082
rect 32362 13030 32414 13082
rect 52962 13030 53014 13082
rect 53026 13030 53078 13082
rect 53090 13030 53142 13082
rect 53154 13030 53206 13082
rect 2412 12767 2464 12776
rect 2412 12733 2421 12767
rect 2421 12733 2455 12767
rect 2455 12733 2464 12767
rect 2412 12724 2464 12733
rect 3884 12792 3936 12844
rect 5724 12792 5776 12844
rect 7380 12792 7432 12844
rect 4988 12767 5040 12776
rect 4988 12733 4997 12767
rect 4997 12733 5031 12767
rect 5031 12733 5040 12767
rect 4988 12724 5040 12733
rect 5172 12767 5224 12776
rect 5172 12733 5181 12767
rect 5181 12733 5215 12767
rect 5215 12733 5224 12767
rect 5172 12724 5224 12733
rect 5448 12767 5500 12776
rect 5448 12733 5457 12767
rect 5457 12733 5491 12767
rect 5491 12733 5500 12767
rect 5448 12724 5500 12733
rect 6920 12724 6972 12776
rect 7288 12724 7340 12776
rect 5264 12656 5316 12708
rect 5356 12699 5408 12708
rect 5356 12665 5365 12699
rect 5365 12665 5399 12699
rect 5399 12665 5408 12699
rect 5356 12656 5408 12665
rect 8116 12767 8168 12776
rect 8116 12733 8125 12767
rect 8125 12733 8159 12767
rect 8159 12733 8168 12767
rect 8116 12724 8168 12733
rect 8484 12928 8536 12980
rect 9772 12971 9824 12980
rect 9772 12937 9781 12971
rect 9781 12937 9815 12971
rect 9815 12937 9824 12971
rect 9772 12928 9824 12937
rect 8760 12835 8812 12844
rect 8760 12801 8769 12835
rect 8769 12801 8803 12835
rect 8803 12801 8812 12835
rect 8760 12792 8812 12801
rect 9956 12835 10008 12844
rect 9956 12801 9965 12835
rect 9965 12801 9999 12835
rect 9999 12801 10008 12835
rect 9956 12792 10008 12801
rect 9128 12767 9180 12776
rect 9128 12733 9137 12767
rect 9137 12733 9171 12767
rect 9171 12733 9180 12767
rect 9128 12724 9180 12733
rect 4160 12588 4212 12640
rect 5816 12588 5868 12640
rect 8668 12588 8720 12640
rect 9496 12631 9548 12640
rect 9496 12597 9505 12631
rect 9505 12597 9539 12631
rect 9539 12597 9548 12631
rect 9496 12588 9548 12597
rect 10232 12792 10284 12844
rect 10324 12699 10376 12708
rect 10324 12665 10333 12699
rect 10333 12665 10367 12699
rect 10367 12665 10376 12699
rect 10324 12656 10376 12665
rect 11244 12656 11296 12708
rect 12532 12860 12584 12912
rect 12716 12903 12768 12912
rect 12716 12869 12725 12903
rect 12725 12869 12759 12903
rect 12759 12869 12768 12903
rect 12716 12860 12768 12869
rect 11980 12792 12032 12844
rect 12808 12835 12860 12844
rect 12808 12801 12817 12835
rect 12817 12801 12851 12835
rect 12851 12801 12860 12835
rect 12808 12792 12860 12801
rect 13636 12928 13688 12980
rect 14096 12903 14148 12912
rect 14096 12869 14105 12903
rect 14105 12869 14139 12903
rect 14139 12869 14148 12903
rect 14096 12860 14148 12869
rect 14464 12928 14516 12980
rect 14924 12928 14976 12980
rect 17408 12971 17460 12980
rect 17408 12937 17417 12971
rect 17417 12937 17451 12971
rect 17451 12937 17460 12971
rect 17408 12928 17460 12937
rect 19432 12928 19484 12980
rect 19524 12928 19576 12980
rect 22928 12971 22980 12980
rect 22928 12937 22937 12971
rect 22937 12937 22971 12971
rect 22971 12937 22980 12971
rect 22928 12928 22980 12937
rect 23388 12971 23440 12980
rect 23388 12937 23397 12971
rect 23397 12937 23431 12971
rect 23431 12937 23440 12971
rect 23388 12928 23440 12937
rect 24216 12971 24268 12980
rect 24216 12937 24225 12971
rect 24225 12937 24259 12971
rect 24259 12937 24268 12971
rect 24216 12928 24268 12937
rect 20812 12860 20864 12912
rect 22468 12860 22520 12912
rect 22652 12860 22704 12912
rect 23296 12860 23348 12912
rect 13084 12724 13136 12776
rect 14740 12767 14792 12776
rect 14740 12733 14749 12767
rect 14749 12733 14783 12767
rect 14783 12733 14792 12767
rect 14740 12724 14792 12733
rect 15292 12767 15344 12776
rect 11888 12656 11940 12708
rect 15292 12733 15301 12767
rect 15301 12733 15335 12767
rect 15335 12733 15344 12767
rect 15292 12724 15344 12733
rect 16948 12767 17000 12776
rect 15200 12656 15252 12708
rect 12256 12588 12308 12640
rect 13728 12588 13780 12640
rect 15476 12588 15528 12640
rect 16028 12588 16080 12640
rect 16948 12733 16957 12767
rect 16957 12733 16991 12767
rect 16991 12733 17000 12767
rect 16948 12724 17000 12733
rect 17500 12724 17552 12776
rect 18236 12767 18288 12776
rect 18236 12733 18245 12767
rect 18245 12733 18279 12767
rect 18279 12733 18288 12767
rect 18236 12724 18288 12733
rect 18328 12724 18380 12776
rect 19524 12792 19576 12844
rect 27712 12928 27764 12980
rect 28172 12928 28224 12980
rect 28816 12928 28868 12980
rect 30932 12971 30984 12980
rect 30932 12937 30941 12971
rect 30941 12937 30975 12971
rect 30975 12937 30984 12971
rect 30932 12928 30984 12937
rect 26056 12860 26108 12912
rect 27160 12860 27212 12912
rect 28356 12860 28408 12912
rect 29828 12860 29880 12912
rect 32588 12928 32640 12980
rect 32680 12971 32732 12980
rect 32680 12937 32689 12971
rect 32689 12937 32723 12971
rect 32723 12937 32732 12971
rect 32680 12928 32732 12937
rect 33508 12928 33560 12980
rect 36176 12928 36228 12980
rect 36360 12928 36412 12980
rect 38108 12971 38160 12980
rect 38108 12937 38117 12971
rect 38117 12937 38151 12971
rect 38151 12937 38160 12971
rect 38108 12928 38160 12937
rect 38844 12928 38896 12980
rect 39396 12928 39448 12980
rect 40408 12928 40460 12980
rect 40868 12928 40920 12980
rect 41512 12971 41564 12980
rect 41512 12937 41521 12971
rect 41521 12937 41555 12971
rect 41555 12937 41564 12971
rect 41512 12928 41564 12937
rect 26332 12835 26384 12844
rect 26332 12801 26341 12835
rect 26341 12801 26375 12835
rect 26375 12801 26384 12835
rect 26332 12792 26384 12801
rect 19623 12767 19675 12776
rect 18696 12656 18748 12708
rect 16948 12588 17000 12640
rect 17684 12588 17736 12640
rect 18880 12588 18932 12640
rect 18972 12588 19024 12640
rect 19623 12733 19625 12767
rect 19625 12733 19659 12767
rect 19659 12733 19675 12767
rect 19623 12724 19675 12733
rect 20904 12724 20956 12776
rect 22836 12724 22888 12776
rect 23664 12767 23716 12776
rect 23664 12733 23673 12767
rect 23673 12733 23707 12767
rect 23707 12733 23716 12767
rect 23664 12724 23716 12733
rect 24860 12724 24912 12776
rect 25964 12724 26016 12776
rect 31668 12792 31720 12844
rect 34980 12860 35032 12912
rect 35256 12860 35308 12912
rect 41328 12860 41380 12912
rect 45192 12971 45244 12980
rect 45192 12937 45201 12971
rect 45201 12937 45235 12971
rect 45235 12937 45244 12971
rect 45192 12928 45244 12937
rect 43536 12903 43588 12912
rect 33140 12835 33192 12844
rect 33140 12801 33149 12835
rect 33149 12801 33183 12835
rect 33183 12801 33192 12835
rect 33140 12792 33192 12801
rect 33416 12792 33468 12844
rect 33784 12792 33836 12844
rect 34244 12792 34296 12844
rect 38752 12792 38804 12844
rect 43536 12869 43545 12903
rect 43545 12869 43579 12903
rect 43579 12869 43588 12903
rect 43536 12860 43588 12869
rect 43720 12860 43772 12912
rect 46940 12928 46992 12980
rect 47216 12971 47268 12980
rect 47216 12937 47225 12971
rect 47225 12937 47259 12971
rect 47259 12937 47268 12971
rect 47216 12928 47268 12937
rect 47584 12971 47636 12980
rect 47584 12937 47593 12971
rect 47593 12937 47627 12971
rect 47627 12937 47636 12971
rect 47584 12928 47636 12937
rect 48044 12928 48096 12980
rect 49608 12928 49660 12980
rect 50712 12971 50764 12980
rect 50712 12937 50721 12971
rect 50721 12937 50755 12971
rect 50755 12937 50764 12971
rect 50712 12928 50764 12937
rect 52552 12928 52604 12980
rect 58256 12971 58308 12980
rect 47124 12860 47176 12912
rect 49240 12860 49292 12912
rect 50252 12860 50304 12912
rect 19524 12699 19576 12708
rect 19524 12665 19533 12699
rect 19533 12665 19567 12699
rect 19567 12665 19576 12699
rect 19524 12656 19576 12665
rect 21180 12631 21232 12640
rect 21180 12597 21189 12631
rect 21189 12597 21223 12631
rect 21223 12597 21232 12631
rect 21824 12699 21876 12708
rect 21824 12665 21833 12699
rect 21833 12665 21867 12699
rect 21867 12665 21876 12699
rect 21824 12656 21876 12665
rect 22192 12656 22244 12708
rect 22468 12656 22520 12708
rect 28540 12724 28592 12776
rect 30196 12767 30248 12776
rect 30196 12733 30205 12767
rect 30205 12733 30239 12767
rect 30239 12733 30248 12767
rect 30196 12724 30248 12733
rect 31392 12767 31444 12776
rect 31392 12733 31401 12767
rect 31401 12733 31435 12767
rect 31435 12733 31444 12767
rect 31392 12724 31444 12733
rect 31576 12724 31628 12776
rect 21180 12588 21232 12597
rect 22560 12588 22612 12640
rect 24768 12588 24820 12640
rect 30012 12656 30064 12708
rect 31208 12699 31260 12708
rect 31208 12665 31217 12699
rect 31217 12665 31251 12699
rect 31251 12665 31260 12699
rect 31208 12656 31260 12665
rect 32128 12699 32180 12708
rect 32128 12665 32137 12699
rect 32137 12665 32171 12699
rect 32171 12665 32180 12699
rect 32128 12656 32180 12665
rect 28724 12631 28776 12640
rect 28724 12597 28733 12631
rect 28733 12597 28767 12631
rect 28767 12597 28776 12631
rect 28724 12588 28776 12597
rect 31392 12588 31444 12640
rect 32036 12588 32088 12640
rect 33048 12724 33100 12776
rect 33968 12724 34020 12776
rect 34520 12724 34572 12776
rect 34060 12699 34112 12708
rect 34060 12665 34069 12699
rect 34069 12665 34103 12699
rect 34103 12665 34112 12699
rect 34060 12656 34112 12665
rect 34796 12656 34848 12708
rect 34612 12631 34664 12640
rect 34612 12597 34621 12631
rect 34621 12597 34655 12631
rect 34655 12597 34664 12631
rect 34612 12588 34664 12597
rect 36176 12724 36228 12776
rect 36728 12767 36780 12776
rect 36728 12733 36737 12767
rect 36737 12733 36771 12767
rect 36771 12733 36780 12767
rect 36728 12724 36780 12733
rect 37004 12767 37056 12776
rect 37004 12733 37013 12767
rect 37013 12733 37047 12767
rect 37047 12733 37056 12767
rect 37004 12724 37056 12733
rect 37188 12767 37240 12776
rect 37188 12733 37197 12767
rect 37197 12733 37231 12767
rect 37231 12733 37240 12767
rect 37188 12724 37240 12733
rect 37740 12767 37792 12776
rect 37740 12733 37749 12767
rect 37749 12733 37783 12767
rect 37783 12733 37792 12767
rect 37740 12724 37792 12733
rect 38660 12724 38712 12776
rect 39212 12724 39264 12776
rect 35348 12656 35400 12708
rect 40868 12724 40920 12776
rect 41420 12724 41472 12776
rect 42984 12792 43036 12844
rect 43352 12792 43404 12844
rect 46848 12792 46900 12844
rect 47308 12835 47360 12844
rect 47308 12801 47317 12835
rect 47317 12801 47351 12835
rect 47351 12801 47360 12835
rect 47308 12792 47360 12801
rect 48688 12792 48740 12844
rect 52368 12860 52420 12912
rect 53656 12860 53708 12912
rect 56048 12903 56100 12912
rect 50528 12792 50580 12844
rect 56048 12869 56057 12903
rect 56057 12869 56091 12903
rect 56091 12869 56100 12903
rect 56048 12860 56100 12869
rect 56784 12903 56836 12912
rect 56784 12869 56793 12903
rect 56793 12869 56827 12903
rect 56827 12869 56836 12903
rect 56784 12860 56836 12869
rect 35808 12631 35860 12640
rect 35808 12597 35817 12631
rect 35817 12597 35851 12631
rect 35851 12597 35860 12631
rect 35808 12588 35860 12597
rect 36452 12588 36504 12640
rect 38108 12588 38160 12640
rect 38844 12588 38896 12640
rect 39028 12588 39080 12640
rect 39488 12588 39540 12640
rect 44548 12724 44600 12776
rect 45560 12724 45612 12776
rect 45836 12767 45888 12776
rect 45836 12733 45845 12767
rect 45845 12733 45879 12767
rect 45879 12733 45888 12767
rect 45836 12724 45888 12733
rect 45928 12724 45980 12776
rect 49424 12724 49476 12776
rect 51908 12767 51960 12776
rect 43352 12656 43404 12708
rect 44272 12699 44324 12708
rect 44272 12665 44281 12699
rect 44281 12665 44315 12699
rect 44315 12665 44324 12699
rect 44272 12656 44324 12665
rect 46940 12699 46992 12708
rect 46940 12665 46949 12699
rect 46949 12665 46983 12699
rect 46983 12665 46992 12699
rect 46940 12656 46992 12665
rect 48504 12699 48556 12708
rect 48504 12665 48513 12699
rect 48513 12665 48547 12699
rect 48547 12665 48556 12699
rect 48504 12656 48556 12665
rect 50068 12699 50120 12708
rect 50068 12665 50077 12699
rect 50077 12665 50111 12699
rect 50111 12665 50120 12699
rect 50068 12656 50120 12665
rect 51908 12733 51917 12767
rect 51917 12733 51951 12767
rect 51951 12733 51960 12767
rect 51908 12724 51960 12733
rect 53288 12767 53340 12776
rect 53288 12733 53297 12767
rect 53297 12733 53331 12767
rect 53331 12733 53340 12767
rect 53288 12724 53340 12733
rect 53472 12724 53524 12776
rect 51540 12656 51592 12708
rect 55220 12792 55272 12844
rect 58256 12937 58265 12971
rect 58265 12937 58299 12971
rect 58299 12937 58308 12971
rect 58256 12928 58308 12937
rect 57796 12792 57848 12844
rect 58900 12835 58952 12844
rect 58900 12801 58909 12835
rect 58909 12801 58943 12835
rect 58943 12801 58952 12835
rect 58900 12792 58952 12801
rect 59268 12792 59320 12844
rect 41972 12588 42024 12640
rect 50252 12588 50304 12640
rect 51632 12588 51684 12640
rect 53288 12588 53340 12640
rect 53380 12588 53432 12640
rect 55128 12656 55180 12708
rect 55680 12631 55732 12640
rect 55680 12597 55689 12631
rect 55689 12597 55723 12631
rect 55723 12597 55732 12631
rect 55680 12588 55732 12597
rect 55864 12656 55916 12708
rect 60004 12631 60056 12640
rect 60004 12597 60013 12631
rect 60013 12597 60047 12631
rect 60047 12597 60056 12631
rect 60004 12588 60056 12597
rect 21774 12486 21826 12538
rect 21838 12486 21890 12538
rect 21902 12486 21954 12538
rect 21966 12486 22018 12538
rect 42566 12486 42618 12538
rect 42630 12486 42682 12538
rect 42694 12486 42746 12538
rect 42758 12486 42810 12538
rect 4068 12384 4120 12436
rect 5908 12384 5960 12436
rect 7012 12384 7064 12436
rect 7564 12384 7616 12436
rect 5356 12316 5408 12368
rect 8300 12316 8352 12368
rect 8760 12384 8812 12436
rect 9864 12384 9916 12436
rect 10324 12384 10376 12436
rect 11152 12384 11204 12436
rect 12072 12427 12124 12436
rect 12072 12393 12081 12427
rect 12081 12393 12115 12427
rect 12115 12393 12124 12427
rect 12072 12384 12124 12393
rect 12164 12384 12216 12436
rect 12808 12384 12860 12436
rect 15476 12384 15528 12436
rect 16304 12384 16356 12436
rect 17776 12384 17828 12436
rect 19340 12384 19392 12436
rect 20260 12384 20312 12436
rect 9128 12316 9180 12368
rect 15200 12316 15252 12368
rect 17316 12316 17368 12368
rect 20904 12359 20956 12368
rect 2688 12248 2740 12300
rect 5080 12291 5132 12300
rect 5080 12257 5089 12291
rect 5089 12257 5123 12291
rect 5123 12257 5132 12291
rect 5080 12248 5132 12257
rect 5448 12291 5500 12300
rect 5448 12257 5457 12291
rect 5457 12257 5491 12291
rect 5491 12257 5500 12291
rect 5448 12248 5500 12257
rect 6552 12248 6604 12300
rect 10692 12291 10744 12300
rect 10692 12257 10701 12291
rect 10701 12257 10735 12291
rect 10735 12257 10744 12291
rect 10692 12248 10744 12257
rect 3332 12180 3384 12232
rect 5540 12223 5592 12232
rect 5540 12189 5549 12223
rect 5549 12189 5583 12223
rect 5583 12189 5592 12223
rect 5540 12180 5592 12189
rect 7564 12223 7616 12232
rect 7564 12189 7570 12223
rect 7570 12189 7616 12223
rect 7564 12180 7616 12189
rect 8208 12180 8260 12232
rect 12164 12248 12216 12300
rect 12532 12248 12584 12300
rect 14280 12248 14332 12300
rect 11888 12180 11940 12232
rect 2872 12112 2924 12164
rect 9404 12112 9456 12164
rect 12164 12112 12216 12164
rect 6920 12087 6972 12096
rect 6920 12053 6929 12087
rect 6929 12053 6963 12087
rect 6963 12053 6972 12087
rect 6920 12044 6972 12053
rect 7564 12044 7616 12096
rect 10600 12087 10652 12096
rect 10600 12053 10609 12087
rect 10609 12053 10643 12087
rect 10643 12053 10652 12087
rect 10600 12044 10652 12053
rect 10968 12087 11020 12096
rect 10968 12053 10977 12087
rect 10977 12053 11011 12087
rect 11011 12053 11020 12087
rect 10968 12044 11020 12053
rect 12716 12044 12768 12096
rect 13084 12044 13136 12096
rect 14096 12180 14148 12232
rect 14924 12180 14976 12232
rect 15660 12248 15712 12300
rect 16212 12248 16264 12300
rect 16672 12291 16724 12300
rect 16672 12257 16681 12291
rect 16681 12257 16715 12291
rect 16715 12257 16724 12291
rect 16672 12248 16724 12257
rect 16856 12291 16908 12300
rect 16856 12257 16865 12291
rect 16865 12257 16899 12291
rect 16899 12257 16908 12291
rect 16856 12248 16908 12257
rect 18696 12248 18748 12300
rect 19524 12248 19576 12300
rect 20628 12291 20680 12300
rect 20628 12257 20637 12291
rect 20637 12257 20671 12291
rect 20671 12257 20680 12291
rect 20628 12248 20680 12257
rect 19156 12180 19208 12232
rect 18328 12112 18380 12164
rect 18420 12112 18472 12164
rect 18972 12112 19024 12164
rect 19616 12112 19668 12164
rect 20536 12112 20588 12164
rect 20904 12325 20913 12359
rect 20913 12325 20947 12359
rect 20947 12325 20956 12359
rect 20904 12316 20956 12325
rect 21088 12384 21140 12436
rect 24492 12427 24544 12436
rect 21456 12248 21508 12300
rect 21732 12291 21784 12300
rect 21732 12257 21741 12291
rect 21741 12257 21775 12291
rect 21775 12257 21784 12291
rect 21732 12248 21784 12257
rect 22100 12248 22152 12300
rect 22928 12291 22980 12300
rect 22928 12257 22937 12291
rect 22937 12257 22971 12291
rect 22971 12257 22980 12291
rect 22928 12248 22980 12257
rect 24492 12393 24501 12427
rect 24501 12393 24535 12427
rect 24535 12393 24544 12427
rect 24492 12384 24544 12393
rect 24860 12384 24912 12436
rect 25780 12384 25832 12436
rect 26056 12384 26108 12436
rect 26240 12427 26292 12436
rect 26240 12393 26249 12427
rect 26249 12393 26283 12427
rect 26283 12393 26292 12427
rect 26240 12384 26292 12393
rect 27712 12427 27764 12436
rect 27712 12393 27721 12427
rect 27721 12393 27755 12427
rect 27755 12393 27764 12427
rect 27712 12384 27764 12393
rect 33140 12384 33192 12436
rect 33324 12384 33376 12436
rect 33508 12427 33560 12436
rect 33508 12393 33517 12427
rect 33517 12393 33551 12427
rect 33551 12393 33560 12427
rect 33508 12384 33560 12393
rect 35256 12427 35308 12436
rect 35256 12393 35265 12427
rect 35265 12393 35299 12427
rect 35299 12393 35308 12427
rect 35256 12384 35308 12393
rect 36268 12384 36320 12436
rect 37188 12427 37240 12436
rect 37188 12393 37197 12427
rect 37197 12393 37231 12427
rect 37231 12393 37240 12427
rect 37188 12384 37240 12393
rect 39580 12384 39632 12436
rect 40684 12427 40736 12436
rect 40684 12393 40693 12427
rect 40693 12393 40727 12427
rect 40727 12393 40736 12427
rect 40684 12384 40736 12393
rect 41788 12427 41840 12436
rect 41788 12393 41797 12427
rect 41797 12393 41831 12427
rect 41831 12393 41840 12427
rect 41788 12384 41840 12393
rect 43076 12427 43128 12436
rect 43076 12393 43085 12427
rect 43085 12393 43119 12427
rect 43119 12393 43128 12427
rect 43076 12384 43128 12393
rect 23112 12316 23164 12368
rect 23940 12316 23992 12368
rect 32496 12316 32548 12368
rect 23848 12248 23900 12300
rect 24952 12291 25004 12300
rect 24952 12257 24961 12291
rect 24961 12257 24995 12291
rect 24995 12257 25004 12291
rect 24952 12248 25004 12257
rect 25320 12291 25372 12300
rect 25320 12257 25329 12291
rect 25329 12257 25363 12291
rect 25363 12257 25372 12291
rect 25320 12248 25372 12257
rect 26240 12248 26292 12300
rect 26792 12291 26844 12300
rect 26792 12257 26801 12291
rect 26801 12257 26835 12291
rect 26835 12257 26844 12291
rect 27252 12291 27304 12300
rect 26792 12248 26844 12257
rect 27252 12257 27261 12291
rect 27261 12257 27295 12291
rect 27295 12257 27304 12291
rect 27252 12248 27304 12257
rect 27344 12248 27396 12300
rect 28540 12248 28592 12300
rect 30104 12291 30156 12300
rect 22560 12180 22612 12232
rect 23296 12180 23348 12232
rect 30104 12257 30113 12291
rect 30113 12257 30147 12291
rect 30147 12257 30156 12291
rect 30104 12248 30156 12257
rect 30288 12248 30340 12300
rect 32588 12248 32640 12300
rect 34152 12316 34204 12368
rect 23112 12112 23164 12164
rect 24216 12112 24268 12164
rect 14464 12044 14516 12096
rect 17316 12044 17368 12096
rect 17500 12087 17552 12096
rect 17500 12053 17509 12087
rect 17509 12053 17543 12087
rect 17543 12053 17552 12087
rect 17500 12044 17552 12053
rect 17684 12044 17736 12096
rect 19524 12044 19576 12096
rect 19800 12044 19852 12096
rect 21456 12044 21508 12096
rect 22192 12044 22244 12096
rect 24124 12087 24176 12096
rect 24124 12053 24133 12087
rect 24133 12053 24167 12087
rect 24167 12053 24176 12087
rect 24124 12044 24176 12053
rect 25780 12044 25832 12096
rect 27160 12112 27212 12164
rect 28908 12180 28960 12232
rect 27712 12112 27764 12164
rect 29184 12112 29236 12164
rect 29460 12112 29512 12164
rect 31576 12112 31628 12164
rect 29000 12087 29052 12096
rect 29000 12053 29009 12087
rect 29009 12053 29043 12087
rect 29043 12053 29052 12087
rect 29000 12044 29052 12053
rect 33968 12248 34020 12300
rect 34336 12291 34388 12300
rect 34336 12257 34345 12291
rect 34345 12257 34379 12291
rect 34379 12257 34388 12291
rect 34336 12248 34388 12257
rect 34520 12248 34572 12300
rect 37740 12359 37792 12368
rect 37740 12325 37749 12359
rect 37749 12325 37783 12359
rect 37783 12325 37792 12359
rect 37740 12316 37792 12325
rect 37832 12316 37884 12368
rect 35716 12291 35768 12300
rect 35716 12257 35725 12291
rect 35725 12257 35759 12291
rect 35759 12257 35768 12291
rect 35716 12248 35768 12257
rect 39764 12316 39816 12368
rect 46112 12359 46164 12368
rect 33692 12180 33744 12232
rect 34796 12180 34848 12232
rect 35532 12112 35584 12164
rect 36084 12223 36136 12232
rect 36084 12189 36093 12223
rect 36093 12189 36127 12223
rect 36127 12189 36136 12223
rect 36084 12180 36136 12189
rect 36820 12180 36872 12232
rect 38292 12223 38344 12232
rect 38292 12189 38301 12223
rect 38301 12189 38335 12223
rect 38335 12189 38344 12223
rect 38292 12180 38344 12189
rect 39948 12248 40000 12300
rect 41880 12248 41932 12300
rect 39856 12180 39908 12232
rect 41512 12180 41564 12232
rect 37832 12112 37884 12164
rect 39672 12112 39724 12164
rect 46112 12325 46121 12359
rect 46121 12325 46155 12359
rect 46155 12325 46164 12359
rect 46112 12316 46164 12325
rect 52552 12384 52604 12436
rect 49240 12316 49292 12368
rect 50252 12316 50304 12368
rect 55404 12316 55456 12368
rect 55864 12359 55916 12368
rect 55864 12325 55873 12359
rect 55873 12325 55907 12359
rect 55907 12325 55916 12359
rect 55864 12316 55916 12325
rect 42984 12248 43036 12300
rect 42156 12180 42208 12232
rect 43444 12180 43496 12232
rect 44272 12248 44324 12300
rect 44916 12248 44968 12300
rect 44180 12223 44232 12232
rect 44180 12189 44189 12223
rect 44189 12189 44223 12223
rect 44223 12189 44232 12223
rect 44180 12180 44232 12189
rect 44456 12223 44508 12232
rect 44456 12189 44465 12223
rect 44465 12189 44499 12223
rect 44499 12189 44508 12223
rect 44456 12180 44508 12189
rect 46848 12248 46900 12300
rect 47032 12248 47084 12300
rect 48320 12248 48372 12300
rect 48872 12248 48924 12300
rect 49056 12291 49108 12300
rect 49056 12257 49065 12291
rect 49065 12257 49099 12291
rect 49099 12257 49108 12291
rect 49056 12248 49108 12257
rect 50712 12291 50764 12300
rect 50712 12257 50721 12291
rect 50721 12257 50755 12291
rect 50755 12257 50764 12291
rect 50712 12248 50764 12257
rect 51448 12248 51500 12300
rect 52828 12248 52880 12300
rect 53472 12248 53524 12300
rect 55128 12291 55180 12300
rect 55128 12257 55137 12291
rect 55137 12257 55171 12291
rect 55171 12257 55180 12291
rect 55128 12248 55180 12257
rect 56876 12248 56928 12300
rect 58072 12316 58124 12368
rect 58440 12384 58492 12436
rect 60004 12316 60056 12368
rect 60556 12248 60608 12300
rect 46572 12180 46624 12232
rect 46664 12223 46716 12232
rect 46664 12189 46673 12223
rect 46673 12189 46707 12223
rect 46707 12189 46716 12223
rect 46664 12180 46716 12189
rect 46940 12180 46992 12232
rect 48964 12223 49016 12232
rect 48964 12189 48973 12223
rect 48973 12189 49007 12223
rect 49007 12189 49016 12223
rect 48964 12180 49016 12189
rect 51264 12223 51316 12232
rect 51264 12189 51273 12223
rect 51273 12189 51307 12223
rect 51307 12189 51316 12223
rect 51264 12180 51316 12189
rect 51724 12223 51776 12232
rect 51724 12189 51733 12223
rect 51733 12189 51767 12223
rect 51767 12189 51776 12223
rect 51724 12180 51776 12189
rect 53288 12180 53340 12232
rect 54116 12180 54168 12232
rect 55496 12223 55548 12232
rect 55496 12189 55505 12223
rect 55505 12189 55539 12223
rect 55539 12189 55548 12223
rect 55496 12180 55548 12189
rect 57888 12180 57940 12232
rect 34796 12044 34848 12096
rect 35624 12087 35676 12096
rect 35624 12053 35633 12087
rect 35633 12053 35667 12087
rect 35667 12053 35676 12087
rect 35624 12044 35676 12053
rect 36452 12044 36504 12096
rect 36820 12087 36872 12096
rect 36820 12053 36829 12087
rect 36829 12053 36863 12087
rect 36863 12053 36872 12087
rect 36820 12044 36872 12053
rect 40868 12044 40920 12096
rect 41788 12044 41840 12096
rect 47032 12112 47084 12164
rect 49056 12112 49108 12164
rect 50252 12112 50304 12164
rect 48504 12044 48556 12096
rect 50068 12087 50120 12096
rect 50068 12053 50077 12087
rect 50077 12053 50111 12087
rect 50111 12053 50120 12087
rect 50068 12044 50120 12053
rect 50528 12044 50580 12096
rect 50620 12044 50672 12096
rect 51080 12044 51132 12096
rect 51632 12112 51684 12164
rect 51908 12112 51960 12164
rect 52276 12112 52328 12164
rect 54208 12112 54260 12164
rect 52368 12087 52420 12096
rect 52368 12053 52377 12087
rect 52377 12053 52411 12087
rect 52411 12053 52420 12087
rect 52368 12044 52420 12053
rect 53932 12087 53984 12096
rect 53932 12053 53941 12087
rect 53941 12053 53975 12087
rect 53975 12053 53984 12087
rect 53932 12044 53984 12053
rect 55220 12044 55272 12096
rect 55404 12087 55456 12096
rect 55404 12053 55413 12087
rect 55413 12053 55447 12087
rect 55447 12053 55456 12087
rect 55404 12044 55456 12053
rect 55956 12044 56008 12096
rect 56692 12044 56744 12096
rect 56876 12087 56928 12096
rect 56876 12053 56885 12087
rect 56885 12053 56919 12087
rect 56919 12053 56928 12087
rect 56876 12044 56928 12053
rect 57796 12112 57848 12164
rect 58164 12044 58216 12096
rect 59176 12087 59228 12096
rect 59176 12053 59185 12087
rect 59185 12053 59219 12087
rect 59219 12053 59228 12087
rect 59176 12044 59228 12053
rect 59728 12087 59780 12096
rect 59728 12053 59737 12087
rect 59737 12053 59771 12087
rect 59771 12053 59780 12087
rect 59728 12044 59780 12053
rect 11378 11942 11430 11994
rect 11442 11942 11494 11994
rect 11506 11942 11558 11994
rect 11570 11942 11622 11994
rect 32170 11942 32222 11994
rect 32234 11942 32286 11994
rect 32298 11942 32350 11994
rect 32362 11942 32414 11994
rect 52962 11942 53014 11994
rect 53026 11942 53078 11994
rect 53090 11942 53142 11994
rect 53154 11942 53206 11994
rect 2872 11883 2924 11892
rect 2872 11849 2881 11883
rect 2881 11849 2915 11883
rect 2915 11849 2924 11883
rect 2872 11840 2924 11849
rect 4712 11840 4764 11892
rect 5448 11840 5500 11892
rect 6552 11883 6604 11892
rect 6552 11849 6561 11883
rect 6561 11849 6595 11883
rect 6595 11849 6604 11883
rect 6552 11840 6604 11849
rect 8024 11840 8076 11892
rect 8392 11840 8444 11892
rect 10968 11840 11020 11892
rect 12164 11883 12216 11892
rect 12164 11849 12173 11883
rect 12173 11849 12207 11883
rect 12207 11849 12216 11883
rect 12164 11840 12216 11849
rect 12532 11840 12584 11892
rect 7564 11815 7616 11824
rect 7564 11781 7573 11815
rect 7573 11781 7607 11815
rect 7607 11781 7616 11815
rect 7564 11772 7616 11781
rect 3332 11747 3384 11756
rect 3332 11713 3341 11747
rect 3341 11713 3375 11747
rect 3375 11713 3384 11747
rect 3332 11704 3384 11713
rect 7656 11747 7708 11756
rect 7656 11713 7665 11747
rect 7665 11713 7699 11747
rect 7699 11713 7708 11747
rect 7656 11704 7708 11713
rect 8208 11704 8260 11756
rect 8484 11704 8536 11756
rect 12624 11772 12676 11824
rect 14464 11840 14516 11892
rect 15660 11883 15712 11892
rect 15660 11849 15669 11883
rect 15669 11849 15703 11883
rect 15703 11849 15712 11883
rect 15660 11840 15712 11849
rect 16856 11840 16908 11892
rect 17500 11840 17552 11892
rect 17592 11840 17644 11892
rect 15844 11772 15896 11824
rect 19156 11772 19208 11824
rect 21088 11815 21140 11824
rect 21088 11781 21097 11815
rect 21097 11781 21131 11815
rect 21131 11781 21140 11815
rect 21088 11772 21140 11781
rect 22100 11840 22152 11892
rect 23848 11883 23900 11892
rect 23848 11849 23857 11883
rect 23857 11849 23891 11883
rect 23891 11849 23900 11883
rect 23848 11840 23900 11849
rect 27252 11840 27304 11892
rect 29000 11883 29052 11892
rect 29000 11849 29009 11883
rect 29009 11849 29043 11883
rect 29043 11849 29052 11883
rect 29000 11840 29052 11849
rect 30196 11840 30248 11892
rect 33324 11840 33376 11892
rect 30748 11772 30800 11824
rect 34152 11840 34204 11892
rect 34336 11883 34388 11892
rect 34336 11849 34345 11883
rect 34345 11849 34379 11883
rect 34379 11849 34388 11883
rect 34336 11840 34388 11849
rect 34520 11840 34572 11892
rect 35532 11883 35584 11892
rect 35532 11849 35541 11883
rect 35541 11849 35575 11883
rect 35575 11849 35584 11883
rect 35532 11840 35584 11849
rect 33692 11772 33744 11824
rect 37004 11840 37056 11892
rect 39764 11883 39816 11892
rect 39764 11849 39773 11883
rect 39773 11849 39807 11883
rect 39807 11849 39816 11883
rect 39764 11840 39816 11849
rect 39948 11840 40000 11892
rect 40868 11883 40920 11892
rect 40868 11849 40877 11883
rect 40877 11849 40911 11883
rect 40911 11849 40920 11883
rect 40868 11840 40920 11849
rect 41512 11840 41564 11892
rect 43352 11840 43404 11892
rect 43444 11840 43496 11892
rect 48412 11883 48464 11892
rect 36452 11772 36504 11824
rect 41972 11772 42024 11824
rect 44456 11815 44508 11824
rect 44456 11781 44465 11815
rect 44465 11781 44499 11815
rect 44499 11781 44508 11815
rect 44456 11772 44508 11781
rect 48412 11849 48421 11883
rect 48421 11849 48455 11883
rect 48455 11849 48464 11883
rect 48412 11840 48464 11849
rect 48780 11883 48832 11892
rect 48780 11849 48789 11883
rect 48789 11849 48823 11883
rect 48823 11849 48832 11883
rect 48780 11840 48832 11849
rect 49056 11840 49108 11892
rect 50528 11883 50580 11892
rect 50528 11849 50537 11883
rect 50537 11849 50571 11883
rect 50571 11849 50580 11883
rect 50528 11840 50580 11849
rect 51724 11840 51776 11892
rect 51908 11840 51960 11892
rect 52368 11883 52420 11892
rect 52368 11849 52377 11883
rect 52377 11849 52411 11883
rect 52411 11849 52420 11883
rect 52368 11840 52420 11849
rect 52460 11840 52512 11892
rect 53472 11883 53524 11892
rect 53472 11849 53481 11883
rect 53481 11849 53515 11883
rect 53515 11849 53524 11883
rect 53472 11840 53524 11849
rect 54576 11883 54628 11892
rect 54576 11849 54585 11883
rect 54585 11849 54619 11883
rect 54619 11849 54628 11883
rect 54576 11840 54628 11849
rect 55496 11840 55548 11892
rect 50896 11772 50948 11824
rect 52000 11815 52052 11824
rect 52000 11781 52009 11815
rect 52009 11781 52043 11815
rect 52043 11781 52052 11815
rect 52000 11772 52052 11781
rect 53564 11772 53616 11824
rect 55404 11772 55456 11824
rect 4252 11636 4304 11688
rect 8668 11636 8720 11688
rect 8852 11679 8904 11688
rect 8852 11645 8861 11679
rect 8861 11645 8895 11679
rect 8895 11645 8904 11679
rect 8852 11636 8904 11645
rect 9772 11636 9824 11688
rect 10600 11636 10652 11688
rect 23940 11704 23992 11756
rect 25780 11747 25832 11756
rect 25780 11713 25789 11747
rect 25789 11713 25823 11747
rect 25823 11713 25832 11747
rect 25780 11704 25832 11713
rect 27160 11747 27212 11756
rect 27160 11713 27169 11747
rect 27169 11713 27203 11747
rect 27203 11713 27212 11747
rect 27160 11704 27212 11713
rect 27436 11704 27488 11756
rect 31668 11704 31720 11756
rect 31760 11704 31812 11756
rect 2872 11500 2924 11552
rect 2964 11500 3016 11552
rect 6920 11568 6972 11620
rect 11244 11636 11296 11688
rect 4620 11500 4672 11552
rect 5080 11543 5132 11552
rect 5080 11509 5089 11543
rect 5089 11509 5123 11543
rect 5123 11509 5132 11543
rect 5080 11500 5132 11509
rect 5540 11543 5592 11552
rect 5540 11509 5549 11543
rect 5549 11509 5583 11543
rect 5583 11509 5592 11543
rect 5540 11500 5592 11509
rect 7012 11500 7064 11552
rect 7196 11500 7248 11552
rect 9772 11543 9824 11552
rect 9772 11509 9781 11543
rect 9781 11509 9815 11543
rect 9815 11509 9824 11543
rect 9772 11500 9824 11509
rect 9956 11500 10008 11552
rect 12348 11568 12400 11620
rect 13728 11568 13780 11620
rect 14280 11636 14332 11688
rect 14464 11679 14516 11688
rect 14464 11645 14473 11679
rect 14473 11645 14507 11679
rect 14507 11645 14516 11679
rect 14464 11636 14516 11645
rect 15200 11636 15252 11688
rect 16396 11636 16448 11688
rect 17960 11636 18012 11688
rect 18328 11679 18380 11688
rect 18328 11645 18337 11679
rect 18337 11645 18371 11679
rect 18371 11645 18380 11679
rect 18328 11636 18380 11645
rect 15292 11568 15344 11620
rect 14464 11500 14516 11552
rect 15108 11500 15160 11552
rect 18052 11568 18104 11620
rect 18236 11568 18288 11620
rect 19616 11636 19668 11688
rect 19800 11636 19852 11688
rect 21088 11636 21140 11688
rect 22192 11679 22244 11688
rect 22192 11645 22201 11679
rect 22201 11645 22235 11679
rect 22235 11645 22244 11679
rect 22192 11636 22244 11645
rect 23020 11636 23072 11688
rect 23296 11636 23348 11688
rect 24492 11636 24544 11688
rect 18880 11611 18932 11620
rect 18880 11577 18889 11611
rect 18889 11577 18923 11611
rect 18923 11577 18932 11611
rect 18880 11568 18932 11577
rect 20904 11568 20956 11620
rect 24124 11611 24176 11620
rect 24124 11577 24133 11611
rect 24133 11577 24167 11611
rect 24167 11577 24176 11611
rect 24124 11568 24176 11577
rect 25136 11568 25188 11620
rect 16396 11543 16448 11552
rect 16396 11509 16405 11543
rect 16405 11509 16439 11543
rect 16439 11509 16448 11543
rect 16396 11500 16448 11509
rect 17776 11543 17828 11552
rect 17776 11509 17785 11543
rect 17785 11509 17819 11543
rect 17819 11509 17828 11543
rect 17776 11500 17828 11509
rect 19156 11500 19208 11552
rect 23020 11543 23072 11552
rect 23020 11509 23029 11543
rect 23029 11509 23063 11543
rect 23063 11509 23072 11543
rect 23020 11500 23072 11509
rect 24952 11500 25004 11552
rect 25412 11500 25464 11552
rect 27804 11636 27856 11688
rect 28908 11636 28960 11688
rect 29000 11636 29052 11688
rect 25872 11500 25924 11552
rect 26792 11500 26844 11552
rect 27528 11500 27580 11552
rect 29092 11568 29144 11620
rect 32404 11704 32456 11756
rect 33876 11747 33928 11756
rect 32864 11636 32916 11688
rect 33416 11679 33468 11688
rect 33416 11645 33425 11679
rect 33425 11645 33459 11679
rect 33459 11645 33468 11679
rect 33416 11636 33468 11645
rect 33876 11713 33885 11747
rect 33885 11713 33919 11747
rect 33919 11713 33928 11747
rect 33876 11704 33928 11713
rect 36820 11704 36872 11756
rect 28264 11500 28316 11552
rect 30196 11543 30248 11552
rect 30196 11509 30205 11543
rect 30205 11509 30239 11543
rect 30239 11509 30248 11543
rect 30196 11500 30248 11509
rect 31484 11500 31536 11552
rect 31760 11611 31812 11620
rect 31760 11577 31769 11611
rect 31769 11577 31803 11611
rect 31803 11577 31812 11611
rect 31760 11568 31812 11577
rect 33508 11568 33560 11620
rect 33600 11568 33652 11620
rect 35164 11568 35216 11620
rect 32496 11500 32548 11552
rect 32588 11500 32640 11552
rect 33048 11500 33100 11552
rect 33140 11500 33192 11552
rect 35348 11500 35400 11552
rect 37832 11704 37884 11756
rect 37464 11679 37516 11688
rect 35624 11568 35676 11620
rect 37464 11645 37473 11679
rect 37473 11645 37507 11679
rect 37507 11645 37516 11679
rect 37464 11636 37516 11645
rect 37280 11611 37332 11620
rect 37280 11577 37289 11611
rect 37289 11577 37323 11611
rect 37323 11577 37332 11611
rect 37280 11568 37332 11577
rect 38660 11611 38712 11620
rect 38660 11577 38669 11611
rect 38669 11577 38703 11611
rect 38703 11577 38712 11611
rect 38660 11568 38712 11577
rect 40408 11568 40460 11620
rect 41696 11704 41748 11756
rect 41788 11679 41840 11688
rect 41788 11645 41797 11679
rect 41797 11645 41831 11679
rect 41831 11645 41840 11679
rect 41788 11636 41840 11645
rect 41972 11636 42024 11688
rect 45284 11704 45336 11756
rect 48320 11704 48372 11756
rect 50620 11704 50672 11756
rect 52460 11747 52512 11756
rect 52460 11713 52469 11747
rect 52469 11713 52503 11747
rect 52503 11713 52512 11747
rect 52460 11704 52512 11713
rect 43444 11568 43496 11620
rect 44548 11568 44600 11620
rect 44916 11636 44968 11688
rect 46848 11679 46900 11688
rect 46848 11645 46857 11679
rect 46857 11645 46891 11679
rect 46891 11645 46900 11679
rect 46848 11636 46900 11645
rect 47032 11636 47084 11688
rect 48412 11636 48464 11688
rect 50252 11679 50304 11688
rect 50252 11645 50261 11679
rect 50261 11645 50295 11679
rect 50295 11645 50304 11679
rect 50252 11636 50304 11645
rect 47492 11568 47544 11620
rect 38292 11543 38344 11552
rect 38292 11509 38301 11543
rect 38301 11509 38335 11543
rect 38335 11509 38344 11543
rect 38292 11500 38344 11509
rect 43904 11500 43956 11552
rect 48964 11568 49016 11620
rect 49424 11568 49476 11620
rect 52000 11636 52052 11688
rect 52276 11636 52328 11688
rect 55496 11747 55548 11756
rect 55496 11713 55505 11747
rect 55505 11713 55539 11747
rect 55539 11713 55548 11747
rect 55496 11704 55548 11713
rect 54116 11679 54168 11688
rect 54116 11645 54125 11679
rect 54125 11645 54159 11679
rect 54159 11645 54168 11679
rect 54116 11636 54168 11645
rect 52828 11568 52880 11620
rect 55772 11772 55824 11824
rect 55956 11815 56008 11824
rect 55956 11781 55965 11815
rect 55965 11781 55999 11815
rect 55999 11781 56008 11815
rect 55956 11772 56008 11781
rect 56232 11840 56284 11892
rect 58900 11840 58952 11892
rect 59544 11815 59596 11824
rect 59544 11781 59553 11815
rect 59553 11781 59587 11815
rect 59587 11781 59596 11815
rect 59544 11772 59596 11781
rect 56784 11704 56836 11756
rect 56140 11636 56192 11688
rect 57428 11679 57480 11688
rect 57428 11645 57437 11679
rect 57437 11645 57471 11679
rect 57471 11645 57480 11679
rect 57428 11636 57480 11645
rect 57796 11679 57848 11688
rect 57796 11645 57805 11679
rect 57805 11645 57839 11679
rect 57839 11645 57848 11679
rect 57796 11636 57848 11645
rect 58164 11679 58216 11688
rect 58164 11645 58173 11679
rect 58173 11645 58207 11679
rect 58207 11645 58216 11679
rect 58164 11636 58216 11645
rect 59728 11679 59780 11688
rect 59728 11645 59737 11679
rect 59737 11645 59771 11679
rect 59771 11645 59780 11679
rect 59728 11636 59780 11645
rect 61108 11704 61160 11756
rect 57612 11568 57664 11620
rect 59268 11568 59320 11620
rect 54852 11500 54904 11552
rect 55036 11500 55088 11552
rect 60832 11568 60884 11620
rect 60556 11543 60608 11552
rect 60556 11509 60565 11543
rect 60565 11509 60599 11543
rect 60599 11509 60608 11543
rect 60556 11500 60608 11509
rect 61108 11500 61160 11552
rect 21774 11398 21826 11450
rect 21838 11398 21890 11450
rect 21902 11398 21954 11450
rect 21966 11398 22018 11450
rect 42566 11398 42618 11450
rect 42630 11398 42682 11450
rect 42694 11398 42746 11450
rect 42758 11398 42810 11450
rect 5632 11296 5684 11348
rect 7104 11296 7156 11348
rect 8392 11339 8444 11348
rect 8392 11305 8401 11339
rect 8401 11305 8435 11339
rect 8435 11305 8444 11339
rect 8392 11296 8444 11305
rect 9772 11296 9824 11348
rect 10692 11339 10744 11348
rect 10692 11305 10701 11339
rect 10701 11305 10735 11339
rect 10735 11305 10744 11339
rect 10692 11296 10744 11305
rect 11244 11296 11296 11348
rect 14004 11296 14056 11348
rect 15108 11339 15160 11348
rect 15108 11305 15117 11339
rect 15117 11305 15151 11339
rect 15151 11305 15160 11339
rect 15108 11296 15160 11305
rect 17040 11339 17092 11348
rect 17040 11305 17049 11339
rect 17049 11305 17083 11339
rect 17083 11305 17092 11339
rect 17040 11296 17092 11305
rect 18880 11296 18932 11348
rect 8852 11271 8904 11280
rect 8852 11237 8861 11271
rect 8861 11237 8895 11271
rect 8895 11237 8904 11271
rect 8852 11228 8904 11237
rect 2872 11160 2924 11212
rect 11980 11203 12032 11212
rect 4988 11092 5040 11144
rect 5356 11092 5408 11144
rect 7196 11092 7248 11144
rect 7472 11135 7524 11144
rect 7472 11101 7478 11135
rect 7478 11101 7524 11135
rect 7472 11092 7524 11101
rect 7656 11135 7708 11144
rect 7656 11101 7665 11135
rect 7665 11101 7699 11135
rect 7699 11101 7708 11135
rect 7656 11092 7708 11101
rect 11980 11169 11989 11203
rect 11989 11169 12023 11203
rect 12023 11169 12032 11203
rect 11980 11160 12032 11169
rect 12072 11160 12124 11212
rect 12256 11160 12308 11212
rect 14924 11228 14976 11280
rect 15292 11271 15344 11280
rect 15292 11237 15301 11271
rect 15301 11237 15335 11271
rect 15335 11237 15344 11271
rect 15292 11228 15344 11237
rect 16120 11228 16172 11280
rect 16856 11228 16908 11280
rect 21180 11296 21232 11348
rect 22744 11296 22796 11348
rect 22928 11339 22980 11348
rect 22928 11305 22937 11339
rect 22937 11305 22971 11339
rect 22971 11305 22980 11339
rect 22928 11296 22980 11305
rect 23204 11296 23256 11348
rect 23480 11296 23532 11348
rect 19984 11271 20036 11280
rect 19984 11237 19993 11271
rect 19993 11237 20027 11271
rect 20027 11237 20036 11271
rect 19984 11228 20036 11237
rect 20904 11271 20956 11280
rect 20904 11237 20913 11271
rect 20913 11237 20947 11271
rect 20947 11237 20956 11271
rect 20904 11228 20956 11237
rect 23572 11228 23624 11280
rect 24768 11228 24820 11280
rect 25780 11228 25832 11280
rect 29000 11296 29052 11348
rect 29368 11296 29420 11348
rect 30748 11296 30800 11348
rect 33232 11339 33284 11348
rect 32404 11228 32456 11280
rect 14188 11160 14240 11212
rect 14280 11160 14332 11212
rect 16212 11160 16264 11212
rect 17684 11160 17736 11212
rect 17776 11160 17828 11212
rect 18696 11160 18748 11212
rect 9956 11092 10008 11144
rect 4252 10999 4304 11008
rect 4252 10965 4261 10999
rect 4261 10965 4295 10999
rect 4295 10965 4304 10999
rect 4252 10956 4304 10965
rect 7104 10999 7156 11008
rect 7104 10965 7113 10999
rect 7113 10965 7147 10999
rect 7147 10965 7156 10999
rect 7104 10956 7156 10965
rect 8300 11024 8352 11076
rect 11796 11067 11848 11076
rect 7380 10956 7432 11008
rect 8392 10956 8444 11008
rect 8760 10956 8812 11008
rect 11796 11033 11805 11067
rect 11805 11033 11839 11067
rect 11839 11033 11848 11067
rect 11796 11024 11848 11033
rect 15844 11092 15896 11144
rect 16672 11092 16724 11144
rect 17868 11135 17920 11144
rect 17592 11024 17644 11076
rect 17868 11101 17877 11135
rect 17877 11101 17911 11135
rect 17911 11101 17920 11135
rect 17868 11092 17920 11101
rect 18880 11092 18932 11144
rect 22468 11203 22520 11212
rect 22468 11169 22477 11203
rect 22477 11169 22511 11203
rect 22511 11169 22520 11203
rect 23480 11203 23532 11212
rect 22468 11160 22520 11169
rect 23480 11169 23489 11203
rect 23489 11169 23523 11203
rect 23523 11169 23532 11203
rect 23480 11160 23532 11169
rect 23664 11203 23716 11212
rect 23664 11169 23673 11203
rect 23673 11169 23707 11203
rect 23707 11169 23716 11203
rect 23664 11160 23716 11169
rect 24860 11160 24912 11212
rect 25136 11203 25188 11212
rect 25136 11169 25145 11203
rect 25145 11169 25179 11203
rect 25179 11169 25188 11203
rect 25136 11160 25188 11169
rect 26332 11160 26384 11212
rect 27160 11160 27212 11212
rect 21272 11135 21324 11144
rect 21272 11101 21281 11135
rect 21281 11101 21315 11135
rect 21315 11101 21324 11135
rect 21272 11092 21324 11101
rect 25320 11092 25372 11144
rect 25872 11092 25924 11144
rect 29460 11160 29512 11212
rect 31576 11160 31628 11212
rect 33232 11305 33241 11339
rect 33241 11305 33275 11339
rect 33275 11305 33284 11339
rect 33232 11296 33284 11305
rect 33692 11339 33744 11348
rect 33692 11305 33701 11339
rect 33701 11305 33735 11339
rect 33735 11305 33744 11339
rect 33692 11296 33744 11305
rect 35900 11296 35952 11348
rect 36084 11339 36136 11348
rect 36084 11305 36093 11339
rect 36093 11305 36127 11339
rect 36127 11305 36136 11339
rect 36084 11296 36136 11305
rect 37464 11339 37516 11348
rect 35440 11271 35492 11280
rect 35440 11237 35449 11271
rect 35449 11237 35483 11271
rect 35483 11237 35492 11271
rect 35440 11228 35492 11237
rect 32588 11160 32640 11212
rect 32864 11160 32916 11212
rect 27804 11092 27856 11144
rect 18328 11024 18380 11076
rect 19064 11067 19116 11076
rect 12808 10999 12860 11008
rect 12808 10965 12817 10999
rect 12817 10965 12851 10999
rect 12851 10965 12860 10999
rect 12808 10956 12860 10965
rect 13820 10999 13872 11008
rect 13820 10965 13844 10999
rect 13844 10965 13872 10999
rect 13820 10956 13872 10965
rect 15200 10956 15252 11008
rect 15476 10999 15528 11008
rect 15476 10965 15500 10999
rect 15500 10965 15528 10999
rect 15476 10956 15528 10965
rect 15568 10999 15620 11008
rect 15568 10965 15577 10999
rect 15577 10965 15611 10999
rect 15611 10965 15620 10999
rect 15568 10956 15620 10965
rect 16212 10956 16264 11008
rect 16304 10999 16356 11008
rect 16304 10965 16313 10999
rect 16313 10965 16347 10999
rect 16347 10965 16356 10999
rect 16304 10956 16356 10965
rect 17960 10956 18012 11008
rect 18696 10956 18748 11008
rect 19064 11033 19073 11067
rect 19073 11033 19107 11067
rect 19107 11033 19116 11067
rect 19064 11024 19116 11033
rect 19248 10956 19300 11008
rect 19524 10999 19576 11008
rect 19524 10965 19533 10999
rect 19533 10965 19567 10999
rect 19567 10965 19576 10999
rect 24952 11024 25004 11076
rect 20352 10999 20404 11008
rect 19524 10956 19576 10965
rect 20352 10965 20361 10999
rect 20361 10965 20395 10999
rect 20395 10965 20404 10999
rect 20352 10956 20404 10965
rect 20444 10956 20496 11008
rect 21732 10956 21784 11008
rect 22100 10956 22152 11008
rect 24676 10956 24728 11008
rect 25780 10956 25832 11008
rect 25964 10999 26016 11008
rect 25964 10965 25973 10999
rect 25973 10965 26007 10999
rect 26007 10965 26016 10999
rect 25964 10956 26016 10965
rect 26056 10956 26108 11008
rect 27160 10999 27212 11008
rect 27160 10965 27169 10999
rect 27169 10965 27203 10999
rect 27203 10965 27212 10999
rect 30104 11024 30156 11076
rect 31760 11024 31812 11076
rect 31944 11067 31996 11076
rect 31944 11033 31953 11067
rect 31953 11033 31987 11067
rect 31987 11033 31996 11067
rect 32772 11092 32824 11144
rect 33140 11092 33192 11144
rect 33784 11135 33836 11144
rect 33784 11101 33793 11135
rect 33793 11101 33827 11135
rect 33827 11101 33836 11135
rect 33784 11092 33836 11101
rect 34336 11160 34388 11212
rect 35348 11160 35400 11212
rect 37464 11305 37473 11339
rect 37473 11305 37507 11339
rect 37507 11305 37516 11339
rect 37464 11296 37516 11305
rect 38476 11296 38528 11348
rect 39764 11296 39816 11348
rect 39856 11296 39908 11348
rect 36820 11271 36872 11280
rect 36360 11092 36412 11144
rect 36820 11237 36829 11271
rect 36829 11237 36863 11271
rect 36863 11237 36872 11271
rect 36820 11228 36872 11237
rect 37372 11228 37424 11280
rect 40500 11228 40552 11280
rect 40592 11228 40644 11280
rect 43444 11296 43496 11348
rect 51264 11339 51316 11348
rect 38844 11160 38896 11212
rect 39396 11160 39448 11212
rect 40408 11203 40460 11212
rect 40408 11169 40417 11203
rect 40417 11169 40451 11203
rect 40451 11169 40460 11203
rect 40408 11160 40460 11169
rect 41512 11160 41564 11212
rect 41696 11160 41748 11212
rect 38292 11092 38344 11144
rect 38752 11135 38804 11144
rect 31944 11024 31996 11033
rect 32496 11024 32548 11076
rect 33600 11024 33652 11076
rect 35716 11067 35768 11076
rect 27160 10956 27212 10965
rect 30472 10956 30524 11008
rect 30932 10956 30984 11008
rect 34428 10956 34480 11008
rect 35716 11033 35725 11067
rect 35725 11033 35759 11067
rect 35759 11033 35768 11067
rect 35716 11024 35768 11033
rect 36452 11024 36504 11076
rect 38016 11024 38068 11076
rect 38752 11101 38761 11135
rect 38761 11101 38795 11135
rect 38795 11101 38804 11135
rect 38752 11092 38804 11101
rect 46664 11228 46716 11280
rect 48044 11271 48096 11280
rect 48044 11237 48053 11271
rect 48053 11237 48087 11271
rect 48087 11237 48096 11271
rect 48044 11228 48096 11237
rect 48780 11228 48832 11280
rect 50896 11271 50948 11280
rect 50896 11237 50905 11271
rect 50905 11237 50939 11271
rect 50939 11237 50948 11271
rect 50896 11228 50948 11237
rect 51264 11305 51273 11339
rect 51273 11305 51307 11339
rect 51307 11305 51316 11339
rect 51264 11296 51316 11305
rect 52552 11296 52604 11348
rect 53564 11296 53616 11348
rect 54116 11296 54168 11348
rect 55220 11296 55272 11348
rect 58072 11296 58124 11348
rect 59544 11339 59596 11348
rect 59544 11305 59553 11339
rect 59553 11305 59587 11339
rect 59587 11305 59596 11339
rect 59544 11296 59596 11305
rect 51632 11228 51684 11280
rect 52368 11228 52420 11280
rect 43352 11203 43404 11212
rect 43352 11169 43361 11203
rect 43361 11169 43395 11203
rect 43395 11169 43404 11203
rect 43352 11160 43404 11169
rect 44180 11160 44232 11212
rect 47584 11203 47636 11212
rect 37096 10999 37148 11008
rect 37096 10965 37105 10999
rect 37105 10965 37139 10999
rect 37139 10965 37148 10999
rect 37096 10956 37148 10965
rect 41880 11024 41932 11076
rect 43168 11092 43220 11144
rect 47584 11169 47593 11203
rect 47593 11169 47627 11203
rect 47627 11169 47636 11203
rect 47584 11160 47636 11169
rect 49332 11160 49384 11212
rect 52276 11160 52328 11212
rect 45376 11092 45428 11144
rect 45560 11092 45612 11144
rect 46848 11135 46900 11144
rect 46848 11101 46857 11135
rect 46857 11101 46891 11135
rect 46891 11101 46900 11135
rect 46848 11092 46900 11101
rect 47860 11092 47912 11144
rect 48504 11092 48556 11144
rect 50344 11135 50396 11144
rect 48872 11024 48924 11076
rect 42064 10956 42116 11008
rect 43904 10999 43956 11008
rect 43904 10965 43913 10999
rect 43913 10965 43947 10999
rect 43947 10965 43956 10999
rect 43904 10956 43956 10965
rect 44364 10999 44416 11008
rect 44364 10965 44373 10999
rect 44373 10965 44407 10999
rect 44407 10965 44416 10999
rect 44364 10956 44416 10965
rect 48780 10999 48832 11008
rect 48780 10965 48789 10999
rect 48789 10965 48823 10999
rect 48823 10965 48832 10999
rect 48780 10956 48832 10965
rect 50344 11101 50353 11135
rect 50353 11101 50387 11135
rect 50387 11101 50396 11135
rect 50344 11092 50396 11101
rect 51448 11092 51500 11144
rect 55036 11228 55088 11280
rect 59176 11228 59228 11280
rect 53196 11135 53248 11144
rect 53196 11101 53205 11135
rect 53205 11101 53239 11135
rect 53239 11101 53248 11135
rect 53196 11092 53248 11101
rect 53472 11092 53524 11144
rect 54944 11160 54996 11212
rect 56416 11203 56468 11212
rect 56416 11169 56425 11203
rect 56425 11169 56459 11203
rect 56459 11169 56468 11203
rect 56416 11160 56468 11169
rect 57428 11160 57480 11212
rect 58808 11160 58860 11212
rect 60464 11203 60516 11212
rect 56784 11135 56836 11144
rect 51356 11024 51408 11076
rect 56784 11101 56793 11135
rect 56793 11101 56827 11135
rect 56827 11101 56836 11135
rect 56784 11092 56836 11101
rect 57336 11092 57388 11144
rect 59176 11135 59228 11144
rect 59176 11101 59185 11135
rect 59185 11101 59219 11135
rect 59219 11101 59228 11135
rect 59176 11092 59228 11101
rect 55772 11024 55824 11076
rect 60464 11169 60473 11203
rect 60473 11169 60507 11203
rect 60507 11169 60516 11203
rect 60464 11160 60516 11169
rect 51080 10956 51132 11008
rect 51724 10999 51776 11008
rect 51724 10965 51733 10999
rect 51733 10965 51767 10999
rect 51767 10965 51776 10999
rect 51724 10956 51776 10965
rect 55956 10999 56008 11008
rect 55956 10965 55965 10999
rect 55965 10965 55999 10999
rect 55999 10965 56008 10999
rect 55956 10956 56008 10965
rect 56600 10999 56652 11008
rect 56600 10965 56624 10999
rect 56624 10965 56652 10999
rect 56600 10956 56652 10965
rect 56692 10999 56744 11008
rect 56692 10965 56701 10999
rect 56701 10965 56735 10999
rect 56735 10965 56744 10999
rect 56692 10956 56744 10965
rect 57244 10956 57296 11008
rect 59268 10956 59320 11008
rect 11378 10854 11430 10906
rect 11442 10854 11494 10906
rect 11506 10854 11558 10906
rect 11570 10854 11622 10906
rect 32170 10854 32222 10906
rect 32234 10854 32286 10906
rect 32298 10854 32350 10906
rect 32362 10854 32414 10906
rect 52962 10854 53014 10906
rect 53026 10854 53078 10906
rect 53090 10854 53142 10906
rect 53154 10854 53206 10906
rect 5264 10752 5316 10804
rect 5448 10752 5500 10804
rect 7656 10752 7708 10804
rect 8300 10752 8352 10804
rect 8668 10752 8720 10804
rect 9956 10795 10008 10804
rect 9956 10761 9965 10795
rect 9965 10761 9999 10795
rect 9999 10761 10008 10795
rect 9956 10752 10008 10761
rect 11888 10752 11940 10804
rect 7288 10684 7340 10736
rect 9772 10684 9824 10736
rect 10692 10684 10744 10736
rect 12072 10684 12124 10736
rect 12624 10752 12676 10804
rect 14188 10752 14240 10804
rect 15292 10752 15344 10804
rect 18328 10752 18380 10804
rect 15844 10727 15896 10736
rect 15844 10693 15853 10727
rect 15853 10693 15887 10727
rect 15887 10693 15896 10727
rect 15844 10684 15896 10693
rect 16212 10727 16264 10736
rect 16212 10693 16221 10727
rect 16221 10693 16255 10727
rect 16255 10693 16264 10727
rect 16212 10684 16264 10693
rect 17868 10684 17920 10736
rect 19156 10752 19208 10804
rect 21272 10752 21324 10804
rect 21732 10752 21784 10804
rect 22284 10752 22336 10804
rect 30104 10752 30156 10804
rect 30196 10795 30248 10804
rect 30196 10761 30205 10795
rect 30205 10761 30239 10795
rect 30239 10761 30248 10795
rect 30472 10795 30524 10804
rect 30196 10752 30248 10761
rect 30472 10761 30481 10795
rect 30481 10761 30515 10795
rect 30515 10761 30524 10795
rect 30472 10752 30524 10761
rect 31208 10752 31260 10804
rect 34520 10752 34572 10804
rect 36360 10795 36412 10804
rect 36360 10761 36369 10795
rect 36369 10761 36403 10795
rect 36403 10761 36412 10795
rect 36360 10752 36412 10761
rect 36636 10752 36688 10804
rect 37924 10752 37976 10804
rect 38568 10752 38620 10804
rect 44548 10795 44600 10804
rect 4252 10591 4304 10600
rect 4252 10557 4261 10591
rect 4261 10557 4295 10591
rect 4295 10557 4304 10591
rect 4252 10548 4304 10557
rect 7380 10548 7432 10600
rect 12808 10616 12860 10668
rect 12900 10616 12952 10668
rect 14280 10616 14332 10668
rect 14924 10659 14976 10668
rect 14924 10625 14933 10659
rect 14933 10625 14967 10659
rect 14967 10625 14976 10659
rect 14924 10616 14976 10625
rect 18604 10659 18656 10668
rect 7104 10480 7156 10532
rect 7840 10548 7892 10600
rect 8668 10591 8720 10600
rect 8668 10557 8677 10591
rect 8677 10557 8711 10591
rect 8711 10557 8720 10591
rect 8668 10548 8720 10557
rect 4988 10412 5040 10464
rect 6368 10412 6420 10464
rect 7472 10412 7524 10464
rect 9772 10412 9824 10464
rect 13452 10548 13504 10600
rect 15108 10548 15160 10600
rect 15200 10480 15252 10532
rect 15568 10480 15620 10532
rect 18604 10625 18613 10659
rect 18613 10625 18647 10659
rect 18647 10625 18656 10659
rect 18604 10616 18656 10625
rect 19616 10684 19668 10736
rect 20720 10684 20772 10736
rect 22928 10727 22980 10736
rect 19616 10591 19668 10600
rect 19616 10557 19625 10591
rect 19625 10557 19659 10591
rect 19659 10557 19668 10591
rect 19616 10548 19668 10557
rect 20352 10548 20404 10600
rect 18236 10480 18288 10532
rect 18788 10480 18840 10532
rect 18972 10523 19024 10532
rect 18972 10489 18981 10523
rect 18981 10489 19015 10523
rect 19015 10489 19024 10523
rect 18972 10480 19024 10489
rect 22928 10693 22937 10727
rect 22937 10693 22971 10727
rect 22971 10693 22980 10727
rect 22928 10684 22980 10693
rect 23480 10727 23532 10736
rect 23480 10693 23489 10727
rect 23489 10693 23523 10727
rect 23523 10693 23532 10727
rect 23480 10684 23532 10693
rect 25044 10684 25096 10736
rect 22652 10659 22704 10668
rect 22652 10625 22661 10659
rect 22661 10625 22695 10659
rect 22695 10625 22704 10659
rect 22652 10616 22704 10625
rect 23204 10548 23256 10600
rect 24676 10548 24728 10600
rect 22100 10523 22152 10532
rect 22100 10489 22109 10523
rect 22109 10489 22143 10523
rect 22143 10489 22152 10523
rect 22100 10480 22152 10489
rect 17408 10455 17460 10464
rect 17408 10421 17417 10455
rect 17417 10421 17451 10455
rect 17451 10421 17460 10455
rect 17408 10412 17460 10421
rect 17776 10412 17828 10464
rect 24952 10591 25004 10600
rect 24952 10557 24961 10591
rect 24961 10557 24995 10591
rect 24995 10557 25004 10591
rect 27804 10616 27856 10668
rect 24952 10548 25004 10557
rect 25596 10548 25648 10600
rect 25780 10548 25832 10600
rect 27160 10591 27212 10600
rect 26148 10523 26200 10532
rect 26148 10489 26157 10523
rect 26157 10489 26191 10523
rect 26191 10489 26200 10523
rect 27160 10557 27169 10591
rect 27169 10557 27203 10591
rect 27203 10557 27212 10591
rect 27160 10548 27212 10557
rect 27252 10548 27304 10600
rect 27528 10548 27580 10600
rect 29092 10616 29144 10668
rect 33784 10684 33836 10736
rect 29368 10591 29420 10600
rect 29368 10557 29377 10591
rect 29377 10557 29411 10591
rect 29411 10557 29420 10591
rect 29368 10548 29420 10557
rect 26148 10480 26200 10489
rect 27620 10480 27672 10532
rect 28264 10480 28316 10532
rect 30932 10548 30984 10600
rect 32312 10591 32364 10600
rect 35992 10616 36044 10668
rect 39028 10684 39080 10736
rect 40500 10684 40552 10736
rect 43168 10727 43220 10736
rect 43168 10693 43177 10727
rect 43177 10693 43211 10727
rect 43211 10693 43220 10727
rect 43168 10684 43220 10693
rect 43352 10684 43404 10736
rect 44548 10761 44557 10795
rect 44557 10761 44591 10795
rect 44591 10761 44600 10795
rect 44548 10752 44600 10761
rect 45100 10752 45152 10804
rect 46664 10752 46716 10804
rect 47584 10752 47636 10804
rect 47860 10795 47912 10804
rect 47860 10761 47869 10795
rect 47869 10761 47903 10795
rect 47903 10761 47912 10795
rect 47860 10752 47912 10761
rect 48228 10752 48280 10804
rect 51448 10795 51500 10804
rect 51448 10761 51457 10795
rect 51457 10761 51491 10795
rect 51491 10761 51500 10795
rect 51448 10752 51500 10761
rect 54944 10752 54996 10804
rect 56140 10795 56192 10804
rect 36452 10659 36504 10668
rect 36452 10625 36461 10659
rect 36461 10625 36495 10659
rect 36495 10625 36504 10659
rect 36452 10616 36504 10625
rect 36728 10659 36780 10668
rect 36728 10625 36737 10659
rect 36737 10625 36771 10659
rect 36771 10625 36780 10659
rect 36728 10616 36780 10625
rect 37096 10616 37148 10668
rect 39396 10659 39448 10668
rect 32312 10557 32328 10591
rect 32328 10557 32362 10591
rect 32362 10557 32364 10591
rect 32312 10548 32364 10557
rect 33692 10548 33744 10600
rect 34152 10548 34204 10600
rect 34704 10548 34756 10600
rect 27068 10412 27120 10464
rect 27160 10412 27212 10464
rect 32036 10480 32088 10532
rect 35072 10523 35124 10532
rect 28908 10412 28960 10464
rect 30840 10455 30892 10464
rect 30840 10421 30849 10455
rect 30849 10421 30883 10455
rect 30883 10421 30892 10455
rect 30840 10412 30892 10421
rect 31576 10412 31628 10464
rect 35072 10489 35081 10523
rect 35081 10489 35115 10523
rect 35115 10489 35124 10523
rect 35072 10480 35124 10489
rect 35808 10480 35860 10532
rect 38292 10548 38344 10600
rect 38844 10548 38896 10600
rect 39028 10548 39080 10600
rect 39396 10625 39405 10659
rect 39405 10625 39439 10659
rect 39439 10625 39448 10659
rect 39396 10616 39448 10625
rect 41696 10616 41748 10668
rect 42064 10659 42116 10668
rect 42064 10625 42073 10659
rect 42073 10625 42107 10659
rect 42107 10625 42116 10659
rect 42064 10616 42116 10625
rect 44916 10616 44968 10668
rect 40684 10591 40736 10600
rect 40684 10557 40693 10591
rect 40693 10557 40727 10591
rect 40727 10557 40736 10591
rect 40684 10548 40736 10557
rect 42984 10548 43036 10600
rect 44364 10591 44416 10600
rect 44364 10557 44373 10591
rect 44373 10557 44407 10591
rect 44407 10557 44416 10591
rect 44364 10548 44416 10557
rect 47952 10684 48004 10736
rect 48320 10727 48372 10736
rect 48320 10693 48329 10727
rect 48329 10693 48363 10727
rect 48363 10693 48372 10727
rect 48320 10684 48372 10693
rect 46940 10616 46992 10668
rect 51356 10684 51408 10736
rect 51908 10727 51960 10736
rect 51908 10693 51917 10727
rect 51917 10693 51951 10727
rect 51951 10693 51960 10727
rect 51908 10684 51960 10693
rect 56140 10761 56149 10795
rect 56149 10761 56183 10795
rect 56183 10761 56192 10795
rect 56140 10752 56192 10761
rect 56784 10795 56836 10804
rect 56784 10761 56793 10795
rect 56793 10761 56827 10795
rect 56827 10761 56836 10795
rect 56784 10752 56836 10761
rect 57612 10795 57664 10804
rect 57612 10761 57621 10795
rect 57621 10761 57655 10795
rect 57655 10761 57664 10795
rect 57612 10752 57664 10761
rect 60464 10752 60516 10804
rect 60832 10727 60884 10736
rect 49332 10659 49384 10668
rect 49332 10625 49341 10659
rect 49341 10625 49375 10659
rect 49375 10625 49384 10659
rect 49332 10616 49384 10625
rect 34336 10455 34388 10464
rect 34336 10421 34345 10455
rect 34345 10421 34379 10455
rect 34379 10421 34388 10455
rect 34336 10412 34388 10421
rect 36820 10412 36872 10464
rect 37924 10412 37976 10464
rect 38660 10480 38712 10532
rect 48596 10548 48648 10600
rect 48780 10548 48832 10600
rect 48872 10591 48924 10600
rect 48872 10557 48881 10591
rect 48881 10557 48915 10591
rect 48915 10557 48924 10591
rect 48872 10548 48924 10557
rect 49424 10548 49476 10600
rect 50344 10616 50396 10668
rect 51816 10616 51868 10668
rect 53932 10616 53984 10668
rect 57336 10659 57388 10668
rect 57336 10625 57345 10659
rect 57345 10625 57379 10659
rect 57379 10625 57388 10659
rect 57336 10616 57388 10625
rect 38752 10455 38804 10464
rect 38752 10421 38761 10455
rect 38761 10421 38795 10455
rect 38795 10421 38804 10455
rect 38752 10412 38804 10421
rect 38936 10412 38988 10464
rect 40868 10455 40920 10464
rect 40868 10421 40877 10455
rect 40877 10421 40911 10455
rect 40911 10421 40920 10455
rect 40868 10412 40920 10421
rect 43536 10412 43588 10464
rect 43904 10412 43956 10464
rect 44088 10455 44140 10464
rect 44088 10421 44097 10455
rect 44097 10421 44131 10455
rect 44131 10421 44140 10455
rect 44088 10412 44140 10421
rect 45468 10455 45520 10464
rect 45468 10421 45477 10455
rect 45477 10421 45511 10455
rect 45511 10421 45520 10455
rect 45468 10412 45520 10421
rect 45836 10455 45888 10464
rect 45836 10421 45845 10455
rect 45845 10421 45879 10455
rect 45879 10421 45888 10455
rect 45836 10412 45888 10421
rect 47400 10455 47452 10464
rect 47400 10421 47409 10455
rect 47409 10421 47443 10455
rect 47443 10421 47452 10455
rect 47400 10412 47452 10421
rect 47584 10412 47636 10464
rect 49608 10480 49660 10532
rect 47952 10412 48004 10464
rect 49516 10412 49568 10464
rect 51724 10591 51776 10600
rect 51724 10557 51733 10591
rect 51733 10557 51767 10591
rect 51767 10557 51776 10591
rect 51724 10548 51776 10557
rect 54484 10548 54536 10600
rect 55496 10548 55548 10600
rect 55956 10591 56008 10600
rect 55956 10557 55965 10591
rect 55965 10557 55999 10591
rect 55999 10557 56008 10591
rect 60832 10693 60841 10727
rect 60841 10693 60875 10727
rect 60875 10693 60884 10727
rect 60832 10684 60884 10693
rect 59544 10659 59596 10668
rect 59544 10625 59553 10659
rect 59553 10625 59587 10659
rect 59587 10625 59596 10659
rect 59544 10616 59596 10625
rect 55956 10548 56008 10557
rect 58348 10548 58400 10600
rect 59268 10591 59320 10600
rect 59268 10557 59277 10591
rect 59277 10557 59311 10591
rect 59311 10557 59320 10591
rect 59268 10548 59320 10557
rect 51172 10412 51224 10464
rect 52276 10455 52328 10464
rect 52276 10421 52285 10455
rect 52285 10421 52319 10455
rect 52319 10421 52328 10455
rect 52276 10412 52328 10421
rect 52828 10455 52880 10464
rect 52828 10421 52837 10455
rect 52837 10421 52871 10455
rect 52871 10421 52880 10455
rect 55404 10480 55456 10532
rect 56508 10480 56560 10532
rect 54392 10455 54444 10464
rect 52828 10412 52880 10421
rect 54392 10421 54401 10455
rect 54401 10421 54435 10455
rect 54435 10421 54444 10455
rect 54392 10412 54444 10421
rect 56600 10412 56652 10464
rect 58808 10455 58860 10464
rect 58808 10421 58817 10455
rect 58817 10421 58851 10455
rect 58851 10421 58860 10455
rect 58808 10412 58860 10421
rect 59084 10455 59136 10464
rect 59084 10421 59093 10455
rect 59093 10421 59127 10455
rect 59127 10421 59136 10455
rect 59084 10412 59136 10421
rect 61292 10412 61344 10464
rect 21774 10310 21826 10362
rect 21838 10310 21890 10362
rect 21902 10310 21954 10362
rect 21966 10310 22018 10362
rect 42566 10310 42618 10362
rect 42630 10310 42682 10362
rect 42694 10310 42746 10362
rect 42758 10310 42810 10362
rect 5448 10208 5500 10260
rect 8852 10208 8904 10260
rect 13820 10251 13872 10260
rect 13820 10217 13829 10251
rect 13829 10217 13863 10251
rect 13863 10217 13872 10251
rect 13820 10208 13872 10217
rect 14188 10251 14240 10260
rect 14188 10217 14197 10251
rect 14197 10217 14231 10251
rect 14231 10217 14240 10251
rect 14188 10208 14240 10217
rect 14924 10251 14976 10260
rect 14924 10217 14933 10251
rect 14933 10217 14967 10251
rect 14967 10217 14976 10251
rect 14924 10208 14976 10217
rect 15476 10208 15528 10260
rect 16396 10208 16448 10260
rect 20076 10208 20128 10260
rect 20444 10208 20496 10260
rect 21180 10208 21232 10260
rect 7472 10140 7524 10192
rect 15108 10140 15160 10192
rect 4252 10072 4304 10124
rect 4804 10072 4856 10124
rect 4988 10072 5040 10124
rect 9772 10115 9824 10124
rect 4712 10047 4764 10056
rect 4712 10013 4721 10047
rect 4721 10013 4755 10047
rect 4755 10013 4764 10047
rect 4712 10004 4764 10013
rect 5724 10004 5776 10056
rect 7288 10004 7340 10056
rect 9772 10081 9781 10115
rect 9781 10081 9815 10115
rect 9815 10081 9824 10115
rect 9772 10072 9824 10081
rect 10876 10072 10928 10124
rect 11796 10072 11848 10124
rect 14372 10072 14424 10124
rect 16028 10072 16080 10124
rect 17408 10072 17460 10124
rect 17776 10072 17828 10124
rect 7840 10047 7892 10056
rect 7840 10013 7849 10047
rect 7849 10013 7883 10047
rect 7883 10013 7892 10047
rect 7840 10004 7892 10013
rect 9680 10047 9732 10056
rect 8944 9936 8996 9988
rect 9680 10013 9689 10047
rect 9689 10013 9723 10047
rect 9723 10013 9732 10047
rect 9680 10004 9732 10013
rect 9956 10004 10008 10056
rect 12072 10004 12124 10056
rect 12716 10004 12768 10056
rect 13728 10004 13780 10056
rect 10692 9936 10744 9988
rect 15568 9936 15620 9988
rect 17960 10004 18012 10056
rect 18236 10140 18288 10192
rect 18328 10115 18380 10124
rect 18328 10081 18337 10115
rect 18337 10081 18371 10115
rect 18371 10081 18380 10115
rect 18328 10072 18380 10081
rect 20352 10140 20404 10192
rect 23020 10208 23072 10260
rect 24216 10208 24268 10260
rect 24860 10251 24912 10260
rect 24860 10217 24869 10251
rect 24869 10217 24903 10251
rect 24903 10217 24912 10251
rect 24860 10208 24912 10217
rect 26332 10251 26384 10260
rect 26332 10217 26341 10251
rect 26341 10217 26375 10251
rect 26375 10217 26384 10251
rect 26332 10208 26384 10217
rect 27620 10208 27672 10260
rect 27712 10208 27764 10260
rect 30840 10208 30892 10260
rect 32588 10251 32640 10260
rect 32588 10217 32597 10251
rect 32597 10217 32631 10251
rect 32631 10217 32640 10251
rect 32588 10208 32640 10217
rect 35072 10208 35124 10260
rect 20812 10072 20864 10124
rect 20996 10004 21048 10056
rect 22100 10072 22152 10124
rect 23204 10072 23256 10124
rect 26056 10140 26108 10192
rect 27896 10140 27948 10192
rect 29184 10183 29236 10192
rect 27436 10072 27488 10124
rect 22192 10047 22244 10056
rect 22192 10013 22201 10047
rect 22201 10013 22235 10047
rect 22235 10013 22244 10047
rect 22192 10004 22244 10013
rect 27252 10047 27304 10056
rect 27252 10013 27261 10047
rect 27261 10013 27295 10047
rect 27295 10013 27304 10047
rect 27252 10004 27304 10013
rect 17592 9936 17644 9988
rect 4160 9868 4212 9920
rect 6368 9911 6420 9920
rect 6368 9877 6377 9911
rect 6377 9877 6411 9911
rect 6411 9877 6420 9911
rect 6368 9868 6420 9877
rect 9312 9868 9364 9920
rect 10508 9911 10560 9920
rect 10508 9877 10517 9911
rect 10517 9877 10551 9911
rect 10551 9877 10560 9911
rect 10508 9868 10560 9877
rect 10876 9868 10928 9920
rect 12900 9868 12952 9920
rect 15200 9868 15252 9920
rect 16304 9911 16356 9920
rect 16304 9877 16313 9911
rect 16313 9877 16347 9911
rect 16347 9877 16356 9911
rect 16304 9868 16356 9877
rect 16672 9911 16724 9920
rect 16672 9877 16681 9911
rect 16681 9877 16715 9911
rect 16715 9877 16724 9911
rect 16672 9868 16724 9877
rect 17776 9911 17828 9920
rect 17776 9877 17785 9911
rect 17785 9877 17819 9911
rect 17819 9877 17828 9911
rect 17776 9868 17828 9877
rect 18052 9868 18104 9920
rect 21180 9936 21232 9988
rect 22468 9936 22520 9988
rect 26332 9936 26384 9988
rect 19340 9868 19392 9920
rect 19708 9911 19760 9920
rect 19708 9877 19717 9911
rect 19717 9877 19751 9911
rect 19751 9877 19760 9911
rect 19708 9868 19760 9877
rect 20720 9911 20772 9920
rect 20720 9877 20729 9911
rect 20729 9877 20763 9911
rect 20763 9877 20772 9911
rect 20720 9868 20772 9877
rect 21364 9868 21416 9920
rect 21732 9868 21784 9920
rect 23940 9868 23992 9920
rect 25320 9911 25372 9920
rect 25320 9877 25329 9911
rect 25329 9877 25363 9911
rect 25363 9877 25372 9911
rect 25320 9868 25372 9877
rect 25596 9868 25648 9920
rect 27528 9868 27580 9920
rect 28356 9868 28408 9920
rect 29184 10149 29193 10183
rect 29193 10149 29227 10183
rect 29227 10149 29236 10183
rect 29184 10140 29236 10149
rect 34336 10140 34388 10192
rect 30288 10072 30340 10124
rect 31576 10004 31628 10056
rect 28724 9936 28776 9988
rect 33232 10072 33284 10124
rect 36084 10115 36136 10124
rect 36084 10081 36093 10115
rect 36093 10081 36127 10115
rect 36127 10081 36136 10115
rect 36084 10072 36136 10081
rect 38660 10115 38712 10124
rect 32312 10004 32364 10056
rect 33140 10047 33192 10056
rect 33140 10013 33149 10047
rect 33149 10013 33183 10047
rect 33183 10013 33192 10047
rect 33140 10004 33192 10013
rect 33508 10004 33560 10056
rect 35440 10004 35492 10056
rect 38660 10081 38669 10115
rect 38669 10081 38703 10115
rect 38703 10081 38712 10115
rect 38660 10072 38712 10081
rect 38936 10140 38988 10192
rect 39856 10183 39908 10192
rect 39856 10149 39865 10183
rect 39865 10149 39899 10183
rect 39899 10149 39908 10183
rect 39856 10140 39908 10149
rect 39028 10115 39080 10124
rect 39028 10081 39037 10115
rect 39037 10081 39071 10115
rect 39071 10081 39080 10115
rect 39028 10072 39080 10081
rect 36544 10047 36596 10056
rect 36544 10013 36553 10047
rect 36553 10013 36587 10047
rect 36587 10013 36596 10047
rect 36544 10004 36596 10013
rect 36820 10004 36872 10056
rect 41604 10140 41656 10192
rect 41972 10140 42024 10192
rect 45836 10208 45888 10260
rect 47308 10208 47360 10260
rect 47768 10208 47820 10260
rect 48320 10251 48372 10260
rect 48320 10217 48329 10251
rect 48329 10217 48363 10251
rect 48363 10217 48372 10251
rect 48320 10208 48372 10217
rect 49608 10208 49660 10260
rect 50436 10208 50488 10260
rect 51080 10208 51132 10260
rect 52000 10208 52052 10260
rect 53932 10251 53984 10260
rect 53932 10217 53941 10251
rect 53941 10217 53975 10251
rect 53975 10217 53984 10251
rect 53932 10208 53984 10217
rect 54484 10208 54536 10260
rect 54944 10208 54996 10260
rect 55772 10251 55824 10260
rect 55772 10217 55781 10251
rect 55781 10217 55815 10251
rect 55815 10217 55824 10251
rect 55772 10208 55824 10217
rect 46020 10183 46072 10192
rect 40316 10047 40368 10056
rect 40316 10013 40325 10047
rect 40325 10013 40359 10047
rect 40359 10013 40368 10047
rect 40316 10004 40368 10013
rect 41788 10115 41840 10124
rect 41788 10081 41797 10115
rect 41797 10081 41831 10115
rect 41831 10081 41840 10115
rect 41788 10072 41840 10081
rect 43904 10072 43956 10124
rect 44824 10115 44876 10124
rect 44824 10081 44833 10115
rect 44833 10081 44867 10115
rect 44867 10081 44876 10115
rect 44824 10072 44876 10081
rect 46020 10149 46029 10183
rect 46029 10149 46063 10183
rect 46063 10149 46072 10183
rect 46020 10140 46072 10149
rect 47400 10140 47452 10192
rect 45560 10072 45612 10124
rect 46664 10115 46716 10124
rect 46664 10081 46673 10115
rect 46673 10081 46707 10115
rect 46707 10081 46716 10115
rect 46664 10072 46716 10081
rect 41052 10004 41104 10056
rect 45284 10047 45336 10056
rect 32956 9936 33008 9988
rect 38752 9936 38804 9988
rect 41420 9936 41472 9988
rect 45284 10013 45293 10047
rect 45293 10013 45327 10047
rect 45327 10013 45336 10047
rect 45284 10004 45336 10013
rect 47584 10072 47636 10124
rect 47768 10115 47820 10124
rect 47768 10081 47777 10115
rect 47777 10081 47811 10115
rect 47811 10081 47820 10115
rect 47768 10072 47820 10081
rect 47860 10072 47912 10124
rect 48688 10072 48740 10124
rect 49332 10072 49384 10124
rect 29092 9868 29144 9920
rect 30104 9868 30156 9920
rect 30288 9868 30340 9920
rect 31208 9868 31260 9920
rect 31760 9911 31812 9920
rect 31760 9877 31769 9911
rect 31769 9877 31803 9911
rect 31803 9877 31812 9911
rect 31760 9868 31812 9877
rect 33876 9868 33928 9920
rect 34336 9868 34388 9920
rect 35532 9868 35584 9920
rect 36176 9868 36228 9920
rect 36912 9911 36964 9920
rect 36912 9877 36921 9911
rect 36921 9877 36955 9911
rect 36955 9877 36964 9911
rect 36912 9868 36964 9877
rect 37924 9911 37976 9920
rect 37924 9877 37933 9911
rect 37933 9877 37967 9911
rect 37967 9877 37976 9911
rect 37924 9868 37976 9877
rect 41512 9911 41564 9920
rect 41512 9877 41521 9911
rect 41521 9877 41555 9911
rect 41555 9877 41564 9911
rect 41512 9868 41564 9877
rect 42892 9911 42944 9920
rect 42892 9877 42901 9911
rect 42901 9877 42935 9911
rect 42935 9877 42944 9911
rect 42892 9868 42944 9877
rect 43076 9868 43128 9920
rect 43536 9911 43588 9920
rect 43536 9877 43545 9911
rect 43545 9877 43579 9911
rect 43579 9877 43588 9911
rect 43536 9868 43588 9877
rect 43904 9911 43956 9920
rect 43904 9877 43913 9911
rect 43913 9877 43947 9911
rect 43947 9877 43956 9911
rect 43904 9868 43956 9877
rect 45468 9936 45520 9988
rect 47216 10004 47268 10056
rect 47124 9936 47176 9988
rect 51540 10140 51592 10192
rect 51264 10115 51316 10124
rect 51264 10081 51273 10115
rect 51273 10081 51307 10115
rect 51307 10081 51316 10115
rect 51264 10072 51316 10081
rect 52736 10072 52788 10124
rect 51540 10004 51592 10056
rect 51632 10004 51684 10056
rect 53564 10072 53616 10124
rect 55404 10140 55456 10192
rect 56416 10208 56468 10260
rect 57244 10251 57296 10260
rect 57244 10217 57253 10251
rect 57253 10217 57287 10251
rect 57287 10217 57296 10251
rect 57244 10208 57296 10217
rect 57336 10208 57388 10260
rect 61844 10208 61896 10260
rect 53840 10004 53892 10056
rect 46480 9911 46532 9920
rect 46480 9877 46489 9911
rect 46489 9877 46523 9911
rect 46523 9877 46532 9911
rect 47216 9911 47268 9920
rect 46480 9868 46532 9877
rect 47216 9877 47225 9911
rect 47225 9877 47259 9911
rect 47259 9877 47268 9911
rect 47216 9868 47268 9877
rect 48412 9868 48464 9920
rect 48688 9911 48740 9920
rect 48688 9877 48697 9911
rect 48697 9877 48731 9911
rect 48731 9877 48740 9911
rect 48688 9868 48740 9877
rect 52828 9979 52880 9988
rect 52828 9945 52837 9979
rect 52837 9945 52871 9979
rect 52871 9945 52880 9979
rect 52828 9936 52880 9945
rect 49608 9868 49660 9920
rect 50252 9868 50304 9920
rect 51816 9868 51868 9920
rect 56508 10115 56560 10124
rect 56508 10081 56517 10115
rect 56517 10081 56551 10115
rect 56551 10081 56560 10115
rect 56508 10072 56560 10081
rect 58440 10115 58492 10124
rect 58440 10081 58449 10115
rect 58449 10081 58483 10115
rect 58483 10081 58492 10115
rect 58440 10072 58492 10081
rect 54760 10004 54812 10056
rect 56416 10047 56468 10056
rect 56416 10013 56425 10047
rect 56425 10013 56459 10047
rect 56459 10013 56468 10047
rect 56416 10004 56468 10013
rect 57796 10004 57848 10056
rect 59084 9936 59136 9988
rect 55220 9911 55272 9920
rect 55220 9877 55229 9911
rect 55229 9877 55263 9911
rect 55263 9877 55272 9911
rect 55220 9868 55272 9877
rect 56600 9868 56652 9920
rect 58164 9868 58216 9920
rect 59452 9868 59504 9920
rect 61292 10072 61344 10124
rect 60464 10047 60516 10056
rect 60464 10013 60473 10047
rect 60473 10013 60507 10047
rect 60507 10013 60516 10047
rect 60464 10004 60516 10013
rect 59820 9868 59872 9920
rect 61844 9868 61896 9920
rect 11378 9766 11430 9818
rect 11442 9766 11494 9818
rect 11506 9766 11558 9818
rect 11570 9766 11622 9818
rect 32170 9766 32222 9818
rect 32234 9766 32286 9818
rect 32298 9766 32350 9818
rect 32362 9766 32414 9818
rect 52962 9766 53014 9818
rect 53026 9766 53078 9818
rect 53090 9766 53142 9818
rect 53154 9766 53206 9818
rect 4804 9664 4856 9716
rect 6368 9664 6420 9716
rect 2964 9639 3016 9648
rect 2964 9605 2973 9639
rect 2973 9605 3007 9639
rect 3007 9605 3016 9639
rect 2964 9596 3016 9605
rect 5356 9596 5408 9648
rect 4252 9528 4304 9580
rect 9956 9664 10008 9716
rect 11796 9707 11848 9716
rect 11796 9673 11805 9707
rect 11805 9673 11839 9707
rect 11839 9673 11848 9707
rect 11796 9664 11848 9673
rect 12256 9707 12308 9716
rect 12256 9673 12265 9707
rect 12265 9673 12299 9707
rect 12299 9673 12308 9707
rect 12256 9664 12308 9673
rect 14280 9664 14332 9716
rect 16028 9707 16080 9716
rect 9680 9596 9732 9648
rect 12808 9596 12860 9648
rect 13544 9596 13596 9648
rect 16028 9673 16037 9707
rect 16037 9673 16071 9707
rect 16071 9673 16080 9707
rect 16028 9664 16080 9673
rect 17960 9664 18012 9716
rect 10508 9528 10560 9580
rect 12164 9528 12216 9580
rect 12624 9528 12676 9580
rect 4160 9503 4212 9512
rect 4160 9469 4169 9503
rect 4169 9469 4203 9503
rect 4203 9469 4212 9503
rect 4160 9460 4212 9469
rect 7104 9503 7156 9512
rect 7104 9469 7113 9503
rect 7113 9469 7147 9503
rect 7147 9469 7156 9503
rect 7104 9460 7156 9469
rect 9312 9503 9364 9512
rect 9312 9469 9321 9503
rect 9321 9469 9355 9503
rect 9355 9469 9364 9503
rect 9312 9460 9364 9469
rect 9864 9435 9916 9444
rect 9864 9401 9873 9435
rect 9873 9401 9907 9435
rect 9907 9401 9916 9435
rect 9864 9392 9916 9401
rect 10692 9460 10744 9512
rect 12900 9503 12952 9512
rect 10876 9392 10928 9444
rect 12900 9469 12909 9503
rect 12909 9469 12943 9503
rect 12943 9469 12952 9503
rect 12900 9460 12952 9469
rect 18328 9596 18380 9648
rect 18788 9664 18840 9716
rect 20812 9664 20864 9716
rect 23204 9707 23256 9716
rect 23204 9673 23213 9707
rect 23213 9673 23247 9707
rect 23247 9673 23256 9707
rect 23204 9664 23256 9673
rect 27436 9707 27488 9716
rect 27436 9673 27445 9707
rect 27445 9673 27479 9707
rect 27479 9673 27488 9707
rect 27436 9664 27488 9673
rect 27620 9664 27672 9716
rect 19156 9596 19208 9648
rect 19800 9639 19852 9648
rect 19800 9605 19809 9639
rect 19809 9605 19843 9639
rect 19843 9605 19852 9639
rect 19800 9596 19852 9605
rect 16396 9528 16448 9580
rect 14280 9460 14332 9512
rect 14740 9460 14792 9512
rect 15200 9460 15252 9512
rect 16028 9460 16080 9512
rect 16672 9503 16724 9512
rect 16672 9469 16681 9503
rect 16681 9469 16715 9503
rect 16715 9469 16724 9503
rect 16672 9460 16724 9469
rect 16948 9528 17000 9580
rect 18512 9528 18564 9580
rect 19064 9528 19116 9580
rect 19248 9528 19300 9580
rect 20720 9528 20772 9580
rect 21916 9571 21968 9580
rect 18052 9460 18104 9512
rect 18236 9503 18288 9512
rect 18236 9469 18245 9503
rect 18245 9469 18279 9503
rect 18279 9469 18288 9503
rect 19984 9503 20036 9512
rect 18236 9460 18288 9469
rect 19984 9469 19993 9503
rect 19993 9469 20027 9503
rect 20027 9469 20036 9503
rect 19984 9460 20036 9469
rect 17224 9392 17276 9444
rect 18696 9392 18748 9444
rect 19248 9392 19300 9444
rect 21088 9460 21140 9512
rect 20260 9392 20312 9444
rect 20812 9435 20864 9444
rect 20812 9401 20821 9435
rect 20821 9401 20855 9435
rect 20855 9401 20864 9435
rect 20812 9392 20864 9401
rect 3056 9324 3108 9376
rect 8944 9324 8996 9376
rect 10692 9324 10744 9376
rect 11060 9324 11112 9376
rect 17592 9324 17644 9376
rect 18144 9324 18196 9376
rect 21088 9324 21140 9376
rect 21272 9367 21324 9376
rect 21272 9333 21281 9367
rect 21281 9333 21315 9367
rect 21315 9333 21324 9367
rect 21272 9324 21324 9333
rect 21916 9537 21925 9571
rect 21925 9537 21959 9571
rect 21959 9537 21968 9571
rect 21916 9528 21968 9537
rect 23388 9596 23440 9648
rect 23112 9460 23164 9512
rect 25044 9596 25096 9648
rect 26792 9596 26844 9648
rect 27252 9596 27304 9648
rect 28908 9664 28960 9716
rect 35900 9664 35952 9716
rect 36544 9664 36596 9716
rect 37096 9664 37148 9716
rect 26148 9528 26200 9580
rect 27068 9528 27120 9580
rect 30288 9596 30340 9648
rect 31944 9596 31996 9648
rect 34336 9596 34388 9648
rect 36728 9639 36780 9648
rect 36728 9605 36737 9639
rect 36737 9605 36771 9639
rect 36771 9605 36780 9639
rect 36728 9596 36780 9605
rect 37832 9596 37884 9648
rect 38476 9639 38528 9648
rect 38476 9605 38485 9639
rect 38485 9605 38519 9639
rect 38519 9605 38528 9639
rect 38476 9596 38528 9605
rect 39028 9664 39080 9716
rect 41604 9664 41656 9716
rect 38844 9596 38896 9648
rect 38936 9596 38988 9648
rect 27988 9528 28040 9580
rect 33508 9571 33560 9580
rect 33508 9537 33517 9571
rect 33517 9537 33551 9571
rect 33551 9537 33560 9571
rect 33508 9528 33560 9537
rect 41420 9596 41472 9648
rect 44180 9639 44232 9648
rect 44180 9605 44189 9639
rect 44189 9605 44223 9639
rect 44223 9605 44232 9639
rect 44180 9596 44232 9605
rect 45284 9639 45336 9648
rect 45284 9605 45293 9639
rect 45293 9605 45327 9639
rect 45327 9605 45336 9639
rect 45284 9596 45336 9605
rect 45560 9639 45612 9648
rect 45560 9605 45569 9639
rect 45569 9605 45603 9639
rect 45603 9605 45612 9639
rect 45560 9596 45612 9605
rect 46664 9639 46716 9648
rect 46664 9605 46673 9639
rect 46673 9605 46707 9639
rect 46707 9605 46716 9639
rect 46664 9596 46716 9605
rect 47032 9639 47084 9648
rect 47032 9605 47041 9639
rect 47041 9605 47075 9639
rect 47075 9605 47084 9639
rect 47032 9596 47084 9605
rect 42892 9571 42944 9580
rect 24952 9460 25004 9512
rect 27620 9503 27672 9512
rect 27620 9469 27629 9503
rect 27629 9469 27663 9503
rect 27663 9469 27672 9503
rect 27620 9460 27672 9469
rect 28448 9460 28500 9512
rect 28724 9503 28776 9512
rect 28724 9469 28733 9503
rect 28733 9469 28767 9503
rect 28767 9469 28776 9503
rect 28724 9460 28776 9469
rect 23020 9324 23072 9376
rect 24860 9367 24912 9376
rect 24860 9333 24869 9367
rect 24869 9333 24903 9367
rect 24903 9333 24912 9367
rect 24860 9324 24912 9333
rect 25320 9324 25372 9376
rect 29092 9392 29144 9444
rect 30288 9460 30340 9512
rect 30656 9392 30708 9444
rect 30840 9392 30892 9444
rect 31760 9392 31812 9444
rect 33324 9460 33376 9512
rect 33968 9503 34020 9512
rect 33968 9469 33977 9503
rect 33977 9469 34011 9503
rect 34011 9469 34020 9503
rect 33968 9460 34020 9469
rect 34152 9503 34204 9512
rect 34152 9469 34161 9503
rect 34161 9469 34195 9503
rect 34195 9469 34204 9503
rect 34152 9460 34204 9469
rect 34336 9503 34388 9512
rect 34336 9469 34345 9503
rect 34345 9469 34379 9503
rect 34379 9469 34388 9503
rect 34336 9460 34388 9469
rect 35532 9460 35584 9512
rect 36176 9460 36228 9512
rect 36912 9503 36964 9512
rect 36912 9469 36921 9503
rect 36921 9469 36955 9503
rect 36955 9469 36964 9503
rect 36912 9460 36964 9469
rect 37096 9503 37148 9512
rect 37096 9469 37105 9503
rect 37105 9469 37139 9503
rect 37139 9469 37148 9503
rect 37096 9460 37148 9469
rect 37924 9460 37976 9512
rect 36544 9392 36596 9444
rect 27436 9324 27488 9376
rect 29920 9324 29972 9376
rect 30012 9324 30064 9376
rect 31116 9324 31168 9376
rect 35992 9324 36044 9376
rect 36176 9324 36228 9376
rect 38660 9392 38712 9444
rect 42892 9537 42901 9571
rect 42901 9537 42935 9571
rect 42935 9537 42944 9571
rect 42892 9528 42944 9537
rect 42984 9528 43036 9580
rect 40408 9460 40460 9512
rect 41236 9503 41288 9512
rect 41236 9469 41245 9503
rect 41245 9469 41279 9503
rect 41279 9469 41288 9503
rect 41236 9460 41288 9469
rect 41420 9503 41472 9512
rect 41420 9469 41429 9503
rect 41429 9469 41463 9503
rect 41463 9469 41472 9503
rect 41604 9503 41656 9512
rect 41420 9460 41472 9469
rect 41604 9469 41613 9503
rect 41613 9469 41647 9503
rect 41647 9469 41656 9503
rect 41604 9460 41656 9469
rect 42340 9460 42392 9512
rect 43904 9460 43956 9512
rect 45652 9528 45704 9580
rect 44088 9392 44140 9444
rect 40040 9324 40092 9376
rect 41604 9324 41656 9376
rect 41696 9324 41748 9376
rect 42984 9324 43036 9376
rect 44824 9367 44876 9376
rect 44824 9333 44833 9367
rect 44833 9333 44867 9367
rect 44867 9333 44876 9367
rect 44824 9324 44876 9333
rect 46020 9460 46072 9512
rect 47860 9596 47912 9648
rect 49608 9707 49660 9716
rect 49608 9673 49617 9707
rect 49617 9673 49651 9707
rect 49651 9673 49660 9707
rect 49608 9664 49660 9673
rect 50436 9639 50488 9648
rect 50436 9605 50445 9639
rect 50445 9605 50479 9639
rect 50479 9605 50488 9639
rect 50436 9596 50488 9605
rect 51264 9596 51316 9648
rect 53840 9664 53892 9716
rect 54392 9707 54444 9716
rect 54392 9673 54401 9707
rect 54401 9673 54435 9707
rect 54435 9673 54444 9707
rect 54392 9664 54444 9673
rect 55404 9707 55456 9716
rect 55404 9673 55413 9707
rect 55413 9673 55447 9707
rect 55447 9673 55456 9707
rect 55404 9664 55456 9673
rect 56048 9664 56100 9716
rect 56416 9707 56468 9716
rect 56416 9673 56425 9707
rect 56425 9673 56459 9707
rect 56459 9673 56468 9707
rect 56416 9664 56468 9673
rect 58164 9707 58216 9716
rect 58164 9673 58173 9707
rect 58173 9673 58207 9707
rect 58207 9673 58216 9707
rect 58164 9664 58216 9673
rect 48320 9571 48372 9580
rect 48320 9537 48329 9571
rect 48329 9537 48363 9571
rect 48363 9537 48372 9571
rect 48320 9528 48372 9537
rect 49240 9528 49292 9580
rect 49700 9460 49752 9512
rect 50252 9460 50304 9512
rect 50528 9503 50580 9512
rect 50528 9469 50537 9503
rect 50537 9469 50571 9503
rect 50571 9469 50580 9503
rect 51724 9503 51776 9512
rect 50528 9460 50580 9469
rect 47216 9392 47268 9444
rect 50068 9435 50120 9444
rect 47768 9324 47820 9376
rect 48044 9324 48096 9376
rect 50068 9401 50077 9435
rect 50077 9401 50111 9435
rect 50111 9401 50120 9435
rect 50068 9392 50120 9401
rect 50344 9392 50396 9444
rect 51724 9469 51733 9503
rect 51733 9469 51767 9503
rect 51767 9469 51776 9503
rect 51724 9460 51776 9469
rect 51816 9460 51868 9512
rect 52368 9528 52420 9580
rect 53288 9528 53340 9580
rect 53564 9528 53616 9580
rect 56508 9596 56560 9648
rect 55128 9571 55180 9580
rect 55128 9537 55137 9571
rect 55137 9537 55171 9571
rect 55171 9537 55180 9571
rect 55128 9528 55180 9537
rect 52644 9460 52696 9512
rect 54944 9460 54996 9512
rect 48780 9324 48832 9376
rect 50896 9324 50948 9376
rect 51448 9324 51500 9376
rect 55680 9324 55732 9376
rect 56140 9460 56192 9512
rect 58348 9503 58400 9512
rect 58348 9469 58357 9503
rect 58357 9469 58391 9503
rect 58391 9469 58400 9503
rect 58348 9460 58400 9469
rect 60556 9460 60608 9512
rect 57336 9324 57388 9376
rect 57796 9367 57848 9376
rect 57796 9333 57805 9367
rect 57805 9333 57839 9367
rect 57839 9333 57848 9367
rect 57796 9324 57848 9333
rect 59820 9324 59872 9376
rect 60464 9367 60516 9376
rect 60464 9333 60473 9367
rect 60473 9333 60507 9367
rect 60507 9333 60516 9367
rect 60464 9324 60516 9333
rect 61292 9367 61344 9376
rect 61292 9333 61301 9367
rect 61301 9333 61335 9367
rect 61335 9333 61344 9367
rect 61292 9324 61344 9333
rect 21774 9222 21826 9274
rect 21838 9222 21890 9274
rect 21902 9222 21954 9274
rect 21966 9222 22018 9274
rect 42566 9222 42618 9274
rect 42630 9222 42682 9274
rect 42694 9222 42746 9274
rect 42758 9222 42810 9274
rect 2596 9027 2648 9036
rect 2596 8993 2605 9027
rect 2605 8993 2639 9027
rect 2639 8993 2648 9027
rect 2596 8984 2648 8993
rect 2872 8984 2924 9036
rect 3056 9027 3108 9036
rect 3056 8993 3065 9027
rect 3065 8993 3099 9027
rect 3099 8993 3108 9027
rect 17224 9120 17276 9172
rect 4712 9052 4764 9104
rect 7104 9052 7156 9104
rect 18420 9052 18472 9104
rect 18604 9095 18656 9104
rect 18604 9061 18613 9095
rect 18613 9061 18647 9095
rect 18647 9061 18656 9095
rect 18604 9052 18656 9061
rect 18696 9052 18748 9104
rect 21640 9052 21692 9104
rect 3056 8984 3108 8993
rect 6552 8984 6604 9036
rect 7196 9027 7248 9036
rect 7196 8993 7205 9027
rect 7205 8993 7239 9027
rect 7239 8993 7248 9027
rect 7196 8984 7248 8993
rect 7288 8984 7340 9036
rect 8024 8984 8076 9036
rect 8760 9027 8812 9036
rect 8760 8993 8769 9027
rect 8769 8993 8803 9027
rect 8803 8993 8812 9027
rect 8760 8984 8812 8993
rect 10140 9027 10192 9036
rect 10140 8993 10149 9027
rect 10149 8993 10183 9027
rect 10183 8993 10192 9027
rect 10140 8984 10192 8993
rect 10508 9027 10560 9036
rect 10508 8993 10517 9027
rect 10517 8993 10551 9027
rect 10551 8993 10560 9027
rect 10508 8984 10560 8993
rect 10876 8984 10928 9036
rect 12348 9027 12400 9036
rect 4344 8916 4396 8968
rect 5448 8959 5500 8968
rect 5448 8925 5457 8959
rect 5457 8925 5491 8959
rect 5491 8925 5500 8959
rect 5448 8916 5500 8925
rect 4160 8848 4212 8900
rect 10600 8959 10652 8968
rect 10600 8925 10609 8959
rect 10609 8925 10643 8959
rect 10643 8925 10652 8959
rect 10600 8916 10652 8925
rect 10784 8916 10836 8968
rect 12348 8993 12357 9027
rect 12357 8993 12391 9027
rect 12391 8993 12400 9027
rect 12348 8984 12400 8993
rect 12992 8984 13044 9036
rect 13544 9027 13596 9036
rect 13544 8993 13553 9027
rect 13553 8993 13587 9027
rect 13587 8993 13596 9027
rect 13544 8984 13596 8993
rect 13728 9027 13780 9036
rect 13728 8993 13737 9027
rect 13737 8993 13771 9027
rect 13771 8993 13780 9027
rect 13728 8984 13780 8993
rect 15936 8984 15988 9036
rect 16028 8984 16080 9036
rect 16764 8984 16816 9036
rect 12532 8959 12584 8968
rect 8208 8848 8260 8900
rect 11152 8891 11204 8900
rect 11152 8857 11161 8891
rect 11161 8857 11195 8891
rect 11195 8857 11204 8891
rect 11152 8848 11204 8857
rect 12532 8925 12541 8959
rect 12541 8925 12575 8959
rect 12575 8925 12584 8959
rect 12532 8916 12584 8925
rect 4068 8780 4120 8832
rect 4804 8780 4856 8832
rect 6276 8823 6328 8832
rect 6276 8789 6285 8823
rect 6285 8789 6319 8823
rect 6319 8789 6328 8823
rect 6276 8780 6328 8789
rect 6368 8780 6420 8832
rect 10508 8780 10560 8832
rect 12256 8780 12308 8832
rect 13636 8959 13688 8968
rect 13636 8925 13645 8959
rect 13645 8925 13679 8959
rect 13679 8925 13688 8959
rect 13636 8916 13688 8925
rect 16120 8916 16172 8968
rect 16396 8916 16448 8968
rect 17316 9027 17368 9036
rect 17316 8993 17325 9027
rect 17325 8993 17359 9027
rect 17359 8993 17368 9027
rect 17316 8984 17368 8993
rect 19156 8984 19208 9036
rect 19248 9027 19300 9036
rect 19248 8993 19257 9027
rect 19257 8993 19291 9027
rect 19291 8993 19300 9027
rect 19248 8984 19300 8993
rect 21456 9027 21508 9036
rect 17224 8959 17276 8968
rect 17224 8925 17233 8959
rect 17233 8925 17267 8959
rect 17267 8925 17276 8959
rect 17224 8916 17276 8925
rect 17500 8916 17552 8968
rect 19340 8916 19392 8968
rect 19708 8916 19760 8968
rect 20904 8959 20956 8968
rect 20904 8925 20913 8959
rect 20913 8925 20947 8959
rect 20947 8925 20956 8959
rect 20904 8916 20956 8925
rect 21456 8993 21465 9027
rect 21465 8993 21499 9027
rect 21499 8993 21508 9027
rect 21456 8984 21508 8993
rect 21548 8984 21600 9036
rect 23112 9120 23164 9172
rect 22376 9027 22428 9036
rect 21272 8916 21324 8968
rect 22376 8993 22385 9027
rect 22385 8993 22419 9027
rect 22419 8993 22428 9027
rect 22376 8984 22428 8993
rect 22284 8959 22336 8968
rect 22284 8925 22293 8959
rect 22293 8925 22327 8959
rect 22327 8925 22336 8959
rect 22284 8916 22336 8925
rect 22560 8916 22612 8968
rect 23940 8916 23992 8968
rect 24860 9052 24912 9104
rect 24400 8984 24452 9036
rect 25044 9027 25096 9036
rect 25044 8993 25053 9027
rect 25053 8993 25087 9027
rect 25087 8993 25096 9027
rect 25044 8984 25096 8993
rect 25412 9027 25464 9036
rect 25412 8993 25421 9027
rect 25421 8993 25455 9027
rect 25455 8993 25464 9027
rect 25412 8984 25464 8993
rect 30288 9052 30340 9104
rect 30380 9052 30432 9104
rect 33324 9120 33376 9172
rect 33508 9163 33560 9172
rect 33508 9129 33517 9163
rect 33517 9129 33551 9163
rect 33551 9129 33560 9163
rect 33508 9120 33560 9129
rect 34520 9120 34572 9172
rect 36452 9120 36504 9172
rect 36544 9120 36596 9172
rect 33692 9095 33744 9104
rect 33692 9061 33701 9095
rect 33701 9061 33735 9095
rect 33735 9061 33744 9095
rect 33692 9052 33744 9061
rect 26148 8984 26200 9036
rect 28448 9027 28500 9036
rect 28448 8993 28457 9027
rect 28457 8993 28491 9027
rect 28491 8993 28500 9027
rect 28448 8984 28500 8993
rect 30012 9027 30064 9036
rect 30012 8993 30021 9027
rect 30021 8993 30055 9027
rect 30055 8993 30064 9027
rect 30012 8984 30064 8993
rect 30104 8984 30156 9036
rect 32404 9027 32456 9036
rect 32404 8993 32413 9027
rect 32413 8993 32447 9027
rect 32447 8993 32456 9027
rect 32404 8984 32456 8993
rect 34612 9052 34664 9104
rect 34888 9052 34940 9104
rect 34520 9027 34572 9036
rect 34520 8993 34529 9027
rect 34529 8993 34563 9027
rect 34563 8993 34572 9027
rect 34520 8984 34572 8993
rect 34704 8984 34756 9036
rect 37280 9052 37332 9104
rect 38292 9095 38344 9104
rect 38292 9061 38301 9095
rect 38301 9061 38335 9095
rect 38335 9061 38344 9095
rect 38292 9052 38344 9061
rect 39488 9052 39540 9104
rect 44824 9052 44876 9104
rect 48688 9052 48740 9104
rect 49332 9120 49384 9172
rect 49976 9120 50028 9172
rect 60648 9120 60700 9172
rect 14004 8848 14056 8900
rect 27160 8916 27212 8968
rect 28356 8959 28408 8968
rect 26608 8848 26660 8900
rect 27436 8848 27488 8900
rect 28356 8925 28365 8959
rect 28365 8925 28399 8959
rect 28399 8925 28408 8959
rect 28356 8916 28408 8925
rect 28816 8916 28868 8968
rect 29460 8916 29512 8968
rect 30748 8959 30800 8968
rect 30748 8925 30757 8959
rect 30757 8925 30791 8959
rect 30791 8925 30800 8959
rect 30748 8916 30800 8925
rect 32772 8916 32824 8968
rect 27620 8848 27672 8900
rect 34796 8916 34848 8968
rect 35532 8959 35584 8968
rect 35532 8925 35541 8959
rect 35541 8925 35575 8959
rect 35575 8925 35584 8959
rect 35532 8916 35584 8925
rect 35716 8916 35768 8968
rect 36268 8848 36320 8900
rect 12992 8780 13044 8832
rect 13820 8780 13872 8832
rect 15200 8780 15252 8832
rect 15476 8780 15528 8832
rect 16120 8823 16172 8832
rect 16120 8789 16129 8823
rect 16129 8789 16163 8823
rect 16163 8789 16172 8823
rect 16120 8780 16172 8789
rect 16764 8823 16816 8832
rect 16764 8789 16773 8823
rect 16773 8789 16807 8823
rect 16807 8789 16816 8823
rect 16764 8780 16816 8789
rect 16856 8823 16908 8832
rect 16856 8789 16865 8823
rect 16865 8789 16899 8823
rect 16899 8789 16908 8823
rect 16856 8780 16908 8789
rect 17408 8780 17460 8832
rect 18144 8780 18196 8832
rect 18512 8780 18564 8832
rect 19892 8780 19944 8832
rect 20260 8780 20312 8832
rect 20352 8823 20404 8832
rect 20352 8789 20361 8823
rect 20361 8789 20395 8823
rect 20395 8789 20404 8823
rect 20352 8780 20404 8789
rect 21548 8780 21600 8832
rect 21824 8780 21876 8832
rect 23480 8780 23532 8832
rect 24400 8823 24452 8832
rect 24400 8789 24409 8823
rect 24409 8789 24443 8823
rect 24443 8789 24452 8823
rect 24400 8780 24452 8789
rect 25872 8823 25924 8832
rect 25872 8789 25881 8823
rect 25881 8789 25915 8823
rect 25915 8789 25924 8823
rect 25872 8780 25924 8789
rect 26240 8823 26292 8832
rect 26240 8789 26249 8823
rect 26249 8789 26283 8823
rect 26283 8789 26292 8823
rect 26240 8780 26292 8789
rect 27712 8780 27764 8832
rect 28632 8823 28684 8832
rect 28632 8789 28641 8823
rect 28641 8789 28675 8823
rect 28675 8789 28684 8823
rect 28632 8780 28684 8789
rect 29276 8823 29328 8832
rect 29276 8789 29285 8823
rect 29285 8789 29319 8823
rect 29319 8789 29328 8823
rect 29276 8780 29328 8789
rect 29368 8780 29420 8832
rect 31208 8780 31260 8832
rect 33416 8780 33468 8832
rect 33876 8780 33928 8832
rect 34888 8780 34940 8832
rect 35072 8823 35124 8832
rect 35072 8789 35081 8823
rect 35081 8789 35115 8823
rect 35115 8789 35124 8823
rect 35072 8780 35124 8789
rect 36728 8823 36780 8832
rect 36728 8789 36737 8823
rect 36737 8789 36771 8823
rect 36771 8789 36780 8823
rect 36728 8780 36780 8789
rect 37188 8823 37240 8832
rect 37188 8789 37197 8823
rect 37197 8789 37231 8823
rect 37231 8789 37240 8823
rect 37188 8780 37240 8789
rect 40040 8984 40092 9036
rect 38476 8959 38528 8968
rect 38476 8925 38485 8959
rect 38485 8925 38519 8959
rect 38519 8925 38528 8959
rect 38476 8916 38528 8925
rect 38752 8959 38804 8968
rect 38752 8925 38761 8959
rect 38761 8925 38795 8959
rect 38795 8925 38804 8959
rect 38752 8916 38804 8925
rect 38844 8916 38896 8968
rect 41696 8984 41748 9036
rect 41972 8984 42024 9036
rect 43536 8984 43588 9036
rect 44364 8984 44416 9036
rect 47400 8984 47452 9036
rect 50528 9052 50580 9104
rect 51172 9052 51224 9104
rect 52368 9052 52420 9104
rect 52460 9052 52512 9104
rect 54208 9052 54260 9104
rect 41604 8959 41656 8968
rect 41604 8925 41613 8959
rect 41613 8925 41647 8959
rect 41647 8925 41656 8959
rect 41604 8916 41656 8925
rect 42248 8916 42300 8968
rect 43352 8959 43404 8968
rect 43352 8925 43361 8959
rect 43361 8925 43395 8959
rect 43395 8925 43404 8959
rect 43352 8916 43404 8925
rect 44088 8916 44140 8968
rect 45100 8916 45152 8968
rect 47768 8916 47820 8968
rect 49792 8916 49844 8968
rect 50896 9027 50948 9036
rect 50896 8993 50905 9027
rect 50905 8993 50939 9027
rect 50939 8993 50948 9027
rect 50896 8984 50948 8993
rect 51356 8984 51408 9036
rect 51448 8984 51500 9036
rect 52736 8984 52788 9036
rect 53564 8984 53616 9036
rect 55220 8984 55272 9036
rect 55404 8984 55456 9036
rect 59268 8984 59320 9036
rect 40316 8848 40368 8900
rect 42340 8848 42392 8900
rect 43076 8848 43128 8900
rect 46112 8848 46164 8900
rect 49976 8848 50028 8900
rect 51816 8848 51868 8900
rect 53288 8916 53340 8968
rect 54300 8916 54352 8968
rect 55128 8916 55180 8968
rect 56140 8959 56192 8968
rect 56140 8925 56149 8959
rect 56149 8925 56183 8959
rect 56183 8925 56192 8959
rect 56140 8916 56192 8925
rect 56416 8959 56468 8968
rect 56416 8925 56425 8959
rect 56425 8925 56459 8959
rect 56459 8925 56468 8959
rect 56416 8916 56468 8925
rect 56508 8916 56560 8968
rect 57060 8916 57112 8968
rect 58624 8959 58676 8968
rect 58624 8925 58633 8959
rect 58633 8925 58667 8959
rect 58667 8925 58676 8959
rect 58624 8916 58676 8925
rect 54760 8848 54812 8900
rect 58256 8848 58308 8900
rect 60464 8891 60516 8900
rect 40592 8823 40644 8832
rect 40592 8789 40601 8823
rect 40601 8789 40635 8823
rect 40635 8789 40644 8823
rect 40592 8780 40644 8789
rect 41052 8780 41104 8832
rect 41236 8823 41288 8832
rect 41236 8789 41245 8823
rect 41245 8789 41279 8823
rect 41279 8789 41288 8823
rect 41236 8780 41288 8789
rect 41972 8780 42024 8832
rect 44272 8823 44324 8832
rect 44272 8789 44281 8823
rect 44281 8789 44315 8823
rect 44315 8789 44324 8823
rect 44272 8780 44324 8789
rect 44640 8823 44692 8832
rect 44640 8789 44649 8823
rect 44649 8789 44683 8823
rect 44683 8789 44692 8823
rect 44640 8780 44692 8789
rect 46296 8823 46348 8832
rect 46296 8789 46305 8823
rect 46305 8789 46339 8823
rect 46339 8789 46348 8823
rect 46296 8780 46348 8789
rect 47032 8823 47084 8832
rect 47032 8789 47041 8823
rect 47041 8789 47075 8823
rect 47075 8789 47084 8823
rect 47032 8780 47084 8789
rect 47400 8780 47452 8832
rect 50068 8823 50120 8832
rect 50068 8789 50077 8823
rect 50077 8789 50111 8823
rect 50111 8789 50120 8823
rect 50068 8780 50120 8789
rect 51540 8823 51592 8832
rect 51540 8789 51549 8823
rect 51549 8789 51583 8823
rect 51583 8789 51592 8823
rect 51540 8780 51592 8789
rect 51724 8780 51776 8832
rect 52276 8780 52328 8832
rect 52828 8780 52880 8832
rect 54852 8823 54904 8832
rect 54852 8789 54861 8823
rect 54861 8789 54895 8823
rect 54895 8789 54904 8823
rect 54852 8780 54904 8789
rect 56324 8780 56376 8832
rect 56508 8780 56560 8832
rect 58440 8823 58492 8832
rect 58440 8789 58449 8823
rect 58449 8789 58483 8823
rect 58483 8789 58492 8823
rect 58440 8780 58492 8789
rect 60464 8857 60473 8891
rect 60473 8857 60507 8891
rect 60507 8857 60516 8891
rect 60464 8848 60516 8857
rect 61844 8984 61896 9036
rect 61108 8959 61160 8968
rect 61108 8925 61117 8959
rect 61117 8925 61151 8959
rect 61151 8925 61160 8959
rect 61108 8916 61160 8925
rect 61384 8916 61436 8968
rect 59084 8780 59136 8832
rect 59820 8823 59872 8832
rect 59820 8789 59829 8823
rect 59829 8789 59863 8823
rect 59863 8789 59872 8823
rect 59820 8780 59872 8789
rect 11378 8678 11430 8730
rect 11442 8678 11494 8730
rect 11506 8678 11558 8730
rect 11570 8678 11622 8730
rect 32170 8678 32222 8730
rect 32234 8678 32286 8730
rect 32298 8678 32350 8730
rect 32362 8678 32414 8730
rect 52962 8678 53014 8730
rect 53026 8678 53078 8730
rect 53090 8678 53142 8730
rect 53154 8678 53206 8730
rect 3056 8619 3108 8628
rect 3056 8585 3065 8619
rect 3065 8585 3099 8619
rect 3099 8585 3108 8619
rect 3056 8576 3108 8585
rect 2872 8508 2924 8560
rect 2596 8440 2648 8492
rect 6368 8576 6420 8628
rect 8760 8576 8812 8628
rect 11152 8576 11204 8628
rect 11888 8619 11940 8628
rect 11888 8585 11897 8619
rect 11897 8585 11931 8619
rect 11931 8585 11940 8619
rect 11888 8576 11940 8585
rect 12348 8576 12400 8628
rect 12532 8576 12584 8628
rect 15108 8619 15160 8628
rect 15108 8585 15117 8619
rect 15117 8585 15151 8619
rect 15151 8585 15160 8619
rect 15108 8576 15160 8585
rect 15936 8576 15988 8628
rect 19984 8576 20036 8628
rect 20260 8576 20312 8628
rect 20904 8576 20956 8628
rect 21640 8576 21692 8628
rect 22376 8576 22428 8628
rect 25412 8576 25464 8628
rect 26516 8576 26568 8628
rect 28448 8619 28500 8628
rect 28448 8585 28457 8619
rect 28457 8585 28491 8619
rect 28491 8585 28500 8619
rect 28448 8576 28500 8585
rect 28540 8576 28592 8628
rect 32496 8576 32548 8628
rect 34796 8576 34848 8628
rect 35900 8576 35952 8628
rect 36452 8576 36504 8628
rect 38752 8619 38804 8628
rect 38752 8585 38761 8619
rect 38761 8585 38795 8619
rect 38795 8585 38804 8619
rect 38752 8576 38804 8585
rect 11060 8508 11112 8560
rect 4068 8372 4120 8424
rect 7288 8440 7340 8492
rect 5448 8304 5500 8356
rect 6644 8347 6696 8356
rect 6644 8313 6653 8347
rect 6653 8313 6687 8347
rect 6687 8313 6696 8347
rect 6644 8304 6696 8313
rect 5816 8279 5868 8288
rect 5816 8245 5825 8279
rect 5825 8245 5859 8279
rect 5859 8245 5868 8279
rect 5816 8236 5868 8245
rect 6092 8236 6144 8288
rect 8208 8304 8260 8356
rect 10876 8440 10928 8492
rect 18052 8551 18104 8560
rect 18052 8517 18061 8551
rect 18061 8517 18095 8551
rect 18095 8517 18104 8551
rect 18052 8508 18104 8517
rect 18328 8508 18380 8560
rect 19340 8508 19392 8560
rect 20352 8508 20404 8560
rect 24952 8508 25004 8560
rect 26700 8508 26752 8560
rect 27344 8508 27396 8560
rect 28908 8508 28960 8560
rect 30012 8508 30064 8560
rect 38844 8508 38896 8560
rect 12072 8440 12124 8492
rect 8852 8347 8904 8356
rect 8852 8313 8861 8347
rect 8861 8313 8895 8347
rect 8895 8313 8904 8347
rect 8852 8304 8904 8313
rect 11244 8415 11296 8424
rect 11244 8381 11253 8415
rect 11253 8381 11287 8415
rect 11287 8381 11296 8415
rect 14004 8415 14056 8424
rect 11244 8372 11296 8381
rect 14004 8381 14013 8415
rect 14013 8381 14047 8415
rect 14047 8381 14056 8415
rect 14004 8372 14056 8381
rect 15016 8440 15068 8492
rect 16120 8440 16172 8492
rect 15108 8372 15160 8424
rect 15200 8372 15252 8424
rect 15752 8372 15804 8424
rect 16764 8372 16816 8424
rect 17224 8372 17276 8424
rect 17500 8440 17552 8492
rect 22008 8440 22060 8492
rect 22100 8440 22152 8492
rect 20352 8415 20404 8424
rect 20352 8381 20361 8415
rect 20361 8381 20395 8415
rect 20395 8381 20404 8415
rect 20352 8372 20404 8381
rect 20720 8415 20772 8424
rect 20720 8381 20729 8415
rect 20729 8381 20763 8415
rect 20763 8381 20772 8415
rect 20720 8372 20772 8381
rect 21548 8372 21600 8424
rect 21732 8415 21784 8424
rect 21732 8381 21741 8415
rect 21741 8381 21775 8415
rect 21775 8381 21784 8415
rect 21732 8372 21784 8381
rect 22192 8415 22244 8424
rect 22192 8381 22201 8415
rect 22201 8381 22235 8415
rect 22235 8381 22244 8415
rect 22192 8372 22244 8381
rect 23480 8372 23532 8424
rect 25228 8372 25280 8424
rect 25872 8372 25924 8424
rect 26240 8372 26292 8424
rect 26516 8372 26568 8424
rect 27160 8415 27212 8424
rect 27160 8381 27169 8415
rect 27169 8381 27203 8415
rect 27203 8381 27212 8415
rect 27160 8372 27212 8381
rect 27344 8372 27396 8424
rect 27620 8415 27672 8424
rect 27620 8381 27629 8415
rect 27629 8381 27663 8415
rect 27663 8381 27672 8415
rect 27620 8372 27672 8381
rect 27896 8415 27948 8424
rect 27896 8381 27905 8415
rect 27905 8381 27939 8415
rect 27939 8381 27948 8415
rect 28540 8440 28592 8492
rect 29276 8483 29328 8492
rect 29276 8449 29285 8483
rect 29285 8449 29319 8483
rect 29319 8449 29328 8483
rect 29276 8440 29328 8449
rect 30564 8440 30616 8492
rect 27896 8372 27948 8381
rect 28724 8372 28776 8424
rect 29368 8415 29420 8424
rect 29368 8381 29377 8415
rect 29377 8381 29411 8415
rect 29411 8381 29420 8415
rect 29368 8372 29420 8381
rect 30656 8415 30708 8424
rect 11520 8304 11572 8356
rect 13452 8347 13504 8356
rect 13452 8313 13461 8347
rect 13461 8313 13495 8347
rect 13495 8313 13504 8347
rect 13452 8304 13504 8313
rect 15936 8304 15988 8356
rect 17408 8347 17460 8356
rect 13176 8236 13228 8288
rect 13728 8236 13780 8288
rect 16580 8236 16632 8288
rect 17408 8313 17417 8347
rect 17417 8313 17451 8347
rect 17451 8313 17460 8347
rect 17408 8304 17460 8313
rect 18144 8236 18196 8288
rect 18880 8304 18932 8356
rect 19708 8304 19760 8356
rect 22008 8304 22060 8356
rect 22284 8304 22336 8356
rect 22744 8304 22796 8356
rect 19800 8236 19852 8288
rect 23296 8236 23348 8288
rect 24952 8236 25004 8288
rect 25044 8279 25096 8288
rect 25044 8245 25053 8279
rect 25053 8245 25087 8279
rect 25087 8245 25096 8279
rect 25044 8236 25096 8245
rect 25320 8236 25372 8288
rect 26976 8236 27028 8288
rect 27528 8279 27580 8288
rect 27528 8245 27537 8279
rect 27537 8245 27571 8279
rect 27571 8245 27580 8279
rect 27528 8236 27580 8245
rect 27712 8236 27764 8288
rect 28172 8236 28224 8288
rect 30656 8381 30665 8415
rect 30665 8381 30699 8415
rect 30699 8381 30708 8415
rect 30656 8372 30708 8381
rect 31300 8372 31352 8424
rect 31852 8415 31904 8424
rect 31852 8381 31861 8415
rect 31861 8381 31895 8415
rect 31895 8381 31904 8415
rect 31852 8372 31904 8381
rect 36084 8440 36136 8492
rect 36728 8440 36780 8492
rect 36820 8440 36872 8492
rect 32036 8372 32088 8424
rect 32312 8304 32364 8356
rect 30656 8236 30708 8288
rect 31300 8279 31352 8288
rect 31300 8245 31309 8279
rect 31309 8245 31343 8279
rect 31343 8245 31352 8279
rect 31300 8236 31352 8245
rect 31852 8236 31904 8288
rect 33048 8236 33100 8288
rect 33692 8372 33744 8424
rect 35072 8372 35124 8424
rect 35164 8372 35216 8424
rect 35440 8415 35492 8424
rect 35440 8381 35449 8415
rect 35449 8381 35483 8415
rect 35483 8381 35492 8415
rect 35440 8372 35492 8381
rect 37188 8415 37240 8424
rect 35532 8236 35584 8288
rect 37188 8381 37197 8415
rect 37197 8381 37231 8415
rect 37231 8381 37240 8415
rect 37188 8372 37240 8381
rect 38660 8440 38712 8492
rect 41420 8576 41472 8628
rect 41880 8576 41932 8628
rect 45560 8576 45612 8628
rect 46296 8576 46348 8628
rect 47308 8508 47360 8560
rect 48504 8551 48556 8560
rect 48504 8517 48513 8551
rect 48513 8517 48547 8551
rect 48547 8517 48556 8551
rect 48504 8508 48556 8517
rect 52736 8619 52788 8628
rect 50252 8508 50304 8560
rect 41236 8440 41288 8492
rect 41972 8483 42024 8492
rect 41972 8449 41981 8483
rect 41981 8449 42015 8483
rect 42015 8449 42024 8483
rect 41972 8440 42024 8449
rect 44272 8440 44324 8492
rect 46296 8440 46348 8492
rect 50068 8483 50120 8492
rect 38384 8347 38436 8356
rect 38384 8313 38393 8347
rect 38393 8313 38427 8347
rect 38427 8313 38436 8347
rect 39948 8372 40000 8424
rect 40316 8415 40368 8424
rect 40316 8381 40325 8415
rect 40325 8381 40359 8415
rect 40359 8381 40368 8415
rect 40316 8372 40368 8381
rect 40500 8415 40552 8424
rect 40500 8381 40509 8415
rect 40509 8381 40543 8415
rect 40543 8381 40552 8415
rect 40500 8372 40552 8381
rect 40592 8415 40644 8424
rect 40592 8381 40601 8415
rect 40601 8381 40635 8415
rect 40635 8381 40644 8415
rect 40592 8372 40644 8381
rect 41512 8372 41564 8424
rect 38384 8304 38436 8313
rect 36268 8279 36320 8288
rect 36268 8245 36277 8279
rect 36277 8245 36311 8279
rect 36311 8245 36320 8279
rect 36268 8236 36320 8245
rect 41604 8236 41656 8288
rect 41696 8236 41748 8288
rect 43260 8372 43312 8424
rect 44456 8372 44508 8424
rect 44640 8415 44692 8424
rect 44640 8381 44649 8415
rect 44649 8381 44683 8415
rect 44683 8381 44692 8415
rect 44640 8372 44692 8381
rect 46848 8372 46900 8424
rect 44732 8304 44784 8356
rect 45468 8347 45520 8356
rect 41880 8236 41932 8288
rect 45100 8279 45152 8288
rect 45100 8245 45109 8279
rect 45109 8245 45143 8279
rect 45143 8245 45152 8279
rect 45100 8236 45152 8245
rect 45468 8313 45477 8347
rect 45477 8313 45511 8347
rect 45511 8313 45520 8347
rect 45468 8304 45520 8313
rect 45744 8304 45796 8356
rect 47308 8372 47360 8424
rect 47492 8415 47544 8424
rect 47492 8381 47501 8415
rect 47501 8381 47535 8415
rect 47535 8381 47544 8415
rect 47492 8372 47544 8381
rect 47768 8372 47820 8424
rect 48504 8372 48556 8424
rect 50068 8449 50077 8483
rect 50077 8449 50111 8483
rect 50111 8449 50120 8483
rect 50068 8440 50120 8449
rect 50160 8440 50212 8492
rect 50620 8440 50672 8492
rect 50896 8440 50948 8492
rect 51264 8440 51316 8492
rect 52736 8585 52745 8619
rect 52745 8585 52779 8619
rect 52779 8585 52788 8619
rect 52736 8576 52788 8585
rect 53564 8619 53616 8628
rect 53564 8585 53573 8619
rect 53573 8585 53607 8619
rect 53607 8585 53616 8619
rect 53564 8576 53616 8585
rect 55864 8576 55916 8628
rect 56140 8576 56192 8628
rect 56600 8576 56652 8628
rect 57704 8576 57756 8628
rect 58624 8619 58676 8628
rect 58624 8585 58633 8619
rect 58633 8585 58667 8619
rect 58667 8585 58676 8619
rect 58624 8576 58676 8585
rect 61844 8619 61896 8628
rect 61844 8585 61853 8619
rect 61853 8585 61887 8619
rect 61887 8585 61896 8619
rect 61844 8576 61896 8585
rect 52828 8508 52880 8560
rect 61108 8551 61160 8560
rect 52184 8440 52236 8492
rect 52276 8440 52328 8492
rect 48872 8372 48924 8424
rect 51172 8372 51224 8424
rect 54208 8415 54260 8424
rect 54208 8381 54217 8415
rect 54217 8381 54251 8415
rect 54251 8381 54260 8415
rect 54208 8372 54260 8381
rect 55220 8372 55272 8424
rect 48044 8304 48096 8356
rect 49240 8304 49292 8356
rect 50252 8347 50304 8356
rect 49516 8279 49568 8288
rect 49516 8245 49525 8279
rect 49525 8245 49559 8279
rect 49559 8245 49568 8279
rect 49516 8236 49568 8245
rect 50252 8313 50261 8347
rect 50261 8313 50295 8347
rect 50295 8313 50304 8347
rect 50252 8304 50304 8313
rect 50620 8304 50672 8356
rect 50804 8347 50856 8356
rect 50804 8313 50813 8347
rect 50813 8313 50847 8347
rect 50847 8313 50856 8347
rect 50804 8304 50856 8313
rect 51080 8304 51132 8356
rect 51632 8304 51684 8356
rect 52460 8347 52512 8356
rect 52460 8313 52469 8347
rect 52469 8313 52503 8347
rect 52503 8313 52512 8347
rect 52460 8304 52512 8313
rect 53840 8347 53892 8356
rect 53840 8313 53849 8347
rect 53849 8313 53883 8347
rect 53883 8313 53892 8347
rect 53840 8304 53892 8313
rect 55312 8304 55364 8356
rect 55404 8347 55456 8356
rect 55404 8313 55413 8347
rect 55413 8313 55447 8347
rect 55447 8313 55456 8347
rect 55404 8304 55456 8313
rect 55864 8415 55916 8424
rect 55864 8381 55873 8415
rect 55873 8381 55907 8415
rect 55907 8381 55916 8415
rect 56508 8440 56560 8492
rect 61108 8517 61117 8551
rect 61117 8517 61151 8551
rect 61151 8517 61160 8551
rect 61108 8508 61160 8517
rect 61292 8508 61344 8560
rect 55864 8372 55916 8381
rect 56140 8372 56192 8424
rect 56324 8415 56376 8424
rect 56324 8381 56333 8415
rect 56333 8381 56367 8415
rect 56367 8381 56376 8415
rect 56324 8372 56376 8381
rect 59820 8440 59872 8492
rect 58348 8372 58400 8424
rect 58532 8372 58584 8424
rect 59084 8415 59136 8424
rect 59084 8381 59093 8415
rect 59093 8381 59127 8415
rect 59127 8381 59136 8415
rect 59084 8372 59136 8381
rect 60648 8372 60700 8424
rect 55956 8304 56008 8356
rect 56416 8304 56468 8356
rect 49884 8236 49936 8288
rect 50712 8236 50764 8288
rect 52000 8236 52052 8288
rect 52184 8236 52236 8288
rect 55772 8236 55824 8288
rect 57612 8279 57664 8288
rect 57612 8245 57621 8279
rect 57621 8245 57655 8279
rect 57655 8245 57664 8279
rect 57612 8236 57664 8245
rect 57704 8236 57756 8288
rect 60924 8236 60976 8288
rect 21774 8134 21826 8186
rect 21838 8134 21890 8186
rect 21902 8134 21954 8186
rect 21966 8134 22018 8186
rect 42566 8134 42618 8186
rect 42630 8134 42682 8186
rect 42694 8134 42746 8186
rect 42758 8134 42810 8186
rect 5816 8032 5868 8084
rect 6092 8007 6144 8016
rect 6092 7973 6101 8007
rect 6101 7973 6135 8007
rect 6135 7973 6144 8007
rect 6092 7964 6144 7973
rect 4344 7939 4396 7948
rect 4344 7905 4353 7939
rect 4353 7905 4387 7939
rect 4387 7905 4396 7939
rect 4344 7896 4396 7905
rect 8208 8032 8260 8084
rect 11520 8075 11572 8084
rect 11520 8041 11529 8075
rect 11529 8041 11563 8075
rect 11563 8041 11572 8075
rect 11520 8032 11572 8041
rect 7288 7896 7340 7948
rect 7564 7939 7616 7948
rect 7564 7905 7573 7939
rect 7573 7905 7607 7939
rect 7607 7905 7616 7939
rect 7564 7896 7616 7905
rect 9956 7939 10008 7948
rect 4068 7871 4120 7880
rect 4068 7837 4077 7871
rect 4077 7837 4111 7871
rect 4111 7837 4120 7871
rect 4068 7828 4120 7837
rect 6828 7828 6880 7880
rect 6552 7760 6604 7812
rect 9956 7905 9965 7939
rect 9965 7905 9999 7939
rect 9999 7905 10008 7939
rect 9956 7896 10008 7905
rect 11244 7939 11296 7948
rect 11244 7905 11253 7939
rect 11253 7905 11287 7939
rect 11287 7905 11296 7939
rect 11244 7896 11296 7905
rect 11888 7896 11940 7948
rect 8024 7828 8076 7880
rect 10600 7828 10652 7880
rect 12072 7871 12124 7880
rect 12072 7837 12081 7871
rect 12081 7837 12115 7871
rect 12115 7837 12124 7871
rect 12072 7828 12124 7837
rect 8208 7760 8260 7812
rect 17224 8032 17276 8084
rect 17316 8075 17368 8084
rect 17316 8041 17325 8075
rect 17325 8041 17359 8075
rect 17359 8041 17368 8075
rect 17316 8032 17368 8041
rect 17960 8032 18012 8084
rect 18328 8032 18380 8084
rect 12532 7964 12584 8016
rect 13176 7896 13228 7948
rect 14188 7896 14240 7948
rect 15016 7939 15068 7948
rect 15016 7905 15025 7939
rect 15025 7905 15059 7939
rect 15059 7905 15068 7939
rect 15016 7896 15068 7905
rect 17500 7964 17552 8016
rect 19524 8032 19576 8084
rect 21088 8032 21140 8084
rect 29644 8032 29696 8084
rect 30748 8032 30800 8084
rect 32312 8032 32364 8084
rect 34612 8075 34664 8084
rect 34612 8041 34621 8075
rect 34621 8041 34655 8075
rect 34655 8041 34664 8075
rect 34612 8032 34664 8041
rect 35256 8075 35308 8084
rect 35256 8041 35265 8075
rect 35265 8041 35299 8075
rect 35299 8041 35308 8075
rect 35256 8032 35308 8041
rect 35440 8032 35492 8084
rect 35808 8032 35860 8084
rect 36268 8032 36320 8084
rect 39120 8032 39172 8084
rect 43536 8075 43588 8084
rect 16580 7896 16632 7948
rect 16948 7896 17000 7948
rect 20168 7896 20220 7948
rect 20904 7939 20956 7948
rect 20904 7905 20913 7939
rect 20913 7905 20947 7939
rect 20947 7905 20956 7939
rect 20904 7896 20956 7905
rect 21088 7939 21140 7948
rect 21088 7905 21097 7939
rect 21097 7905 21131 7939
rect 21131 7905 21140 7939
rect 21088 7896 21140 7905
rect 24400 7964 24452 8016
rect 24492 7964 24544 8016
rect 25872 7964 25924 8016
rect 26516 7964 26568 8016
rect 27896 7964 27948 8016
rect 28908 7964 28960 8016
rect 29368 8007 29420 8016
rect 29368 7973 29377 8007
rect 29377 7973 29411 8007
rect 29411 7973 29420 8007
rect 29368 7964 29420 7973
rect 30196 7964 30248 8016
rect 32772 7964 32824 8016
rect 34244 7964 34296 8016
rect 35624 7964 35676 8016
rect 24308 7896 24360 7948
rect 26332 7896 26384 7948
rect 27436 7896 27488 7948
rect 28816 7939 28868 7948
rect 28816 7905 28825 7939
rect 28825 7905 28859 7939
rect 28859 7905 28868 7939
rect 28816 7896 28868 7905
rect 29092 7896 29144 7948
rect 13360 7828 13412 7880
rect 13912 7828 13964 7880
rect 16212 7828 16264 7880
rect 17500 7828 17552 7880
rect 18236 7828 18288 7880
rect 19708 7871 19760 7880
rect 19708 7837 19717 7871
rect 19717 7837 19751 7871
rect 19751 7837 19760 7871
rect 19708 7828 19760 7837
rect 25228 7871 25280 7880
rect 25228 7837 25237 7871
rect 25237 7837 25271 7871
rect 25271 7837 25280 7871
rect 25228 7828 25280 7837
rect 26700 7828 26752 7880
rect 26976 7828 27028 7880
rect 12440 7760 12492 7812
rect 6276 7692 6328 7744
rect 6736 7692 6788 7744
rect 7564 7692 7616 7744
rect 8760 7692 8812 7744
rect 10968 7692 11020 7744
rect 13084 7735 13136 7744
rect 13084 7701 13093 7735
rect 13093 7701 13127 7735
rect 13127 7701 13136 7735
rect 13084 7692 13136 7701
rect 13268 7692 13320 7744
rect 13636 7735 13688 7744
rect 13636 7701 13645 7735
rect 13645 7701 13679 7735
rect 13679 7701 13688 7735
rect 13636 7692 13688 7701
rect 14464 7735 14516 7744
rect 14464 7701 14473 7735
rect 14473 7701 14507 7735
rect 14507 7701 14516 7735
rect 14464 7692 14516 7701
rect 15752 7760 15804 7812
rect 16672 7735 16724 7744
rect 16672 7701 16681 7735
rect 16681 7701 16715 7735
rect 16715 7701 16724 7735
rect 16672 7692 16724 7701
rect 18880 7760 18932 7812
rect 22284 7692 22336 7744
rect 22468 7735 22520 7744
rect 22468 7701 22477 7735
rect 22477 7701 22511 7735
rect 22511 7701 22520 7735
rect 22468 7692 22520 7701
rect 23296 7735 23348 7744
rect 23296 7701 23305 7735
rect 23305 7701 23339 7735
rect 23339 7701 23348 7735
rect 23296 7692 23348 7701
rect 24860 7760 24912 7812
rect 26240 7803 26292 7812
rect 26240 7769 26249 7803
rect 26249 7769 26283 7803
rect 26283 7769 26292 7803
rect 26240 7760 26292 7769
rect 25320 7692 25372 7744
rect 25780 7692 25832 7744
rect 25872 7692 25924 7744
rect 27988 7692 28040 7744
rect 28448 7735 28500 7744
rect 28448 7701 28457 7735
rect 28457 7701 28491 7735
rect 28491 7701 28500 7735
rect 28448 7692 28500 7701
rect 29092 7760 29144 7812
rect 29920 7896 29972 7948
rect 31208 7896 31260 7948
rect 32496 7896 32548 7948
rect 34704 7896 34756 7948
rect 29460 7828 29512 7880
rect 29828 7828 29880 7880
rect 33692 7828 33744 7880
rect 33784 7871 33836 7880
rect 33784 7837 33793 7871
rect 33793 7837 33827 7871
rect 33827 7837 33836 7871
rect 33784 7828 33836 7837
rect 34244 7828 34296 7880
rect 38016 7964 38068 8016
rect 38476 7964 38528 8016
rect 43536 8041 43545 8075
rect 43545 8041 43579 8075
rect 43579 8041 43588 8075
rect 43536 8032 43588 8041
rect 44272 8032 44324 8084
rect 44456 8032 44508 8084
rect 45468 8032 45520 8084
rect 45744 8075 45796 8084
rect 45744 8041 45753 8075
rect 45753 8041 45787 8075
rect 45787 8041 45796 8075
rect 45744 8032 45796 8041
rect 39120 7896 39172 7948
rect 40316 7896 40368 7948
rect 41696 7896 41748 7948
rect 43628 7964 43680 8016
rect 45100 7964 45152 8016
rect 45652 7964 45704 8016
rect 44824 7939 44876 7948
rect 44824 7905 44833 7939
rect 44833 7905 44867 7939
rect 44867 7905 44876 7939
rect 44824 7896 44876 7905
rect 45192 7939 45244 7948
rect 45192 7905 45201 7939
rect 45201 7905 45235 7939
rect 45235 7905 45244 7939
rect 45192 7896 45244 7905
rect 47032 8032 47084 8084
rect 47308 8032 47360 8084
rect 50344 8032 50396 8084
rect 51080 8032 51132 8084
rect 51356 8075 51408 8084
rect 51356 8041 51365 8075
rect 51365 8041 51399 8075
rect 51399 8041 51408 8075
rect 51356 8032 51408 8041
rect 52184 8032 52236 8084
rect 53380 8032 53432 8084
rect 53932 8075 53984 8084
rect 53932 8041 53941 8075
rect 53941 8041 53975 8075
rect 53975 8041 53984 8075
rect 53932 8032 53984 8041
rect 55128 8075 55180 8084
rect 55128 8041 55137 8075
rect 55137 8041 55171 8075
rect 55171 8041 55180 8075
rect 55128 8032 55180 8041
rect 55312 8032 55364 8084
rect 53840 7964 53892 8016
rect 57612 8032 57664 8084
rect 58164 8032 58216 8084
rect 58440 8032 58492 8084
rect 59268 8032 59320 8084
rect 47400 7896 47452 7948
rect 47676 7939 47728 7948
rect 47676 7905 47685 7939
rect 47685 7905 47719 7939
rect 47719 7905 47728 7939
rect 47676 7896 47728 7905
rect 34980 7828 35032 7880
rect 35716 7828 35768 7880
rect 35900 7871 35952 7880
rect 35900 7837 35909 7871
rect 35909 7837 35943 7871
rect 35943 7837 35952 7871
rect 35900 7828 35952 7837
rect 39304 7871 39356 7880
rect 39304 7837 39313 7871
rect 39313 7837 39347 7871
rect 39347 7837 39356 7871
rect 39304 7828 39356 7837
rect 39672 7871 39724 7880
rect 39672 7837 39681 7871
rect 39681 7837 39715 7871
rect 39715 7837 39724 7871
rect 39672 7828 39724 7837
rect 41972 7828 42024 7880
rect 42248 7871 42300 7880
rect 42248 7837 42257 7871
rect 42257 7837 42291 7871
rect 42291 7837 42300 7871
rect 42248 7828 42300 7837
rect 44272 7828 44324 7880
rect 44732 7871 44784 7880
rect 44732 7837 44741 7871
rect 44741 7837 44775 7871
rect 44775 7837 44784 7871
rect 44732 7828 44784 7837
rect 46940 7828 46992 7880
rect 48780 7896 48832 7948
rect 49148 7939 49200 7948
rect 49148 7905 49157 7939
rect 49157 7905 49191 7939
rect 49191 7905 49200 7939
rect 49148 7896 49200 7905
rect 48136 7828 48188 7880
rect 52000 7939 52052 7948
rect 49792 7828 49844 7880
rect 49884 7828 49936 7880
rect 50252 7828 50304 7880
rect 38292 7760 38344 7812
rect 38752 7760 38804 7812
rect 39212 7760 39264 7812
rect 29368 7692 29420 7744
rect 29920 7692 29972 7744
rect 31208 7735 31260 7744
rect 31208 7701 31217 7735
rect 31217 7701 31251 7735
rect 31251 7701 31260 7735
rect 31208 7692 31260 7701
rect 31484 7735 31536 7744
rect 31484 7701 31493 7735
rect 31493 7701 31527 7735
rect 31527 7701 31536 7735
rect 31484 7692 31536 7701
rect 33968 7692 34020 7744
rect 34520 7692 34572 7744
rect 39764 7692 39816 7744
rect 40868 7735 40920 7744
rect 40868 7701 40877 7735
rect 40877 7701 40911 7735
rect 40911 7701 40920 7735
rect 40868 7692 40920 7701
rect 41604 7760 41656 7812
rect 47492 7760 47544 7812
rect 47676 7760 47728 7812
rect 47952 7760 48004 7812
rect 48412 7760 48464 7812
rect 48596 7760 48648 7812
rect 50712 7871 50764 7880
rect 50712 7837 50721 7871
rect 50721 7837 50755 7871
rect 50755 7837 50764 7871
rect 52000 7905 52009 7939
rect 52009 7905 52043 7939
rect 52043 7905 52052 7939
rect 52000 7896 52052 7905
rect 52460 7896 52512 7948
rect 53748 7896 53800 7948
rect 56140 7939 56192 7948
rect 56140 7905 56149 7939
rect 56149 7905 56183 7939
rect 56183 7905 56192 7939
rect 56140 7896 56192 7905
rect 59084 7964 59136 8016
rect 50712 7828 50764 7837
rect 51908 7871 51960 7880
rect 51908 7837 51917 7871
rect 51917 7837 51951 7871
rect 51951 7837 51960 7871
rect 51908 7828 51960 7837
rect 55404 7828 55456 7880
rect 56692 7896 56744 7948
rect 58164 7939 58216 7948
rect 58164 7905 58173 7939
rect 58173 7905 58207 7939
rect 58207 7905 58216 7939
rect 58164 7896 58216 7905
rect 58256 7939 58308 7948
rect 58256 7905 58265 7939
rect 58265 7905 58299 7939
rect 58299 7905 58308 7939
rect 58256 7896 58308 7905
rect 58716 7939 58768 7948
rect 57520 7828 57572 7880
rect 58716 7905 58725 7939
rect 58725 7905 58759 7939
rect 58759 7905 58768 7939
rect 58716 7896 58768 7905
rect 60924 7939 60976 7948
rect 60924 7905 60933 7939
rect 60933 7905 60967 7939
rect 60967 7905 60976 7939
rect 60924 7896 60976 7905
rect 55956 7803 56008 7812
rect 55956 7769 55965 7803
rect 55965 7769 55999 7803
rect 55999 7769 56008 7803
rect 55956 7760 56008 7769
rect 56324 7760 56376 7812
rect 59452 7760 59504 7812
rect 41880 7692 41932 7744
rect 42432 7692 42484 7744
rect 43076 7735 43128 7744
rect 43076 7701 43085 7735
rect 43085 7701 43119 7735
rect 43119 7701 43128 7735
rect 43076 7692 43128 7701
rect 46204 7735 46256 7744
rect 46204 7701 46213 7735
rect 46213 7701 46247 7735
rect 46247 7701 46256 7735
rect 46204 7692 46256 7701
rect 46664 7692 46716 7744
rect 48228 7735 48280 7744
rect 48228 7701 48237 7735
rect 48237 7701 48271 7735
rect 48271 7701 48280 7735
rect 48228 7692 48280 7701
rect 49608 7692 49660 7744
rect 50620 7735 50672 7744
rect 50620 7701 50629 7735
rect 50629 7701 50663 7735
rect 50663 7701 50672 7735
rect 50620 7692 50672 7701
rect 51172 7692 51224 7744
rect 53288 7692 53340 7744
rect 54300 7692 54352 7744
rect 55864 7692 55916 7744
rect 59636 7692 59688 7744
rect 11378 7590 11430 7642
rect 11442 7590 11494 7642
rect 11506 7590 11558 7642
rect 11570 7590 11622 7642
rect 32170 7590 32222 7642
rect 32234 7590 32286 7642
rect 32298 7590 32350 7642
rect 32362 7590 32414 7642
rect 52962 7590 53014 7642
rect 53026 7590 53078 7642
rect 53090 7590 53142 7642
rect 53154 7590 53206 7642
rect 4344 7531 4396 7540
rect 4344 7497 4353 7531
rect 4353 7497 4387 7531
rect 4387 7497 4396 7531
rect 4344 7488 4396 7497
rect 8852 7488 8904 7540
rect 7748 7420 7800 7472
rect 8760 7463 8812 7472
rect 8760 7429 8769 7463
rect 8769 7429 8803 7463
rect 8803 7429 8812 7463
rect 8760 7420 8812 7429
rect 5448 7395 5500 7404
rect 5448 7361 5457 7395
rect 5457 7361 5491 7395
rect 5491 7361 5500 7395
rect 5448 7352 5500 7361
rect 6276 7395 6328 7404
rect 6276 7361 6285 7395
rect 6285 7361 6319 7395
rect 6319 7361 6328 7395
rect 6276 7352 6328 7361
rect 6736 7352 6788 7404
rect 6552 7284 6604 7336
rect 7104 7284 7156 7336
rect 4896 7259 4948 7268
rect 4896 7225 4905 7259
rect 4905 7225 4939 7259
rect 4939 7225 4948 7259
rect 4896 7216 4948 7225
rect 7748 7284 7800 7336
rect 7932 7327 7984 7336
rect 7932 7293 7941 7327
rect 7941 7293 7975 7327
rect 7975 7293 7984 7327
rect 7932 7284 7984 7293
rect 8208 7216 8260 7268
rect 3700 7191 3752 7200
rect 3700 7157 3709 7191
rect 3709 7157 3743 7191
rect 3743 7157 3752 7191
rect 3700 7148 3752 7157
rect 4068 7148 4120 7200
rect 5540 7148 5592 7200
rect 6828 7148 6880 7200
rect 12532 7488 12584 7540
rect 13360 7463 13412 7472
rect 12532 7352 12584 7404
rect 13084 7395 13136 7404
rect 13084 7361 13093 7395
rect 13093 7361 13127 7395
rect 13127 7361 13136 7395
rect 13084 7352 13136 7361
rect 10232 7284 10284 7336
rect 12348 7284 12400 7336
rect 12440 7327 12492 7336
rect 12440 7293 12449 7327
rect 12449 7293 12483 7327
rect 12483 7293 12492 7327
rect 12440 7284 12492 7293
rect 9956 7148 10008 7200
rect 13360 7429 13369 7463
rect 13369 7429 13403 7463
rect 13403 7429 13412 7463
rect 13360 7420 13412 7429
rect 16764 7488 16816 7540
rect 18236 7531 18288 7540
rect 18236 7497 18245 7531
rect 18245 7497 18279 7531
rect 18279 7497 18288 7531
rect 18236 7488 18288 7497
rect 20904 7488 20956 7540
rect 23480 7531 23532 7540
rect 23480 7497 23489 7531
rect 23489 7497 23523 7531
rect 23523 7497 23532 7531
rect 23480 7488 23532 7497
rect 25320 7488 25372 7540
rect 26516 7488 26568 7540
rect 28724 7531 28776 7540
rect 28724 7497 28733 7531
rect 28733 7497 28767 7531
rect 28767 7497 28776 7531
rect 28724 7488 28776 7497
rect 28816 7488 28868 7540
rect 24768 7420 24820 7472
rect 13544 7352 13596 7404
rect 15292 7352 15344 7404
rect 15752 7395 15804 7404
rect 15752 7361 15761 7395
rect 15761 7361 15795 7395
rect 15795 7361 15804 7395
rect 15752 7352 15804 7361
rect 17224 7352 17276 7404
rect 29828 7420 29880 7472
rect 30196 7488 30248 7540
rect 31024 7531 31076 7540
rect 31024 7497 31033 7531
rect 31033 7497 31067 7531
rect 31067 7497 31076 7531
rect 31024 7488 31076 7497
rect 33876 7531 33928 7540
rect 33876 7497 33885 7531
rect 33885 7497 33919 7531
rect 33919 7497 33928 7531
rect 33876 7488 33928 7497
rect 34612 7488 34664 7540
rect 41696 7531 41748 7540
rect 41696 7497 41705 7531
rect 41705 7497 41739 7531
rect 41739 7497 41748 7531
rect 41696 7488 41748 7497
rect 41972 7488 42024 7540
rect 42800 7488 42852 7540
rect 44732 7531 44784 7540
rect 44732 7497 44741 7531
rect 44741 7497 44775 7531
rect 44775 7497 44784 7531
rect 44732 7488 44784 7497
rect 44824 7488 44876 7540
rect 35900 7420 35952 7472
rect 39672 7420 39724 7472
rect 45560 7420 45612 7472
rect 46480 7463 46532 7472
rect 46480 7429 46489 7463
rect 46489 7429 46523 7463
rect 46523 7429 46532 7463
rect 46480 7420 46532 7429
rect 46664 7488 46716 7540
rect 47492 7488 47544 7540
rect 47676 7488 47728 7540
rect 51632 7488 51684 7540
rect 52000 7488 52052 7540
rect 53748 7531 53800 7540
rect 52552 7420 52604 7472
rect 28448 7352 28500 7404
rect 29000 7352 29052 7404
rect 14188 7284 14240 7336
rect 14464 7284 14516 7336
rect 16304 7284 16356 7336
rect 16672 7327 16724 7336
rect 16672 7293 16681 7327
rect 16681 7293 16715 7327
rect 16715 7293 16724 7327
rect 16672 7284 16724 7293
rect 17684 7284 17736 7336
rect 18144 7284 18196 7336
rect 18880 7284 18932 7336
rect 19708 7284 19760 7336
rect 10876 7148 10928 7200
rect 11888 7191 11940 7200
rect 11888 7157 11897 7191
rect 11897 7157 11931 7191
rect 11931 7157 11940 7191
rect 11888 7148 11940 7157
rect 12256 7191 12308 7200
rect 12256 7157 12265 7191
rect 12265 7157 12299 7191
rect 12299 7157 12308 7191
rect 12256 7148 12308 7157
rect 16212 7191 16264 7200
rect 16212 7157 16221 7191
rect 16221 7157 16255 7191
rect 16255 7157 16264 7191
rect 16212 7148 16264 7157
rect 17500 7216 17552 7268
rect 19524 7216 19576 7268
rect 20076 7284 20128 7336
rect 21180 7327 21232 7336
rect 21180 7293 21189 7327
rect 21189 7293 21223 7327
rect 21223 7293 21232 7327
rect 21180 7284 21232 7293
rect 21548 7284 21600 7336
rect 22100 7284 22152 7336
rect 23848 7284 23900 7336
rect 24308 7327 24360 7336
rect 24308 7293 24317 7327
rect 24317 7293 24351 7327
rect 24351 7293 24360 7327
rect 24308 7284 24360 7293
rect 18604 7148 18656 7200
rect 18788 7191 18840 7200
rect 18788 7157 18797 7191
rect 18797 7157 18831 7191
rect 18831 7157 18840 7191
rect 18788 7148 18840 7157
rect 18880 7148 18932 7200
rect 20076 7148 20128 7200
rect 20260 7216 20312 7268
rect 20812 7191 20864 7200
rect 20812 7157 20821 7191
rect 20821 7157 20855 7191
rect 20855 7157 20864 7191
rect 20812 7148 20864 7157
rect 22284 7216 22336 7268
rect 24492 7327 24544 7336
rect 24492 7293 24501 7327
rect 24501 7293 24535 7327
rect 24535 7293 24544 7327
rect 24492 7284 24544 7293
rect 25320 7284 25372 7336
rect 25964 7284 26016 7336
rect 26240 7216 26292 7268
rect 26884 7327 26936 7336
rect 26884 7293 26893 7327
rect 26893 7293 26927 7327
rect 26927 7293 26936 7327
rect 26884 7284 26936 7293
rect 27160 7284 27212 7336
rect 27896 7284 27948 7336
rect 28080 7284 28132 7336
rect 31484 7352 31536 7404
rect 32036 7352 32088 7404
rect 27068 7216 27120 7268
rect 23112 7148 23164 7200
rect 23940 7191 23992 7200
rect 23940 7157 23949 7191
rect 23949 7157 23983 7191
rect 23983 7157 23992 7191
rect 23940 7148 23992 7157
rect 25320 7191 25372 7200
rect 25320 7157 25329 7191
rect 25329 7157 25363 7191
rect 25363 7157 25372 7191
rect 25320 7148 25372 7157
rect 25964 7148 26016 7200
rect 27804 7259 27856 7268
rect 27804 7225 27813 7259
rect 27813 7225 27847 7259
rect 27847 7225 27856 7259
rect 27804 7216 27856 7225
rect 29276 7259 29328 7268
rect 29276 7225 29285 7259
rect 29285 7225 29319 7259
rect 29319 7225 29328 7259
rect 29276 7216 29328 7225
rect 28264 7148 28316 7200
rect 29552 7259 29604 7268
rect 29552 7225 29561 7259
rect 29561 7225 29595 7259
rect 29595 7225 29604 7259
rect 29552 7216 29604 7225
rect 30748 7284 30800 7336
rect 31300 7284 31352 7336
rect 33784 7352 33836 7404
rect 34704 7395 34756 7404
rect 34704 7361 34713 7395
rect 34713 7361 34747 7395
rect 34747 7361 34756 7395
rect 34704 7352 34756 7361
rect 30012 7259 30064 7268
rect 30012 7225 30021 7259
rect 30021 7225 30055 7259
rect 30055 7225 30064 7259
rect 30012 7216 30064 7225
rect 30656 7148 30708 7200
rect 31760 7191 31812 7200
rect 31760 7157 31769 7191
rect 31769 7157 31803 7191
rect 31803 7157 31812 7191
rect 31760 7148 31812 7157
rect 32404 7191 32456 7200
rect 32404 7157 32413 7191
rect 32413 7157 32447 7191
rect 32447 7157 32456 7191
rect 32404 7148 32456 7157
rect 34612 7284 34664 7336
rect 34980 7327 35032 7336
rect 34980 7293 34989 7327
rect 34989 7293 35023 7327
rect 35023 7293 35032 7327
rect 34980 7284 35032 7293
rect 39212 7327 39264 7336
rect 33508 7148 33560 7200
rect 35992 7148 36044 7200
rect 36636 7191 36688 7200
rect 36636 7157 36645 7191
rect 36645 7157 36679 7191
rect 36679 7157 36688 7191
rect 36636 7148 36688 7157
rect 39212 7293 39221 7327
rect 39221 7293 39255 7327
rect 39255 7293 39264 7327
rect 39212 7284 39264 7293
rect 39396 7327 39448 7336
rect 39396 7293 39405 7327
rect 39405 7293 39439 7327
rect 39439 7293 39448 7327
rect 39396 7284 39448 7293
rect 40408 7284 40460 7336
rect 42340 7327 42392 7336
rect 42340 7293 42349 7327
rect 42349 7293 42383 7327
rect 42383 7293 42392 7327
rect 42340 7284 42392 7293
rect 42432 7284 42484 7336
rect 38384 7216 38436 7268
rect 39764 7216 39816 7268
rect 41052 7259 41104 7268
rect 41052 7225 41061 7259
rect 41061 7225 41095 7259
rect 41095 7225 41104 7259
rect 41052 7216 41104 7225
rect 46112 7352 46164 7404
rect 37280 7148 37332 7200
rect 38660 7148 38712 7200
rect 39120 7148 39172 7200
rect 40592 7148 40644 7200
rect 43352 7216 43404 7268
rect 41328 7148 41380 7200
rect 44456 7148 44508 7200
rect 44732 7148 44784 7200
rect 45192 7216 45244 7268
rect 46480 7284 46532 7336
rect 46204 7259 46256 7268
rect 46204 7225 46213 7259
rect 46213 7225 46247 7259
rect 46247 7225 46256 7259
rect 46204 7216 46256 7225
rect 46296 7216 46348 7268
rect 48688 7352 48740 7404
rect 49608 7352 49660 7404
rect 50160 7352 50212 7404
rect 51908 7352 51960 7404
rect 46664 7284 46716 7336
rect 46940 7259 46992 7268
rect 46940 7225 46949 7259
rect 46949 7225 46983 7259
rect 46983 7225 46992 7259
rect 46940 7216 46992 7225
rect 47676 7216 47728 7268
rect 47952 7259 48004 7268
rect 47216 7148 47268 7200
rect 47952 7225 47961 7259
rect 47961 7225 47995 7259
rect 47995 7225 48004 7259
rect 47952 7216 48004 7225
rect 48136 7259 48188 7268
rect 48136 7225 48145 7259
rect 48145 7225 48179 7259
rect 48179 7225 48188 7259
rect 48136 7216 48188 7225
rect 48504 7259 48556 7268
rect 48504 7225 48513 7259
rect 48513 7225 48547 7259
rect 48547 7225 48556 7259
rect 48504 7216 48556 7225
rect 48780 7259 48832 7268
rect 48780 7225 48789 7259
rect 48789 7225 48823 7259
rect 48823 7225 48832 7259
rect 48780 7216 48832 7225
rect 48596 7148 48648 7200
rect 50068 7284 50120 7336
rect 50344 7327 50396 7336
rect 50344 7293 50353 7327
rect 50353 7293 50387 7327
rect 50387 7293 50396 7327
rect 50344 7284 50396 7293
rect 50988 7284 51040 7336
rect 53748 7497 53757 7531
rect 53757 7497 53791 7531
rect 53791 7497 53800 7531
rect 53748 7488 53800 7497
rect 55404 7488 55456 7540
rect 56140 7488 56192 7540
rect 57060 7531 57112 7540
rect 57060 7497 57069 7531
rect 57069 7497 57103 7531
rect 57103 7497 57112 7531
rect 57060 7488 57112 7497
rect 53012 7463 53064 7472
rect 53012 7429 53021 7463
rect 53021 7429 53055 7463
rect 53055 7429 53064 7463
rect 59912 7488 59964 7540
rect 60924 7488 60976 7540
rect 53012 7420 53064 7429
rect 57612 7420 57664 7472
rect 57704 7420 57756 7472
rect 56324 7352 56376 7404
rect 55772 7327 55824 7336
rect 49148 7259 49200 7268
rect 49148 7225 49157 7259
rect 49157 7225 49191 7259
rect 49191 7225 49200 7259
rect 49148 7216 49200 7225
rect 49884 7216 49936 7268
rect 50712 7148 50764 7200
rect 51632 7148 51684 7200
rect 52736 7216 52788 7268
rect 55772 7293 55781 7327
rect 55781 7293 55815 7327
rect 55815 7293 55824 7327
rect 55772 7284 55824 7293
rect 55864 7284 55916 7336
rect 57060 7284 57112 7336
rect 57796 7284 57848 7336
rect 58072 7327 58124 7336
rect 58072 7293 58081 7327
rect 58081 7293 58115 7327
rect 58115 7293 58124 7327
rect 58072 7284 58124 7293
rect 59636 7327 59688 7336
rect 57980 7216 58032 7268
rect 59636 7293 59645 7327
rect 59645 7293 59679 7327
rect 59679 7293 59688 7327
rect 59636 7284 59688 7293
rect 59820 7284 59872 7336
rect 58716 7259 58768 7268
rect 58716 7225 58725 7259
rect 58725 7225 58759 7259
rect 58759 7225 58768 7259
rect 58716 7216 58768 7225
rect 52184 7148 52236 7200
rect 53564 7148 53616 7200
rect 54116 7191 54168 7200
rect 54116 7157 54125 7191
rect 54125 7157 54159 7191
rect 54159 7157 54168 7191
rect 54116 7148 54168 7157
rect 56600 7148 56652 7200
rect 58072 7148 58124 7200
rect 21774 7046 21826 7098
rect 21838 7046 21890 7098
rect 21902 7046 21954 7098
rect 21966 7046 22018 7098
rect 42566 7046 42618 7098
rect 42630 7046 42682 7098
rect 42694 7046 42746 7098
rect 42758 7046 42810 7098
rect 7288 6944 7340 6996
rect 7932 6987 7984 6996
rect 7932 6953 7941 6987
rect 7941 6953 7975 6987
rect 7975 6953 7984 6987
rect 7932 6944 7984 6953
rect 9956 6987 10008 6996
rect 9956 6953 9965 6987
rect 9965 6953 9999 6987
rect 9999 6953 10008 6987
rect 9956 6944 10008 6953
rect 12256 6944 12308 6996
rect 13636 6944 13688 6996
rect 18512 6944 18564 6996
rect 18604 6944 18656 6996
rect 20720 6944 20772 6996
rect 6552 6919 6604 6928
rect 6552 6885 6561 6919
rect 6561 6885 6595 6919
rect 6595 6885 6604 6919
rect 6552 6876 6604 6885
rect 6736 6919 6788 6928
rect 6736 6885 6745 6919
rect 6745 6885 6779 6919
rect 6779 6885 6788 6919
rect 6736 6876 6788 6885
rect 6920 6919 6972 6928
rect 6920 6885 6929 6919
rect 6929 6885 6963 6919
rect 6963 6885 6972 6919
rect 6920 6876 6972 6885
rect 8208 6851 8260 6860
rect 8208 6817 8217 6851
rect 8217 6817 8251 6851
rect 8251 6817 8260 6851
rect 12532 6876 12584 6928
rect 8208 6808 8260 6817
rect 3700 6740 3752 6792
rect 4804 6740 4856 6792
rect 8300 6740 8352 6792
rect 7196 6672 7248 6724
rect 3240 6647 3292 6656
rect 3240 6613 3249 6647
rect 3249 6613 3283 6647
rect 3283 6613 3292 6647
rect 3240 6604 3292 6613
rect 3516 6647 3568 6656
rect 3516 6613 3525 6647
rect 3525 6613 3559 6647
rect 3559 6613 3568 6647
rect 3516 6604 3568 6613
rect 8208 6604 8260 6656
rect 12992 6808 13044 6860
rect 10232 6740 10284 6792
rect 10784 6740 10836 6792
rect 14740 6876 14792 6928
rect 16304 6919 16356 6928
rect 16304 6885 16313 6919
rect 16313 6885 16347 6919
rect 16347 6885 16356 6919
rect 16304 6876 16356 6885
rect 13820 6851 13872 6860
rect 13820 6817 13829 6851
rect 13829 6817 13863 6851
rect 13863 6817 13872 6851
rect 13820 6808 13872 6817
rect 14372 6851 14424 6860
rect 13912 6740 13964 6792
rect 14372 6817 14381 6851
rect 14381 6817 14415 6851
rect 14415 6817 14424 6851
rect 14372 6808 14424 6817
rect 15660 6808 15712 6860
rect 15200 6740 15252 6792
rect 16212 6808 16264 6860
rect 17224 6808 17276 6860
rect 17500 6851 17552 6860
rect 17500 6817 17509 6851
rect 17509 6817 17543 6851
rect 17543 6817 17552 6851
rect 17500 6808 17552 6817
rect 18236 6876 18288 6928
rect 21272 6944 21324 6996
rect 21364 6944 21416 6996
rect 23296 6944 23348 6996
rect 24124 6944 24176 6996
rect 24308 6944 24360 6996
rect 28080 6944 28132 6996
rect 28448 6944 28500 6996
rect 29920 6944 29972 6996
rect 31208 6987 31260 6996
rect 31208 6953 31217 6987
rect 31217 6953 31251 6987
rect 31251 6953 31260 6987
rect 31208 6944 31260 6953
rect 18052 6808 18104 6860
rect 17040 6783 17092 6792
rect 17040 6749 17049 6783
rect 17049 6749 17083 6783
rect 17083 6749 17092 6783
rect 17040 6740 17092 6749
rect 17132 6740 17184 6792
rect 11244 6604 11296 6656
rect 11704 6604 11756 6656
rect 15936 6672 15988 6724
rect 18144 6672 18196 6724
rect 14188 6604 14240 6656
rect 16120 6647 16172 6656
rect 16120 6613 16129 6647
rect 16129 6613 16163 6647
rect 16163 6613 16172 6647
rect 16120 6604 16172 6613
rect 16212 6604 16264 6656
rect 17132 6604 17184 6656
rect 17224 6604 17276 6656
rect 18236 6647 18288 6656
rect 18236 6613 18245 6647
rect 18245 6613 18279 6647
rect 18279 6613 18288 6647
rect 18236 6604 18288 6613
rect 19064 6851 19116 6860
rect 19064 6817 19073 6851
rect 19073 6817 19107 6851
rect 19107 6817 19116 6851
rect 19064 6808 19116 6817
rect 19248 6808 19300 6860
rect 19524 6851 19576 6860
rect 19524 6817 19533 6851
rect 19533 6817 19567 6851
rect 19567 6817 19576 6851
rect 19524 6808 19576 6817
rect 20076 6808 20128 6860
rect 20628 6808 20680 6860
rect 22560 6851 22612 6860
rect 22560 6817 22569 6851
rect 22569 6817 22603 6851
rect 22603 6817 22612 6851
rect 22560 6808 22612 6817
rect 22652 6851 22704 6860
rect 22652 6817 22661 6851
rect 22661 6817 22695 6851
rect 22695 6817 22704 6851
rect 22652 6808 22704 6817
rect 24032 6808 24084 6860
rect 24308 6808 24360 6860
rect 26516 6876 26568 6928
rect 21824 6783 21876 6792
rect 19340 6672 19392 6724
rect 21824 6749 21833 6783
rect 21833 6749 21867 6783
rect 21867 6749 21876 6783
rect 21824 6740 21876 6749
rect 24860 6740 24912 6792
rect 25320 6808 25372 6860
rect 26700 6851 26752 6860
rect 26700 6817 26709 6851
rect 26709 6817 26743 6851
rect 26743 6817 26752 6851
rect 26700 6808 26752 6817
rect 23756 6672 23808 6724
rect 24676 6672 24728 6724
rect 25412 6740 25464 6792
rect 25780 6740 25832 6792
rect 26332 6783 26384 6792
rect 26332 6749 26341 6783
rect 26341 6749 26375 6783
rect 26375 6749 26384 6783
rect 27068 6808 27120 6860
rect 27160 6851 27212 6860
rect 27160 6817 27169 6851
rect 27169 6817 27203 6851
rect 27203 6817 27212 6851
rect 28264 6876 28316 6928
rect 28540 6876 28592 6928
rect 29000 6876 29052 6928
rect 29092 6876 29144 6928
rect 33416 6944 33468 6996
rect 38752 6944 38804 6996
rect 39028 6944 39080 6996
rect 39672 6987 39724 6996
rect 39672 6953 39681 6987
rect 39681 6953 39715 6987
rect 39715 6953 39724 6987
rect 39672 6944 39724 6953
rect 39856 6944 39908 6996
rect 45192 6944 45244 6996
rect 34520 6876 34572 6928
rect 27160 6808 27212 6817
rect 27436 6808 27488 6860
rect 28724 6808 28776 6860
rect 29460 6851 29512 6860
rect 26332 6740 26384 6749
rect 28264 6740 28316 6792
rect 29460 6817 29469 6851
rect 29469 6817 29503 6851
rect 29503 6817 29512 6851
rect 29460 6808 29512 6817
rect 30012 6808 30064 6860
rect 30564 6808 30616 6860
rect 31300 6808 31352 6860
rect 29092 6740 29144 6792
rect 32956 6808 33008 6860
rect 32496 6740 32548 6792
rect 33416 6740 33468 6792
rect 33692 6740 33744 6792
rect 34244 6740 34296 6792
rect 36912 6851 36964 6860
rect 36912 6817 36921 6851
rect 36921 6817 36955 6851
rect 36955 6817 36964 6851
rect 36912 6808 36964 6817
rect 38384 6851 38436 6860
rect 38384 6817 38393 6851
rect 38393 6817 38427 6851
rect 38427 6817 38436 6851
rect 38384 6808 38436 6817
rect 38752 6851 38804 6860
rect 38752 6817 38761 6851
rect 38761 6817 38795 6851
rect 38795 6817 38804 6851
rect 38752 6808 38804 6817
rect 25136 6672 25188 6724
rect 26240 6672 26292 6724
rect 26884 6672 26936 6724
rect 28816 6672 28868 6724
rect 19892 6604 19944 6656
rect 20168 6647 20220 6656
rect 20168 6613 20177 6647
rect 20177 6613 20211 6647
rect 20211 6613 20220 6647
rect 20168 6604 20220 6613
rect 20536 6604 20588 6656
rect 22468 6604 22520 6656
rect 22836 6647 22888 6656
rect 22836 6613 22845 6647
rect 22845 6613 22879 6647
rect 22879 6613 22888 6647
rect 22836 6604 22888 6613
rect 22928 6604 22980 6656
rect 24308 6647 24360 6656
rect 24308 6613 24317 6647
rect 24317 6613 24351 6647
rect 24351 6613 24360 6647
rect 24308 6604 24360 6613
rect 24860 6647 24912 6656
rect 24860 6613 24869 6647
rect 24869 6613 24903 6647
rect 24903 6613 24912 6647
rect 24860 6604 24912 6613
rect 28632 6604 28684 6656
rect 29552 6672 29604 6724
rect 31668 6672 31720 6724
rect 35900 6740 35952 6792
rect 37280 6783 37332 6792
rect 37280 6749 37289 6783
rect 37289 6749 37323 6783
rect 37323 6749 37332 6783
rect 37280 6740 37332 6749
rect 38476 6740 38528 6792
rect 39764 6876 39816 6928
rect 39396 6808 39448 6860
rect 43076 6876 43128 6928
rect 46940 6944 46992 6996
rect 48596 6944 48648 6996
rect 50988 6944 51040 6996
rect 51632 6944 51684 6996
rect 54208 6944 54260 6996
rect 45560 6876 45612 6928
rect 45652 6876 45704 6928
rect 41604 6851 41656 6860
rect 41604 6817 41613 6851
rect 41613 6817 41647 6851
rect 41647 6817 41656 6851
rect 41604 6808 41656 6817
rect 41788 6808 41840 6860
rect 43352 6808 43404 6860
rect 44640 6808 44692 6860
rect 46204 6808 46256 6860
rect 47400 6876 47452 6928
rect 54116 6876 54168 6928
rect 55036 6876 55088 6928
rect 42984 6740 43036 6792
rect 36452 6672 36504 6724
rect 36544 6672 36596 6724
rect 38660 6672 38712 6724
rect 38752 6672 38804 6724
rect 39212 6715 39264 6724
rect 39212 6681 39221 6715
rect 39221 6681 39255 6715
rect 39255 6681 39264 6715
rect 39212 6672 39264 6681
rect 39304 6672 39356 6724
rect 44732 6740 44784 6792
rect 46388 6740 46440 6792
rect 46664 6740 46716 6792
rect 48412 6808 48464 6860
rect 48596 6851 48648 6860
rect 48596 6817 48605 6851
rect 48605 6817 48639 6851
rect 48639 6817 48648 6851
rect 48596 6808 48648 6817
rect 49700 6808 49752 6860
rect 49884 6808 49936 6860
rect 50344 6808 50396 6860
rect 50712 6808 50764 6860
rect 50988 6808 51040 6860
rect 52460 6851 52512 6860
rect 52460 6817 52469 6851
rect 52469 6817 52503 6851
rect 52503 6817 52512 6851
rect 52460 6808 52512 6817
rect 30380 6604 30432 6656
rect 30932 6604 30984 6656
rect 31944 6647 31996 6656
rect 31944 6613 31953 6647
rect 31953 6613 31987 6647
rect 31987 6613 31996 6647
rect 31944 6604 31996 6613
rect 32588 6604 32640 6656
rect 35624 6647 35676 6656
rect 35624 6613 35633 6647
rect 35633 6613 35667 6647
rect 35667 6613 35676 6647
rect 35624 6604 35676 6613
rect 39764 6647 39816 6656
rect 39764 6613 39773 6647
rect 39773 6613 39807 6647
rect 39807 6613 39816 6647
rect 39764 6604 39816 6613
rect 45100 6672 45152 6724
rect 47216 6783 47268 6792
rect 47216 6749 47225 6783
rect 47225 6749 47259 6783
rect 47259 6749 47268 6783
rect 47216 6740 47268 6749
rect 47400 6740 47452 6792
rect 52184 6783 52236 6792
rect 52184 6749 52193 6783
rect 52193 6749 52227 6783
rect 52227 6749 52236 6783
rect 52184 6740 52236 6749
rect 46940 6672 46992 6724
rect 41880 6604 41932 6656
rect 42524 6647 42576 6656
rect 42524 6613 42533 6647
rect 42533 6613 42567 6647
rect 42567 6613 42576 6647
rect 42524 6604 42576 6613
rect 44180 6604 44232 6656
rect 46112 6604 46164 6656
rect 47492 6604 47544 6656
rect 47952 6604 48004 6656
rect 49608 6647 49660 6656
rect 49608 6613 49617 6647
rect 49617 6613 49651 6647
rect 49651 6613 49660 6647
rect 49608 6604 49660 6613
rect 51172 6672 51224 6724
rect 53288 6808 53340 6860
rect 54944 6851 54996 6860
rect 53840 6740 53892 6792
rect 54944 6817 54953 6851
rect 54953 6817 54987 6851
rect 54987 6817 54996 6851
rect 54944 6808 54996 6817
rect 56600 6944 56652 6996
rect 57704 6944 57756 6996
rect 57612 6876 57664 6928
rect 55956 6740 56008 6792
rect 57336 6808 57388 6860
rect 57520 6851 57572 6860
rect 57520 6817 57529 6851
rect 57529 6817 57563 6851
rect 57563 6817 57572 6851
rect 57520 6808 57572 6817
rect 57796 6808 57848 6860
rect 59728 6876 59780 6928
rect 57980 6740 58032 6792
rect 58256 6740 58308 6792
rect 59636 6808 59688 6860
rect 59912 6851 59964 6860
rect 59912 6817 59921 6851
rect 59921 6817 59955 6851
rect 59955 6817 59964 6851
rect 59912 6808 59964 6817
rect 60648 6808 60700 6860
rect 60004 6740 60056 6792
rect 61292 6740 61344 6792
rect 61568 6783 61620 6792
rect 61568 6749 61577 6783
rect 61577 6749 61611 6783
rect 61611 6749 61620 6783
rect 61568 6740 61620 6749
rect 58532 6672 58584 6724
rect 53288 6647 53340 6656
rect 53288 6613 53297 6647
rect 53297 6613 53331 6647
rect 53331 6613 53340 6647
rect 53288 6604 53340 6613
rect 54024 6647 54076 6656
rect 54024 6613 54033 6647
rect 54033 6613 54067 6647
rect 54067 6613 54076 6647
rect 54024 6604 54076 6613
rect 55588 6604 55640 6656
rect 55864 6647 55916 6656
rect 55864 6613 55873 6647
rect 55873 6613 55907 6647
rect 55907 6613 55916 6647
rect 55864 6604 55916 6613
rect 55956 6604 56008 6656
rect 56140 6604 56192 6656
rect 57612 6604 57664 6656
rect 58808 6604 58860 6656
rect 11378 6502 11430 6554
rect 11442 6502 11494 6554
rect 11506 6502 11558 6554
rect 11570 6502 11622 6554
rect 32170 6502 32222 6554
rect 32234 6502 32286 6554
rect 32298 6502 32350 6554
rect 32362 6502 32414 6554
rect 52962 6502 53014 6554
rect 53026 6502 53078 6554
rect 53090 6502 53142 6554
rect 53154 6502 53206 6554
rect 4896 6400 4948 6452
rect 6920 6400 6972 6452
rect 7380 6400 7432 6452
rect 9312 6400 9364 6452
rect 13912 6400 13964 6452
rect 3516 6307 3568 6316
rect 3516 6273 3525 6307
rect 3525 6273 3559 6307
rect 3559 6273 3568 6307
rect 3516 6264 3568 6273
rect 6736 6264 6788 6316
rect 12716 6332 12768 6384
rect 16028 6332 16080 6384
rect 16304 6332 16356 6384
rect 20168 6400 20220 6452
rect 20720 6400 20772 6452
rect 18052 6332 18104 6384
rect 19984 6375 20036 6384
rect 19984 6341 19993 6375
rect 19993 6341 20027 6375
rect 20027 6341 20036 6375
rect 19984 6332 20036 6341
rect 3240 6239 3292 6248
rect 2320 6060 2372 6112
rect 3240 6205 3249 6239
rect 3249 6205 3283 6239
rect 3283 6205 3292 6239
rect 3240 6196 3292 6205
rect 10140 6307 10192 6316
rect 8116 6196 8168 6248
rect 7196 6128 7248 6180
rect 8208 6128 8260 6180
rect 9220 6196 9272 6248
rect 10140 6273 10149 6307
rect 10149 6273 10183 6307
rect 10183 6273 10192 6307
rect 10140 6264 10192 6273
rect 10784 6307 10836 6316
rect 10784 6273 10793 6307
rect 10793 6273 10827 6307
rect 10827 6273 10836 6307
rect 10784 6264 10836 6273
rect 9772 6196 9824 6248
rect 11060 6239 11112 6248
rect 11060 6205 11069 6239
rect 11069 6205 11103 6239
rect 11103 6205 11112 6239
rect 11060 6196 11112 6205
rect 11980 6196 12032 6248
rect 6644 6060 6696 6112
rect 8300 6060 8352 6112
rect 9312 6060 9364 6112
rect 9496 6060 9548 6112
rect 12440 6128 12492 6180
rect 14372 6264 14424 6316
rect 15016 6239 15068 6248
rect 13544 6128 13596 6180
rect 15016 6205 15025 6239
rect 15025 6205 15059 6239
rect 15059 6205 15068 6239
rect 15016 6196 15068 6205
rect 15752 6196 15804 6248
rect 16120 6239 16172 6248
rect 16120 6205 16129 6239
rect 16129 6205 16163 6239
rect 16163 6205 16172 6239
rect 16120 6196 16172 6205
rect 15200 6128 15252 6180
rect 15936 6128 15988 6180
rect 16764 6196 16816 6248
rect 18236 6264 18288 6316
rect 19432 6264 19484 6316
rect 20536 6332 20588 6384
rect 25780 6400 25832 6452
rect 31944 6400 31996 6452
rect 33876 6443 33928 6452
rect 33876 6409 33885 6443
rect 33885 6409 33919 6443
rect 33919 6409 33928 6443
rect 33876 6400 33928 6409
rect 22928 6332 22980 6384
rect 24032 6332 24084 6384
rect 12532 6060 12584 6112
rect 13176 6060 13228 6112
rect 13820 6060 13872 6112
rect 14648 6060 14700 6112
rect 15016 6060 15068 6112
rect 16120 6060 16172 6112
rect 17132 6060 17184 6112
rect 17408 6103 17460 6112
rect 17408 6069 17417 6103
rect 17417 6069 17451 6103
rect 17451 6069 17460 6103
rect 17408 6060 17460 6069
rect 17960 6196 18012 6248
rect 18696 6196 18748 6248
rect 19064 6239 19116 6248
rect 19064 6205 19073 6239
rect 19073 6205 19107 6239
rect 19107 6205 19116 6239
rect 19064 6196 19116 6205
rect 19340 6196 19392 6248
rect 22652 6264 22704 6316
rect 24860 6332 24912 6384
rect 28356 6332 28408 6384
rect 31484 6332 31536 6384
rect 20168 6196 20220 6248
rect 20536 6239 20588 6248
rect 20536 6205 20545 6239
rect 20545 6205 20579 6239
rect 20579 6205 20588 6239
rect 20536 6196 20588 6205
rect 20628 6196 20680 6248
rect 21640 6239 21692 6248
rect 21640 6205 21649 6239
rect 21649 6205 21683 6239
rect 21683 6205 21692 6239
rect 21640 6196 21692 6205
rect 23756 6196 23808 6248
rect 18052 6171 18104 6180
rect 18052 6137 18061 6171
rect 18061 6137 18095 6171
rect 18095 6137 18104 6171
rect 18052 6128 18104 6137
rect 18236 6128 18288 6180
rect 20904 6060 20956 6112
rect 21824 6128 21876 6180
rect 24584 6264 24636 6316
rect 25136 6264 25188 6316
rect 26516 6264 26568 6316
rect 25320 6239 25372 6248
rect 25320 6205 25329 6239
rect 25329 6205 25363 6239
rect 25363 6205 25372 6239
rect 25320 6196 25372 6205
rect 25596 6196 25648 6248
rect 25872 6196 25924 6248
rect 27620 6264 27672 6316
rect 27068 6196 27120 6248
rect 28448 6264 28500 6316
rect 28724 6307 28776 6316
rect 28724 6273 28733 6307
rect 28733 6273 28767 6307
rect 28767 6273 28776 6307
rect 28724 6264 28776 6273
rect 29552 6307 29604 6316
rect 29552 6273 29561 6307
rect 29561 6273 29595 6307
rect 29595 6273 29604 6307
rect 29552 6264 29604 6273
rect 31668 6264 31720 6316
rect 34888 6375 34940 6384
rect 34888 6341 34897 6375
rect 34897 6341 34931 6375
rect 34931 6341 34940 6375
rect 37924 6375 37976 6384
rect 34888 6332 34940 6341
rect 35532 6264 35584 6316
rect 27804 6196 27856 6248
rect 30012 6196 30064 6248
rect 31300 6239 31352 6248
rect 31300 6205 31309 6239
rect 31309 6205 31343 6239
rect 31343 6205 31352 6239
rect 31300 6196 31352 6205
rect 32036 6239 32088 6248
rect 24860 6128 24912 6180
rect 28264 6171 28316 6180
rect 28264 6137 28273 6171
rect 28273 6137 28307 6171
rect 28307 6137 28316 6171
rect 28264 6128 28316 6137
rect 28816 6128 28868 6180
rect 29092 6171 29144 6180
rect 29092 6137 29101 6171
rect 29101 6137 29135 6171
rect 29135 6137 29144 6171
rect 29092 6128 29144 6137
rect 31668 6128 31720 6180
rect 23664 6060 23716 6112
rect 24492 6060 24544 6112
rect 26792 6060 26844 6112
rect 27712 6060 27764 6112
rect 31392 6060 31444 6112
rect 31484 6060 31536 6112
rect 32036 6205 32045 6239
rect 32045 6205 32079 6239
rect 32079 6205 32088 6239
rect 32036 6196 32088 6205
rect 31944 6128 31996 6180
rect 34244 6239 34296 6248
rect 34244 6205 34253 6239
rect 34253 6205 34287 6239
rect 34287 6205 34296 6239
rect 34244 6196 34296 6205
rect 35624 6239 35676 6248
rect 35624 6205 35633 6239
rect 35633 6205 35667 6239
rect 35667 6205 35676 6239
rect 35624 6196 35676 6205
rect 35992 6239 36044 6248
rect 35992 6205 36001 6239
rect 36001 6205 36035 6239
rect 36035 6205 36044 6239
rect 35992 6196 36044 6205
rect 37924 6341 37933 6375
rect 37933 6341 37967 6375
rect 37967 6341 37976 6375
rect 37924 6332 37976 6341
rect 39396 6307 39448 6316
rect 35256 6171 35308 6180
rect 35256 6137 35265 6171
rect 35265 6137 35299 6171
rect 35299 6137 35308 6171
rect 35256 6128 35308 6137
rect 35716 6128 35768 6180
rect 31852 6060 31904 6112
rect 32496 6060 32548 6112
rect 33508 6103 33560 6112
rect 33508 6069 33517 6103
rect 33517 6069 33551 6103
rect 33551 6069 33560 6103
rect 33508 6060 33560 6069
rect 34612 6060 34664 6112
rect 38660 6239 38712 6248
rect 38660 6205 38669 6239
rect 38669 6205 38703 6239
rect 38703 6205 38712 6239
rect 38660 6196 38712 6205
rect 38936 6196 38988 6248
rect 39396 6273 39405 6307
rect 39405 6273 39439 6307
rect 39439 6273 39448 6307
rect 39396 6264 39448 6273
rect 40500 6332 40552 6384
rect 42432 6400 42484 6452
rect 42892 6400 42944 6452
rect 45560 6443 45612 6452
rect 45560 6409 45569 6443
rect 45569 6409 45603 6443
rect 45603 6409 45612 6443
rect 45560 6400 45612 6409
rect 46204 6400 46256 6452
rect 47308 6400 47360 6452
rect 47952 6443 48004 6452
rect 47952 6409 47961 6443
rect 47961 6409 47995 6443
rect 47995 6409 48004 6443
rect 47952 6400 48004 6409
rect 48504 6400 48556 6452
rect 50344 6400 50396 6452
rect 52184 6400 52236 6452
rect 42064 6264 42116 6316
rect 41880 6196 41932 6248
rect 42432 6239 42484 6248
rect 42432 6205 42455 6239
rect 42455 6205 42484 6239
rect 42432 6196 42484 6205
rect 40500 6171 40552 6180
rect 39488 6060 39540 6112
rect 40500 6137 40509 6171
rect 40509 6137 40543 6171
rect 40543 6137 40552 6171
rect 40500 6128 40552 6137
rect 42892 6239 42944 6248
rect 42892 6205 42901 6239
rect 42901 6205 42935 6239
rect 42935 6205 42944 6239
rect 42892 6196 42944 6205
rect 43352 6196 43404 6248
rect 44088 6264 44140 6316
rect 44640 6264 44692 6316
rect 50620 6332 50672 6384
rect 54760 6400 54812 6452
rect 54944 6443 54996 6452
rect 54944 6409 54953 6443
rect 54953 6409 54987 6443
rect 54987 6409 54996 6443
rect 54944 6400 54996 6409
rect 55496 6400 55548 6452
rect 55772 6400 55824 6452
rect 57704 6400 57756 6452
rect 57796 6400 57848 6452
rect 56600 6332 56652 6384
rect 44364 6196 44416 6248
rect 44732 6239 44784 6248
rect 42984 6128 43036 6180
rect 43720 6171 43772 6180
rect 43720 6137 43729 6171
rect 43729 6137 43763 6171
rect 43763 6137 43772 6171
rect 44732 6205 44741 6239
rect 44741 6205 44775 6239
rect 44775 6205 44784 6239
rect 44732 6196 44784 6205
rect 46112 6196 46164 6248
rect 46296 6196 46348 6248
rect 47400 6196 47452 6248
rect 48504 6264 48556 6316
rect 53288 6307 53340 6316
rect 47952 6196 48004 6248
rect 49976 6196 50028 6248
rect 50436 6196 50488 6248
rect 51908 6239 51960 6248
rect 51908 6205 51917 6239
rect 51917 6205 51951 6239
rect 51951 6205 51960 6239
rect 51908 6196 51960 6205
rect 53012 6239 53064 6248
rect 53012 6205 53021 6239
rect 53021 6205 53055 6239
rect 53055 6205 53064 6239
rect 53012 6196 53064 6205
rect 53288 6273 53297 6307
rect 53297 6273 53331 6307
rect 53331 6273 53340 6307
rect 53288 6264 53340 6273
rect 53380 6264 53432 6316
rect 55864 6264 55916 6316
rect 57520 6264 57572 6316
rect 58256 6264 58308 6316
rect 43720 6128 43772 6137
rect 44916 6128 44968 6180
rect 46756 6128 46808 6180
rect 46848 6128 46900 6180
rect 46664 6060 46716 6112
rect 49056 6060 49108 6112
rect 55588 6128 55640 6180
rect 49700 6060 49752 6112
rect 50068 6060 50120 6112
rect 50804 6103 50856 6112
rect 50804 6069 50813 6103
rect 50813 6069 50847 6103
rect 50847 6069 50856 6103
rect 50804 6060 50856 6069
rect 50896 6060 50948 6112
rect 52368 6060 52420 6112
rect 52552 6060 52604 6112
rect 58348 6239 58400 6248
rect 57980 6103 58032 6112
rect 57980 6069 57989 6103
rect 57989 6069 58023 6103
rect 58023 6069 58032 6103
rect 57980 6060 58032 6069
rect 58348 6205 58357 6239
rect 58357 6205 58391 6239
rect 58391 6205 58400 6239
rect 58348 6196 58400 6205
rect 58440 6060 58492 6112
rect 60004 6103 60056 6112
rect 60004 6069 60013 6103
rect 60013 6069 60047 6103
rect 60047 6069 60056 6103
rect 60004 6060 60056 6069
rect 60280 6060 60332 6112
rect 61384 6264 61436 6316
rect 60648 6239 60700 6248
rect 60648 6205 60657 6239
rect 60657 6205 60691 6239
rect 60691 6205 60700 6239
rect 60648 6196 60700 6205
rect 61568 6103 61620 6112
rect 61568 6069 61577 6103
rect 61577 6069 61611 6103
rect 61611 6069 61620 6103
rect 61568 6060 61620 6069
rect 21774 5958 21826 6010
rect 21838 5958 21890 6010
rect 21902 5958 21954 6010
rect 21966 5958 22018 6010
rect 42566 5958 42618 6010
rect 42630 5958 42682 6010
rect 42694 5958 42746 6010
rect 42758 5958 42810 6010
rect 3516 5788 3568 5840
rect 2688 5763 2740 5772
rect 2688 5729 2697 5763
rect 2697 5729 2731 5763
rect 2731 5729 2740 5763
rect 2688 5720 2740 5729
rect 4620 5720 4672 5772
rect 2596 5695 2648 5704
rect 2596 5661 2605 5695
rect 2605 5661 2639 5695
rect 2639 5661 2648 5695
rect 2596 5652 2648 5661
rect 5172 5720 5224 5772
rect 6920 5856 6972 5908
rect 7196 5856 7248 5908
rect 9404 5899 9456 5908
rect 6552 5788 6604 5840
rect 6184 5720 6236 5772
rect 8208 5788 8260 5840
rect 9404 5865 9413 5899
rect 9413 5865 9447 5899
rect 9447 5865 9456 5899
rect 9404 5856 9456 5865
rect 16764 5856 16816 5908
rect 17040 5856 17092 5908
rect 20720 5899 20772 5908
rect 8392 5788 8444 5840
rect 11704 5788 11756 5840
rect 12900 5788 12952 5840
rect 18788 5788 18840 5840
rect 8300 5720 8352 5772
rect 9772 5763 9824 5772
rect 9772 5729 9781 5763
rect 9781 5729 9815 5763
rect 9815 5729 9824 5763
rect 9772 5720 9824 5729
rect 11060 5720 11112 5772
rect 11888 5720 11940 5772
rect 13636 5720 13688 5772
rect 15016 5720 15068 5772
rect 16120 5720 16172 5772
rect 16304 5763 16356 5772
rect 16304 5729 16313 5763
rect 16313 5729 16347 5763
rect 16347 5729 16356 5763
rect 16304 5720 16356 5729
rect 17776 5720 17828 5772
rect 18144 5720 18196 5772
rect 18696 5720 18748 5772
rect 19340 5788 19392 5840
rect 19800 5788 19852 5840
rect 20720 5865 20729 5899
rect 20729 5865 20763 5899
rect 20763 5865 20772 5899
rect 20720 5856 20772 5865
rect 22100 5856 22152 5908
rect 22836 5856 22888 5908
rect 23112 5899 23164 5908
rect 23112 5865 23121 5899
rect 23121 5865 23155 5899
rect 23155 5865 23164 5899
rect 23112 5856 23164 5865
rect 23664 5899 23716 5908
rect 23664 5865 23673 5899
rect 23673 5865 23707 5899
rect 23707 5865 23716 5899
rect 23664 5856 23716 5865
rect 24032 5856 24084 5908
rect 28264 5856 28316 5908
rect 31392 5856 31444 5908
rect 20904 5788 20956 5840
rect 21272 5788 21324 5840
rect 19616 5720 19668 5772
rect 21548 5763 21600 5772
rect 21548 5729 21557 5763
rect 21557 5729 21591 5763
rect 21591 5729 21600 5763
rect 21548 5720 21600 5729
rect 22652 5720 22704 5772
rect 22928 5763 22980 5772
rect 22928 5729 22937 5763
rect 22937 5729 22971 5763
rect 22971 5729 22980 5763
rect 22928 5720 22980 5729
rect 4988 5652 5040 5704
rect 5448 5652 5500 5704
rect 7748 5652 7800 5704
rect 9680 5695 9732 5704
rect 9680 5661 9689 5695
rect 9689 5661 9723 5695
rect 9723 5661 9732 5695
rect 9680 5652 9732 5661
rect 10232 5652 10284 5704
rect 11704 5652 11756 5704
rect 5172 5584 5224 5636
rect 8116 5584 8168 5636
rect 11060 5627 11112 5636
rect 11060 5593 11069 5627
rect 11069 5593 11103 5627
rect 11103 5593 11112 5627
rect 11060 5584 11112 5593
rect 12532 5584 12584 5636
rect 14096 5627 14148 5636
rect 14096 5593 14105 5627
rect 14105 5593 14139 5627
rect 14139 5593 14148 5627
rect 14096 5584 14148 5593
rect 14924 5584 14976 5636
rect 16580 5652 16632 5704
rect 18052 5652 18104 5704
rect 2320 5516 2372 5568
rect 3516 5559 3568 5568
rect 3516 5525 3525 5559
rect 3525 5525 3559 5559
rect 3559 5525 3568 5559
rect 3516 5516 3568 5525
rect 3792 5559 3844 5568
rect 3792 5525 3801 5559
rect 3801 5525 3835 5559
rect 3835 5525 3844 5559
rect 3792 5516 3844 5525
rect 5632 5516 5684 5568
rect 5724 5516 5776 5568
rect 7012 5559 7064 5568
rect 7012 5525 7021 5559
rect 7021 5525 7055 5559
rect 7055 5525 7064 5559
rect 7012 5516 7064 5525
rect 8852 5516 8904 5568
rect 8944 5516 8996 5568
rect 10416 5516 10468 5568
rect 12808 5559 12860 5568
rect 12808 5525 12817 5559
rect 12817 5525 12851 5559
rect 12851 5525 12860 5559
rect 12808 5516 12860 5525
rect 15108 5559 15160 5568
rect 15108 5525 15117 5559
rect 15117 5525 15151 5559
rect 15151 5525 15160 5559
rect 15108 5516 15160 5525
rect 15936 5584 15988 5636
rect 22376 5584 22428 5636
rect 24032 5720 24084 5772
rect 24860 5788 24912 5840
rect 25320 5788 25372 5840
rect 25596 5788 25648 5840
rect 26424 5788 26476 5840
rect 24400 5763 24452 5772
rect 24400 5729 24409 5763
rect 24409 5729 24443 5763
rect 24443 5729 24452 5763
rect 24400 5720 24452 5729
rect 24676 5720 24728 5772
rect 23204 5652 23256 5704
rect 18696 5516 18748 5568
rect 19340 5516 19392 5568
rect 21732 5516 21784 5568
rect 24400 5584 24452 5636
rect 25044 5652 25096 5704
rect 26700 5652 26752 5704
rect 26976 5695 27028 5704
rect 26976 5661 26985 5695
rect 26985 5661 27019 5695
rect 27019 5661 27028 5695
rect 29092 5720 29144 5772
rect 29460 5763 29512 5772
rect 29460 5729 29469 5763
rect 29469 5729 29503 5763
rect 29503 5729 29512 5763
rect 29460 5720 29512 5729
rect 29552 5763 29604 5772
rect 29552 5729 29561 5763
rect 29561 5729 29595 5763
rect 29595 5729 29604 5763
rect 30012 5763 30064 5772
rect 29552 5720 29604 5729
rect 30012 5729 30021 5763
rect 30021 5729 30055 5763
rect 30055 5729 30064 5763
rect 30012 5720 30064 5729
rect 31024 5763 31076 5772
rect 31024 5729 31033 5763
rect 31033 5729 31067 5763
rect 31067 5729 31076 5763
rect 31024 5720 31076 5729
rect 31300 5720 31352 5772
rect 32956 5788 33008 5840
rect 26976 5652 27028 5661
rect 28632 5652 28684 5704
rect 29828 5652 29880 5704
rect 31484 5695 31536 5704
rect 31484 5661 31493 5695
rect 31493 5661 31527 5695
rect 31527 5661 31536 5695
rect 31484 5652 31536 5661
rect 32496 5720 32548 5772
rect 35256 5856 35308 5908
rect 41328 5856 41380 5908
rect 41604 5899 41656 5908
rect 41604 5865 41613 5899
rect 41613 5865 41647 5899
rect 41647 5865 41656 5899
rect 41604 5856 41656 5865
rect 42248 5856 42300 5908
rect 42984 5899 43036 5908
rect 42984 5865 42993 5899
rect 42993 5865 43027 5899
rect 43027 5865 43036 5899
rect 42984 5856 43036 5865
rect 34152 5788 34204 5840
rect 38384 5831 38436 5840
rect 33600 5720 33652 5772
rect 34888 5763 34940 5772
rect 34888 5729 34897 5763
rect 34897 5729 34931 5763
rect 34931 5729 34940 5763
rect 34888 5720 34940 5729
rect 34980 5763 35032 5772
rect 34980 5729 34989 5763
rect 34989 5729 35023 5763
rect 35023 5729 35032 5763
rect 35164 5763 35216 5772
rect 34980 5720 35032 5729
rect 35164 5729 35173 5763
rect 35173 5729 35207 5763
rect 35207 5729 35216 5763
rect 35164 5720 35216 5729
rect 35348 5763 35400 5772
rect 35348 5729 35357 5763
rect 35357 5729 35391 5763
rect 35391 5729 35400 5763
rect 35348 5720 35400 5729
rect 35440 5720 35492 5772
rect 37004 5720 37056 5772
rect 37280 5720 37332 5772
rect 37740 5763 37792 5772
rect 37740 5729 37749 5763
rect 37749 5729 37783 5763
rect 37783 5729 37792 5763
rect 37740 5720 37792 5729
rect 38384 5797 38393 5831
rect 38393 5797 38427 5831
rect 38427 5797 38436 5831
rect 38384 5788 38436 5797
rect 41880 5788 41932 5840
rect 48228 5856 48280 5908
rect 49148 5899 49200 5908
rect 49148 5865 49157 5899
rect 49157 5865 49191 5899
rect 49191 5865 49200 5899
rect 49148 5856 49200 5865
rect 49976 5899 50028 5908
rect 49976 5865 49985 5899
rect 49985 5865 50019 5899
rect 50019 5865 50028 5899
rect 49976 5856 50028 5865
rect 43444 5831 43496 5840
rect 43444 5797 43453 5831
rect 43453 5797 43487 5831
rect 43487 5797 43496 5831
rect 43444 5788 43496 5797
rect 46296 5788 46348 5840
rect 52184 5856 52236 5908
rect 52276 5856 52328 5908
rect 41696 5720 41748 5772
rect 41972 5763 42024 5772
rect 41972 5729 41981 5763
rect 41981 5729 42015 5763
rect 42015 5729 42024 5763
rect 41972 5720 42024 5729
rect 43904 5720 43956 5772
rect 44088 5720 44140 5772
rect 44364 5720 44416 5772
rect 45008 5763 45060 5772
rect 45008 5729 45017 5763
rect 45017 5729 45051 5763
rect 45051 5729 45060 5763
rect 45008 5720 45060 5729
rect 45100 5763 45152 5772
rect 45100 5729 45109 5763
rect 45109 5729 45143 5763
rect 45143 5729 45152 5763
rect 45100 5720 45152 5729
rect 29368 5584 29420 5636
rect 29460 5584 29512 5636
rect 30104 5584 30156 5636
rect 31208 5584 31260 5636
rect 35164 5584 35216 5636
rect 35992 5584 36044 5636
rect 36176 5584 36228 5636
rect 39028 5652 39080 5704
rect 39304 5695 39356 5704
rect 39304 5661 39313 5695
rect 39313 5661 39347 5695
rect 39347 5661 39356 5695
rect 39304 5652 39356 5661
rect 39580 5695 39632 5704
rect 39580 5661 39589 5695
rect 39589 5661 39623 5695
rect 39623 5661 39632 5695
rect 39580 5652 39632 5661
rect 40224 5652 40276 5704
rect 40868 5652 40920 5704
rect 41144 5652 41196 5704
rect 43720 5652 43772 5704
rect 44456 5652 44508 5704
rect 52828 5788 52880 5840
rect 46664 5763 46716 5772
rect 46664 5729 46673 5763
rect 46673 5729 46707 5763
rect 46707 5729 46716 5763
rect 46664 5720 46716 5729
rect 48044 5720 48096 5772
rect 48228 5720 48280 5772
rect 49700 5720 49752 5772
rect 50252 5763 50304 5772
rect 50252 5729 50261 5763
rect 50261 5729 50295 5763
rect 50295 5729 50304 5763
rect 50252 5720 50304 5729
rect 50436 5720 50488 5772
rect 50896 5763 50948 5772
rect 50896 5729 50905 5763
rect 50905 5729 50939 5763
rect 50939 5729 50948 5763
rect 50896 5720 50948 5729
rect 51816 5720 51868 5772
rect 53380 5763 53432 5772
rect 53380 5729 53389 5763
rect 53389 5729 53423 5763
rect 53423 5729 53432 5763
rect 54760 5788 54812 5840
rect 55128 5788 55180 5840
rect 55864 5856 55916 5908
rect 57796 5856 57848 5908
rect 57980 5856 58032 5908
rect 58348 5856 58400 5908
rect 58716 5856 58768 5908
rect 55772 5788 55824 5840
rect 57336 5788 57388 5840
rect 57612 5788 57664 5840
rect 53380 5720 53432 5729
rect 56508 5720 56560 5772
rect 57796 5720 57848 5772
rect 58072 5720 58124 5772
rect 58256 5720 58308 5772
rect 58900 5720 58952 5772
rect 46756 5695 46808 5704
rect 46756 5661 46765 5695
rect 46765 5661 46799 5695
rect 46799 5661 46808 5695
rect 46756 5652 46808 5661
rect 49148 5652 49200 5704
rect 39120 5584 39172 5636
rect 40776 5584 40828 5636
rect 42892 5584 42944 5636
rect 44732 5584 44784 5636
rect 44824 5627 44876 5636
rect 44824 5593 44833 5627
rect 44833 5593 44867 5627
rect 44867 5593 44876 5627
rect 44824 5584 44876 5593
rect 23940 5559 23992 5568
rect 23940 5525 23949 5559
rect 23949 5525 23983 5559
rect 23983 5525 23992 5559
rect 23940 5516 23992 5525
rect 24032 5516 24084 5568
rect 26608 5516 26660 5568
rect 26792 5516 26844 5568
rect 27804 5559 27856 5568
rect 27804 5525 27813 5559
rect 27813 5525 27847 5559
rect 27847 5525 27856 5559
rect 27804 5516 27856 5525
rect 27988 5516 28040 5568
rect 29276 5516 29328 5568
rect 29552 5516 29604 5568
rect 30288 5516 30340 5568
rect 31116 5559 31168 5568
rect 31116 5525 31125 5559
rect 31125 5525 31159 5559
rect 31159 5525 31168 5559
rect 31116 5516 31168 5525
rect 31852 5559 31904 5568
rect 31852 5525 31861 5559
rect 31861 5525 31895 5559
rect 31895 5525 31904 5559
rect 31852 5516 31904 5525
rect 32588 5516 32640 5568
rect 32772 5516 32824 5568
rect 33508 5516 33560 5568
rect 34520 5516 34572 5568
rect 34980 5516 35032 5568
rect 35256 5516 35308 5568
rect 35716 5516 35768 5568
rect 35900 5516 35952 5568
rect 36360 5516 36412 5568
rect 36728 5559 36780 5568
rect 36728 5525 36737 5559
rect 36737 5525 36771 5559
rect 36771 5525 36780 5559
rect 36728 5516 36780 5525
rect 37924 5559 37976 5568
rect 37924 5525 37933 5559
rect 37933 5525 37967 5559
rect 37967 5525 37976 5559
rect 37924 5516 37976 5525
rect 38384 5516 38436 5568
rect 38752 5559 38804 5568
rect 38752 5525 38761 5559
rect 38761 5525 38795 5559
rect 38795 5525 38804 5559
rect 38752 5516 38804 5525
rect 40592 5516 40644 5568
rect 41788 5516 41840 5568
rect 48688 5584 48740 5636
rect 49332 5584 49384 5636
rect 50252 5584 50304 5636
rect 50988 5584 51040 5636
rect 53288 5584 53340 5636
rect 53840 5652 53892 5704
rect 54944 5652 54996 5704
rect 55588 5584 55640 5636
rect 55772 5627 55824 5636
rect 55772 5593 55796 5627
rect 55796 5593 55824 5627
rect 55772 5584 55824 5593
rect 56140 5652 56192 5704
rect 57152 5695 57204 5704
rect 57152 5661 57161 5695
rect 57161 5661 57195 5695
rect 57195 5661 57204 5695
rect 57152 5652 57204 5661
rect 58164 5695 58216 5704
rect 58164 5661 58173 5695
rect 58173 5661 58207 5695
rect 58207 5661 58216 5695
rect 58164 5652 58216 5661
rect 46112 5516 46164 5568
rect 46664 5516 46716 5568
rect 47768 5516 47820 5568
rect 47952 5516 48004 5568
rect 48412 5516 48464 5568
rect 50160 5516 50212 5568
rect 50344 5559 50396 5568
rect 50344 5525 50353 5559
rect 50353 5525 50387 5559
rect 50387 5525 50396 5559
rect 50344 5516 50396 5525
rect 51448 5516 51500 5568
rect 54668 5559 54720 5568
rect 54668 5525 54677 5559
rect 54677 5525 54711 5559
rect 54711 5525 54720 5559
rect 54668 5516 54720 5525
rect 55496 5559 55548 5568
rect 55496 5525 55505 5559
rect 55505 5525 55539 5559
rect 55539 5525 55548 5559
rect 55496 5516 55548 5525
rect 56048 5516 56100 5568
rect 56232 5559 56284 5568
rect 56232 5525 56241 5559
rect 56241 5525 56275 5559
rect 56275 5525 56284 5559
rect 56232 5516 56284 5525
rect 56600 5516 56652 5568
rect 59636 5584 59688 5636
rect 59268 5516 59320 5568
rect 59728 5516 59780 5568
rect 61292 5720 61344 5772
rect 60464 5695 60516 5704
rect 60464 5661 60473 5695
rect 60473 5661 60507 5695
rect 60507 5661 60516 5695
rect 60464 5652 60516 5661
rect 61752 5559 61804 5568
rect 61752 5525 61761 5559
rect 61761 5525 61795 5559
rect 61795 5525 61804 5559
rect 61752 5516 61804 5525
rect 11378 5414 11430 5466
rect 11442 5414 11494 5466
rect 11506 5414 11558 5466
rect 11570 5414 11622 5466
rect 32170 5414 32222 5466
rect 32234 5414 32286 5466
rect 32298 5414 32350 5466
rect 32362 5414 32414 5466
rect 52962 5414 53014 5466
rect 53026 5414 53078 5466
rect 53090 5414 53142 5466
rect 53154 5414 53206 5466
rect 2688 5312 2740 5364
rect 4068 5312 4120 5364
rect 14096 5312 14148 5364
rect 15016 5312 15068 5364
rect 16304 5312 16356 5364
rect 4988 5287 5040 5296
rect 4988 5253 4997 5287
rect 4997 5253 5031 5287
rect 5031 5253 5040 5287
rect 4988 5244 5040 5253
rect 5172 5244 5224 5296
rect 6184 5287 6236 5296
rect 6184 5253 6193 5287
rect 6193 5253 6227 5287
rect 6227 5253 6236 5287
rect 6184 5244 6236 5253
rect 7748 5244 7800 5296
rect 8300 5287 8352 5296
rect 8300 5253 8309 5287
rect 8309 5253 8343 5287
rect 8343 5253 8352 5287
rect 8300 5244 8352 5253
rect 9496 5244 9548 5296
rect 11888 5287 11940 5296
rect 11888 5253 11897 5287
rect 11897 5253 11931 5287
rect 11931 5253 11940 5287
rect 11888 5244 11940 5253
rect 7932 5176 7984 5228
rect 9404 5219 9456 5228
rect 9404 5185 9413 5219
rect 9413 5185 9447 5219
rect 9447 5185 9456 5219
rect 9404 5176 9456 5185
rect 9772 5176 9824 5228
rect 2320 5108 2372 5160
rect 3516 5108 3568 5160
rect 4068 5108 4120 5160
rect 5632 5151 5684 5160
rect 5632 5117 5641 5151
rect 5641 5117 5675 5151
rect 5675 5117 5684 5151
rect 5632 5108 5684 5117
rect 7012 5151 7064 5160
rect 7012 5117 7021 5151
rect 7021 5117 7055 5151
rect 7055 5117 7064 5151
rect 7012 5108 7064 5117
rect 8024 5108 8076 5160
rect 8852 5108 8904 5160
rect 9312 5151 9364 5160
rect 9312 5117 9321 5151
rect 9321 5117 9355 5151
rect 9355 5117 9364 5151
rect 9312 5108 9364 5117
rect 10324 5151 10376 5160
rect 2596 4972 2648 5024
rect 8300 5040 8352 5092
rect 8576 5083 8628 5092
rect 8576 5049 8585 5083
rect 8585 5049 8619 5083
rect 8619 5049 8628 5083
rect 8576 5040 8628 5049
rect 10324 5117 10333 5151
rect 10333 5117 10367 5151
rect 10367 5117 10376 5151
rect 10324 5108 10376 5117
rect 10508 5176 10560 5228
rect 12348 5176 12400 5228
rect 12808 5176 12860 5228
rect 15844 5244 15896 5296
rect 18144 5312 18196 5364
rect 19064 5355 19116 5364
rect 19064 5321 19073 5355
rect 19073 5321 19107 5355
rect 19107 5321 19116 5355
rect 19064 5312 19116 5321
rect 19156 5312 19208 5364
rect 20812 5312 20864 5364
rect 18604 5244 18656 5296
rect 20260 5244 20312 5296
rect 19340 5176 19392 5228
rect 21916 5244 21968 5296
rect 22192 5312 22244 5364
rect 24216 5355 24268 5364
rect 24216 5321 24225 5355
rect 24225 5321 24259 5355
rect 24259 5321 24268 5355
rect 24216 5312 24268 5321
rect 27252 5312 27304 5364
rect 28172 5312 28224 5364
rect 24676 5287 24728 5296
rect 24676 5253 24685 5287
rect 24685 5253 24719 5287
rect 24719 5253 24728 5287
rect 24676 5244 24728 5253
rect 26792 5244 26844 5296
rect 29092 5244 29144 5296
rect 32496 5312 32548 5364
rect 32864 5312 32916 5364
rect 35348 5312 35400 5364
rect 35992 5355 36044 5364
rect 35992 5321 36001 5355
rect 36001 5321 36035 5355
rect 36035 5321 36044 5355
rect 35992 5312 36044 5321
rect 36452 5312 36504 5364
rect 37740 5312 37792 5364
rect 38016 5312 38068 5364
rect 39580 5355 39632 5364
rect 39580 5321 39589 5355
rect 39589 5321 39623 5355
rect 39623 5321 39632 5355
rect 39580 5312 39632 5321
rect 39764 5312 39816 5364
rect 40868 5312 40920 5364
rect 41788 5355 41840 5364
rect 41788 5321 41797 5355
rect 41797 5321 41831 5355
rect 41831 5321 41840 5355
rect 41788 5312 41840 5321
rect 41972 5312 42024 5364
rect 42892 5312 42944 5364
rect 43352 5312 43404 5364
rect 44456 5312 44508 5364
rect 44732 5312 44784 5364
rect 45008 5312 45060 5364
rect 31668 5244 31720 5296
rect 31944 5244 31996 5296
rect 35256 5287 35308 5296
rect 35256 5253 35265 5287
rect 35265 5253 35299 5287
rect 35299 5253 35308 5287
rect 35256 5244 35308 5253
rect 39028 5244 39080 5296
rect 39120 5244 39172 5296
rect 40776 5287 40828 5296
rect 40776 5253 40785 5287
rect 40785 5253 40819 5287
rect 40819 5253 40828 5287
rect 40776 5244 40828 5253
rect 40960 5244 41012 5296
rect 43904 5287 43956 5296
rect 43904 5253 43913 5287
rect 43913 5253 43947 5287
rect 43947 5253 43956 5287
rect 43904 5244 43956 5253
rect 11704 5108 11756 5160
rect 14556 5108 14608 5160
rect 14648 5108 14700 5160
rect 15568 5151 15620 5160
rect 15568 5117 15577 5151
rect 15577 5117 15611 5151
rect 15611 5117 15620 5151
rect 15568 5108 15620 5117
rect 15936 5151 15988 5160
rect 15936 5117 15945 5151
rect 15945 5117 15979 5151
rect 15979 5117 15988 5151
rect 15936 5108 15988 5117
rect 16028 5151 16080 5160
rect 16028 5117 16037 5151
rect 16037 5117 16071 5151
rect 16071 5117 16080 5151
rect 16028 5108 16080 5117
rect 17776 5108 17828 5160
rect 18512 5108 18564 5160
rect 21548 5176 21600 5228
rect 22284 5176 22336 5228
rect 22836 5176 22888 5228
rect 22928 5176 22980 5228
rect 20352 5108 20404 5160
rect 20720 5108 20772 5160
rect 20996 5108 21048 5160
rect 5356 4972 5408 5024
rect 5816 5015 5868 5024
rect 5816 4981 5825 5015
rect 5825 4981 5859 5015
rect 5859 4981 5868 5015
rect 5816 4972 5868 4981
rect 7840 4972 7892 5024
rect 12072 5040 12124 5092
rect 13636 5040 13688 5092
rect 18236 5083 18288 5092
rect 18236 5049 18245 5083
rect 18245 5049 18279 5083
rect 18279 5049 18288 5083
rect 18236 5040 18288 5049
rect 10048 4972 10100 5024
rect 10232 5015 10284 5024
rect 10232 4981 10241 5015
rect 10241 4981 10275 5015
rect 10275 4981 10284 5015
rect 10232 4972 10284 4981
rect 10968 4972 11020 5024
rect 15752 4972 15804 5024
rect 18328 4972 18380 5024
rect 22192 5040 22244 5092
rect 22468 5151 22520 5160
rect 22468 5117 22477 5151
rect 22477 5117 22511 5151
rect 22511 5117 22520 5151
rect 22468 5108 22520 5117
rect 22652 5108 22704 5160
rect 24124 5176 24176 5228
rect 24216 5108 24268 5160
rect 25044 5219 25096 5228
rect 25044 5185 25053 5219
rect 25053 5185 25087 5219
rect 25087 5185 25096 5219
rect 25044 5176 25096 5185
rect 25228 5176 25280 5228
rect 25964 5108 26016 5160
rect 19524 4972 19576 5024
rect 20352 4972 20404 5024
rect 20904 4972 20956 5024
rect 22284 5015 22336 5024
rect 22284 4981 22293 5015
rect 22293 4981 22327 5015
rect 22327 4981 22336 5015
rect 22284 4972 22336 4981
rect 22560 4972 22612 5024
rect 26056 4972 26108 5024
rect 26240 5176 26292 5228
rect 26976 5176 27028 5228
rect 31852 5176 31904 5228
rect 32128 5176 32180 5228
rect 26700 5108 26752 5160
rect 27896 5108 27948 5160
rect 28080 5151 28132 5160
rect 28080 5117 28089 5151
rect 28089 5117 28123 5151
rect 28123 5117 28132 5151
rect 28080 5108 28132 5117
rect 28264 5151 28316 5160
rect 28264 5117 28273 5151
rect 28273 5117 28307 5151
rect 28307 5117 28316 5151
rect 28264 5108 28316 5117
rect 28356 5108 28408 5160
rect 29828 5151 29880 5160
rect 29828 5117 29837 5151
rect 29837 5117 29871 5151
rect 29871 5117 29880 5151
rect 29828 5108 29880 5117
rect 29920 5151 29972 5160
rect 29920 5117 29929 5151
rect 29929 5117 29963 5151
rect 29963 5117 29972 5151
rect 30104 5151 30156 5160
rect 29920 5108 29972 5117
rect 30104 5117 30113 5151
rect 30113 5117 30147 5151
rect 30147 5117 30156 5151
rect 30104 5108 30156 5117
rect 30288 5151 30340 5160
rect 30288 5117 30297 5151
rect 30297 5117 30331 5151
rect 30331 5117 30340 5151
rect 30288 5108 30340 5117
rect 31392 5151 31444 5160
rect 31392 5117 31401 5151
rect 31401 5117 31435 5151
rect 31435 5117 31444 5151
rect 31392 5108 31444 5117
rect 27160 5040 27212 5092
rect 29000 5083 29052 5092
rect 29000 5049 29009 5083
rect 29009 5049 29043 5083
rect 29043 5049 29052 5083
rect 29000 5040 29052 5049
rect 30196 5040 30248 5092
rect 32588 5108 32640 5160
rect 33508 5176 33560 5228
rect 37924 5176 37976 5228
rect 41144 5219 41196 5228
rect 33232 5108 33284 5160
rect 34244 5151 34296 5160
rect 34244 5117 34253 5151
rect 34253 5117 34287 5151
rect 34287 5117 34296 5151
rect 34244 5108 34296 5117
rect 36084 5108 36136 5160
rect 36176 5151 36228 5160
rect 36176 5117 36185 5151
rect 36185 5117 36219 5151
rect 36219 5117 36228 5151
rect 36360 5151 36412 5160
rect 36176 5108 36228 5117
rect 36360 5117 36369 5151
rect 36369 5117 36403 5151
rect 36403 5117 36412 5151
rect 36360 5108 36412 5117
rect 38016 5151 38068 5160
rect 38016 5117 38025 5151
rect 38025 5117 38059 5151
rect 38059 5117 38068 5151
rect 38016 5108 38068 5117
rect 38384 5151 38436 5160
rect 38384 5117 38393 5151
rect 38393 5117 38427 5151
rect 38427 5117 38436 5151
rect 38384 5108 38436 5117
rect 29736 4972 29788 5024
rect 29920 4972 29972 5024
rect 31668 5040 31720 5092
rect 31024 5015 31076 5024
rect 31024 4981 31033 5015
rect 31033 4981 31067 5015
rect 31067 4981 31076 5015
rect 31024 4972 31076 4981
rect 34520 5040 34572 5092
rect 36544 5040 36596 5092
rect 37556 5040 37608 5092
rect 32680 4972 32732 5024
rect 33324 4972 33376 5024
rect 33600 5015 33652 5024
rect 33600 4981 33609 5015
rect 33609 4981 33643 5015
rect 33643 4981 33652 5015
rect 33600 4972 33652 4981
rect 37004 5015 37056 5024
rect 37004 4981 37013 5015
rect 37013 4981 37047 5015
rect 37047 4981 37056 5015
rect 37004 4972 37056 4981
rect 37372 5015 37424 5024
rect 37372 4981 37381 5015
rect 37381 4981 37415 5015
rect 37415 4981 37424 5015
rect 37372 4972 37424 4981
rect 37464 4972 37516 5024
rect 38936 5151 38988 5160
rect 38936 5117 38945 5151
rect 38945 5117 38979 5151
rect 38979 5117 38988 5151
rect 38936 5108 38988 5117
rect 39304 5108 39356 5160
rect 40500 5108 40552 5160
rect 41144 5185 41153 5219
rect 41153 5185 41187 5219
rect 41187 5185 41196 5219
rect 41144 5176 41196 5185
rect 44088 5176 44140 5228
rect 41972 5151 42024 5160
rect 41972 5117 41981 5151
rect 41981 5117 42015 5151
rect 42015 5117 42024 5151
rect 41972 5108 42024 5117
rect 42892 5108 42944 5160
rect 43628 5108 43680 5160
rect 46112 5244 46164 5296
rect 44824 5176 44876 5228
rect 48872 5312 48924 5364
rect 50252 5312 50304 5364
rect 50436 5312 50488 5364
rect 51816 5312 51868 5364
rect 46296 5287 46348 5296
rect 46296 5253 46305 5287
rect 46305 5253 46339 5287
rect 46339 5253 46348 5287
rect 46296 5244 46348 5253
rect 47124 5244 47176 5296
rect 53380 5287 53432 5296
rect 53380 5253 53389 5287
rect 53389 5253 53423 5287
rect 53423 5253 53432 5287
rect 53380 5244 53432 5253
rect 53840 5312 53892 5364
rect 55220 5312 55272 5364
rect 55772 5312 55824 5364
rect 56048 5312 56100 5364
rect 58900 5355 58952 5364
rect 58900 5321 58909 5355
rect 58909 5321 58943 5355
rect 58943 5321 58952 5355
rect 58900 5312 58952 5321
rect 61292 5312 61344 5364
rect 54024 5244 54076 5296
rect 39028 5040 39080 5092
rect 44548 5108 44600 5160
rect 45008 5108 45060 5160
rect 48136 5176 48188 5228
rect 49516 5176 49568 5228
rect 50620 5176 50672 5228
rect 52736 5176 52788 5228
rect 43812 5040 43864 5092
rect 47860 5108 47912 5160
rect 49332 5151 49384 5160
rect 49332 5117 49341 5151
rect 49341 5117 49375 5151
rect 49375 5117 49384 5151
rect 49332 5108 49384 5117
rect 49700 5151 49752 5160
rect 49700 5117 49709 5151
rect 49709 5117 49743 5151
rect 49743 5117 49752 5151
rect 49700 5108 49752 5117
rect 50896 5151 50948 5160
rect 50896 5117 50905 5151
rect 50905 5117 50939 5151
rect 50939 5117 50948 5151
rect 50896 5108 50948 5117
rect 52644 5151 52696 5160
rect 52644 5117 52653 5151
rect 52653 5117 52687 5151
rect 52687 5117 52696 5151
rect 52644 5108 52696 5117
rect 52828 5108 52880 5160
rect 39212 5015 39264 5024
rect 39212 4981 39221 5015
rect 39221 4981 39255 5015
rect 39255 4981 39264 5015
rect 39212 4972 39264 4981
rect 40224 4972 40276 5024
rect 40868 4972 40920 5024
rect 41972 4972 42024 5024
rect 46572 5015 46624 5024
rect 46572 4981 46581 5015
rect 46581 4981 46615 5015
rect 46615 4981 46624 5015
rect 46572 4972 46624 4981
rect 47952 5040 48004 5092
rect 54668 5108 54720 5160
rect 55220 5108 55272 5160
rect 55404 5151 55456 5160
rect 55404 5117 55413 5151
rect 55413 5117 55447 5151
rect 55447 5117 55456 5151
rect 55404 5108 55456 5117
rect 55496 5108 55548 5160
rect 56416 5176 56468 5228
rect 57980 5219 58032 5228
rect 54576 5083 54628 5092
rect 54576 5049 54585 5083
rect 54585 5049 54619 5083
rect 54619 5049 54628 5083
rect 54576 5040 54628 5049
rect 48044 4972 48096 5024
rect 49516 4972 49568 5024
rect 51540 4972 51592 5024
rect 52552 4972 52604 5024
rect 57152 5108 57204 5160
rect 57980 5185 57989 5219
rect 57989 5185 58023 5219
rect 58023 5185 58032 5219
rect 57980 5176 58032 5185
rect 58624 5108 58676 5160
rect 59084 5151 59136 5160
rect 59084 5117 59093 5151
rect 59093 5117 59127 5151
rect 59127 5117 59136 5151
rect 59084 5108 59136 5117
rect 59268 5151 59320 5160
rect 59268 5117 59277 5151
rect 59277 5117 59311 5151
rect 59311 5117 59320 5151
rect 59268 5108 59320 5117
rect 59728 5151 59780 5160
rect 59728 5117 59737 5151
rect 59737 5117 59771 5151
rect 59771 5117 59780 5151
rect 59728 5108 59780 5117
rect 59820 5151 59872 5160
rect 59820 5117 59829 5151
rect 59829 5117 59863 5151
rect 59863 5117 59872 5151
rect 59820 5108 59872 5117
rect 61016 5108 61068 5160
rect 61200 5040 61252 5092
rect 56508 4972 56560 5024
rect 57060 5015 57112 5024
rect 57060 4981 57069 5015
rect 57069 4981 57103 5015
rect 57103 4981 57112 5015
rect 57060 4972 57112 4981
rect 60004 4972 60056 5024
rect 60464 4972 60516 5024
rect 61016 4972 61068 5024
rect 21774 4870 21826 4922
rect 21838 4870 21890 4922
rect 21902 4870 21954 4922
rect 21966 4870 22018 4922
rect 42566 4870 42618 4922
rect 42630 4870 42682 4922
rect 42694 4870 42746 4922
rect 42758 4870 42810 4922
rect 2504 4700 2556 4752
rect 12164 4768 12216 4820
rect 14924 4811 14976 4820
rect 14924 4777 14933 4811
rect 14933 4777 14967 4811
rect 14967 4777 14976 4811
rect 14924 4768 14976 4777
rect 15568 4768 15620 4820
rect 17224 4768 17276 4820
rect 17776 4768 17828 4820
rect 18052 4768 18104 4820
rect 21548 4768 21600 4820
rect 4068 4743 4120 4752
rect 4068 4709 4077 4743
rect 4077 4709 4111 4743
rect 4111 4709 4120 4743
rect 4068 4700 4120 4709
rect 2872 4632 2924 4684
rect 4528 4675 4580 4684
rect 4528 4641 4537 4675
rect 4537 4641 4571 4675
rect 4571 4641 4580 4675
rect 4528 4632 4580 4641
rect 5172 4632 5224 4684
rect 8760 4700 8812 4752
rect 8852 4700 8904 4752
rect 7840 4632 7892 4684
rect 8668 4632 8720 4684
rect 4804 4564 4856 4616
rect 7288 4607 7340 4616
rect 7288 4573 7297 4607
rect 7297 4573 7331 4607
rect 7331 4573 7340 4607
rect 9680 4632 9732 4684
rect 9772 4632 9824 4684
rect 10140 4632 10192 4684
rect 7288 4564 7340 4573
rect 8852 4564 8904 4616
rect 9588 4564 9640 4616
rect 11704 4632 11756 4684
rect 11888 4632 11940 4684
rect 12072 4700 12124 4752
rect 23940 4768 23992 4820
rect 24216 4768 24268 4820
rect 24400 4811 24452 4820
rect 24400 4777 24409 4811
rect 24409 4777 24443 4811
rect 24443 4777 24452 4811
rect 24400 4768 24452 4777
rect 24860 4811 24912 4820
rect 24860 4777 24869 4811
rect 24869 4777 24903 4811
rect 24903 4777 24912 4811
rect 24860 4768 24912 4777
rect 26056 4768 26108 4820
rect 22192 4700 22244 4752
rect 29828 4743 29880 4752
rect 29828 4709 29837 4743
rect 29837 4709 29871 4743
rect 29871 4709 29880 4743
rect 29828 4700 29880 4709
rect 11060 4564 11112 4616
rect 13912 4632 13964 4684
rect 10784 4496 10836 4548
rect 13084 4539 13136 4548
rect 13084 4505 13093 4539
rect 13093 4505 13127 4539
rect 13127 4505 13136 4539
rect 13084 4496 13136 4505
rect 14096 4564 14148 4616
rect 14740 4632 14792 4684
rect 16580 4675 16632 4684
rect 16212 4564 16264 4616
rect 16580 4641 16589 4675
rect 16589 4641 16623 4675
rect 16623 4641 16632 4675
rect 16580 4632 16632 4641
rect 16672 4632 16724 4684
rect 17408 4607 17460 4616
rect 17408 4573 17417 4607
rect 17417 4573 17451 4607
rect 17451 4573 17460 4607
rect 18144 4632 18196 4684
rect 18604 4675 18656 4684
rect 18604 4641 18613 4675
rect 18613 4641 18647 4675
rect 18647 4641 18656 4675
rect 18604 4632 18656 4641
rect 19340 4632 19392 4684
rect 19984 4632 20036 4684
rect 20904 4675 20956 4684
rect 20904 4641 20913 4675
rect 20913 4641 20947 4675
rect 20947 4641 20956 4675
rect 20904 4632 20956 4641
rect 21180 4675 21232 4684
rect 21180 4641 21189 4675
rect 21189 4641 21223 4675
rect 21223 4641 21232 4675
rect 21180 4632 21232 4641
rect 22928 4632 22980 4684
rect 23848 4675 23900 4684
rect 23848 4641 23857 4675
rect 23857 4641 23891 4675
rect 23891 4641 23900 4675
rect 23848 4632 23900 4641
rect 24492 4632 24544 4684
rect 25136 4675 25188 4684
rect 25136 4641 25145 4675
rect 25145 4641 25179 4675
rect 25179 4641 25188 4675
rect 25136 4632 25188 4641
rect 25320 4675 25372 4684
rect 25320 4641 25329 4675
rect 25329 4641 25363 4675
rect 25363 4641 25372 4675
rect 25320 4632 25372 4641
rect 27160 4675 27212 4684
rect 27160 4641 27169 4675
rect 27169 4641 27203 4675
rect 27203 4641 27212 4675
rect 27160 4632 27212 4641
rect 27436 4675 27488 4684
rect 27436 4641 27445 4675
rect 27445 4641 27479 4675
rect 27479 4641 27488 4675
rect 27436 4632 27488 4641
rect 17408 4564 17460 4573
rect 18328 4564 18380 4616
rect 18972 4564 19024 4616
rect 20720 4564 20772 4616
rect 21272 4564 21324 4616
rect 16672 4496 16724 4548
rect 25780 4564 25832 4616
rect 28632 4632 28684 4684
rect 28908 4632 28960 4684
rect 29000 4632 29052 4684
rect 29460 4632 29512 4684
rect 30472 4700 30524 4752
rect 30656 4700 30708 4752
rect 31760 4743 31812 4752
rect 31760 4709 31769 4743
rect 31769 4709 31803 4743
rect 31803 4709 31812 4743
rect 31760 4700 31812 4709
rect 38660 4700 38712 4752
rect 39580 4700 39632 4752
rect 39764 4768 39816 4820
rect 46572 4768 46624 4820
rect 47216 4768 47268 4820
rect 48136 4768 48188 4820
rect 49792 4811 49844 4820
rect 49792 4777 49801 4811
rect 49801 4777 49835 4811
rect 49835 4777 49844 4811
rect 49792 4768 49844 4777
rect 50068 4768 50120 4820
rect 50896 4768 50948 4820
rect 21548 4496 21600 4548
rect 3516 4471 3568 4480
rect 3516 4437 3525 4471
rect 3525 4437 3559 4471
rect 3559 4437 3568 4471
rect 3516 4428 3568 4437
rect 5356 4428 5408 4480
rect 7840 4428 7892 4480
rect 8024 4428 8076 4480
rect 8668 4428 8720 4480
rect 9496 4428 9548 4480
rect 10692 4428 10744 4480
rect 11244 4471 11296 4480
rect 11244 4437 11253 4471
rect 11253 4437 11287 4471
rect 11287 4437 11296 4471
rect 11244 4428 11296 4437
rect 11980 4428 12032 4480
rect 12532 4471 12584 4480
rect 12532 4437 12541 4471
rect 12541 4437 12575 4471
rect 12575 4437 12584 4471
rect 12532 4428 12584 4437
rect 12716 4428 12768 4480
rect 13360 4428 13412 4480
rect 13636 4428 13688 4480
rect 15200 4428 15252 4480
rect 15476 4471 15528 4480
rect 15476 4437 15485 4471
rect 15485 4437 15519 4471
rect 15519 4437 15528 4471
rect 15476 4428 15528 4437
rect 16120 4428 16172 4480
rect 17500 4428 17552 4480
rect 17960 4428 18012 4480
rect 19800 4471 19852 4480
rect 19800 4437 19809 4471
rect 19809 4437 19843 4471
rect 19843 4437 19852 4471
rect 19800 4428 19852 4437
rect 20260 4471 20312 4480
rect 20260 4437 20269 4471
rect 20269 4437 20303 4471
rect 20303 4437 20312 4471
rect 20260 4428 20312 4437
rect 20536 4428 20588 4480
rect 20720 4471 20772 4480
rect 20720 4437 20729 4471
rect 20729 4437 20763 4471
rect 20763 4437 20772 4471
rect 20720 4428 20772 4437
rect 22192 4471 22244 4480
rect 22192 4437 22201 4471
rect 22201 4437 22235 4471
rect 22235 4437 22244 4471
rect 22192 4428 22244 4437
rect 22652 4428 22704 4480
rect 23020 4428 23072 4480
rect 23664 4471 23716 4480
rect 23664 4437 23673 4471
rect 23673 4437 23707 4471
rect 23707 4437 23716 4471
rect 23664 4428 23716 4437
rect 24492 4428 24544 4480
rect 25780 4428 25832 4480
rect 26608 4496 26660 4548
rect 32772 4632 32824 4684
rect 30196 4564 30248 4616
rect 34428 4632 34480 4684
rect 34980 4675 35032 4684
rect 33508 4564 33560 4616
rect 34520 4564 34572 4616
rect 34980 4641 34989 4675
rect 34989 4641 35023 4675
rect 35023 4641 35032 4675
rect 34980 4632 35032 4641
rect 35440 4675 35492 4684
rect 35440 4641 35449 4675
rect 35449 4641 35483 4675
rect 35483 4641 35492 4675
rect 35440 4632 35492 4641
rect 36452 4675 36504 4684
rect 36452 4641 36461 4675
rect 36461 4641 36495 4675
rect 36495 4641 36504 4675
rect 36452 4632 36504 4641
rect 37924 4675 37976 4684
rect 37924 4641 37933 4675
rect 37933 4641 37967 4675
rect 37967 4641 37976 4675
rect 37924 4632 37976 4641
rect 39028 4632 39080 4684
rect 39856 4675 39908 4684
rect 39856 4641 39865 4675
rect 39865 4641 39899 4675
rect 39899 4641 39908 4675
rect 39856 4632 39908 4641
rect 40224 4675 40276 4684
rect 40224 4641 40233 4675
rect 40233 4641 40267 4675
rect 40267 4641 40276 4675
rect 40224 4632 40276 4641
rect 40316 4632 40368 4684
rect 27896 4428 27948 4480
rect 29644 4471 29696 4480
rect 29644 4437 29653 4471
rect 29653 4437 29687 4471
rect 29687 4437 29696 4471
rect 29644 4428 29696 4437
rect 30288 4496 30340 4548
rect 30472 4428 30524 4480
rect 31852 4496 31904 4548
rect 32312 4496 32364 4548
rect 32496 4496 32548 4548
rect 32956 4496 33008 4548
rect 33140 4539 33192 4548
rect 33140 4505 33149 4539
rect 33149 4505 33183 4539
rect 33183 4505 33192 4539
rect 33140 4496 33192 4505
rect 35808 4564 35860 4616
rect 35992 4564 36044 4616
rect 37188 4564 37240 4616
rect 37556 4564 37608 4616
rect 37924 4496 37976 4548
rect 38568 4496 38620 4548
rect 38752 4496 38804 4548
rect 39580 4564 39632 4616
rect 42156 4632 42208 4684
rect 43812 4700 43864 4752
rect 44088 4700 44140 4752
rect 47124 4743 47176 4752
rect 47124 4709 47133 4743
rect 47133 4709 47167 4743
rect 47167 4709 47176 4743
rect 47124 4700 47176 4709
rect 47492 4743 47544 4752
rect 47492 4709 47501 4743
rect 47501 4709 47535 4743
rect 47535 4709 47544 4743
rect 47492 4700 47544 4709
rect 48964 4700 49016 4752
rect 49608 4700 49660 4752
rect 41972 4564 42024 4616
rect 40040 4496 40092 4548
rect 43628 4632 43680 4684
rect 46112 4675 46164 4684
rect 45652 4607 45704 4616
rect 45652 4573 45661 4607
rect 45661 4573 45695 4607
rect 45695 4573 45704 4607
rect 45652 4564 45704 4573
rect 42432 4496 42484 4548
rect 46112 4641 46121 4675
rect 46121 4641 46155 4675
rect 46155 4641 46164 4675
rect 46112 4632 46164 4641
rect 46296 4675 46348 4684
rect 46296 4641 46305 4675
rect 46305 4641 46339 4675
rect 46339 4641 46348 4675
rect 46296 4632 46348 4641
rect 47584 4632 47636 4684
rect 48136 4632 48188 4684
rect 49700 4632 49752 4684
rect 50344 4700 50396 4752
rect 57060 4768 57112 4820
rect 57336 4811 57388 4820
rect 57336 4777 57345 4811
rect 57345 4777 57379 4811
rect 57379 4777 57388 4811
rect 57336 4768 57388 4777
rect 58072 4811 58124 4820
rect 58072 4777 58081 4811
rect 58081 4777 58115 4811
rect 58115 4777 58124 4811
rect 58072 4768 58124 4777
rect 51540 4743 51592 4752
rect 51540 4709 51549 4743
rect 51549 4709 51583 4743
rect 51583 4709 51592 4743
rect 51540 4700 51592 4709
rect 51816 4700 51868 4752
rect 52276 4743 52328 4752
rect 52276 4709 52285 4743
rect 52285 4709 52319 4743
rect 52319 4709 52328 4743
rect 52276 4700 52328 4709
rect 52368 4700 52420 4752
rect 53656 4700 53708 4752
rect 55404 4743 55456 4752
rect 52000 4632 52052 4684
rect 53196 4632 53248 4684
rect 55404 4709 55413 4743
rect 55413 4709 55447 4743
rect 55447 4709 55456 4743
rect 55404 4700 55456 4709
rect 54484 4632 54536 4684
rect 54760 4632 54812 4684
rect 61568 4768 61620 4820
rect 59820 4700 59872 4752
rect 58348 4632 58400 4684
rect 59084 4675 59136 4684
rect 59084 4641 59093 4675
rect 59093 4641 59127 4675
rect 59127 4641 59136 4675
rect 59084 4632 59136 4641
rect 61016 4675 61068 4684
rect 61016 4641 61025 4675
rect 61025 4641 61059 4675
rect 61059 4641 61068 4675
rect 61016 4632 61068 4641
rect 61200 4675 61252 4684
rect 61200 4641 61209 4675
rect 61209 4641 61243 4675
rect 61243 4641 61252 4675
rect 61200 4632 61252 4641
rect 47860 4607 47912 4616
rect 47860 4573 47869 4607
rect 47869 4573 47903 4607
rect 47903 4573 47912 4607
rect 47860 4564 47912 4573
rect 48872 4564 48924 4616
rect 50620 4564 50672 4616
rect 33324 4428 33376 4480
rect 33968 4471 34020 4480
rect 33968 4437 33977 4471
rect 33977 4437 34011 4471
rect 34011 4437 34020 4471
rect 33968 4428 34020 4437
rect 35440 4428 35492 4480
rect 36452 4428 36504 4480
rect 37372 4471 37424 4480
rect 37372 4437 37381 4471
rect 37381 4437 37415 4471
rect 37415 4437 37424 4471
rect 37372 4428 37424 4437
rect 40868 4428 40920 4480
rect 43628 4471 43680 4480
rect 43628 4437 43637 4471
rect 43637 4437 43671 4471
rect 43671 4437 43680 4471
rect 43628 4428 43680 4437
rect 44180 4471 44232 4480
rect 44180 4437 44189 4471
rect 44189 4437 44223 4471
rect 44223 4437 44232 4471
rect 44180 4428 44232 4437
rect 45560 4428 45612 4480
rect 51172 4496 51224 4548
rect 48136 4428 48188 4480
rect 48688 4428 48740 4480
rect 49148 4471 49200 4480
rect 49148 4437 49157 4471
rect 49157 4437 49191 4471
rect 49191 4437 49200 4471
rect 49148 4428 49200 4437
rect 50988 4428 51040 4480
rect 51448 4496 51500 4548
rect 52368 4496 52420 4548
rect 51540 4428 51592 4480
rect 51908 4428 51960 4480
rect 52184 4428 52236 4480
rect 52736 4428 52788 4480
rect 54024 4564 54076 4616
rect 56048 4607 56100 4616
rect 54300 4539 54352 4548
rect 54300 4505 54309 4539
rect 54309 4505 54343 4539
rect 54343 4505 54352 4539
rect 54300 4496 54352 4505
rect 54668 4496 54720 4548
rect 55128 4428 55180 4480
rect 56048 4573 56057 4607
rect 56057 4573 56091 4607
rect 56091 4573 56100 4607
rect 56048 4564 56100 4573
rect 58900 4564 58952 4616
rect 59268 4607 59320 4616
rect 59268 4573 59277 4607
rect 59277 4573 59311 4607
rect 59311 4573 59320 4607
rect 59268 4564 59320 4573
rect 59360 4564 59412 4616
rect 61752 4564 61804 4616
rect 59452 4496 59504 4548
rect 58440 4428 58492 4480
rect 59544 4471 59596 4480
rect 59544 4437 59553 4471
rect 59553 4437 59587 4471
rect 59587 4437 59596 4471
rect 59544 4428 59596 4437
rect 61476 4471 61528 4480
rect 61476 4437 61485 4471
rect 61485 4437 61519 4471
rect 61519 4437 61528 4471
rect 61476 4428 61528 4437
rect 11378 4326 11430 4378
rect 11442 4326 11494 4378
rect 11506 4326 11558 4378
rect 11570 4326 11622 4378
rect 32170 4326 32222 4378
rect 32234 4326 32286 4378
rect 32298 4326 32350 4378
rect 32362 4326 32414 4378
rect 52962 4326 53014 4378
rect 53026 4326 53078 4378
rect 53090 4326 53142 4378
rect 53154 4326 53206 4378
rect 2504 4267 2556 4276
rect 2504 4233 2513 4267
rect 2513 4233 2547 4267
rect 2547 4233 2556 4267
rect 2504 4224 2556 4233
rect 3608 4267 3660 4276
rect 3608 4233 3617 4267
rect 3617 4233 3651 4267
rect 3651 4233 3660 4267
rect 3608 4224 3660 4233
rect 4528 4224 4580 4276
rect 7288 4267 7340 4276
rect 7288 4233 7297 4267
rect 7297 4233 7331 4267
rect 7331 4233 7340 4267
rect 7288 4224 7340 4233
rect 8760 4267 8812 4276
rect 8760 4233 8769 4267
rect 8769 4233 8803 4267
rect 8803 4233 8812 4267
rect 8760 4224 8812 4233
rect 9588 4224 9640 4276
rect 11704 4224 11756 4276
rect 12256 4267 12308 4276
rect 12256 4233 12265 4267
rect 12265 4233 12299 4267
rect 12299 4233 12308 4267
rect 12256 4224 12308 4233
rect 12440 4224 12492 4276
rect 12716 4267 12768 4276
rect 12716 4233 12725 4267
rect 12725 4233 12759 4267
rect 12759 4233 12768 4267
rect 12716 4224 12768 4233
rect 13912 4267 13964 4276
rect 5172 4199 5224 4208
rect 5172 4165 5181 4199
rect 5181 4165 5215 4199
rect 5215 4165 5224 4199
rect 5172 4156 5224 4165
rect 8852 4156 8904 4208
rect 9496 4156 9548 4208
rect 3700 4131 3752 4140
rect 3700 4097 3709 4131
rect 3709 4097 3743 4131
rect 3743 4097 3752 4131
rect 3700 4088 3752 4097
rect 7012 4088 7064 4140
rect 10416 4156 10468 4208
rect 11888 4199 11940 4208
rect 3056 4020 3108 4072
rect 3516 4063 3568 4072
rect 3516 4029 3522 4063
rect 3522 4029 3568 4063
rect 4068 4063 4120 4072
rect 3516 4020 3568 4029
rect 4068 4029 4077 4063
rect 4077 4029 4111 4063
rect 4111 4029 4120 4063
rect 4068 4020 4120 4029
rect 5356 4063 5408 4072
rect 5356 4029 5365 4063
rect 5365 4029 5399 4063
rect 5399 4029 5408 4063
rect 5356 4020 5408 4029
rect 8024 4020 8076 4072
rect 9864 4063 9916 4072
rect 9864 4029 9870 4063
rect 9870 4029 9916 4063
rect 9864 4020 9916 4029
rect 11060 4088 11112 4140
rect 11888 4165 11897 4199
rect 11897 4165 11931 4199
rect 11931 4165 11940 4199
rect 11888 4156 11940 4165
rect 13912 4233 13921 4267
rect 13921 4233 13955 4267
rect 13955 4233 13964 4267
rect 13912 4224 13964 4233
rect 16580 4224 16632 4276
rect 16672 4224 16724 4276
rect 17500 4224 17552 4276
rect 20812 4224 20864 4276
rect 22192 4224 22244 4276
rect 23572 4224 23624 4276
rect 23848 4267 23900 4276
rect 23848 4233 23857 4267
rect 23857 4233 23891 4267
rect 23891 4233 23900 4267
rect 23848 4224 23900 4233
rect 23940 4224 23992 4276
rect 27436 4267 27488 4276
rect 14832 4199 14884 4208
rect 3332 3995 3384 4004
rect 3332 3961 3341 3995
rect 3341 3961 3375 3995
rect 3375 3961 3384 3995
rect 3332 3952 3384 3961
rect 3608 3952 3660 4004
rect 5632 3952 5684 4004
rect 9496 3952 9548 4004
rect 10784 4020 10836 4072
rect 11244 4063 11296 4072
rect 11244 4029 11253 4063
rect 11253 4029 11287 4063
rect 11287 4029 11296 4063
rect 13360 4088 13412 4140
rect 13728 4088 13780 4140
rect 14832 4165 14841 4199
rect 14841 4165 14875 4199
rect 14875 4165 14884 4199
rect 14832 4156 14884 4165
rect 14924 4156 14976 4208
rect 17408 4156 17460 4208
rect 19248 4156 19300 4208
rect 25596 4156 25648 4208
rect 20904 4088 20956 4140
rect 21088 4088 21140 4140
rect 21180 4088 21232 4140
rect 22008 4088 22060 4140
rect 22100 4088 22152 4140
rect 11244 4020 11296 4029
rect 13176 4020 13228 4072
rect 14188 4020 14240 4072
rect 14372 4063 14424 4072
rect 14372 4029 14381 4063
rect 14381 4029 14415 4063
rect 14415 4029 14424 4063
rect 14372 4020 14424 4029
rect 14464 4020 14516 4072
rect 12532 3952 12584 4004
rect 2872 3927 2924 3936
rect 2872 3893 2881 3927
rect 2881 3893 2915 3927
rect 2915 3893 2924 3927
rect 2872 3884 2924 3893
rect 6552 3884 6604 3936
rect 7104 3884 7156 3936
rect 7472 3884 7524 3936
rect 7840 3884 7892 3936
rect 8024 3884 8076 3936
rect 9772 3884 9824 3936
rect 10692 3927 10744 3936
rect 10692 3893 10701 3927
rect 10701 3893 10735 3927
rect 10735 3893 10744 3927
rect 10692 3884 10744 3893
rect 10784 3884 10836 3936
rect 13636 3952 13688 4004
rect 15200 4020 15252 4072
rect 18788 4063 18840 4072
rect 15660 3952 15712 4004
rect 15936 3952 15988 4004
rect 18788 4029 18797 4063
rect 18797 4029 18831 4063
rect 18831 4029 18840 4063
rect 18788 4020 18840 4029
rect 20536 4063 20588 4072
rect 18236 3952 18288 4004
rect 20168 3952 20220 4004
rect 20536 4029 20545 4063
rect 20545 4029 20579 4063
rect 20579 4029 20588 4063
rect 20536 4020 20588 4029
rect 20628 4020 20680 4072
rect 22192 3995 22244 4004
rect 22192 3961 22201 3995
rect 22201 3961 22235 3995
rect 22235 3961 22244 3995
rect 22192 3952 22244 3961
rect 22652 4020 22704 4072
rect 24308 4020 24360 4072
rect 25320 4088 25372 4140
rect 25412 4088 25464 4140
rect 27436 4233 27445 4267
rect 27445 4233 27479 4267
rect 27479 4233 27488 4267
rect 27436 4224 27488 4233
rect 29460 4224 29512 4276
rect 31024 4224 31076 4276
rect 25780 4088 25832 4140
rect 29368 4156 29420 4208
rect 30288 4156 30340 4208
rect 24676 4063 24728 4072
rect 24676 4029 24685 4063
rect 24685 4029 24719 4063
rect 24719 4029 24728 4063
rect 24676 4020 24728 4029
rect 24768 4020 24820 4072
rect 26332 4063 26384 4072
rect 26332 4029 26341 4063
rect 26341 4029 26375 4063
rect 26375 4029 26384 4063
rect 26332 4020 26384 4029
rect 27252 4020 27304 4072
rect 27620 4020 27672 4072
rect 29644 4088 29696 4140
rect 32036 4224 32088 4276
rect 33968 4224 34020 4276
rect 34244 4267 34296 4276
rect 34244 4233 34253 4267
rect 34253 4233 34287 4267
rect 34287 4233 34296 4267
rect 34244 4224 34296 4233
rect 34520 4224 34572 4276
rect 35808 4224 35860 4276
rect 36268 4224 36320 4276
rect 39028 4224 39080 4276
rect 40316 4267 40368 4276
rect 40316 4233 40325 4267
rect 40325 4233 40359 4267
rect 40359 4233 40368 4267
rect 40316 4224 40368 4233
rect 40408 4224 40460 4276
rect 41972 4224 42024 4276
rect 31300 4156 31352 4208
rect 32220 4131 32272 4140
rect 27896 4063 27948 4072
rect 27896 4029 27905 4063
rect 27905 4029 27939 4063
rect 27939 4029 27948 4063
rect 27896 4020 27948 4029
rect 28172 4020 28224 4072
rect 30012 4020 30064 4072
rect 30472 4020 30524 4072
rect 30748 4063 30800 4072
rect 30748 4029 30757 4063
rect 30757 4029 30791 4063
rect 30791 4029 30800 4063
rect 30748 4020 30800 4029
rect 31392 4020 31444 4072
rect 32220 4097 32229 4131
rect 32229 4097 32263 4131
rect 32263 4097 32272 4131
rect 32220 4088 32272 4097
rect 34428 4156 34480 4208
rect 39764 4156 39816 4208
rect 39856 4156 39908 4208
rect 42432 4156 42484 4208
rect 43628 4156 43680 4208
rect 44180 4224 44232 4276
rect 46756 4224 46808 4276
rect 47032 4224 47084 4276
rect 47952 4224 48004 4276
rect 49148 4199 49200 4208
rect 49148 4165 49157 4199
rect 49157 4165 49191 4199
rect 49191 4165 49200 4199
rect 49148 4156 49200 4165
rect 52552 4156 52604 4208
rect 53288 4156 53340 4208
rect 54484 4199 54536 4208
rect 54484 4165 54493 4199
rect 54493 4165 54527 4199
rect 54527 4165 54536 4199
rect 54484 4156 54536 4165
rect 55036 4156 55088 4208
rect 32588 4020 32640 4072
rect 36084 4088 36136 4140
rect 37188 4088 37240 4140
rect 39580 4131 39632 4140
rect 33508 4063 33560 4072
rect 33508 4029 33517 4063
rect 33517 4029 33551 4063
rect 33551 4029 33560 4063
rect 33508 4020 33560 4029
rect 34244 4020 34296 4072
rect 34520 4020 34572 4072
rect 35992 4063 36044 4072
rect 35992 4029 36001 4063
rect 36001 4029 36035 4063
rect 36035 4029 36044 4063
rect 35992 4020 36044 4029
rect 36268 4063 36320 4072
rect 36268 4029 36277 4063
rect 36277 4029 36311 4063
rect 36311 4029 36320 4063
rect 36268 4020 36320 4029
rect 36452 4020 36504 4072
rect 37924 4020 37976 4072
rect 38936 4020 38988 4072
rect 39580 4097 39589 4131
rect 39589 4097 39623 4131
rect 39623 4097 39632 4131
rect 39580 4088 39632 4097
rect 40960 4020 41012 4072
rect 42064 4063 42116 4072
rect 13452 3884 13504 3936
rect 15108 3884 15160 3936
rect 16488 3927 16540 3936
rect 16488 3893 16497 3927
rect 16497 3893 16531 3927
rect 16531 3893 16540 3927
rect 16488 3884 16540 3893
rect 16580 3927 16632 3936
rect 16580 3893 16589 3927
rect 16589 3893 16623 3927
rect 16623 3893 16632 3927
rect 16580 3884 16632 3893
rect 22376 3884 22428 3936
rect 22652 3884 22704 3936
rect 23388 3927 23440 3936
rect 23388 3893 23397 3927
rect 23397 3893 23431 3927
rect 23431 3893 23440 3927
rect 23388 3884 23440 3893
rect 24952 3927 25004 3936
rect 24952 3893 24961 3927
rect 24961 3893 24995 3927
rect 24995 3893 25004 3927
rect 24952 3884 25004 3893
rect 25136 3952 25188 4004
rect 26516 3952 26568 4004
rect 27804 3995 27856 4004
rect 27804 3961 27813 3995
rect 27813 3961 27847 3995
rect 27847 3961 27856 3995
rect 27804 3952 27856 3961
rect 28356 3995 28408 4004
rect 28356 3961 28365 3995
rect 28365 3961 28399 3995
rect 28399 3961 28408 3995
rect 28356 3952 28408 3961
rect 25596 3884 25648 3936
rect 27160 3927 27212 3936
rect 27160 3893 27169 3927
rect 27169 3893 27203 3927
rect 27203 3893 27212 3927
rect 28632 3927 28684 3936
rect 27160 3884 27212 3893
rect 28632 3893 28641 3927
rect 28641 3893 28675 3927
rect 28675 3893 28684 3927
rect 28632 3884 28684 3893
rect 30196 3952 30248 4004
rect 31944 3952 31996 4004
rect 30656 3884 30708 3936
rect 31484 3884 31536 3936
rect 32772 3927 32824 3936
rect 32772 3893 32781 3927
rect 32781 3893 32815 3927
rect 32815 3893 32824 3927
rect 32772 3884 32824 3893
rect 34980 3952 35032 4004
rect 37740 3952 37792 4004
rect 38752 3952 38804 4004
rect 42064 4029 42073 4063
rect 42073 4029 42107 4063
rect 42107 4029 42116 4063
rect 42064 4020 42116 4029
rect 45652 4088 45704 4140
rect 44180 3995 44232 4004
rect 44180 3961 44189 3995
rect 44189 3961 44223 3995
rect 44223 3961 44232 3995
rect 44180 3952 44232 3961
rect 35992 3884 36044 3936
rect 36176 3884 36228 3936
rect 41604 3927 41656 3936
rect 41604 3893 41613 3927
rect 41613 3893 41647 3927
rect 41647 3893 41656 3927
rect 41604 3884 41656 3893
rect 42156 3884 42208 3936
rect 44732 3884 44784 3936
rect 44824 3884 44876 3936
rect 45100 3952 45152 4004
rect 46940 4020 46992 4072
rect 47032 4063 47084 4072
rect 47032 4029 47041 4063
rect 47041 4029 47075 4063
rect 47075 4029 47084 4063
rect 47952 4088 48004 4140
rect 49240 4088 49292 4140
rect 50620 4088 50672 4140
rect 52184 4088 52236 4140
rect 52828 4088 52880 4140
rect 47032 4020 47084 4029
rect 46296 3995 46348 4004
rect 46296 3961 46305 3995
rect 46305 3961 46339 3995
rect 46339 3961 46348 3995
rect 46296 3952 46348 3961
rect 48412 4020 48464 4072
rect 48504 4020 48556 4072
rect 48688 4020 48740 4072
rect 49792 4020 49844 4072
rect 51724 4063 51776 4072
rect 46020 3884 46072 3936
rect 46204 3884 46256 3936
rect 47492 3884 47544 3936
rect 48320 3884 48372 3936
rect 48872 3884 48924 3936
rect 50068 3884 50120 3936
rect 50252 3884 50304 3936
rect 51080 3927 51132 3936
rect 51080 3893 51089 3927
rect 51089 3893 51123 3927
rect 51123 3893 51132 3927
rect 51724 4029 51733 4063
rect 51733 4029 51767 4063
rect 51767 4029 51776 4063
rect 51724 4020 51776 4029
rect 51816 4063 51868 4072
rect 51816 4029 51825 4063
rect 51825 4029 51859 4063
rect 51859 4029 51868 4063
rect 51816 4020 51868 4029
rect 52552 4020 52604 4072
rect 53380 4063 53432 4072
rect 53380 4029 53389 4063
rect 53389 4029 53423 4063
rect 53423 4029 53432 4063
rect 53380 4020 53432 4029
rect 53564 4020 53616 4072
rect 53656 4063 53708 4072
rect 53656 4029 53665 4063
rect 53665 4029 53699 4063
rect 53699 4029 53708 4063
rect 54116 4088 54168 4140
rect 54760 4088 54812 4140
rect 55220 4088 55272 4140
rect 53656 4020 53708 4029
rect 52000 3952 52052 4004
rect 53932 3952 53984 4004
rect 54668 3995 54720 4004
rect 54668 3961 54677 3995
rect 54677 3961 54711 3995
rect 54711 3961 54720 3995
rect 54668 3952 54720 3961
rect 55128 4020 55180 4072
rect 56140 4156 56192 4208
rect 59268 4224 59320 4276
rect 61200 4224 61252 4276
rect 59544 4088 59596 4140
rect 61016 4088 61068 4140
rect 51080 3884 51132 3893
rect 53288 3884 53340 3936
rect 53380 3884 53432 3936
rect 54852 3884 54904 3936
rect 55036 3995 55088 4004
rect 55036 3961 55045 3995
rect 55045 3961 55079 3995
rect 55079 3961 55088 3995
rect 55036 3952 55088 3961
rect 55220 3952 55272 4004
rect 58072 4020 58124 4072
rect 58440 4020 58492 4072
rect 57612 3952 57664 4004
rect 55588 3884 55640 3936
rect 55680 3884 55732 3936
rect 56048 3927 56100 3936
rect 56048 3893 56057 3927
rect 56057 3893 56091 3927
rect 56091 3893 56100 3927
rect 56048 3884 56100 3893
rect 57336 3884 57388 3936
rect 61476 4020 61528 4072
rect 61752 4088 61804 4140
rect 21774 3782 21826 3834
rect 21838 3782 21890 3834
rect 21902 3782 21954 3834
rect 21966 3782 22018 3834
rect 42566 3782 42618 3834
rect 42630 3782 42682 3834
rect 42694 3782 42746 3834
rect 42758 3782 42810 3834
rect 3332 3680 3384 3732
rect 4804 3680 4856 3732
rect 5724 3680 5776 3732
rect 7472 3680 7524 3732
rect 7840 3680 7892 3732
rect 8576 3680 8628 3732
rect 9588 3680 9640 3732
rect 9864 3680 9916 3732
rect 14096 3723 14148 3732
rect 2228 3612 2280 3664
rect 2872 3544 2924 3596
rect 3424 3544 3476 3596
rect 3792 3544 3844 3596
rect 7932 3612 7984 3664
rect 8944 3612 8996 3664
rect 5908 3587 5960 3596
rect 5908 3553 5917 3587
rect 5917 3553 5951 3587
rect 5951 3553 5960 3587
rect 5908 3544 5960 3553
rect 6644 3544 6696 3596
rect 7748 3544 7800 3596
rect 8300 3544 8352 3596
rect 10140 3587 10192 3596
rect 10140 3553 10149 3587
rect 10149 3553 10183 3587
rect 10183 3553 10192 3587
rect 10140 3544 10192 3553
rect 14096 3689 14105 3723
rect 14105 3689 14139 3723
rect 14139 3689 14148 3723
rect 14096 3680 14148 3689
rect 16580 3680 16632 3732
rect 12256 3587 12308 3596
rect 2780 3476 2832 3528
rect 6184 3476 6236 3528
rect 5724 3408 5776 3460
rect 5356 3383 5408 3392
rect 5356 3349 5365 3383
rect 5365 3349 5399 3383
rect 5399 3349 5408 3383
rect 5356 3340 5408 3349
rect 9312 3476 9364 3528
rect 7012 3408 7064 3460
rect 7656 3408 7708 3460
rect 9036 3408 9088 3460
rect 9404 3408 9456 3460
rect 9680 3408 9732 3460
rect 12256 3553 12265 3587
rect 12265 3553 12299 3587
rect 12299 3553 12308 3587
rect 12256 3544 12308 3553
rect 12624 3544 12676 3596
rect 12808 3587 12860 3596
rect 12808 3553 12817 3587
rect 12817 3553 12851 3587
rect 12851 3553 12860 3587
rect 12808 3544 12860 3553
rect 12900 3544 12952 3596
rect 17684 3612 17736 3664
rect 15660 3587 15712 3596
rect 15660 3553 15669 3587
rect 15669 3553 15703 3587
rect 15703 3553 15712 3587
rect 16212 3587 16264 3596
rect 15660 3544 15712 3553
rect 16212 3553 16221 3587
rect 16221 3553 16255 3587
rect 16255 3553 16264 3587
rect 16212 3544 16264 3553
rect 17408 3587 17460 3596
rect 17408 3553 17417 3587
rect 17417 3553 17451 3587
rect 17451 3553 17460 3587
rect 17408 3544 17460 3553
rect 17868 3544 17920 3596
rect 18052 3680 18104 3732
rect 19524 3680 19576 3732
rect 18236 3612 18288 3664
rect 20444 3680 20496 3732
rect 20812 3680 20864 3732
rect 22376 3680 22428 3732
rect 23020 3680 23072 3732
rect 23112 3680 23164 3732
rect 23848 3680 23900 3732
rect 25044 3680 25096 3732
rect 25596 3680 25648 3732
rect 26332 3680 26384 3732
rect 26424 3680 26476 3732
rect 31852 3680 31904 3732
rect 32036 3680 32088 3732
rect 32772 3680 32824 3732
rect 23664 3612 23716 3664
rect 23756 3612 23808 3664
rect 25228 3612 25280 3664
rect 11244 3519 11296 3528
rect 11244 3485 11253 3519
rect 11253 3485 11287 3519
rect 11287 3485 11296 3519
rect 11244 3476 11296 3485
rect 11612 3451 11664 3460
rect 11612 3417 11621 3451
rect 11621 3417 11655 3451
rect 11655 3417 11664 3451
rect 11612 3408 11664 3417
rect 6828 3383 6880 3392
rect 6828 3349 6837 3383
rect 6837 3349 6871 3383
rect 6871 3349 6880 3383
rect 6828 3340 6880 3349
rect 7196 3383 7248 3392
rect 7196 3349 7205 3383
rect 7205 3349 7239 3383
rect 7239 3349 7248 3383
rect 7196 3340 7248 3349
rect 7288 3340 7340 3392
rect 10876 3340 10928 3392
rect 13452 3476 13504 3528
rect 15016 3519 15068 3528
rect 15016 3485 15025 3519
rect 15025 3485 15059 3519
rect 15059 3485 15068 3519
rect 15016 3476 15068 3485
rect 15936 3476 15988 3528
rect 18328 3476 18380 3528
rect 18696 3544 18748 3596
rect 20996 3544 21048 3596
rect 21272 3544 21324 3596
rect 23572 3544 23624 3596
rect 24860 3544 24912 3596
rect 25320 3587 25372 3596
rect 25320 3553 25329 3587
rect 25329 3553 25363 3587
rect 25363 3553 25372 3587
rect 25320 3544 25372 3553
rect 26516 3587 26568 3596
rect 26516 3553 26525 3587
rect 26525 3553 26559 3587
rect 26559 3553 26568 3587
rect 26516 3544 26568 3553
rect 26792 3544 26844 3596
rect 28080 3587 28132 3596
rect 28080 3553 28089 3587
rect 28089 3553 28123 3587
rect 28123 3553 28132 3587
rect 28080 3544 28132 3553
rect 28264 3587 28316 3596
rect 28264 3553 28273 3587
rect 28273 3553 28307 3587
rect 28307 3553 28316 3587
rect 28264 3544 28316 3553
rect 29092 3612 29144 3664
rect 30472 3612 30524 3664
rect 33508 3612 33560 3664
rect 28908 3544 28960 3596
rect 29920 3544 29972 3596
rect 30288 3544 30340 3596
rect 30564 3587 30616 3596
rect 30564 3553 30573 3587
rect 30573 3553 30607 3587
rect 30607 3553 30616 3587
rect 30564 3544 30616 3553
rect 30656 3544 30708 3596
rect 33968 3544 34020 3596
rect 36728 3680 36780 3732
rect 37740 3680 37792 3732
rect 36268 3612 36320 3664
rect 38016 3680 38068 3732
rect 38844 3680 38896 3732
rect 38936 3680 38988 3732
rect 41236 3680 41288 3732
rect 41972 3723 42024 3732
rect 41972 3689 41981 3723
rect 41981 3689 42015 3723
rect 42015 3689 42024 3723
rect 41972 3680 42024 3689
rect 41420 3612 41472 3664
rect 41604 3655 41656 3664
rect 41604 3621 41613 3655
rect 41613 3621 41647 3655
rect 41647 3621 41656 3655
rect 46204 3680 46256 3732
rect 46296 3680 46348 3732
rect 48044 3680 48096 3732
rect 48964 3680 49016 3732
rect 49056 3680 49108 3732
rect 49884 3723 49936 3732
rect 49884 3689 49893 3723
rect 49893 3689 49927 3723
rect 49927 3689 49936 3723
rect 49884 3680 49936 3689
rect 50068 3680 50120 3732
rect 41604 3612 41656 3621
rect 44824 3612 44876 3664
rect 46940 3612 46992 3664
rect 47216 3655 47268 3664
rect 47216 3621 47225 3655
rect 47225 3621 47259 3655
rect 47259 3621 47268 3655
rect 47216 3612 47268 3621
rect 47400 3612 47452 3664
rect 34428 3544 34480 3596
rect 34704 3587 34756 3596
rect 34704 3553 34713 3587
rect 34713 3553 34747 3587
rect 34747 3553 34756 3587
rect 34704 3544 34756 3553
rect 19616 3519 19668 3528
rect 12348 3408 12400 3460
rect 14096 3408 14148 3460
rect 19616 3485 19625 3519
rect 19625 3485 19659 3519
rect 19659 3485 19668 3519
rect 19616 3476 19668 3485
rect 20076 3476 20128 3528
rect 21364 3476 21416 3528
rect 23388 3519 23440 3528
rect 23388 3485 23397 3519
rect 23397 3485 23431 3519
rect 23431 3485 23440 3519
rect 23388 3476 23440 3485
rect 23756 3476 23808 3528
rect 24584 3476 24636 3528
rect 24768 3476 24820 3528
rect 27620 3519 27672 3528
rect 27620 3485 27629 3519
rect 27629 3485 27663 3519
rect 27663 3485 27672 3519
rect 27620 3476 27672 3485
rect 12900 3340 12952 3392
rect 13268 3383 13320 3392
rect 13268 3349 13277 3383
rect 13277 3349 13311 3383
rect 13311 3349 13320 3383
rect 13268 3340 13320 3349
rect 13820 3383 13872 3392
rect 13820 3349 13829 3383
rect 13829 3349 13863 3383
rect 13863 3349 13872 3383
rect 13820 3340 13872 3349
rect 14372 3340 14424 3392
rect 15936 3340 15988 3392
rect 16120 3340 16172 3392
rect 18604 3340 18656 3392
rect 19248 3340 19300 3392
rect 20260 3408 20312 3460
rect 20444 3408 20496 3460
rect 22468 3408 22520 3460
rect 21824 3340 21876 3392
rect 22744 3340 22796 3392
rect 24492 3340 24544 3392
rect 24584 3340 24636 3392
rect 26516 3408 26568 3460
rect 26792 3408 26844 3460
rect 27896 3408 27948 3460
rect 26148 3340 26200 3392
rect 26332 3383 26384 3392
rect 26332 3349 26341 3383
rect 26341 3349 26375 3383
rect 26375 3349 26384 3383
rect 26332 3340 26384 3349
rect 26976 3340 27028 3392
rect 27252 3340 27304 3392
rect 27436 3383 27488 3392
rect 27436 3349 27445 3383
rect 27445 3349 27479 3383
rect 27479 3349 27488 3383
rect 27436 3340 27488 3349
rect 31760 3476 31812 3528
rect 31944 3476 31996 3528
rect 32680 3476 32732 3528
rect 31024 3408 31076 3460
rect 34336 3408 34388 3460
rect 35900 3544 35952 3596
rect 36360 3544 36412 3596
rect 38476 3544 38528 3596
rect 38752 3544 38804 3596
rect 40316 3544 40368 3596
rect 40684 3587 40736 3596
rect 40684 3553 40693 3587
rect 40693 3553 40727 3587
rect 40727 3553 40736 3587
rect 40684 3544 40736 3553
rect 42064 3587 42116 3596
rect 42064 3553 42073 3587
rect 42073 3553 42107 3587
rect 42107 3553 42116 3587
rect 42064 3544 42116 3553
rect 43076 3544 43128 3596
rect 43720 3587 43772 3596
rect 43720 3553 43729 3587
rect 43729 3553 43763 3587
rect 43763 3553 43772 3587
rect 43720 3544 43772 3553
rect 39212 3519 39264 3528
rect 39212 3485 39221 3519
rect 39221 3485 39255 3519
rect 39255 3485 39264 3519
rect 39212 3476 39264 3485
rect 40592 3519 40644 3528
rect 40592 3485 40601 3519
rect 40601 3485 40635 3519
rect 40635 3485 40644 3519
rect 40592 3476 40644 3485
rect 36636 3408 36688 3460
rect 45192 3544 45244 3596
rect 45560 3587 45612 3596
rect 45560 3553 45569 3587
rect 45569 3553 45603 3587
rect 45603 3553 45612 3587
rect 45560 3544 45612 3553
rect 46204 3544 46256 3596
rect 46756 3544 46808 3596
rect 47860 3544 47912 3596
rect 48872 3544 48924 3596
rect 50804 3612 50856 3664
rect 50068 3587 50120 3596
rect 50068 3553 50077 3587
rect 50077 3553 50111 3587
rect 50111 3553 50120 3587
rect 50068 3544 50120 3553
rect 51080 3587 51132 3596
rect 51080 3553 51089 3587
rect 51089 3553 51123 3587
rect 51123 3553 51132 3587
rect 51080 3544 51132 3553
rect 51724 3544 51776 3596
rect 52000 3587 52052 3596
rect 52000 3553 52009 3587
rect 52009 3553 52043 3587
rect 52043 3553 52052 3587
rect 52000 3544 52052 3553
rect 52184 3544 52236 3596
rect 52368 3680 52420 3732
rect 54024 3680 54076 3732
rect 54852 3680 54904 3732
rect 56232 3723 56284 3732
rect 52368 3544 52420 3596
rect 53380 3587 53432 3596
rect 33048 3340 33100 3392
rect 33232 3383 33284 3392
rect 33232 3349 33241 3383
rect 33241 3349 33275 3383
rect 33275 3349 33284 3383
rect 33232 3340 33284 3349
rect 33508 3383 33560 3392
rect 33508 3349 33517 3383
rect 33517 3349 33551 3383
rect 33551 3349 33560 3383
rect 33508 3340 33560 3349
rect 34520 3340 34572 3392
rect 36452 3340 36504 3392
rect 38476 3340 38528 3392
rect 39488 3383 39540 3392
rect 39488 3349 39497 3383
rect 39497 3349 39531 3383
rect 39531 3349 39540 3383
rect 39488 3340 39540 3349
rect 40132 3383 40184 3392
rect 40132 3349 40141 3383
rect 40141 3349 40175 3383
rect 40175 3349 40184 3383
rect 40132 3340 40184 3349
rect 44640 3476 44692 3528
rect 44824 3451 44876 3460
rect 44824 3417 44833 3451
rect 44833 3417 44867 3451
rect 44867 3417 44876 3451
rect 44824 3408 44876 3417
rect 45100 3451 45152 3460
rect 45100 3417 45109 3451
rect 45109 3417 45143 3451
rect 45143 3417 45152 3451
rect 45100 3408 45152 3417
rect 42800 3340 42852 3392
rect 42984 3383 43036 3392
rect 42984 3349 42993 3383
rect 42993 3349 43027 3383
rect 43027 3349 43036 3383
rect 42984 3340 43036 3349
rect 43996 3383 44048 3392
rect 43996 3349 44005 3383
rect 44005 3349 44039 3383
rect 44039 3349 44048 3383
rect 43996 3340 44048 3349
rect 44272 3340 44324 3392
rect 45468 3476 45520 3528
rect 53380 3553 53389 3587
rect 53389 3553 53423 3587
rect 53423 3553 53432 3587
rect 53380 3544 53432 3553
rect 54668 3612 54720 3664
rect 53748 3544 53800 3596
rect 54576 3544 54628 3596
rect 54944 3587 54996 3596
rect 54944 3553 54953 3587
rect 54953 3553 54987 3587
rect 54987 3553 54996 3587
rect 54944 3544 54996 3553
rect 55036 3587 55088 3596
rect 55036 3553 55045 3587
rect 55045 3553 55079 3587
rect 55079 3553 55088 3587
rect 55036 3544 55088 3553
rect 55312 3544 55364 3596
rect 55680 3655 55732 3664
rect 55680 3621 55689 3655
rect 55689 3621 55723 3655
rect 55723 3621 55732 3655
rect 56232 3689 56241 3723
rect 56241 3689 56275 3723
rect 56275 3689 56284 3723
rect 56232 3680 56284 3689
rect 59912 3680 59964 3732
rect 57336 3655 57388 3664
rect 55680 3612 55732 3621
rect 57336 3621 57345 3655
rect 57345 3621 57379 3655
rect 57379 3621 57388 3655
rect 57336 3612 57388 3621
rect 60464 3612 60516 3664
rect 56508 3587 56560 3596
rect 56508 3553 56517 3587
rect 56517 3553 56551 3587
rect 56551 3553 56560 3587
rect 56508 3544 56560 3553
rect 57244 3544 57296 3596
rect 58348 3587 58400 3596
rect 58348 3553 58357 3587
rect 58357 3553 58391 3587
rect 58391 3553 58400 3587
rect 58348 3544 58400 3553
rect 58532 3587 58584 3596
rect 58532 3553 58541 3587
rect 58541 3553 58575 3587
rect 58575 3553 58584 3587
rect 58532 3544 58584 3553
rect 58716 3544 58768 3596
rect 59452 3544 59504 3596
rect 59636 3544 59688 3596
rect 60280 3544 60332 3596
rect 46388 3408 46440 3460
rect 46848 3408 46900 3460
rect 50252 3408 50304 3460
rect 50620 3408 50672 3460
rect 51172 3408 51224 3460
rect 52092 3408 52144 3460
rect 57060 3476 57112 3528
rect 57980 3476 58032 3528
rect 59360 3476 59412 3528
rect 59820 3476 59872 3528
rect 62304 3476 62356 3528
rect 53840 3451 53892 3460
rect 53840 3417 53849 3451
rect 53849 3417 53883 3451
rect 53883 3417 53892 3451
rect 53840 3408 53892 3417
rect 53932 3408 53984 3460
rect 61292 3408 61344 3460
rect 47308 3340 47360 3392
rect 48688 3340 48740 3392
rect 49332 3340 49384 3392
rect 51540 3383 51592 3392
rect 51540 3349 51549 3383
rect 51549 3349 51583 3383
rect 51583 3349 51592 3383
rect 51540 3340 51592 3349
rect 51816 3340 51868 3392
rect 52460 3340 52512 3392
rect 52644 3340 52696 3392
rect 53288 3340 53340 3392
rect 58532 3340 58584 3392
rect 59820 3340 59872 3392
rect 60556 3340 60608 3392
rect 62212 3340 62264 3392
rect 11378 3238 11430 3290
rect 11442 3238 11494 3290
rect 11506 3238 11558 3290
rect 11570 3238 11622 3290
rect 32170 3238 32222 3290
rect 32234 3238 32286 3290
rect 32298 3238 32350 3290
rect 32362 3238 32414 3290
rect 52962 3238 53014 3290
rect 53026 3238 53078 3290
rect 53090 3238 53142 3290
rect 53154 3238 53206 3290
rect 2780 3136 2832 3188
rect 2872 3136 2924 3188
rect 3884 3136 3936 3188
rect 5908 3179 5960 3188
rect 5908 3145 5917 3179
rect 5917 3145 5951 3179
rect 5951 3145 5960 3179
rect 5908 3136 5960 3145
rect 6644 3136 6696 3188
rect 7748 3136 7800 3188
rect 11244 3136 11296 3188
rect 12532 3136 12584 3188
rect 14464 3179 14516 3188
rect 14464 3145 14473 3179
rect 14473 3145 14507 3179
rect 14507 3145 14516 3179
rect 14464 3136 14516 3145
rect 15660 3136 15712 3188
rect 17776 3179 17828 3188
rect 3608 3068 3660 3120
rect 6828 3068 6880 3120
rect 13268 3068 13320 3120
rect 2320 2975 2372 2984
rect 2320 2941 2329 2975
rect 2329 2941 2363 2975
rect 2363 2941 2372 2975
rect 2320 2932 2372 2941
rect 5356 3000 5408 3052
rect 7196 3000 7248 3052
rect 7748 3000 7800 3052
rect 7932 3043 7984 3052
rect 7932 3009 7941 3043
rect 7941 3009 7975 3043
rect 7975 3009 7984 3043
rect 7932 3000 7984 3009
rect 8392 3000 8444 3052
rect 9312 3000 9364 3052
rect 9588 3000 9640 3052
rect 10416 3043 10468 3052
rect 5908 2932 5960 2984
rect 7656 2932 7708 2984
rect 7840 2975 7892 2984
rect 7840 2941 7849 2975
rect 7849 2941 7883 2975
rect 7883 2941 7892 2975
rect 7840 2932 7892 2941
rect 9036 2932 9088 2984
rect 9772 2932 9824 2984
rect 10416 3009 10425 3043
rect 10425 3009 10459 3043
rect 10459 3009 10468 3043
rect 10416 3000 10468 3009
rect 12348 3000 12400 3052
rect 12808 3000 12860 3052
rect 13820 3068 13872 3120
rect 16212 3068 16264 3120
rect 17776 3145 17785 3179
rect 17785 3145 17819 3179
rect 17819 3145 17828 3179
rect 17776 3136 17828 3145
rect 18052 3179 18104 3188
rect 18052 3145 18061 3179
rect 18061 3145 18095 3179
rect 18095 3145 18104 3179
rect 18052 3136 18104 3145
rect 18144 3136 18196 3188
rect 21272 3179 21324 3188
rect 18696 3068 18748 3120
rect 18972 3068 19024 3120
rect 13728 3043 13780 3052
rect 11152 2975 11204 2984
rect 4712 2864 4764 2916
rect 8116 2864 8168 2916
rect 9588 2864 9640 2916
rect 11152 2941 11161 2975
rect 11161 2941 11195 2975
rect 11195 2941 11204 2975
rect 11152 2932 11204 2941
rect 12256 2975 12308 2984
rect 12256 2941 12265 2975
rect 12265 2941 12299 2975
rect 12299 2941 12308 2975
rect 12256 2932 12308 2941
rect 13728 3009 13737 3043
rect 13737 3009 13771 3043
rect 13771 3009 13780 3043
rect 13728 3000 13780 3009
rect 19064 3000 19116 3052
rect 20352 3000 20404 3052
rect 2136 2796 2188 2848
rect 8300 2796 8352 2848
rect 10324 2796 10376 2848
rect 13452 2864 13504 2916
rect 15016 2932 15068 2984
rect 15936 2975 15988 2984
rect 15936 2941 15945 2975
rect 15945 2941 15979 2975
rect 15979 2941 15988 2975
rect 15936 2932 15988 2941
rect 16120 2975 16172 2984
rect 16120 2941 16129 2975
rect 16129 2941 16163 2975
rect 16163 2941 16172 2975
rect 16120 2932 16172 2941
rect 16396 2932 16448 2984
rect 18052 2932 18104 2984
rect 18328 2975 18380 2984
rect 18328 2941 18337 2975
rect 18337 2941 18371 2975
rect 18371 2941 18380 2975
rect 18328 2932 18380 2941
rect 20076 2975 20128 2984
rect 14096 2864 14148 2916
rect 15200 2864 15252 2916
rect 15384 2864 15436 2916
rect 17408 2907 17460 2916
rect 14556 2796 14608 2848
rect 17408 2873 17417 2907
rect 17417 2873 17451 2907
rect 17451 2873 17460 2907
rect 17408 2864 17460 2873
rect 17684 2864 17736 2916
rect 17868 2864 17920 2916
rect 20076 2941 20085 2975
rect 20085 2941 20119 2975
rect 20119 2941 20128 2975
rect 20076 2932 20128 2941
rect 20168 2975 20220 2984
rect 20168 2941 20177 2975
rect 20177 2941 20211 2975
rect 20211 2941 20220 2975
rect 20720 3000 20772 3052
rect 21272 3145 21281 3179
rect 21281 3145 21315 3179
rect 21315 3145 21324 3179
rect 21272 3136 21324 3145
rect 22652 3136 22704 3188
rect 23480 3136 23532 3188
rect 25320 3179 25372 3188
rect 21548 3068 21600 3120
rect 21824 3068 21876 3120
rect 22100 3000 22152 3052
rect 22376 3000 22428 3052
rect 20168 2932 20220 2941
rect 23112 3000 23164 3052
rect 23572 3000 23624 3052
rect 25320 3145 25329 3179
rect 25329 3145 25363 3179
rect 25363 3145 25372 3179
rect 25320 3136 25372 3145
rect 24492 3068 24544 3120
rect 27436 3136 27488 3188
rect 28172 3136 28224 3188
rect 28264 3136 28316 3188
rect 28724 3136 28776 3188
rect 32036 3136 32088 3188
rect 32680 3136 32732 3188
rect 34520 3136 34572 3188
rect 34704 3179 34756 3188
rect 34704 3145 34713 3179
rect 34713 3145 34747 3179
rect 34747 3145 34756 3179
rect 34704 3136 34756 3145
rect 38016 3136 38068 3188
rect 41236 3136 41288 3188
rect 42064 3179 42116 3188
rect 42064 3145 42073 3179
rect 42073 3145 42107 3179
rect 42107 3145 42116 3179
rect 42064 3136 42116 3145
rect 43444 3136 43496 3188
rect 43628 3136 43680 3188
rect 43996 3136 44048 3188
rect 46112 3136 46164 3188
rect 48596 3136 48648 3188
rect 50068 3136 50120 3188
rect 52368 3136 52420 3188
rect 52644 3136 52696 3188
rect 53840 3179 53892 3188
rect 53840 3145 53849 3179
rect 53849 3145 53883 3179
rect 53883 3145 53892 3179
rect 53840 3136 53892 3145
rect 54668 3136 54720 3188
rect 55128 3136 55180 3188
rect 56324 3179 56376 3188
rect 56324 3145 56333 3179
rect 56333 3145 56367 3179
rect 56367 3145 56376 3179
rect 56324 3136 56376 3145
rect 56508 3136 56560 3188
rect 57244 3136 57296 3188
rect 57612 3179 57664 3188
rect 57612 3145 57621 3179
rect 57621 3145 57655 3179
rect 57655 3145 57664 3179
rect 57612 3136 57664 3145
rect 57980 3179 58032 3188
rect 57980 3145 57989 3179
rect 57989 3145 58023 3179
rect 58023 3145 58032 3179
rect 58624 3179 58676 3188
rect 57980 3136 58032 3145
rect 58624 3145 58633 3179
rect 58633 3145 58667 3179
rect 58667 3145 58676 3179
rect 58624 3136 58676 3145
rect 59544 3136 59596 3188
rect 60556 3136 60608 3188
rect 61292 3179 61344 3188
rect 61292 3145 61301 3179
rect 61301 3145 61335 3179
rect 61335 3145 61344 3179
rect 61292 3136 61344 3145
rect 62304 3179 62356 3188
rect 62304 3145 62313 3179
rect 62313 3145 62347 3179
rect 62347 3145 62356 3179
rect 62304 3136 62356 3145
rect 27804 3068 27856 3120
rect 25228 3000 25280 3052
rect 28356 3000 28408 3052
rect 28448 3000 28500 3052
rect 30748 3068 30800 3120
rect 31852 3068 31904 3120
rect 32128 3068 32180 3120
rect 33324 3068 33376 3120
rect 37464 3068 37516 3120
rect 39764 3068 39816 3120
rect 39948 3111 40000 3120
rect 39948 3077 39957 3111
rect 39957 3077 39991 3111
rect 39991 3077 40000 3111
rect 39948 3068 40000 3077
rect 40316 3111 40368 3120
rect 40316 3077 40325 3111
rect 40325 3077 40359 3111
rect 40359 3077 40368 3111
rect 40316 3068 40368 3077
rect 41972 3068 42024 3120
rect 22560 2975 22612 2984
rect 22560 2941 22569 2975
rect 22569 2941 22603 2975
rect 22603 2941 22612 2975
rect 22744 2975 22796 2984
rect 22560 2932 22612 2941
rect 22744 2941 22753 2975
rect 22753 2941 22787 2975
rect 22787 2941 22796 2975
rect 22744 2932 22796 2941
rect 24584 2975 24636 2984
rect 20444 2864 20496 2916
rect 22836 2864 22888 2916
rect 18696 2796 18748 2848
rect 20720 2796 20772 2848
rect 22192 2796 22244 2848
rect 22560 2796 22612 2848
rect 24584 2941 24593 2975
rect 24593 2941 24627 2975
rect 24627 2941 24636 2975
rect 24584 2932 24636 2941
rect 24860 2932 24912 2984
rect 26976 2932 27028 2984
rect 24308 2864 24360 2916
rect 26608 2907 26660 2916
rect 26608 2873 26617 2907
rect 26617 2873 26651 2907
rect 26651 2873 26660 2907
rect 26608 2864 26660 2873
rect 27712 2975 27764 2984
rect 27712 2941 27721 2975
rect 27721 2941 27755 2975
rect 27755 2941 27764 2975
rect 29276 2975 29328 2984
rect 27712 2932 27764 2941
rect 29276 2941 29285 2975
rect 29285 2941 29319 2975
rect 29319 2941 29328 2975
rect 29276 2932 29328 2941
rect 29460 2975 29512 2984
rect 29460 2941 29469 2975
rect 29469 2941 29503 2975
rect 29503 2941 29512 2975
rect 29460 2932 29512 2941
rect 30196 3000 30248 3052
rect 32496 3000 32548 3052
rect 33968 3043 34020 3052
rect 33968 3009 33977 3043
rect 33977 3009 34011 3043
rect 34011 3009 34020 3043
rect 33968 3000 34020 3009
rect 36728 3000 36780 3052
rect 36912 3000 36964 3052
rect 31024 2975 31076 2984
rect 31024 2941 31033 2975
rect 31033 2941 31067 2975
rect 31067 2941 31076 2975
rect 31024 2932 31076 2941
rect 31208 2932 31260 2984
rect 31484 2975 31536 2984
rect 31484 2941 31493 2975
rect 31493 2941 31527 2975
rect 31527 2941 31536 2975
rect 31484 2932 31536 2941
rect 23388 2796 23440 2848
rect 26516 2796 26568 2848
rect 30564 2864 30616 2916
rect 33232 2932 33284 2984
rect 33508 2975 33560 2984
rect 33508 2941 33517 2975
rect 33517 2941 33551 2975
rect 33551 2941 33560 2975
rect 33508 2932 33560 2941
rect 34796 2932 34848 2984
rect 36268 2975 36320 2984
rect 29460 2796 29512 2848
rect 32680 2864 32732 2916
rect 33416 2907 33468 2916
rect 33416 2873 33425 2907
rect 33425 2873 33459 2907
rect 33459 2873 33468 2907
rect 33416 2864 33468 2873
rect 36268 2941 36277 2975
rect 36277 2941 36311 2975
rect 36311 2941 36320 2975
rect 36268 2932 36320 2941
rect 36360 2975 36412 2984
rect 36360 2941 36369 2975
rect 36369 2941 36403 2975
rect 36403 2941 36412 2975
rect 36360 2932 36412 2941
rect 36544 2932 36596 2984
rect 37740 2932 37792 2984
rect 38016 2932 38068 2984
rect 38844 2932 38896 2984
rect 32956 2839 33008 2848
rect 32956 2805 32965 2839
rect 32965 2805 32999 2839
rect 32999 2805 33008 2839
rect 32956 2796 33008 2805
rect 36176 2864 36228 2916
rect 38476 2907 38528 2916
rect 35900 2796 35952 2848
rect 38476 2873 38485 2907
rect 38485 2873 38519 2907
rect 38519 2873 38528 2907
rect 38476 2864 38528 2873
rect 40040 3000 40092 3052
rect 40132 3000 40184 3052
rect 40776 3043 40828 3052
rect 40776 3009 40785 3043
rect 40785 3009 40819 3043
rect 40819 3009 40828 3043
rect 40776 3000 40828 3009
rect 39304 2932 39356 2984
rect 39948 2932 40000 2984
rect 40500 2975 40552 2984
rect 40500 2941 40509 2975
rect 40509 2941 40543 2975
rect 40543 2941 40552 2975
rect 40500 2932 40552 2941
rect 42892 3068 42944 3120
rect 45008 3068 45060 3120
rect 46296 3068 46348 3120
rect 47032 3068 47084 3120
rect 49056 3068 49108 3120
rect 52184 3068 52236 3120
rect 53472 3068 53524 3120
rect 56140 3068 56192 3120
rect 42984 2975 43036 2984
rect 37280 2796 37332 2848
rect 38752 2796 38804 2848
rect 40316 2796 40368 2848
rect 42984 2941 42993 2975
rect 42993 2941 43027 2975
rect 43027 2941 43036 2975
rect 42984 2932 43036 2941
rect 50436 3000 50488 3052
rect 51172 3000 51224 3052
rect 51724 3000 51776 3052
rect 44732 2975 44784 2984
rect 44732 2941 44741 2975
rect 44741 2941 44775 2975
rect 44775 2941 44784 2975
rect 45008 2975 45060 2984
rect 44732 2932 44784 2941
rect 45008 2941 45017 2975
rect 45017 2941 45051 2975
rect 45051 2941 45060 2975
rect 45008 2932 45060 2941
rect 45192 2975 45244 2984
rect 45192 2941 45201 2975
rect 45201 2941 45235 2975
rect 45235 2941 45244 2975
rect 45192 2932 45244 2941
rect 42892 2864 42944 2916
rect 43996 2907 44048 2916
rect 43996 2873 44005 2907
rect 44005 2873 44039 2907
rect 44039 2873 44048 2907
rect 43996 2864 44048 2873
rect 45376 2864 45428 2916
rect 43076 2839 43128 2848
rect 43076 2805 43085 2839
rect 43085 2805 43119 2839
rect 43119 2805 43128 2839
rect 43076 2796 43128 2805
rect 43720 2796 43772 2848
rect 45560 2796 45612 2848
rect 46112 2932 46164 2984
rect 46296 2975 46348 2984
rect 46296 2941 46305 2975
rect 46305 2941 46339 2975
rect 46339 2941 46348 2975
rect 47032 2975 47084 2984
rect 46296 2932 46348 2941
rect 47032 2941 47041 2975
rect 47041 2941 47075 2975
rect 47075 2941 47084 2975
rect 47032 2932 47084 2941
rect 46020 2864 46072 2916
rect 48228 2932 48280 2984
rect 49332 2975 49384 2984
rect 49332 2941 49341 2975
rect 49341 2941 49375 2975
rect 49375 2941 49384 2975
rect 49332 2932 49384 2941
rect 49884 2975 49936 2984
rect 49884 2941 49893 2975
rect 49893 2941 49927 2975
rect 49927 2941 49936 2975
rect 49884 2932 49936 2941
rect 48136 2864 48188 2916
rect 50528 2932 50580 2984
rect 51540 2932 51592 2984
rect 54392 3000 54444 3052
rect 55036 3000 55088 3052
rect 57888 3068 57940 3120
rect 60832 3068 60884 3120
rect 62212 3068 62264 3120
rect 61200 3043 61252 3052
rect 61200 3009 61206 3043
rect 61206 3009 61240 3043
rect 61240 3009 61252 3043
rect 61200 3000 61252 3009
rect 54116 2975 54168 2984
rect 54116 2941 54125 2975
rect 54125 2941 54159 2975
rect 54159 2941 54168 2975
rect 54116 2932 54168 2941
rect 46940 2796 46992 2848
rect 48320 2796 48372 2848
rect 51080 2864 51132 2916
rect 52000 2864 52052 2916
rect 52276 2907 52328 2916
rect 52276 2873 52285 2907
rect 52285 2873 52319 2907
rect 52319 2873 52328 2907
rect 52276 2864 52328 2873
rect 53564 2864 53616 2916
rect 55312 2975 55364 2984
rect 55312 2941 55321 2975
rect 55321 2941 55355 2975
rect 55355 2941 55364 2975
rect 55312 2932 55364 2941
rect 56232 2932 56284 2984
rect 59820 2975 59872 2984
rect 51816 2796 51868 2848
rect 53748 2839 53800 2848
rect 53748 2805 53757 2839
rect 53757 2805 53791 2839
rect 53791 2805 53800 2839
rect 55128 2864 55180 2916
rect 55588 2864 55640 2916
rect 59820 2941 59829 2975
rect 59829 2941 59863 2975
rect 59863 2941 59872 2975
rect 59820 2932 59872 2941
rect 60004 2975 60056 2984
rect 60004 2941 60013 2975
rect 60013 2941 60047 2975
rect 60047 2941 60056 2975
rect 60004 2932 60056 2941
rect 53748 2796 53800 2805
rect 59452 2796 59504 2848
rect 64144 2932 64196 2984
rect 60280 2907 60332 2916
rect 60280 2873 60289 2907
rect 60289 2873 60323 2907
rect 60323 2873 60332 2907
rect 60280 2864 60332 2873
rect 63224 2864 63276 2916
rect 61200 2796 61252 2848
rect 21774 2694 21826 2746
rect 21838 2694 21890 2746
rect 21902 2694 21954 2746
rect 21966 2694 22018 2746
rect 42566 2694 42618 2746
rect 42630 2694 42682 2746
rect 42694 2694 42746 2746
rect 42758 2694 42810 2746
rect 3056 2635 3108 2644
rect 3056 2601 3065 2635
rect 3065 2601 3099 2635
rect 3099 2601 3108 2635
rect 3056 2592 3108 2601
rect 5724 2635 5776 2644
rect 5724 2601 5733 2635
rect 5733 2601 5767 2635
rect 5767 2601 5776 2635
rect 5724 2592 5776 2601
rect 6184 2592 6236 2644
rect 9036 2592 9088 2644
rect 9588 2592 9640 2644
rect 10416 2592 10468 2644
rect 12348 2635 12400 2644
rect 12348 2601 12357 2635
rect 12357 2601 12391 2635
rect 12391 2601 12400 2635
rect 12348 2592 12400 2601
rect 12900 2635 12952 2644
rect 12900 2601 12909 2635
rect 12909 2601 12943 2635
rect 12943 2601 12952 2635
rect 12900 2592 12952 2601
rect 13360 2592 13412 2644
rect 9404 2524 9456 2576
rect 2964 2499 3016 2508
rect 2964 2465 2973 2499
rect 2973 2465 3007 2499
rect 3007 2465 3016 2499
rect 2964 2456 3016 2465
rect 4712 2456 4764 2508
rect 8116 2456 8168 2508
rect 2320 2388 2372 2440
rect 3608 2388 3660 2440
rect 11980 2456 12032 2508
rect 15200 2635 15252 2644
rect 15200 2601 15209 2635
rect 15209 2601 15243 2635
rect 15243 2601 15252 2635
rect 15200 2592 15252 2601
rect 16396 2592 16448 2644
rect 19340 2592 19392 2644
rect 19616 2635 19668 2644
rect 19616 2601 19625 2635
rect 19625 2601 19659 2635
rect 19659 2601 19668 2635
rect 19616 2592 19668 2601
rect 13084 2388 13136 2440
rect 17868 2524 17920 2576
rect 14464 2499 14516 2508
rect 14464 2465 14473 2499
rect 14473 2465 14507 2499
rect 14507 2465 14516 2499
rect 14464 2456 14516 2465
rect 15292 2456 15344 2508
rect 15752 2499 15804 2508
rect 15752 2465 15761 2499
rect 15761 2465 15795 2499
rect 15795 2465 15804 2499
rect 15752 2456 15804 2465
rect 17592 2456 17644 2508
rect 19800 2524 19852 2576
rect 23020 2524 23072 2576
rect 23480 2567 23532 2576
rect 23480 2533 23489 2567
rect 23489 2533 23523 2567
rect 23523 2533 23532 2567
rect 23480 2524 23532 2533
rect 24860 2592 24912 2644
rect 26424 2592 26476 2644
rect 26608 2635 26660 2644
rect 26608 2601 26617 2635
rect 26617 2601 26651 2635
rect 26651 2601 26660 2635
rect 26608 2592 26660 2601
rect 26700 2592 26752 2644
rect 29000 2592 29052 2644
rect 31944 2592 31996 2644
rect 32680 2592 32732 2644
rect 34796 2592 34848 2644
rect 35900 2592 35952 2644
rect 39028 2592 39080 2644
rect 2136 2295 2188 2304
rect 2136 2261 2145 2295
rect 2145 2261 2179 2295
rect 2179 2261 2188 2295
rect 2136 2252 2188 2261
rect 7840 2252 7892 2304
rect 15384 2320 15436 2372
rect 17684 2252 17736 2304
rect 19248 2388 19300 2440
rect 19984 2456 20036 2508
rect 21548 2456 21600 2508
rect 24308 2499 24360 2508
rect 24308 2465 24317 2499
rect 24317 2465 24351 2499
rect 24351 2465 24360 2499
rect 24308 2456 24360 2465
rect 25044 2456 25096 2508
rect 28080 2524 28132 2576
rect 30748 2499 30800 2508
rect 30748 2465 30757 2499
rect 30757 2465 30791 2499
rect 30791 2465 30800 2499
rect 30748 2456 30800 2465
rect 31116 2499 31168 2508
rect 31116 2465 31125 2499
rect 31125 2465 31159 2499
rect 31159 2465 31168 2499
rect 31116 2456 31168 2465
rect 33692 2456 33744 2508
rect 37004 2524 37056 2576
rect 36084 2456 36136 2508
rect 36636 2499 36688 2508
rect 36636 2465 36645 2499
rect 36645 2465 36679 2499
rect 36679 2465 36688 2499
rect 36636 2456 36688 2465
rect 37280 2456 37332 2508
rect 40776 2635 40828 2644
rect 40776 2601 40785 2635
rect 40785 2601 40819 2635
rect 40819 2601 40828 2635
rect 40776 2592 40828 2601
rect 41420 2592 41472 2644
rect 39212 2524 39264 2576
rect 40592 2524 40644 2576
rect 41052 2524 41104 2576
rect 39764 2499 39816 2508
rect 21456 2431 21508 2440
rect 21456 2397 21465 2431
rect 21465 2397 21499 2431
rect 21499 2397 21508 2431
rect 21456 2388 21508 2397
rect 22376 2388 22428 2440
rect 18052 2320 18104 2372
rect 18880 2320 18932 2372
rect 24124 2320 24176 2372
rect 31208 2388 31260 2440
rect 25872 2320 25924 2372
rect 32956 2388 33008 2440
rect 39764 2465 39773 2499
rect 39773 2465 39807 2499
rect 39807 2465 39816 2499
rect 39764 2456 39816 2465
rect 40408 2456 40460 2508
rect 38660 2388 38712 2440
rect 39028 2431 39080 2440
rect 39028 2397 39037 2431
rect 39037 2397 39071 2431
rect 39071 2397 39080 2431
rect 39028 2388 39080 2397
rect 41972 2388 42024 2440
rect 43076 2320 43128 2372
rect 22744 2252 22796 2304
rect 22836 2252 22888 2304
rect 24768 2252 24820 2304
rect 32588 2252 32640 2304
rect 34428 2252 34480 2304
rect 37280 2252 37332 2304
rect 38476 2252 38528 2304
rect 42156 2252 42208 2304
rect 42432 2295 42484 2304
rect 42432 2261 42441 2295
rect 42441 2261 42475 2295
rect 42475 2261 42484 2295
rect 42432 2252 42484 2261
rect 43996 2592 44048 2644
rect 46204 2635 46256 2644
rect 46204 2601 46213 2635
rect 46213 2601 46247 2635
rect 46247 2601 46256 2635
rect 46204 2592 46256 2601
rect 46940 2592 46992 2644
rect 48136 2592 48188 2644
rect 49884 2635 49936 2644
rect 49884 2601 49893 2635
rect 49893 2601 49927 2635
rect 49927 2601 49936 2635
rect 49884 2592 49936 2601
rect 51908 2635 51960 2644
rect 51908 2601 51917 2635
rect 51917 2601 51951 2635
rect 51951 2601 51960 2635
rect 51908 2592 51960 2601
rect 52000 2592 52052 2644
rect 54668 2635 54720 2644
rect 54668 2601 54677 2635
rect 54677 2601 54711 2635
rect 54711 2601 54720 2635
rect 54668 2592 54720 2601
rect 54944 2635 54996 2644
rect 54944 2601 54953 2635
rect 54953 2601 54987 2635
rect 54987 2601 54996 2635
rect 54944 2592 54996 2601
rect 57244 2592 57296 2644
rect 58532 2635 58584 2644
rect 58532 2601 58541 2635
rect 58541 2601 58575 2635
rect 58575 2601 58584 2635
rect 58532 2592 58584 2601
rect 62212 2635 62264 2644
rect 62212 2601 62221 2635
rect 62221 2601 62255 2635
rect 62255 2601 62264 2635
rect 62212 2592 62264 2601
rect 47584 2524 47636 2576
rect 49792 2524 49844 2576
rect 50528 2524 50580 2576
rect 51264 2524 51316 2576
rect 53472 2524 53524 2576
rect 59452 2567 59504 2576
rect 59452 2533 59461 2567
rect 59461 2533 59495 2567
rect 59495 2533 59504 2567
rect 59452 2524 59504 2533
rect 44272 2431 44324 2440
rect 44272 2397 44281 2431
rect 44281 2397 44315 2431
rect 44315 2397 44324 2431
rect 44272 2388 44324 2397
rect 49056 2456 49108 2508
rect 51080 2456 51132 2508
rect 53748 2456 53800 2508
rect 48320 2388 48372 2440
rect 49332 2388 49384 2440
rect 47308 2320 47360 2372
rect 48228 2295 48280 2304
rect 48228 2261 48252 2295
rect 48252 2261 48280 2295
rect 48228 2252 48280 2261
rect 49884 2320 49936 2372
rect 50804 2388 50856 2440
rect 58072 2388 58124 2440
rect 58808 2388 58860 2440
rect 61476 2456 61528 2508
rect 62396 2456 62448 2508
rect 51540 2295 51592 2304
rect 51540 2261 51549 2295
rect 51549 2261 51583 2295
rect 51583 2261 51592 2295
rect 51540 2252 51592 2261
rect 53472 2295 53524 2304
rect 53472 2261 53481 2295
rect 53481 2261 53515 2295
rect 53515 2261 53524 2295
rect 53472 2252 53524 2261
rect 55956 2295 56008 2304
rect 55956 2261 55965 2295
rect 55965 2261 55999 2295
rect 55999 2261 56008 2295
rect 55956 2252 56008 2261
rect 59728 2295 59780 2304
rect 59728 2261 59737 2295
rect 59737 2261 59771 2295
rect 59771 2261 59780 2295
rect 59728 2252 59780 2261
rect 59912 2295 59964 2304
rect 59912 2261 59921 2295
rect 59921 2261 59955 2295
rect 59955 2261 59964 2295
rect 59912 2252 59964 2261
rect 61476 2252 61528 2304
rect 62396 2252 62448 2304
rect 11378 2150 11430 2202
rect 11442 2150 11494 2202
rect 11506 2150 11558 2202
rect 11570 2150 11622 2202
rect 32170 2150 32222 2202
rect 32234 2150 32286 2202
rect 32298 2150 32350 2202
rect 32362 2150 32414 2202
rect 52962 2150 53014 2202
rect 53026 2150 53078 2202
rect 53090 2150 53142 2202
rect 53154 2150 53206 2202
rect 2136 2048 2188 2100
rect 15200 2048 15252 2100
rect 15752 2048 15804 2100
rect 42156 2048 42208 2100
rect 42708 2048 42760 2100
rect 48228 2048 48280 2100
rect 49976 2048 50028 2100
rect 51540 2048 51592 2100
rect 59912 2048 59964 2100
rect 9220 1980 9272 2032
rect 19984 1980 20036 2032
rect 42432 1980 42484 2032
rect 49332 1980 49384 2032
rect 15292 1912 15344 1964
rect 40500 1912 40552 1964
rect 44272 1912 44324 1964
rect 55956 1912 56008 1964
rect 16304 1844 16356 1896
rect 17592 1844 17644 1896
rect 21456 1776 21508 1828
rect 1216 1368 1268 1420
rect 7288 1368 7340 1420
rect 32220 1368 32272 1420
rect 36912 1368 36964 1420
rect 4068 1300 4120 1352
rect 24952 1300 25004 1352
rect 30472 1300 30524 1352
rect 32772 1300 32824 1352
<< metal2 >>
rect 938 19162 994 19962
rect 2870 19162 2926 19962
rect 4802 19162 4858 19962
rect 6734 19162 6790 19962
rect 8758 19162 8814 19962
rect 10690 19162 10746 19962
rect 12622 19162 12678 19962
rect 14646 19162 14702 19962
rect 16578 19162 16634 19962
rect 18510 19162 18566 19962
rect 20534 19162 20590 19962
rect 22466 19162 22522 19962
rect 24398 19162 24454 19962
rect 26330 19162 26386 19962
rect 28354 19162 28410 19962
rect 30286 19162 30342 19962
rect 32218 19162 32274 19962
rect 34242 19162 34298 19962
rect 36174 19162 36230 19962
rect 38106 19162 38162 19962
rect 40130 19162 40186 19962
rect 42062 19162 42118 19962
rect 43994 19162 44050 19962
rect 45926 19162 45982 19962
rect 47950 19162 48006 19962
rect 49882 19162 49938 19962
rect 51814 19162 51870 19962
rect 53838 19162 53894 19962
rect 55770 19162 55826 19962
rect 57702 19162 57758 19962
rect 59726 19162 59782 19962
rect 61658 19162 61714 19962
rect 63590 19162 63646 19962
rect 952 15910 980 19162
rect 940 15904 992 15910
rect 940 15846 992 15852
rect 2884 15094 2912 19162
rect 3974 18864 4030 18873
rect 3974 18799 4030 18808
rect 3608 15904 3660 15910
rect 3608 15846 3660 15852
rect 2872 15088 2924 15094
rect 2872 15030 2924 15036
rect 3146 14512 3202 14521
rect 3146 14447 3202 14456
rect 3160 14006 3188 14447
rect 3148 14000 3200 14006
rect 3148 13942 3200 13948
rect 2412 13184 2464 13190
rect 2412 13126 2464 13132
rect 2424 12782 2452 13126
rect 2412 12776 2464 12782
rect 2412 12718 2464 12724
rect 2688 12300 2740 12306
rect 2688 12242 2740 12248
rect 2700 12186 2728 12242
rect 3332 12232 3384 12238
rect 2700 12158 2820 12186
rect 3332 12174 3384 12180
rect 2792 11778 2820 12158
rect 2872 12164 2924 12170
rect 2872 12106 2924 12112
rect 2884 11898 2912 12106
rect 2872 11892 2924 11898
rect 2872 11834 2924 11840
rect 2792 11750 2912 11778
rect 3344 11762 3372 12174
rect 2884 11558 2912 11750
rect 3332 11756 3384 11762
rect 3332 11698 3384 11704
rect 2872 11552 2924 11558
rect 2872 11494 2924 11500
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 2884 11218 2912 11494
rect 2872 11212 2924 11218
rect 2872 11154 2924 11160
rect 2884 9042 2912 11154
rect 2976 9654 3004 11494
rect 2964 9648 3016 9654
rect 2964 9590 3016 9596
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 3068 9042 3096 9318
rect 2596 9036 2648 9042
rect 2596 8978 2648 8984
rect 2872 9036 2924 9042
rect 2872 8978 2924 8984
rect 3056 9036 3108 9042
rect 3056 8978 3108 8984
rect 2608 8498 2636 8978
rect 2884 8566 2912 8978
rect 3068 8634 3096 8978
rect 3056 8628 3108 8634
rect 3056 8570 3108 8576
rect 2872 8560 2924 8566
rect 2872 8502 2924 8508
rect 2596 8492 2648 8498
rect 2596 8434 2648 8440
rect 3240 6656 3292 6662
rect 3240 6598 3292 6604
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3252 6254 3280 6598
rect 3528 6322 3556 6598
rect 3516 6316 3568 6322
rect 3516 6258 3568 6264
rect 3240 6248 3292 6254
rect 3240 6190 3292 6196
rect 2320 6112 2372 6118
rect 2320 6054 2372 6060
rect 2332 5574 2360 6054
rect 3528 5846 3556 6258
rect 3516 5840 3568 5846
rect 3516 5782 3568 5788
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 2596 5704 2648 5710
rect 2596 5646 2648 5652
rect 2320 5568 2372 5574
rect 2320 5510 2372 5516
rect 2332 5166 2360 5510
rect 2320 5160 2372 5166
rect 2320 5102 2372 5108
rect 2228 3664 2280 3670
rect 2228 3606 2280 3612
rect 386 3088 442 3097
rect 386 3023 442 3032
rect 400 800 428 3023
rect 2136 2848 2188 2854
rect 2136 2790 2188 2796
rect 2148 2310 2176 2790
rect 2136 2304 2188 2310
rect 2136 2246 2188 2252
rect 2148 2106 2176 2246
rect 2136 2100 2188 2106
rect 2136 2042 2188 2048
rect 1216 1420 1268 1426
rect 1216 1362 1268 1368
rect 1228 800 1256 1362
rect 2240 898 2268 3606
rect 2332 2990 2360 5102
rect 2608 5030 2636 5646
rect 2700 5370 2728 5714
rect 3516 5568 3568 5574
rect 3516 5510 3568 5516
rect 2688 5364 2740 5370
rect 2688 5306 2740 5312
rect 3528 5166 3556 5510
rect 3516 5160 3568 5166
rect 3516 5102 3568 5108
rect 2596 5024 2648 5030
rect 2596 4966 2648 4972
rect 2778 4992 2834 5001
rect 2778 4927 2834 4936
rect 2504 4752 2556 4758
rect 2504 4694 2556 4700
rect 2516 4282 2544 4694
rect 2504 4276 2556 4282
rect 2504 4218 2556 4224
rect 2792 3534 2820 4927
rect 2872 4684 2924 4690
rect 2872 4626 2924 4632
rect 2884 3942 2912 4626
rect 3516 4480 3568 4486
rect 3516 4422 3568 4428
rect 3528 4078 3556 4422
rect 3620 4282 3648 15846
rect 3988 13297 4016 18799
rect 4066 16688 4122 16697
rect 4066 16623 4122 16632
rect 4080 15026 4108 16623
rect 4816 16454 4844 19162
rect 4804 16448 4856 16454
rect 4804 16390 4856 16396
rect 6748 15706 6776 19162
rect 8116 16652 8168 16658
rect 8116 16594 8168 16600
rect 7932 16584 7984 16590
rect 7932 16526 7984 16532
rect 7944 15910 7972 16526
rect 8128 16250 8156 16594
rect 8208 16516 8260 16522
rect 8208 16458 8260 16464
rect 8116 16244 8168 16250
rect 8116 16186 8168 16192
rect 7288 15904 7340 15910
rect 7288 15846 7340 15852
rect 7932 15904 7984 15910
rect 7932 15846 7984 15852
rect 6736 15700 6788 15706
rect 6736 15642 6788 15648
rect 7300 15502 7328 15846
rect 7840 15700 7892 15706
rect 7840 15642 7892 15648
rect 5356 15496 5408 15502
rect 5356 15438 5408 15444
rect 5632 15496 5684 15502
rect 5632 15438 5684 15444
rect 7288 15496 7340 15502
rect 7288 15438 7340 15444
rect 5368 15162 5396 15438
rect 5644 15162 5672 15438
rect 7196 15428 7248 15434
rect 7196 15370 7248 15376
rect 7208 15162 7236 15370
rect 5356 15156 5408 15162
rect 5356 15098 5408 15104
rect 5632 15156 5684 15162
rect 5632 15098 5684 15104
rect 6276 15156 6328 15162
rect 6276 15098 6328 15104
rect 7196 15156 7248 15162
rect 7196 15098 7248 15104
rect 5368 15042 5396 15098
rect 4068 15020 4120 15026
rect 5368 15014 5488 15042
rect 4068 14962 4120 14968
rect 5356 14952 5408 14958
rect 5356 14894 5408 14900
rect 4896 14612 4948 14618
rect 4896 14554 4948 14560
rect 4908 14074 4936 14554
rect 5368 14346 5396 14894
rect 5460 14822 5488 15014
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 5448 14816 5500 14822
rect 5448 14758 5500 14764
rect 5356 14340 5408 14346
rect 5356 14282 5408 14288
rect 4896 14068 4948 14074
rect 4896 14010 4948 14016
rect 4908 13938 4936 14010
rect 4896 13932 4948 13938
rect 4896 13874 4948 13880
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 4528 13864 4580 13870
rect 4528 13806 4580 13812
rect 3974 13288 4030 13297
rect 3974 13223 4030 13232
rect 3884 13184 3936 13190
rect 3884 13126 3936 13132
rect 3896 12850 3924 13126
rect 3884 12844 3936 12850
rect 3884 12786 3936 12792
rect 4172 12646 4200 13806
rect 4540 13530 4568 13806
rect 4712 13796 4764 13802
rect 4712 13738 4764 13744
rect 4528 13524 4580 13530
rect 4528 13466 4580 13472
rect 4724 13190 4752 13738
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 4988 13388 5040 13394
rect 4988 13330 5040 13336
rect 4712 13184 4764 13190
rect 4712 13126 4764 13132
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 4080 12209 4108 12378
rect 4066 12200 4122 12209
rect 4066 12135 4122 12144
rect 4724 11898 4752 13126
rect 5000 12782 5028 13330
rect 5172 13184 5224 13190
rect 5172 13126 5224 13132
rect 5184 12782 5212 13126
rect 5460 12782 5488 13466
rect 5552 13462 5580 14894
rect 5908 14884 5960 14890
rect 5908 14826 5960 14832
rect 5724 14272 5776 14278
rect 5724 14214 5776 14220
rect 5632 13932 5684 13938
rect 5632 13874 5684 13880
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 4988 12776 5040 12782
rect 4988 12718 5040 12724
rect 5172 12776 5224 12782
rect 5172 12718 5224 12724
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 5264 12708 5316 12714
rect 5264 12650 5316 12656
rect 5356 12708 5408 12714
rect 5356 12650 5408 12656
rect 5080 12300 5132 12306
rect 5080 12242 5132 12248
rect 4712 11892 4764 11898
rect 4712 11834 4764 11840
rect 4252 11688 4304 11694
rect 4252 11630 4304 11636
rect 4264 11014 4292 11630
rect 5092 11558 5120 12242
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 3974 10704 4030 10713
rect 3974 10639 4030 10648
rect 3882 10024 3938 10033
rect 3882 9959 3938 9968
rect 3896 7857 3924 9959
rect 3882 7848 3938 7857
rect 3882 7783 3938 7792
rect 3700 7200 3752 7206
rect 3700 7142 3752 7148
rect 3712 6798 3740 7142
rect 3700 6792 3752 6798
rect 3700 6734 3752 6740
rect 3792 5568 3844 5574
rect 3792 5510 3844 5516
rect 3608 4276 3660 4282
rect 3608 4218 3660 4224
rect 3056 4072 3108 4078
rect 3056 4014 3108 4020
rect 3516 4072 3568 4078
rect 3516 4014 3568 4020
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2884 3602 2912 3878
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2792 3194 2820 3470
rect 2884 3194 2912 3538
rect 2780 3188 2832 3194
rect 2780 3130 2832 3136
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 2320 2984 2372 2990
rect 2320 2926 2372 2932
rect 2332 2446 2360 2926
rect 3068 2650 3096 4014
rect 3620 4010 3648 4218
rect 3700 4140 3752 4146
rect 3700 4082 3752 4088
rect 3332 4004 3384 4010
rect 3332 3946 3384 3952
rect 3608 4004 3660 4010
rect 3608 3946 3660 3952
rect 3344 3738 3372 3946
rect 3422 3768 3478 3777
rect 3332 3732 3384 3738
rect 3422 3703 3478 3712
rect 3332 3674 3384 3680
rect 3436 3602 3464 3703
rect 3424 3596 3476 3602
rect 3424 3538 3476 3544
rect 3608 3120 3660 3126
rect 3608 3062 3660 3068
rect 3056 2644 3108 2650
rect 3056 2586 3108 2592
rect 2964 2508 3016 2514
rect 2964 2450 3016 2456
rect 2320 2440 2372 2446
rect 2320 2382 2372 2388
rect 2148 870 2268 898
rect 2148 800 2176 870
rect 2976 800 3004 2450
rect 3620 2446 3648 3062
rect 3712 2825 3740 4082
rect 3804 3602 3832 5510
rect 3792 3596 3844 3602
rect 3792 3538 3844 3544
rect 3804 3176 3832 3538
rect 3884 3188 3936 3194
rect 3804 3148 3884 3176
rect 3884 3130 3936 3136
rect 3698 2816 3754 2825
rect 3988 2802 4016 10639
rect 4264 10606 4292 10950
rect 4252 10600 4304 10606
rect 4252 10542 4304 10548
rect 4264 10130 4292 10542
rect 4252 10124 4304 10130
rect 4252 10066 4304 10072
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 4172 9518 4200 9862
rect 4264 9586 4292 10066
rect 4252 9580 4304 9586
rect 4252 9522 4304 9528
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 4172 8906 4200 9454
rect 4344 8968 4396 8974
rect 4344 8910 4396 8916
rect 4160 8900 4212 8906
rect 4160 8842 4212 8848
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 4080 8430 4108 8774
rect 4068 8424 4120 8430
rect 4068 8366 4120 8372
rect 4080 7886 4108 8366
rect 4356 7954 4384 8910
rect 4344 7948 4396 7954
rect 4344 7890 4396 7896
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 4080 7206 4108 7822
rect 4356 7546 4384 7890
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 4068 7200 4120 7206
rect 4068 7142 4120 7148
rect 4632 5778 4660 11494
rect 4988 11144 5040 11150
rect 4988 11086 5040 11092
rect 5000 10470 5028 11086
rect 5276 10810 5304 12650
rect 5368 12374 5396 12650
rect 5356 12368 5408 12374
rect 5356 12310 5408 12316
rect 5448 12300 5500 12306
rect 5448 12242 5500 12248
rect 5460 11898 5488 12242
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5448 11892 5500 11898
rect 5448 11834 5500 11840
rect 5552 11558 5580 12174
rect 5540 11552 5592 11558
rect 5540 11494 5592 11500
rect 5644 11354 5672 13874
rect 5736 13734 5764 14214
rect 5724 13728 5776 13734
rect 5724 13670 5776 13676
rect 5736 13002 5764 13670
rect 5736 12974 5856 13002
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5632 11348 5684 11354
rect 5632 11290 5684 11296
rect 5356 11144 5408 11150
rect 5356 11086 5408 11092
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 4988 10464 5040 10470
rect 4988 10406 5040 10412
rect 5000 10130 5028 10406
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 4988 10124 5040 10130
rect 4988 10066 5040 10072
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4724 9110 4752 9998
rect 4816 9722 4844 10066
rect 4804 9716 4856 9722
rect 4804 9658 4856 9664
rect 4712 9104 4764 9110
rect 4712 9046 4764 9052
rect 4816 8838 4844 9658
rect 5368 9654 5396 11086
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5460 10266 5488 10746
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5736 10062 5764 12786
rect 5828 12646 5856 12974
rect 5816 12640 5868 12646
rect 5816 12582 5868 12588
rect 5920 12442 5948 14826
rect 6000 14476 6052 14482
rect 6000 14418 6052 14424
rect 6012 14074 6040 14418
rect 6288 14278 6316 15098
rect 7300 14958 7328 15438
rect 7472 15428 7524 15434
rect 7472 15370 7524 15376
rect 7288 14952 7340 14958
rect 7116 14912 7288 14940
rect 7116 14822 7144 14912
rect 7288 14894 7340 14900
rect 7104 14816 7156 14822
rect 7104 14758 7156 14764
rect 7484 14550 7512 15370
rect 7656 15360 7708 15366
rect 7656 15302 7708 15308
rect 7668 14958 7696 15302
rect 7748 15020 7800 15026
rect 7748 14962 7800 14968
rect 7656 14952 7708 14958
rect 7656 14894 7708 14900
rect 7472 14544 7524 14550
rect 7472 14486 7524 14492
rect 6276 14272 6328 14278
rect 6276 14214 6328 14220
rect 7104 14272 7156 14278
rect 7104 14214 7156 14220
rect 6000 14068 6052 14074
rect 6000 14010 6052 14016
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 5908 12436 5960 12442
rect 5908 12378 5960 12384
rect 6564 12306 6592 13262
rect 6932 13258 6960 13806
rect 7012 13388 7064 13394
rect 7012 13330 7064 13336
rect 6920 13252 6972 13258
rect 6920 13194 6972 13200
rect 6932 12782 6960 13194
rect 6920 12776 6972 12782
rect 6920 12718 6972 12724
rect 7024 12442 7052 13330
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 6552 12300 6604 12306
rect 6552 12242 6604 12248
rect 6564 11898 6592 12242
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 6552 11892 6604 11898
rect 6552 11834 6604 11840
rect 6932 11626 6960 12038
rect 6920 11620 6972 11626
rect 6920 11562 6972 11568
rect 7012 11552 7064 11558
rect 7012 11494 7064 11500
rect 7024 11234 7052 11494
rect 7116 11354 7144 14214
rect 7484 14074 7512 14486
rect 7472 14068 7524 14074
rect 7472 14010 7524 14016
rect 7760 13870 7788 14962
rect 7852 14482 7880 15642
rect 7944 14550 7972 15846
rect 8220 15638 8248 16458
rect 8208 15632 8260 15638
rect 8208 15574 8260 15580
rect 8300 15564 8352 15570
rect 8300 15506 8352 15512
rect 8024 14952 8076 14958
rect 8024 14894 8076 14900
rect 7932 14544 7984 14550
rect 7932 14486 7984 14492
rect 7840 14476 7892 14482
rect 7840 14418 7892 14424
rect 8036 14074 8064 14894
rect 8312 14890 8340 15506
rect 8772 15094 8800 19162
rect 9496 16652 9548 16658
rect 9496 16594 9548 16600
rect 9508 16454 9536 16594
rect 9036 16448 9088 16454
rect 9036 16390 9088 16396
rect 9496 16448 9548 16454
rect 9496 16390 9548 16396
rect 9048 16114 9076 16390
rect 9036 16108 9088 16114
rect 9036 16050 9088 16056
rect 9048 15638 9076 16050
rect 9036 15632 9088 15638
rect 9036 15574 9088 15580
rect 9508 15366 9536 16390
rect 10704 16250 10732 19162
rect 11352 17436 11648 17456
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11430 17382 11432 17434
rect 11494 17382 11506 17434
rect 11568 17382 11570 17434
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11352 17360 11648 17380
rect 12256 17196 12308 17202
rect 12256 17138 12308 17144
rect 12268 16658 12296 17138
rect 12636 16794 12664 19162
rect 14660 17338 14688 19162
rect 14648 17332 14700 17338
rect 14648 17274 14700 17280
rect 13912 17128 13964 17134
rect 13912 17070 13964 17076
rect 12624 16788 12676 16794
rect 12624 16730 12676 16736
rect 12256 16652 12308 16658
rect 12256 16594 12308 16600
rect 11244 16584 11296 16590
rect 11244 16526 11296 16532
rect 10876 16448 10928 16454
rect 10876 16390 10928 16396
rect 10692 16244 10744 16250
rect 10692 16186 10744 16192
rect 10888 16046 10916 16390
rect 11256 16250 11284 16526
rect 11980 16448 12032 16454
rect 11980 16390 12032 16396
rect 11352 16348 11648 16368
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11430 16294 11432 16346
rect 11494 16294 11506 16346
rect 11568 16294 11570 16346
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11352 16272 11648 16292
rect 11244 16244 11296 16250
rect 11244 16186 11296 16192
rect 10876 16040 10928 16046
rect 10876 15982 10928 15988
rect 10888 15706 10916 15982
rect 11152 15972 11204 15978
rect 11152 15914 11204 15920
rect 10876 15700 10928 15706
rect 10876 15642 10928 15648
rect 10888 15434 10916 15642
rect 10876 15428 10928 15434
rect 10876 15370 10928 15376
rect 8944 15360 8996 15366
rect 8944 15302 8996 15308
rect 9496 15360 9548 15366
rect 9496 15302 9548 15308
rect 10508 15360 10560 15366
rect 10508 15302 10560 15308
rect 8760 15088 8812 15094
rect 8760 15030 8812 15036
rect 8300 14884 8352 14890
rect 8300 14826 8352 14832
rect 8116 14476 8168 14482
rect 8116 14418 8168 14424
rect 8128 14074 8156 14418
rect 8024 14068 8076 14074
rect 8024 14010 8076 14016
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 7748 13864 7800 13870
rect 7748 13806 7800 13812
rect 8024 13864 8076 13870
rect 8024 13806 8076 13812
rect 7760 13530 7788 13806
rect 7748 13524 7800 13530
rect 7748 13466 7800 13472
rect 7288 13388 7340 13394
rect 7288 13330 7340 13336
rect 7300 12782 7328 13330
rect 7380 13320 7432 13326
rect 7380 13262 7432 13268
rect 7392 12850 7420 13262
rect 8036 13190 8064 13806
rect 8116 13524 8168 13530
rect 8116 13466 8168 13472
rect 8024 13184 8076 13190
rect 8024 13126 8076 13132
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 7288 12776 7340 12782
rect 7288 12718 7340 12724
rect 7564 12436 7616 12442
rect 7564 12378 7616 12384
rect 7576 12238 7604 12378
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7564 12096 7616 12102
rect 7564 12038 7616 12044
rect 7576 11830 7604 12038
rect 8036 11898 8064 13126
rect 8128 12782 8156 13466
rect 8116 12776 8168 12782
rect 8116 12718 8168 12724
rect 8312 12374 8340 14826
rect 8956 14414 8984 15302
rect 10520 14958 10548 15302
rect 11164 14958 11192 15914
rect 11244 15496 11296 15502
rect 11244 15438 11296 15444
rect 10416 14952 10468 14958
rect 10416 14894 10468 14900
rect 10508 14952 10560 14958
rect 10508 14894 10560 14900
rect 11152 14952 11204 14958
rect 11152 14894 11204 14900
rect 10428 14482 10456 14894
rect 11256 14822 11284 15438
rect 11992 15366 12020 16390
rect 12268 16250 12296 16594
rect 12256 16244 12308 16250
rect 12176 16204 12256 16232
rect 12176 15570 12204 16204
rect 12256 16186 12308 16192
rect 12256 16040 12308 16046
rect 12256 15982 12308 15988
rect 12164 15564 12216 15570
rect 12164 15506 12216 15512
rect 11980 15360 12032 15366
rect 11980 15302 12032 15308
rect 11352 15260 11648 15280
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11430 15206 11432 15258
rect 11494 15206 11506 15258
rect 11568 15206 11570 15258
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11352 15184 11648 15204
rect 11520 14884 11572 14890
rect 11520 14826 11572 14832
rect 11244 14816 11296 14822
rect 11244 14758 11296 14764
rect 10784 14612 10836 14618
rect 10784 14554 10836 14560
rect 9680 14476 9732 14482
rect 9680 14418 9732 14424
rect 9864 14476 9916 14482
rect 9864 14418 9916 14424
rect 10416 14476 10468 14482
rect 10416 14418 10468 14424
rect 8944 14408 8996 14414
rect 8944 14350 8996 14356
rect 8956 14074 8984 14350
rect 9496 14272 9548 14278
rect 9496 14214 9548 14220
rect 8944 14068 8996 14074
rect 8944 14010 8996 14016
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 8484 13184 8536 13190
rect 8484 13126 8536 13132
rect 8496 12986 8524 13126
rect 8484 12980 8536 12986
rect 8484 12922 8536 12928
rect 8772 12850 8800 13874
rect 9508 13870 9536 14214
rect 9496 13864 9548 13870
rect 9496 13806 9548 13812
rect 9312 13728 9364 13734
rect 9312 13670 9364 13676
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 8668 12640 8720 12646
rect 8668 12582 8720 12588
rect 8300 12368 8352 12374
rect 8300 12310 8352 12316
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 8024 11892 8076 11898
rect 8024 11834 8076 11840
rect 7564 11824 7616 11830
rect 7564 11766 7616 11772
rect 8220 11762 8248 12174
rect 8392 11892 8444 11898
rect 8392 11834 8444 11840
rect 7656 11756 7708 11762
rect 7656 11698 7708 11704
rect 8208 11756 8260 11762
rect 8208 11698 8260 11704
rect 7196 11552 7248 11558
rect 7196 11494 7248 11500
rect 7104 11348 7156 11354
rect 7104 11290 7156 11296
rect 7024 11206 7144 11234
rect 7116 11014 7144 11206
rect 7208 11150 7236 11494
rect 7668 11150 7696 11698
rect 8404 11354 8432 11834
rect 8484 11756 8536 11762
rect 8484 11698 8536 11704
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7656 11144 7708 11150
rect 7656 11086 7708 11092
rect 7104 11008 7156 11014
rect 7104 10950 7156 10956
rect 7380 11008 7432 11014
rect 7380 10950 7432 10956
rect 7116 10538 7144 10950
rect 7288 10736 7340 10742
rect 7288 10678 7340 10684
rect 7104 10532 7156 10538
rect 7104 10474 7156 10480
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 6380 9926 6408 10406
rect 7300 10062 7328 10678
rect 7392 10606 7420 10950
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7288 10056 7340 10062
rect 7288 9998 7340 10004
rect 6368 9920 6420 9926
rect 6368 9862 6420 9868
rect 6380 9722 6408 9862
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 5356 9648 5408 9654
rect 5356 9590 5408 9596
rect 7104 9512 7156 9518
rect 7104 9454 7156 9460
rect 7116 9110 7144 9454
rect 7104 9104 7156 9110
rect 7104 9046 7156 9052
rect 7300 9042 7328 9998
rect 6552 9036 6604 9042
rect 7196 9036 7248 9042
rect 6604 8996 6684 9024
rect 6552 8978 6604 8984
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 5460 8362 5488 8910
rect 6276 8832 6328 8838
rect 6276 8774 6328 8780
rect 6368 8832 6420 8838
rect 6368 8774 6420 8780
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 5460 7410 5488 8298
rect 5816 8288 5868 8294
rect 5816 8230 5868 8236
rect 6092 8288 6144 8294
rect 6092 8230 6144 8236
rect 5828 8090 5856 8230
rect 5816 8084 5868 8090
rect 5816 8026 5868 8032
rect 6104 8022 6132 8230
rect 6092 8016 6144 8022
rect 6092 7958 6144 7964
rect 6288 7750 6316 8774
rect 6380 8634 6408 8774
rect 6368 8628 6420 8634
rect 6368 8570 6420 8576
rect 6656 8401 6684 8996
rect 7196 8978 7248 8984
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 6642 8392 6698 8401
rect 6642 8327 6644 8336
rect 6696 8327 6698 8336
rect 6644 8298 6696 8304
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6552 7812 6604 7818
rect 6552 7754 6604 7760
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 6274 7440 6330 7449
rect 5448 7404 5500 7410
rect 6274 7375 6276 7384
rect 5448 7346 5500 7352
rect 6328 7375 6330 7384
rect 6276 7346 6328 7352
rect 4896 7268 4948 7274
rect 4896 7210 4948 7216
rect 4804 6792 4856 6798
rect 4908 6746 4936 7210
rect 4856 6740 4936 6746
rect 4804 6734 4936 6740
rect 4816 6718 4936 6734
rect 4908 6458 4936 6718
rect 4896 6452 4948 6458
rect 4896 6394 4948 6400
rect 4620 5772 4672 5778
rect 4620 5714 4672 5720
rect 5172 5772 5224 5778
rect 5172 5714 5224 5720
rect 4988 5704 5040 5710
rect 4988 5646 5040 5652
rect 4066 5536 4122 5545
rect 4066 5471 4122 5480
rect 4080 5370 4108 5471
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 5000 5302 5028 5646
rect 5184 5642 5212 5714
rect 5460 5710 5488 7346
rect 6564 7342 6592 7754
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 6748 7410 6776 7686
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 6552 7336 6604 7342
rect 6552 7278 6604 7284
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 5172 5636 5224 5642
rect 5172 5578 5224 5584
rect 5184 5302 5212 5578
rect 4988 5296 5040 5302
rect 4988 5238 5040 5244
rect 5172 5296 5224 5302
rect 5172 5238 5224 5244
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 4080 4758 4108 5102
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 4068 4752 4120 4758
rect 4068 4694 4120 4700
rect 4526 4720 4582 4729
rect 4526 4655 4528 4664
rect 4580 4655 4582 4664
rect 5172 4684 5224 4690
rect 4528 4626 4580 4632
rect 5172 4626 5224 4632
rect 4540 4282 4568 4626
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 4528 4276 4580 4282
rect 4528 4218 4580 4224
rect 4068 4072 4120 4078
rect 4066 4040 4068 4049
rect 4120 4040 4122 4049
rect 4066 3975 4122 3984
rect 4816 3738 4844 4558
rect 5184 4214 5212 4626
rect 5368 4486 5396 4966
rect 5356 4480 5408 4486
rect 5356 4422 5408 4428
rect 5172 4208 5224 4214
rect 5172 4150 5224 4156
rect 5368 4078 5396 4422
rect 5356 4072 5408 4078
rect 5356 4014 5408 4020
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4802 3632 4858 3641
rect 4802 3567 4858 3576
rect 4712 2916 4764 2922
rect 4712 2858 4764 2864
rect 3698 2751 3754 2760
rect 3804 2774 4016 2802
rect 3804 2666 3832 2774
rect 3804 2638 3924 2666
rect 3608 2440 3660 2446
rect 3608 2382 3660 2388
rect 3896 800 3924 2638
rect 4724 2514 4752 2858
rect 4712 2508 4764 2514
rect 4712 2450 4764 2456
rect 4068 1352 4120 1358
rect 4068 1294 4120 1300
rect 4080 1193 4108 1294
rect 4066 1184 4122 1193
rect 4066 1119 4122 1128
rect 4816 800 4844 3567
rect 5356 3392 5408 3398
rect 5356 3334 5408 3340
rect 5368 3058 5396 3334
rect 5356 3052 5408 3058
rect 5356 2994 5408 3000
rect 5552 898 5580 7142
rect 6564 6934 6592 7278
rect 6748 6934 6776 7346
rect 6840 7206 6868 7822
rect 7104 7336 7156 7342
rect 7104 7278 7156 7284
rect 6828 7200 6880 7206
rect 6828 7142 6880 7148
rect 6552 6928 6604 6934
rect 6552 6870 6604 6876
rect 6736 6928 6788 6934
rect 6736 6870 6788 6876
rect 6920 6928 6972 6934
rect 6920 6870 6972 6876
rect 6564 5846 6592 6870
rect 6748 6322 6776 6870
rect 6932 6458 6960 6870
rect 6920 6452 6972 6458
rect 6920 6394 6972 6400
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 6644 6112 6696 6118
rect 6644 6054 6696 6060
rect 6552 5840 6604 5846
rect 6552 5782 6604 5788
rect 6184 5772 6236 5778
rect 6184 5714 6236 5720
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 5724 5568 5776 5574
rect 5724 5510 5776 5516
rect 5644 5166 5672 5510
rect 5632 5160 5684 5166
rect 5632 5102 5684 5108
rect 5644 4010 5672 5102
rect 5632 4004 5684 4010
rect 5632 3946 5684 3952
rect 5736 3738 5764 5510
rect 6196 5302 6224 5714
rect 6184 5296 6236 5302
rect 6184 5238 6236 5244
rect 5816 5024 5868 5030
rect 5814 4992 5816 5001
rect 5868 4992 5870 5001
rect 5814 4927 5870 4936
rect 6552 3936 6604 3942
rect 6552 3878 6604 3884
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5736 3466 5764 3674
rect 5908 3596 5960 3602
rect 5908 3538 5960 3544
rect 5724 3460 5776 3466
rect 5724 3402 5776 3408
rect 5736 2650 5764 3402
rect 5920 3194 5948 3538
rect 6184 3528 6236 3534
rect 6184 3470 6236 3476
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 5920 2990 5948 3130
rect 5908 2984 5960 2990
rect 5908 2926 5960 2932
rect 6196 2650 6224 3470
rect 5724 2644 5776 2650
rect 5724 2586 5776 2592
rect 6184 2644 6236 2650
rect 6184 2586 6236 2592
rect 5552 870 5672 898
rect 5644 800 5672 870
rect 6564 800 6592 3878
rect 6656 3602 6684 6054
rect 6932 5914 6960 6394
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 7024 5166 7052 5510
rect 7012 5160 7064 5166
rect 7012 5102 7064 5108
rect 7024 4146 7052 5102
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 6644 3596 6696 3602
rect 6644 3538 6696 3544
rect 6656 3194 6684 3538
rect 7024 3466 7052 4082
rect 7116 3942 7144 7278
rect 7208 6730 7236 8978
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 7300 7954 7328 8434
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 7300 7002 7328 7890
rect 7288 6996 7340 7002
rect 7288 6938 7340 6944
rect 7196 6724 7248 6730
rect 7196 6666 7248 6672
rect 7392 6458 7420 10542
rect 7484 10470 7512 11086
rect 7668 10810 7696 11086
rect 8300 11076 8352 11082
rect 8300 11018 8352 11024
rect 8312 10810 8340 11018
rect 8404 11014 8432 11290
rect 8392 11008 8444 11014
rect 8392 10950 8444 10956
rect 7656 10804 7708 10810
rect 7656 10746 7708 10752
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 8496 10713 8524 11698
rect 8680 11694 8708 12582
rect 8772 12442 8800 12786
rect 9128 12776 9180 12782
rect 9128 12718 9180 12724
rect 8760 12436 8812 12442
rect 8760 12378 8812 12384
rect 9140 12374 9168 12718
rect 9128 12368 9180 12374
rect 9324 12345 9352 13670
rect 9402 13560 9458 13569
rect 9402 13495 9458 13504
rect 9416 13190 9444 13495
rect 9404 13184 9456 13190
rect 9404 13126 9456 13132
rect 9128 12310 9180 12316
rect 9310 12336 9366 12345
rect 9310 12271 9366 12280
rect 9416 12170 9444 13126
rect 9508 12646 9536 13806
rect 9588 13796 9640 13802
rect 9588 13738 9640 13744
rect 9600 13326 9628 13738
rect 9692 13326 9720 14418
rect 9876 13569 9904 14418
rect 10324 14408 10376 14414
rect 10324 14350 10376 14356
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 9968 13734 9996 13874
rect 9956 13728 10008 13734
rect 9956 13670 10008 13676
rect 9862 13560 9918 13569
rect 9862 13495 9918 13504
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 9588 13320 9640 13326
rect 9588 13262 9640 13268
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9600 12889 9628 13262
rect 9784 12986 9812 13330
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9586 12880 9642 12889
rect 9586 12815 9642 12824
rect 9496 12640 9548 12646
rect 9494 12608 9496 12617
rect 9548 12608 9550 12617
rect 9494 12543 9550 12552
rect 9404 12164 9456 12170
rect 9404 12106 9456 12112
rect 9784 11694 9812 12922
rect 9968 12850 9996 13670
rect 10232 13184 10284 13190
rect 10232 13126 10284 13132
rect 10244 12850 10272 13126
rect 9956 12844 10008 12850
rect 9956 12786 10008 12792
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 10336 12714 10364 14350
rect 10796 14074 10824 14554
rect 11152 14340 11204 14346
rect 11152 14282 11204 14288
rect 10784 14068 10836 14074
rect 10784 14010 10836 14016
rect 11164 13954 11192 14282
rect 11256 14074 11284 14758
rect 11532 14414 11560 14826
rect 11520 14408 11572 14414
rect 11520 14350 11572 14356
rect 11352 14172 11648 14192
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11430 14118 11432 14170
rect 11494 14118 11506 14170
rect 11568 14118 11570 14170
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11352 14096 11648 14116
rect 11244 14068 11296 14074
rect 11244 14010 11296 14016
rect 11164 13938 11284 13954
rect 11164 13932 11296 13938
rect 11164 13926 11244 13932
rect 11244 13874 11296 13880
rect 11152 13864 11204 13870
rect 11152 13806 11204 13812
rect 10600 13728 10652 13734
rect 10600 13670 10652 13676
rect 10612 13462 10640 13670
rect 10600 13456 10652 13462
rect 10600 13398 10652 13404
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 10508 13252 10560 13258
rect 10508 13194 10560 13200
rect 10324 12708 10376 12714
rect 10324 12650 10376 12656
rect 10336 12442 10364 12650
rect 9864 12436 9916 12442
rect 9864 12378 9916 12384
rect 10324 12436 10376 12442
rect 10324 12378 10376 12384
rect 8668 11688 8720 11694
rect 8668 11630 8720 11636
rect 8852 11688 8904 11694
rect 8852 11630 8904 11636
rect 9772 11688 9824 11694
rect 9772 11630 9824 11636
rect 8680 10810 8708 11630
rect 8864 11286 8892 11630
rect 9784 11558 9812 11630
rect 9772 11552 9824 11558
rect 9772 11494 9824 11500
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 8852 11280 8904 11286
rect 8852 11222 8904 11228
rect 8760 11008 8812 11014
rect 8760 10950 8812 10956
rect 8668 10804 8720 10810
rect 8668 10746 8720 10752
rect 8482 10704 8538 10713
rect 8772 10690 8800 10950
rect 8482 10639 8538 10648
rect 8680 10662 8800 10690
rect 8680 10606 8708 10662
rect 7840 10600 7892 10606
rect 7840 10542 7892 10548
rect 8668 10600 8720 10606
rect 8668 10542 8720 10548
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 7484 10198 7512 10406
rect 7472 10192 7524 10198
rect 7472 10134 7524 10140
rect 7852 10062 7880 10542
rect 7840 10056 7892 10062
rect 7840 9998 7892 10004
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 7562 7984 7618 7993
rect 7562 7919 7564 7928
rect 7616 7919 7618 7928
rect 7564 7890 7616 7896
rect 7576 7750 7604 7890
rect 8036 7886 8064 8978
rect 8208 8900 8260 8906
rect 8208 8842 8260 8848
rect 8220 8362 8248 8842
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 8220 8090 8248 8298
rect 8208 8084 8260 8090
rect 8208 8026 8260 8032
rect 8024 7880 8076 7886
rect 8024 7822 8076 7828
rect 8208 7812 8260 7818
rect 8208 7754 8260 7760
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 7196 6180 7248 6186
rect 7196 6122 7248 6128
rect 7208 5914 7236 6122
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 7288 4616 7340 4622
rect 7288 4558 7340 4564
rect 7300 4282 7328 4558
rect 7288 4276 7340 4282
rect 7288 4218 7340 4224
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 7484 3738 7512 3878
rect 7472 3732 7524 3738
rect 7472 3674 7524 3680
rect 7576 3618 7604 7686
rect 7748 7472 7800 7478
rect 7748 7414 7800 7420
rect 7760 7342 7788 7414
rect 7748 7336 7800 7342
rect 7748 7278 7800 7284
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 7760 5710 7788 7278
rect 7944 7002 7972 7278
rect 8220 7274 8248 7754
rect 8208 7268 8260 7274
rect 8208 7210 8260 7216
rect 7932 6996 7984 7002
rect 7932 6938 7984 6944
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 8220 6662 8248 6802
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8208 6656 8260 6662
rect 8208 6598 8260 6604
rect 8116 6248 8168 6254
rect 8116 6190 8168 6196
rect 7748 5704 7800 5710
rect 7748 5646 7800 5652
rect 7760 5302 7788 5646
rect 8128 5642 8156 6190
rect 8220 6186 8248 6598
rect 8208 6180 8260 6186
rect 8208 6122 8260 6128
rect 8220 5846 8248 6122
rect 8312 6118 8340 6734
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8208 5840 8260 5846
rect 8208 5782 8260 5788
rect 8392 5840 8444 5846
rect 8392 5782 8444 5788
rect 8300 5772 8352 5778
rect 8300 5714 8352 5720
rect 8116 5636 8168 5642
rect 8116 5578 8168 5584
rect 8312 5302 8340 5714
rect 7748 5296 7800 5302
rect 7748 5238 7800 5244
rect 8300 5296 8352 5302
rect 8300 5238 8352 5244
rect 7932 5228 7984 5234
rect 7932 5170 7984 5176
rect 7840 5024 7892 5030
rect 7840 4966 7892 4972
rect 7852 4690 7880 4966
rect 7840 4684 7892 4690
rect 7840 4626 7892 4632
rect 7852 4486 7880 4626
rect 7840 4480 7892 4486
rect 7840 4422 7892 4428
rect 7852 3942 7880 4422
rect 7840 3936 7892 3942
rect 7840 3878 7892 3884
rect 7840 3732 7892 3738
rect 7840 3674 7892 3680
rect 7484 3590 7604 3618
rect 7748 3596 7800 3602
rect 7012 3460 7064 3466
rect 7012 3402 7064 3408
rect 6828 3392 6880 3398
rect 6828 3334 6880 3340
rect 7196 3392 7248 3398
rect 7196 3334 7248 3340
rect 7288 3392 7340 3398
rect 7288 3334 7340 3340
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 6840 3126 6868 3334
rect 6828 3120 6880 3126
rect 6828 3062 6880 3068
rect 7208 3058 7236 3334
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 7300 1426 7328 3334
rect 7288 1420 7340 1426
rect 7288 1362 7340 1368
rect 7484 800 7512 3590
rect 7748 3538 7800 3544
rect 7656 3460 7708 3466
rect 7656 3402 7708 3408
rect 7668 2990 7696 3402
rect 7760 3194 7788 3538
rect 7748 3188 7800 3194
rect 7748 3130 7800 3136
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 7656 2984 7708 2990
rect 7656 2926 7708 2932
rect 7760 2666 7788 2994
rect 7852 2990 7880 3674
rect 7944 3670 7972 5170
rect 8024 5160 8076 5166
rect 8024 5102 8076 5108
rect 8298 5128 8354 5137
rect 8036 4486 8064 5102
rect 8298 5063 8300 5072
rect 8352 5063 8354 5072
rect 8300 5034 8352 5040
rect 8024 4480 8076 4486
rect 8024 4422 8076 4428
rect 8036 4078 8064 4422
rect 8024 4072 8076 4078
rect 8024 4014 8076 4020
rect 8036 3942 8064 4014
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 7932 3664 7984 3670
rect 7932 3606 7984 3612
rect 7944 3058 7972 3606
rect 8300 3596 8352 3602
rect 8404 3584 8432 5782
rect 8576 5092 8628 5098
rect 8576 5034 8628 5040
rect 8588 3738 8616 5034
rect 8680 4690 8708 10542
rect 8864 10266 8892 11222
rect 9784 10742 9812 11290
rect 9772 10736 9824 10742
rect 9772 10678 9824 10684
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 8852 10260 8904 10266
rect 8852 10202 8904 10208
rect 9784 10130 9812 10406
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 8944 9988 8996 9994
rect 8944 9930 8996 9936
rect 8956 9382 8984 9930
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 9324 9518 9352 9862
rect 9692 9654 9720 9998
rect 9680 9648 9732 9654
rect 9680 9590 9732 9596
rect 9312 9512 9364 9518
rect 9312 9454 9364 9460
rect 8944 9376 8996 9382
rect 8944 9318 8996 9324
rect 8760 9036 8812 9042
rect 8760 8978 8812 8984
rect 8772 8634 8800 8978
rect 8760 8628 8812 8634
rect 8760 8570 8812 8576
rect 8852 8356 8904 8362
rect 8852 8298 8904 8304
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 8772 7478 8800 7686
rect 8864 7546 8892 8298
rect 8852 7540 8904 7546
rect 8852 7482 8904 7488
rect 8760 7472 8812 7478
rect 8760 7414 8812 7420
rect 8956 5574 8984 9318
rect 9324 6458 9352 9454
rect 9692 8378 9720 9590
rect 9876 9450 9904 12378
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 9968 11150 9996 11494
rect 9956 11144 10008 11150
rect 9956 11086 10008 11092
rect 9968 10810 9996 11086
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 9956 10056 10008 10062
rect 9956 9998 10008 10004
rect 9968 9722 9996 9998
rect 10520 9926 10548 13194
rect 10704 12306 10732 13262
rect 11164 13190 11192 13806
rect 11704 13796 11756 13802
rect 11704 13738 11756 13744
rect 11716 13462 11744 13738
rect 11704 13456 11756 13462
rect 11704 13398 11756 13404
rect 11992 13394 12020 15302
rect 12176 14890 12204 15506
rect 12164 14884 12216 14890
rect 12164 14826 12216 14832
rect 11980 13388 12032 13394
rect 11980 13330 12032 13336
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 11164 12442 11192 13126
rect 11352 13084 11648 13104
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11430 13030 11432 13082
rect 11494 13030 11506 13082
rect 11568 13030 11570 13082
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11352 13008 11648 13028
rect 11992 12850 12020 13330
rect 12072 13184 12124 13190
rect 12072 13126 12124 13132
rect 11980 12844 12032 12850
rect 11980 12786 12032 12792
rect 11244 12708 11296 12714
rect 11244 12650 11296 12656
rect 11888 12708 11940 12714
rect 11888 12650 11940 12656
rect 11152 12436 11204 12442
rect 11152 12378 11204 12384
rect 10692 12300 10744 12306
rect 10692 12242 10744 12248
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 10612 11694 10640 12038
rect 10600 11688 10652 11694
rect 10600 11630 10652 11636
rect 10704 11354 10732 12242
rect 10968 12096 11020 12102
rect 10968 12038 11020 12044
rect 10980 11898 11008 12038
rect 10968 11892 11020 11898
rect 10968 11834 11020 11840
rect 11256 11694 11284 12650
rect 11900 12238 11928 12650
rect 12084 12442 12112 13126
rect 12268 12646 12296 15982
rect 12636 14958 12664 16730
rect 13924 16658 13952 17070
rect 13912 16652 13964 16658
rect 13912 16594 13964 16600
rect 13360 15972 13412 15978
rect 13360 15914 13412 15920
rect 13268 15904 13320 15910
rect 13268 15846 13320 15852
rect 13280 15366 13308 15846
rect 13372 15638 13400 15914
rect 13360 15632 13412 15638
rect 13360 15574 13412 15580
rect 13820 15428 13872 15434
rect 13820 15370 13872 15376
rect 13268 15360 13320 15366
rect 13268 15302 13320 15308
rect 13280 14958 13308 15302
rect 12624 14952 12676 14958
rect 12624 14894 12676 14900
rect 13268 14952 13320 14958
rect 13268 14894 13320 14900
rect 13452 14952 13504 14958
rect 13452 14894 13504 14900
rect 12900 14816 12952 14822
rect 12900 14758 12952 14764
rect 12440 14408 12492 14414
rect 12440 14350 12492 14356
rect 12452 13870 12480 14350
rect 12440 13864 12492 13870
rect 12440 13806 12492 13812
rect 12622 13696 12678 13705
rect 12622 13631 12678 13640
rect 12636 13394 12664 13631
rect 12624 13388 12676 13394
rect 12544 13348 12624 13376
rect 12544 12918 12572 13348
rect 12624 13330 12676 13336
rect 12624 13252 12676 13258
rect 12624 13194 12676 13200
rect 12716 13252 12768 13258
rect 12716 13194 12768 13200
rect 12532 12912 12584 12918
rect 12532 12854 12584 12860
rect 12256 12640 12308 12646
rect 12256 12582 12308 12588
rect 12072 12436 12124 12442
rect 12072 12378 12124 12384
rect 12164 12436 12216 12442
rect 12164 12378 12216 12384
rect 12176 12306 12204 12378
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 12532 12300 12584 12306
rect 12532 12242 12584 12248
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11352 11996 11648 12016
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11430 11942 11432 11994
rect 11494 11942 11506 11994
rect 11568 11942 11570 11994
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11352 11920 11648 11940
rect 11244 11688 11296 11694
rect 11244 11630 11296 11636
rect 11256 11354 11284 11630
rect 10692 11348 10744 11354
rect 10692 11290 10744 11296
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 11796 11076 11848 11082
rect 11796 11018 11848 11024
rect 11352 10908 11648 10928
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11430 10854 11432 10906
rect 11494 10854 11506 10906
rect 11568 10854 11570 10906
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11352 10832 11648 10852
rect 10692 10736 10744 10742
rect 10692 10678 10744 10684
rect 10704 9994 10732 10678
rect 11808 10130 11836 11018
rect 11900 10810 11928 12174
rect 12164 12164 12216 12170
rect 12164 12106 12216 12112
rect 12176 11898 12204 12106
rect 12544 11898 12572 12242
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 12532 11892 12584 11898
rect 12532 11834 12584 11840
rect 11980 11212 12032 11218
rect 11980 11154 12032 11160
rect 12072 11212 12124 11218
rect 12072 11154 12124 11160
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 10876 10124 10928 10130
rect 10876 10066 10928 10072
rect 11796 10124 11848 10130
rect 11796 10066 11848 10072
rect 10692 9988 10744 9994
rect 10692 9930 10744 9936
rect 10888 9926 10916 10066
rect 10508 9920 10560 9926
rect 10508 9862 10560 9868
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 9956 9716 10008 9722
rect 9956 9658 10008 9664
rect 10520 9586 10548 9862
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 9864 9444 9916 9450
rect 9864 9386 9916 9392
rect 10520 9042 10548 9522
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10704 9382 10732 9454
rect 10888 9450 10916 9862
rect 11352 9820 11648 9840
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11430 9766 11432 9818
rect 11494 9766 11506 9818
rect 11568 9766 11570 9818
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11352 9744 11648 9764
rect 11808 9722 11836 10066
rect 11796 9716 11848 9722
rect 11796 9658 11848 9664
rect 10876 9444 10928 9450
rect 10876 9386 10928 9392
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 11060 9376 11112 9382
rect 11060 9318 11112 9324
rect 10140 9036 10192 9042
rect 10140 8978 10192 8984
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 9600 8350 9720 8378
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 8852 5568 8904 5574
rect 8852 5510 8904 5516
rect 8944 5568 8996 5574
rect 8944 5510 8996 5516
rect 8864 5166 8892 5510
rect 8852 5160 8904 5166
rect 8852 5102 8904 5108
rect 8864 4758 8892 5102
rect 8942 4992 8998 5001
rect 8942 4927 8998 4936
rect 8760 4752 8812 4758
rect 8760 4694 8812 4700
rect 8852 4752 8904 4758
rect 8852 4694 8904 4700
rect 8668 4684 8720 4690
rect 8668 4626 8720 4632
rect 8680 4486 8708 4626
rect 8668 4480 8720 4486
rect 8668 4422 8720 4428
rect 8772 4282 8800 4694
rect 8864 4622 8892 4694
rect 8852 4616 8904 4622
rect 8852 4558 8904 4564
rect 8760 4276 8812 4282
rect 8760 4218 8812 4224
rect 8864 4214 8892 4558
rect 8852 4208 8904 4214
rect 8852 4150 8904 4156
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 8956 3670 8984 4927
rect 8944 3664 8996 3670
rect 8944 3606 8996 3612
rect 8352 3556 8432 3584
rect 8300 3538 8352 3544
rect 8404 3058 8432 3556
rect 9036 3460 9088 3466
rect 9036 3402 9088 3408
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 8392 3052 8444 3058
rect 8392 2994 8444 3000
rect 9048 2990 9076 3402
rect 7840 2984 7892 2990
rect 7838 2952 7840 2961
rect 9036 2984 9088 2990
rect 7892 2952 7894 2961
rect 9036 2926 9088 2932
rect 7838 2887 7894 2896
rect 8116 2916 8168 2922
rect 8116 2858 8168 2864
rect 7760 2638 7880 2666
rect 7852 2310 7880 2638
rect 8128 2514 8156 2858
rect 8300 2848 8352 2854
rect 8300 2790 8352 2796
rect 8116 2508 8168 2514
rect 8116 2450 8168 2456
rect 7840 2304 7892 2310
rect 7840 2246 7892 2252
rect 8312 800 8340 2790
rect 9048 2650 9076 2926
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 9232 2038 9260 6190
rect 9312 6112 9364 6118
rect 9312 6054 9364 6060
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9324 5166 9352 6054
rect 9404 5908 9456 5914
rect 9404 5850 9456 5856
rect 9416 5234 9444 5850
rect 9508 5302 9536 6054
rect 9496 5296 9548 5302
rect 9496 5238 9548 5244
rect 9404 5228 9456 5234
rect 9404 5170 9456 5176
rect 9312 5160 9364 5166
rect 9312 5102 9364 5108
rect 9600 4622 9628 8350
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 9968 7206 9996 7890
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 9968 7002 9996 7142
rect 9956 6996 10008 7002
rect 9956 6938 10008 6944
rect 10152 6322 10180 8978
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 10508 8832 10560 8838
rect 10508 8774 10560 8780
rect 10232 7336 10284 7342
rect 10232 7278 10284 7284
rect 10244 6798 10272 7278
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 9784 5778 9812 6190
rect 9772 5772 9824 5778
rect 9772 5714 9824 5720
rect 9680 5704 9732 5710
rect 9680 5646 9732 5652
rect 9692 4690 9720 5646
rect 9784 5234 9812 5714
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 9784 4690 9812 5170
rect 10244 5030 10272 5646
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 10324 5160 10376 5166
rect 10324 5102 10376 5108
rect 10048 5024 10100 5030
rect 10048 4966 10100 4972
rect 10232 5024 10284 5030
rect 10232 4966 10284 4972
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 9588 4616 9640 4622
rect 9588 4558 9640 4564
rect 9496 4480 9548 4486
rect 9496 4422 9548 4428
rect 9508 4214 9536 4422
rect 9600 4282 9628 4558
rect 9588 4276 9640 4282
rect 9588 4218 9640 4224
rect 9496 4208 9548 4214
rect 9496 4150 9548 4156
rect 9496 4004 9548 4010
rect 9600 3992 9628 4218
rect 9864 4072 9916 4078
rect 9864 4014 9916 4020
rect 9548 3964 9628 3992
rect 9496 3946 9548 3952
rect 9600 3890 9628 3964
rect 9772 3936 9824 3942
rect 9600 3862 9720 3890
rect 9772 3878 9824 3884
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 9324 3058 9352 3470
rect 9404 3460 9456 3466
rect 9404 3402 9456 3408
rect 9312 3052 9364 3058
rect 9312 2994 9364 3000
rect 9416 2582 9444 3402
rect 9600 3058 9628 3674
rect 9692 3466 9720 3862
rect 9680 3460 9732 3466
rect 9680 3402 9732 3408
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 9784 2990 9812 3878
rect 9876 3738 9904 4014
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9772 2984 9824 2990
rect 9772 2926 9824 2932
rect 9588 2916 9640 2922
rect 9588 2858 9640 2864
rect 9600 2650 9628 2858
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 9404 2576 9456 2582
rect 9404 2518 9456 2524
rect 9220 2032 9272 2038
rect 9220 1974 9272 1980
rect 9232 800 9260 1974
rect 10060 800 10088 4966
rect 10138 4856 10194 4865
rect 10138 4791 10194 4800
rect 10152 4690 10180 4791
rect 10140 4684 10192 4690
rect 10140 4626 10192 4632
rect 10152 3602 10180 4626
rect 10140 3596 10192 3602
rect 10140 3538 10192 3544
rect 10336 2854 10364 5102
rect 10428 4214 10456 5510
rect 10520 5234 10548 8774
rect 10612 7886 10640 8910
rect 10600 7880 10652 7886
rect 10600 7822 10652 7828
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 10704 4486 10732 9318
rect 10876 9036 10928 9042
rect 10876 8978 10928 8984
rect 10784 8968 10836 8974
rect 10784 8910 10836 8916
rect 10796 6798 10824 8910
rect 10888 8498 10916 8978
rect 11072 8566 11100 9318
rect 11150 8936 11206 8945
rect 11150 8871 11152 8880
rect 11204 8871 11206 8880
rect 11152 8842 11204 8848
rect 11164 8634 11192 8842
rect 11352 8732 11648 8752
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11430 8678 11432 8730
rect 11494 8678 11506 8730
rect 11568 8678 11570 8730
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11352 8656 11648 8676
rect 11886 8664 11942 8673
rect 11152 8628 11204 8634
rect 11886 8599 11888 8608
rect 11152 8570 11204 8576
rect 11940 8599 11942 8608
rect 11888 8570 11940 8576
rect 11060 8560 11112 8566
rect 11060 8502 11112 8508
rect 10876 8492 10928 8498
rect 10876 8434 10928 8440
rect 11164 8412 11192 8570
rect 11244 8424 11296 8430
rect 11164 8384 11244 8412
rect 11244 8366 11296 8372
rect 11520 8356 11572 8362
rect 11520 8298 11572 8304
rect 11532 8090 11560 8298
rect 11520 8084 11572 8090
rect 11520 8026 11572 8032
rect 11244 7948 11296 7954
rect 11244 7890 11296 7896
rect 11888 7948 11940 7954
rect 11888 7890 11940 7896
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 10876 7200 10928 7206
rect 10876 7142 10928 7148
rect 10784 6792 10836 6798
rect 10784 6734 10836 6740
rect 10796 6322 10824 6734
rect 10784 6316 10836 6322
rect 10784 6258 10836 6264
rect 10784 4548 10836 4554
rect 10784 4490 10836 4496
rect 10692 4480 10744 4486
rect 10692 4422 10744 4428
rect 10416 4208 10468 4214
rect 10416 4150 10468 4156
rect 10704 3942 10732 4422
rect 10796 4078 10824 4490
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 10796 3942 10824 4014
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 10784 3936 10836 3942
rect 10784 3878 10836 3884
rect 10416 3052 10468 3058
rect 10416 2994 10468 3000
rect 10324 2848 10376 2854
rect 10324 2790 10376 2796
rect 10428 2650 10456 2994
rect 10704 2689 10732 3878
rect 10888 3398 10916 7142
rect 10980 6089 11008 7686
rect 11256 6662 11284 7890
rect 11352 7644 11648 7664
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11430 7590 11432 7642
rect 11494 7590 11506 7642
rect 11568 7590 11570 7642
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11352 7568 11648 7588
rect 11900 7585 11928 7890
rect 11886 7576 11942 7585
rect 11886 7511 11942 7520
rect 11900 7206 11928 7511
rect 11888 7200 11940 7206
rect 11888 7142 11940 7148
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11352 6556 11648 6576
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11430 6502 11432 6554
rect 11494 6502 11506 6554
rect 11568 6502 11570 6554
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11352 6480 11648 6500
rect 11060 6248 11112 6254
rect 11060 6190 11112 6196
rect 10966 6080 11022 6089
rect 10966 6015 11022 6024
rect 11072 5778 11100 6190
rect 11716 5846 11744 6598
rect 11992 6254 12020 11154
rect 12084 10742 12112 11154
rect 12072 10736 12124 10742
rect 12072 10678 12124 10684
rect 12072 10056 12124 10062
rect 12072 9998 12124 10004
rect 12084 9466 12112 9998
rect 12176 9586 12204 11834
rect 12636 11830 12664 13194
rect 12728 12918 12756 13194
rect 12716 12912 12768 12918
rect 12716 12854 12768 12860
rect 12728 12102 12756 12854
rect 12808 12844 12860 12850
rect 12808 12786 12860 12792
rect 12820 12442 12848 12786
rect 12808 12436 12860 12442
rect 12808 12378 12860 12384
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 12624 11824 12676 11830
rect 12624 11766 12676 11772
rect 12348 11620 12400 11626
rect 12348 11562 12400 11568
rect 12256 11212 12308 11218
rect 12256 11154 12308 11160
rect 12268 9722 12296 11154
rect 12256 9716 12308 9722
rect 12256 9658 12308 9664
rect 12164 9580 12216 9586
rect 12164 9522 12216 9528
rect 12084 9438 12296 9466
rect 12268 8838 12296 9438
rect 12360 9042 12388 11562
rect 12808 11008 12860 11014
rect 12808 10950 12860 10956
rect 12624 10804 12676 10810
rect 12624 10746 12676 10752
rect 12636 9586 12664 10746
rect 12820 10674 12848 10950
rect 12912 10674 12940 14758
rect 13464 14482 13492 14894
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 13280 13938 13492 13954
rect 13268 13932 13504 13938
rect 13320 13926 13452 13932
rect 13268 13874 13320 13880
rect 13452 13874 13504 13880
rect 13832 13870 13860 15370
rect 13924 15366 13952 16594
rect 14280 16448 14332 16454
rect 14280 16390 14332 16396
rect 14292 16046 14320 16390
rect 14660 16250 14688 17274
rect 15752 17196 15804 17202
rect 15752 17138 15804 17144
rect 15764 16590 15792 17138
rect 16592 16810 16620 19162
rect 18524 17134 18552 19162
rect 19156 17264 19208 17270
rect 19156 17206 19208 17212
rect 18512 17128 18564 17134
rect 18512 17070 18564 17076
rect 18328 17060 18380 17066
rect 18328 17002 18380 17008
rect 16592 16794 16712 16810
rect 16592 16788 16724 16794
rect 16592 16782 16672 16788
rect 16672 16730 16724 16736
rect 17132 16788 17184 16794
rect 17132 16730 17184 16736
rect 15752 16584 15804 16590
rect 15752 16526 15804 16532
rect 16028 16584 16080 16590
rect 16028 16526 16080 16532
rect 14648 16244 14700 16250
rect 14648 16186 14700 16192
rect 14660 16114 14688 16186
rect 14648 16108 14700 16114
rect 14648 16050 14700 16056
rect 14280 16040 14332 16046
rect 14280 15982 14332 15988
rect 14292 15706 14320 15982
rect 15764 15910 15792 16526
rect 16040 16250 16068 16526
rect 16028 16244 16080 16250
rect 16028 16186 16080 16192
rect 16764 16108 16816 16114
rect 16764 16050 16816 16056
rect 17040 16108 17092 16114
rect 17040 16050 17092 16056
rect 16396 16040 16448 16046
rect 16396 15982 16448 15988
rect 15568 15904 15620 15910
rect 15568 15846 15620 15852
rect 15752 15904 15804 15910
rect 15752 15846 15804 15852
rect 14280 15700 14332 15706
rect 14200 15660 14280 15688
rect 14004 15564 14056 15570
rect 14004 15506 14056 15512
rect 13912 15360 13964 15366
rect 13912 15302 13964 15308
rect 14016 14278 14044 15506
rect 14096 15496 14148 15502
rect 14096 15438 14148 15444
rect 14108 15094 14136 15438
rect 14096 15088 14148 15094
rect 14096 15030 14148 15036
rect 14200 15026 14228 15660
rect 14280 15642 14332 15648
rect 15200 15564 15252 15570
rect 15200 15506 15252 15512
rect 15212 15026 15240 15506
rect 15580 15094 15608 15846
rect 15764 15502 15792 15846
rect 15752 15496 15804 15502
rect 15752 15438 15804 15444
rect 16408 15434 16436 15982
rect 16120 15428 16172 15434
rect 16120 15370 16172 15376
rect 16396 15428 16448 15434
rect 16396 15370 16448 15376
rect 15568 15088 15620 15094
rect 15568 15030 15620 15036
rect 14188 15020 14240 15026
rect 14188 14962 14240 14968
rect 15200 15020 15252 15026
rect 15200 14962 15252 14968
rect 14280 14952 14332 14958
rect 14280 14894 14332 14900
rect 16028 14952 16080 14958
rect 16028 14894 16080 14900
rect 14096 14544 14148 14550
rect 14096 14486 14148 14492
rect 14004 14272 14056 14278
rect 14004 14214 14056 14220
rect 14108 14226 14136 14486
rect 14292 14482 14320 14894
rect 16040 14822 16068 14894
rect 16028 14816 16080 14822
rect 16028 14758 16080 14764
rect 16040 14482 16068 14758
rect 14280 14476 14332 14482
rect 14280 14418 14332 14424
rect 15936 14476 15988 14482
rect 15936 14418 15988 14424
rect 16028 14476 16080 14482
rect 16028 14418 16080 14424
rect 13912 13932 13964 13938
rect 13912 13874 13964 13880
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 13636 13796 13688 13802
rect 13636 13738 13688 13744
rect 13082 13424 13138 13433
rect 13082 13359 13084 13368
rect 13136 13359 13138 13368
rect 13084 13330 13136 13336
rect 13648 12986 13676 13738
rect 13728 13524 13780 13530
rect 13728 13466 13780 13472
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 13084 12776 13136 12782
rect 13084 12718 13136 12724
rect 13096 12102 13124 12718
rect 13740 12646 13768 13466
rect 13924 13462 13952 13874
rect 13912 13456 13964 13462
rect 13912 13398 13964 13404
rect 13728 12640 13780 12646
rect 13728 12582 13780 12588
rect 13084 12096 13136 12102
rect 13084 12038 13136 12044
rect 12808 10668 12860 10674
rect 12808 10610 12860 10616
rect 12900 10668 12952 10674
rect 12900 10610 12952 10616
rect 12716 10056 12768 10062
rect 12716 9998 12768 10004
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12348 9036 12400 9042
rect 12348 8978 12400 8984
rect 12256 8832 12308 8838
rect 12256 8774 12308 8780
rect 12268 8514 12296 8774
rect 12360 8634 12388 8978
rect 12532 8968 12584 8974
rect 12532 8910 12584 8916
rect 12544 8634 12572 8910
rect 12348 8628 12400 8634
rect 12348 8570 12400 8576
rect 12532 8628 12584 8634
rect 12532 8570 12584 8576
rect 12072 8492 12124 8498
rect 12268 8486 12388 8514
rect 12072 8434 12124 8440
rect 12084 7886 12112 8434
rect 12072 7880 12124 7886
rect 12072 7822 12124 7828
rect 12360 7342 12388 8486
rect 12532 8016 12584 8022
rect 12532 7958 12584 7964
rect 12440 7812 12492 7818
rect 12440 7754 12492 7760
rect 12452 7342 12480 7754
rect 12544 7546 12572 7958
rect 12532 7540 12584 7546
rect 12532 7482 12584 7488
rect 12532 7404 12584 7410
rect 12532 7346 12584 7352
rect 12348 7336 12400 7342
rect 12348 7278 12400 7284
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 12256 7200 12308 7206
rect 12256 7142 12308 7148
rect 12268 7002 12296 7142
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 11980 6248 12032 6254
rect 11980 6190 12032 6196
rect 11704 5840 11756 5846
rect 11704 5782 11756 5788
rect 11060 5772 11112 5778
rect 11060 5714 11112 5720
rect 11888 5772 11940 5778
rect 11888 5714 11940 5720
rect 11072 5642 11100 5714
rect 11704 5704 11756 5710
rect 11704 5646 11756 5652
rect 11060 5636 11112 5642
rect 11060 5578 11112 5584
rect 11352 5468 11648 5488
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11430 5414 11432 5466
rect 11494 5414 11506 5466
rect 11568 5414 11570 5466
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11352 5392 11648 5412
rect 11716 5166 11744 5646
rect 11900 5302 11928 5714
rect 11888 5296 11940 5302
rect 11888 5238 11940 5244
rect 12360 5234 12388 7278
rect 12452 6186 12480 7278
rect 12544 6934 12572 7346
rect 12532 6928 12584 6934
rect 12532 6870 12584 6876
rect 12728 6474 12756 9998
rect 12820 9654 12848 10610
rect 12900 9920 12952 9926
rect 12900 9862 12952 9868
rect 12808 9648 12860 9654
rect 12808 9590 12860 9596
rect 12912 9518 12940 9862
rect 12900 9512 12952 9518
rect 12900 9454 12952 9460
rect 12728 6446 12848 6474
rect 12716 6384 12768 6390
rect 12716 6326 12768 6332
rect 12440 6180 12492 6186
rect 12440 6122 12492 6128
rect 12532 6112 12584 6118
rect 12532 6054 12584 6060
rect 12544 5642 12572 6054
rect 12532 5636 12584 5642
rect 12532 5578 12584 5584
rect 12348 5228 12400 5234
rect 12348 5170 12400 5176
rect 11704 5160 11756 5166
rect 11704 5102 11756 5108
rect 11886 5128 11942 5137
rect 12162 5128 12218 5137
rect 11886 5063 11942 5072
rect 12072 5092 12124 5098
rect 10968 5024 11020 5030
rect 10968 4966 11020 4972
rect 10876 3392 10928 3398
rect 10876 3334 10928 3340
rect 10690 2680 10746 2689
rect 10416 2644 10468 2650
rect 10690 2615 10746 2624
rect 10416 2586 10468 2592
rect 10980 800 11008 4966
rect 11900 4690 11928 5063
rect 12162 5063 12218 5072
rect 12072 5034 12124 5040
rect 12084 4758 12112 5034
rect 12176 4826 12204 5063
rect 12164 4820 12216 4826
rect 12164 4762 12216 4768
rect 12072 4752 12124 4758
rect 12072 4694 12124 4700
rect 11704 4684 11756 4690
rect 11704 4626 11756 4632
rect 11888 4684 11940 4690
rect 11888 4626 11940 4632
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 11072 4146 11100 4558
rect 11244 4480 11296 4486
rect 11244 4422 11296 4428
rect 11150 4176 11206 4185
rect 11060 4140 11112 4146
rect 11150 4111 11206 4120
rect 11060 4082 11112 4088
rect 11164 2990 11192 4111
rect 11256 4078 11284 4422
rect 11352 4380 11648 4400
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11430 4326 11432 4378
rect 11494 4326 11506 4378
rect 11568 4326 11570 4378
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11352 4304 11648 4324
rect 11716 4282 11744 4626
rect 11704 4276 11756 4282
rect 11704 4218 11756 4224
rect 11900 4214 11928 4626
rect 12544 4604 12572 5578
rect 12728 5114 12756 6326
rect 12820 5658 12848 6446
rect 12912 5846 12940 9454
rect 12992 9036 13044 9042
rect 12992 8978 13044 8984
rect 13004 8838 13032 8978
rect 12992 8832 13044 8838
rect 12992 8774 13044 8780
rect 13004 6866 13032 8774
rect 13096 7750 13124 12038
rect 13726 11792 13782 11801
rect 13726 11727 13782 11736
rect 13740 11626 13768 11727
rect 13728 11620 13780 11626
rect 13728 11562 13780 11568
rect 13452 10600 13504 10606
rect 13452 10542 13504 10548
rect 13464 8480 13492 10542
rect 13740 10062 13768 11562
rect 14016 11354 14044 14214
rect 14108 14198 14228 14226
rect 14200 13938 14228 14198
rect 14292 14006 14320 14418
rect 15948 14278 15976 14418
rect 14740 14272 14792 14278
rect 14740 14214 14792 14220
rect 14832 14272 14884 14278
rect 14832 14214 14884 14220
rect 15936 14272 15988 14278
rect 15936 14214 15988 14220
rect 14752 14074 14780 14214
rect 14372 14068 14424 14074
rect 14372 14010 14424 14016
rect 14740 14068 14792 14074
rect 14740 14010 14792 14016
rect 14280 14000 14332 14006
rect 14280 13942 14332 13948
rect 14188 13932 14240 13938
rect 14188 13874 14240 13880
rect 14096 13388 14148 13394
rect 14096 13330 14148 13336
rect 14108 12918 14136 13330
rect 14200 13326 14228 13874
rect 14188 13320 14240 13326
rect 14188 13262 14240 13268
rect 14096 12912 14148 12918
rect 14096 12854 14148 12860
rect 14108 12238 14136 12854
rect 14280 12300 14332 12306
rect 14280 12242 14332 12248
rect 14096 12232 14148 12238
rect 14096 12174 14148 12180
rect 14292 11694 14320 12242
rect 14280 11688 14332 11694
rect 14280 11630 14332 11636
rect 14004 11348 14056 11354
rect 14004 11290 14056 11296
rect 14292 11218 14320 11630
rect 14188 11212 14240 11218
rect 14188 11154 14240 11160
rect 14280 11212 14332 11218
rect 14280 11154 14332 11160
rect 13820 11008 13872 11014
rect 13820 10950 13872 10956
rect 13832 10266 13860 10950
rect 14200 10810 14228 11154
rect 14188 10804 14240 10810
rect 14188 10746 14240 10752
rect 14200 10266 14228 10746
rect 14292 10674 14320 11154
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 14188 10260 14240 10266
rect 14188 10202 14240 10208
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 13544 9648 13596 9654
rect 13544 9590 13596 9596
rect 13556 9042 13584 9590
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 13728 9036 13780 9042
rect 13728 8978 13780 8984
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 13464 8452 13584 8480
rect 13452 8356 13504 8362
rect 13452 8298 13504 8304
rect 13176 8288 13228 8294
rect 13176 8230 13228 8236
rect 13188 7954 13216 8230
rect 13176 7948 13228 7954
rect 13176 7890 13228 7896
rect 13084 7744 13136 7750
rect 13084 7686 13136 7692
rect 13084 7404 13136 7410
rect 13188 7392 13216 7890
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 13268 7744 13320 7750
rect 13268 7686 13320 7692
rect 13136 7364 13216 7392
rect 13084 7346 13136 7352
rect 12992 6860 13044 6866
rect 12992 6802 13044 6808
rect 13176 6112 13228 6118
rect 13280 6100 13308 7686
rect 13372 7478 13400 7822
rect 13360 7472 13412 7478
rect 13360 7414 13412 7420
rect 13228 6072 13308 6100
rect 13176 6054 13228 6060
rect 12900 5840 12952 5846
rect 12900 5782 12952 5788
rect 12820 5630 13032 5658
rect 12808 5568 12860 5574
rect 12808 5510 12860 5516
rect 12820 5234 12848 5510
rect 12808 5228 12860 5234
rect 12808 5170 12860 5176
rect 12728 5086 12940 5114
rect 12452 4576 12572 4604
rect 11980 4480 12032 4486
rect 11980 4422 12032 4428
rect 11888 4208 11940 4214
rect 11888 4150 11940 4156
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 11610 3496 11666 3505
rect 11256 3194 11284 3470
rect 11610 3431 11612 3440
rect 11664 3431 11666 3440
rect 11612 3402 11664 3408
rect 11352 3292 11648 3312
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11430 3238 11432 3290
rect 11494 3238 11506 3290
rect 11568 3238 11570 3290
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11352 3216 11648 3236
rect 11244 3188 11296 3194
rect 11244 3130 11296 3136
rect 11152 2984 11204 2990
rect 11150 2952 11152 2961
rect 11204 2952 11206 2961
rect 11150 2887 11206 2896
rect 11352 2204 11648 2224
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11430 2150 11432 2202
rect 11494 2150 11506 2202
rect 11568 2150 11570 2202
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11352 2128 11648 2148
rect 11900 800 11928 4150
rect 11992 2514 12020 4422
rect 12254 4312 12310 4321
rect 12452 4282 12480 4576
rect 12532 4480 12584 4486
rect 12532 4422 12584 4428
rect 12716 4480 12768 4486
rect 12716 4422 12768 4428
rect 12254 4247 12256 4256
rect 12308 4247 12310 4256
rect 12440 4276 12492 4282
rect 12256 4218 12308 4224
rect 12440 4218 12492 4224
rect 12452 4185 12480 4218
rect 12438 4176 12494 4185
rect 12438 4111 12494 4120
rect 12544 4010 12572 4422
rect 12728 4282 12756 4422
rect 12716 4276 12768 4282
rect 12636 4236 12716 4264
rect 12532 4004 12584 4010
rect 12532 3946 12584 3952
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 12268 2990 12296 3538
rect 12348 3460 12400 3466
rect 12348 3402 12400 3408
rect 12360 3058 12388 3402
rect 12544 3194 12572 3946
rect 12636 3602 12664 4236
rect 12716 4218 12768 4224
rect 12912 4162 12940 5086
rect 12728 4134 12940 4162
rect 12624 3596 12676 3602
rect 12624 3538 12676 3544
rect 12532 3188 12584 3194
rect 12532 3130 12584 3136
rect 12348 3052 12400 3058
rect 12348 2994 12400 3000
rect 12256 2984 12308 2990
rect 12256 2926 12308 2932
rect 12360 2650 12388 2994
rect 12348 2644 12400 2650
rect 12348 2586 12400 2592
rect 11980 2508 12032 2514
rect 11980 2450 12032 2456
rect 12728 800 12756 4134
rect 12808 3596 12860 3602
rect 12808 3538 12860 3544
rect 12900 3596 12952 3602
rect 12900 3538 12952 3544
rect 12820 3058 12848 3538
rect 12912 3398 12940 3538
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 12912 3233 12940 3334
rect 12898 3224 12954 3233
rect 12898 3159 12954 3168
rect 12808 3052 12860 3058
rect 12808 2994 12860 3000
rect 12912 2650 12940 3159
rect 13004 2825 13032 5630
rect 13084 4548 13136 4554
rect 13084 4490 13136 4496
rect 12990 2816 13046 2825
rect 12990 2751 13046 2760
rect 12900 2644 12952 2650
rect 12900 2586 12952 2592
rect 13096 2446 13124 4490
rect 13188 4078 13216 6054
rect 13372 4486 13400 7414
rect 13464 6225 13492 8298
rect 13556 7410 13584 8452
rect 13648 7750 13676 8910
rect 13740 8294 13768 8978
rect 13832 8838 13860 10202
rect 14292 9722 14320 10610
rect 14384 10130 14412 14010
rect 14752 13938 14780 14010
rect 14740 13932 14792 13938
rect 14740 13874 14792 13880
rect 14740 13796 14792 13802
rect 14740 13738 14792 13744
rect 14752 13530 14780 13738
rect 14740 13524 14792 13530
rect 14740 13466 14792 13472
rect 14844 13410 14872 14214
rect 15292 14068 15344 14074
rect 15292 14010 15344 14016
rect 14924 14000 14976 14006
rect 14924 13942 14976 13948
rect 14936 13530 14964 13942
rect 14924 13524 14976 13530
rect 14924 13466 14976 13472
rect 14660 13394 14872 13410
rect 14648 13388 14872 13394
rect 14700 13382 14872 13388
rect 14924 13388 14976 13394
rect 14648 13330 14700 13336
rect 14924 13330 14976 13336
rect 14832 13320 14884 13326
rect 14752 13280 14832 13308
rect 14464 12980 14516 12986
rect 14464 12922 14516 12928
rect 14476 12102 14504 12922
rect 14752 12782 14780 13280
rect 14832 13262 14884 13268
rect 14936 12986 14964 13330
rect 14924 12980 14976 12986
rect 14924 12922 14976 12928
rect 15304 12782 15332 14010
rect 15948 13938 15976 14214
rect 15936 13932 15988 13938
rect 15936 13874 15988 13880
rect 15568 13864 15620 13870
rect 15568 13806 15620 13812
rect 15580 13326 15608 13806
rect 16028 13388 16080 13394
rect 16028 13330 16080 13336
rect 15568 13320 15620 13326
rect 15568 13262 15620 13268
rect 14740 12776 14792 12782
rect 14740 12718 14792 12724
rect 15292 12776 15344 12782
rect 16040 12753 16068 13330
rect 15292 12718 15344 12724
rect 16026 12744 16082 12753
rect 15200 12708 15252 12714
rect 16026 12679 16082 12688
rect 15200 12650 15252 12656
rect 15212 12374 15240 12650
rect 16040 12646 16068 12679
rect 15476 12640 15528 12646
rect 15476 12582 15528 12588
rect 16028 12640 16080 12646
rect 16028 12582 16080 12588
rect 15488 12442 15516 12582
rect 15476 12436 15528 12442
rect 15476 12378 15528 12384
rect 15200 12368 15252 12374
rect 15200 12310 15252 12316
rect 15660 12300 15712 12306
rect 15660 12242 15712 12248
rect 14924 12232 14976 12238
rect 14924 12174 14976 12180
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14476 11898 14504 12038
rect 14464 11892 14516 11898
rect 14464 11834 14516 11840
rect 14464 11688 14516 11694
rect 14464 11630 14516 11636
rect 14476 11558 14504 11630
rect 14464 11552 14516 11558
rect 14464 11494 14516 11500
rect 14936 11286 14964 12174
rect 15672 11898 15700 12242
rect 15660 11892 15712 11898
rect 15660 11834 15712 11840
rect 15844 11824 15896 11830
rect 15212 11750 15424 11778
rect 15844 11766 15896 11772
rect 15212 11694 15240 11750
rect 15200 11688 15252 11694
rect 15200 11630 15252 11636
rect 15292 11620 15344 11626
rect 15292 11562 15344 11568
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 15120 11354 15148 11494
rect 15108 11348 15160 11354
rect 15108 11290 15160 11296
rect 14924 11280 14976 11286
rect 14924 11222 14976 11228
rect 14936 10674 14964 11222
rect 14924 10668 14976 10674
rect 14924 10610 14976 10616
rect 14936 10266 14964 10610
rect 15120 10606 15148 11290
rect 15304 11286 15332 11562
rect 15292 11280 15344 11286
rect 15292 11222 15344 11228
rect 15200 11008 15252 11014
rect 15200 10950 15252 10956
rect 15108 10600 15160 10606
rect 15108 10542 15160 10548
rect 15212 10538 15240 10950
rect 15304 10810 15332 11222
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 15200 10532 15252 10538
rect 15200 10474 15252 10480
rect 14924 10260 14976 10266
rect 14924 10202 14976 10208
rect 15108 10192 15160 10198
rect 15108 10134 15160 10140
rect 14372 10124 14424 10130
rect 14372 10066 14424 10072
rect 14280 9716 14332 9722
rect 14280 9658 14332 9664
rect 14292 9518 14320 9658
rect 14280 9512 14332 9518
rect 14280 9454 14332 9460
rect 14740 9512 14792 9518
rect 14740 9454 14792 9460
rect 14004 8900 14056 8906
rect 14004 8842 14056 8848
rect 13820 8832 13872 8838
rect 13820 8774 13872 8780
rect 14016 8430 14044 8842
rect 14004 8424 14056 8430
rect 14004 8366 14056 8372
rect 13728 8288 13780 8294
rect 13728 8230 13780 8236
rect 14188 7948 14240 7954
rect 14188 7890 14240 7896
rect 13912 7880 13964 7886
rect 13912 7822 13964 7828
rect 13636 7744 13688 7750
rect 13636 7686 13688 7692
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 13636 6996 13688 7002
rect 13636 6938 13688 6944
rect 13450 6216 13506 6225
rect 13450 6151 13506 6160
rect 13544 6180 13596 6186
rect 13544 6122 13596 6128
rect 13360 4480 13412 4486
rect 13360 4422 13412 4428
rect 13372 4146 13400 4422
rect 13556 4185 13584 6122
rect 13648 5778 13676 6938
rect 13820 6860 13872 6866
rect 13820 6802 13872 6808
rect 13832 6118 13860 6802
rect 13924 6798 13952 7822
rect 14200 7342 14228 7890
rect 14464 7744 14516 7750
rect 14464 7686 14516 7692
rect 14476 7342 14504 7686
rect 14188 7336 14240 7342
rect 14188 7278 14240 7284
rect 14464 7336 14516 7342
rect 14464 7278 14516 7284
rect 13912 6792 13964 6798
rect 13912 6734 13964 6740
rect 13924 6458 13952 6734
rect 14200 6662 14228 7278
rect 14752 6934 14780 9454
rect 15120 8634 15148 10134
rect 15200 9920 15252 9926
rect 15200 9862 15252 9868
rect 15212 9518 15240 9862
rect 15200 9512 15252 9518
rect 15200 9454 15252 9460
rect 15200 8832 15252 8838
rect 15200 8774 15252 8780
rect 15108 8628 15160 8634
rect 15108 8570 15160 8576
rect 15016 8492 15068 8498
rect 15016 8434 15068 8440
rect 15028 7954 15056 8434
rect 15120 8430 15148 8570
rect 15212 8430 15240 8774
rect 15108 8424 15160 8430
rect 15108 8366 15160 8372
rect 15200 8424 15252 8430
rect 15200 8366 15252 8372
rect 15016 7948 15068 7954
rect 15016 7890 15068 7896
rect 15290 7712 15346 7721
rect 15290 7647 15346 7656
rect 15304 7410 15332 7647
rect 15292 7404 15344 7410
rect 15292 7346 15344 7352
rect 14740 6928 14792 6934
rect 14740 6870 14792 6876
rect 14372 6860 14424 6866
rect 14372 6802 14424 6808
rect 14188 6656 14240 6662
rect 14188 6598 14240 6604
rect 13912 6452 13964 6458
rect 13912 6394 13964 6400
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13636 5772 13688 5778
rect 13636 5714 13688 5720
rect 13648 5098 13676 5714
rect 14096 5636 14148 5642
rect 14096 5578 14148 5584
rect 14108 5370 14136 5578
rect 14096 5364 14148 5370
rect 14096 5306 14148 5312
rect 13636 5092 13688 5098
rect 13636 5034 13688 5040
rect 13912 4684 13964 4690
rect 13912 4626 13964 4632
rect 13636 4480 13688 4486
rect 13636 4422 13688 4428
rect 13542 4176 13598 4185
rect 13360 4140 13412 4146
rect 13542 4111 13598 4120
rect 13360 4082 13412 4088
rect 13176 4072 13228 4078
rect 13228 4020 13492 4026
rect 13176 4014 13492 4020
rect 13188 3998 13492 4014
rect 13464 3942 13492 3998
rect 13452 3936 13504 3942
rect 13452 3878 13504 3884
rect 13556 3890 13584 4111
rect 13648 4010 13676 4422
rect 13924 4282 13952 4626
rect 14096 4616 14148 4622
rect 14096 4558 14148 4564
rect 13912 4276 13964 4282
rect 13912 4218 13964 4224
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 13636 4004 13688 4010
rect 13636 3946 13688 3952
rect 13556 3862 13676 3890
rect 13358 3768 13414 3777
rect 13358 3703 13414 3712
rect 13268 3392 13320 3398
rect 13268 3334 13320 3340
rect 13280 3126 13308 3334
rect 13268 3120 13320 3126
rect 13268 3062 13320 3068
rect 13372 2650 13400 3703
rect 13452 3528 13504 3534
rect 13452 3470 13504 3476
rect 13464 2922 13492 3470
rect 13452 2916 13504 2922
rect 13452 2858 13504 2864
rect 13360 2644 13412 2650
rect 13360 2586 13412 2592
rect 13084 2440 13136 2446
rect 13084 2382 13136 2388
rect 13648 800 13676 3862
rect 13740 3058 13768 4082
rect 14108 3738 14136 4558
rect 14200 4078 14228 6598
rect 14384 6322 14412 6802
rect 14372 6316 14424 6322
rect 14372 6258 14424 6264
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 14660 5166 14688 6054
rect 14556 5160 14608 5166
rect 14556 5102 14608 5108
rect 14648 5160 14700 5166
rect 14648 5102 14700 5108
rect 14188 4072 14240 4078
rect 14188 4014 14240 4020
rect 14372 4072 14424 4078
rect 14372 4014 14424 4020
rect 14464 4072 14516 4078
rect 14464 4014 14516 4020
rect 14096 3732 14148 3738
rect 14096 3674 14148 3680
rect 14108 3466 14136 3674
rect 14096 3460 14148 3466
rect 14096 3402 14148 3408
rect 13820 3392 13872 3398
rect 13818 3360 13820 3369
rect 13872 3360 13874 3369
rect 13818 3295 13874 3304
rect 13832 3126 13860 3295
rect 13820 3120 13872 3126
rect 13820 3062 13872 3068
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 14108 2922 14136 3402
rect 14384 3398 14412 4014
rect 14372 3392 14424 3398
rect 14372 3334 14424 3340
rect 14476 3194 14504 4014
rect 14464 3188 14516 3194
rect 14464 3130 14516 3136
rect 14096 2916 14148 2922
rect 14096 2858 14148 2864
rect 14476 2514 14504 3130
rect 14568 2854 14596 5102
rect 14752 4690 14780 6870
rect 15200 6792 15252 6798
rect 15200 6734 15252 6740
rect 15016 6248 15068 6254
rect 15016 6190 15068 6196
rect 15028 6118 15056 6190
rect 15212 6186 15240 6734
rect 15200 6180 15252 6186
rect 15200 6122 15252 6128
rect 15016 6112 15068 6118
rect 15016 6054 15068 6060
rect 15028 5778 15056 6054
rect 15016 5772 15068 5778
rect 15016 5714 15068 5720
rect 14924 5636 14976 5642
rect 14924 5578 14976 5584
rect 14936 4826 14964 5578
rect 15028 5370 15056 5714
rect 15108 5568 15160 5574
rect 15108 5510 15160 5516
rect 15016 5364 15068 5370
rect 15016 5306 15068 5312
rect 14924 4820 14976 4826
rect 14924 4762 14976 4768
rect 14740 4684 14792 4690
rect 14740 4626 14792 4632
rect 14936 4214 14964 4762
rect 14832 4208 14884 4214
rect 14832 4150 14884 4156
rect 14924 4208 14976 4214
rect 14924 4150 14976 4156
rect 14844 3913 14872 4150
rect 15120 3942 15148 5510
rect 15200 4480 15252 4486
rect 15200 4422 15252 4428
rect 15212 4078 15240 4422
rect 15200 4072 15252 4078
rect 15200 4014 15252 4020
rect 15108 3936 15160 3942
rect 14830 3904 14886 3913
rect 15108 3878 15160 3884
rect 14830 3839 14886 3848
rect 15016 3528 15068 3534
rect 15016 3470 15068 3476
rect 15028 2990 15056 3470
rect 15016 2984 15068 2990
rect 15016 2926 15068 2932
rect 15200 2916 15252 2922
rect 15200 2858 15252 2864
rect 14556 2848 14608 2854
rect 14556 2790 14608 2796
rect 14464 2508 14516 2514
rect 14464 2450 14516 2456
rect 14568 800 14596 2790
rect 15212 2650 15240 2858
rect 15200 2644 15252 2650
rect 15200 2586 15252 2592
rect 15212 2106 15240 2586
rect 15304 2514 15332 7346
rect 15396 4570 15424 11750
rect 15856 11150 15884 11766
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 15476 11008 15528 11014
rect 15476 10950 15528 10956
rect 15568 11008 15620 11014
rect 15568 10950 15620 10956
rect 15488 10266 15516 10950
rect 15580 10538 15608 10950
rect 15856 10742 15884 11086
rect 15844 10736 15896 10742
rect 15844 10678 15896 10684
rect 15568 10532 15620 10538
rect 15568 10474 15620 10480
rect 15476 10260 15528 10266
rect 15476 10202 15528 10208
rect 15488 8838 15516 10202
rect 15580 9994 15608 10474
rect 16040 10130 16068 12582
rect 16132 11286 16160 15370
rect 16776 15366 16804 16050
rect 16856 15428 16908 15434
rect 16856 15370 16908 15376
rect 16764 15360 16816 15366
rect 16764 15302 16816 15308
rect 16868 14822 16896 15370
rect 17052 15094 17080 16050
rect 17144 16046 17172 16730
rect 18052 16652 18104 16658
rect 18052 16594 18104 16600
rect 18064 16250 18092 16594
rect 18052 16244 18104 16250
rect 18052 16186 18104 16192
rect 18064 16114 18092 16186
rect 18052 16108 18104 16114
rect 18052 16050 18104 16056
rect 17132 16040 17184 16046
rect 17132 15982 17184 15988
rect 18340 15638 18368 17002
rect 18512 16584 18564 16590
rect 18512 16526 18564 16532
rect 18524 15638 18552 16526
rect 19168 16046 19196 17206
rect 19248 17060 19300 17066
rect 19248 17002 19300 17008
rect 19260 16794 19288 17002
rect 20444 16992 20496 16998
rect 20444 16934 20496 16940
rect 19248 16788 19300 16794
rect 19248 16730 19300 16736
rect 19984 16584 20036 16590
rect 19984 16526 20036 16532
rect 19996 16250 20024 16526
rect 20352 16448 20404 16454
rect 20352 16390 20404 16396
rect 19984 16244 20036 16250
rect 19984 16186 20036 16192
rect 19800 16176 19852 16182
rect 19800 16118 19852 16124
rect 19156 16040 19208 16046
rect 19156 15982 19208 15988
rect 19168 15706 19196 15982
rect 19156 15700 19208 15706
rect 19156 15642 19208 15648
rect 18328 15632 18380 15638
rect 18328 15574 18380 15580
rect 18512 15632 18564 15638
rect 18512 15574 18564 15580
rect 19812 15570 19840 16118
rect 20364 16046 20392 16390
rect 20352 16040 20404 16046
rect 20352 15982 20404 15988
rect 19340 15564 19392 15570
rect 19340 15506 19392 15512
rect 19524 15564 19576 15570
rect 19524 15506 19576 15512
rect 19800 15564 19852 15570
rect 19800 15506 19852 15512
rect 18144 15428 18196 15434
rect 18144 15370 18196 15376
rect 17868 15360 17920 15366
rect 17868 15302 17920 15308
rect 17040 15088 17092 15094
rect 17040 15030 17092 15036
rect 17880 14958 17908 15302
rect 18156 15094 18184 15370
rect 18144 15088 18196 15094
rect 18144 15030 18196 15036
rect 17868 14952 17920 14958
rect 17868 14894 17920 14900
rect 18328 14952 18380 14958
rect 18328 14894 18380 14900
rect 17880 14822 17908 14894
rect 16856 14816 16908 14822
rect 16856 14758 16908 14764
rect 17868 14816 17920 14822
rect 17868 14758 17920 14764
rect 16868 14414 16896 14758
rect 16856 14408 16908 14414
rect 16856 14350 16908 14356
rect 17132 14408 17184 14414
rect 17132 14350 17184 14356
rect 16396 14340 16448 14346
rect 16396 14282 16448 14288
rect 16408 14074 16436 14282
rect 16580 14272 16632 14278
rect 16580 14214 16632 14220
rect 16764 14272 16816 14278
rect 16764 14214 16816 14220
rect 16396 14068 16448 14074
rect 16396 14010 16448 14016
rect 16212 13864 16264 13870
rect 16212 13806 16264 13812
rect 16224 12306 16252 13806
rect 16592 13394 16620 14214
rect 16776 13870 16804 14214
rect 16764 13864 16816 13870
rect 16764 13806 16816 13812
rect 16868 13530 16896 14350
rect 17038 13968 17094 13977
rect 17144 13938 17172 14350
rect 18340 14278 18368 14894
rect 18880 14884 18932 14890
rect 18880 14826 18932 14832
rect 18892 14618 18920 14826
rect 18880 14612 18932 14618
rect 18880 14554 18932 14560
rect 18328 14272 18380 14278
rect 18328 14214 18380 14220
rect 17222 14104 17278 14113
rect 17222 14039 17278 14048
rect 17038 13903 17040 13912
rect 17092 13903 17094 13912
rect 17132 13932 17184 13938
rect 17040 13874 17092 13880
rect 17132 13874 17184 13880
rect 17236 13682 17264 14039
rect 17684 14000 17736 14006
rect 17684 13942 17736 13948
rect 18696 14000 18748 14006
rect 18696 13942 18748 13948
rect 17052 13654 17264 13682
rect 17408 13728 17460 13734
rect 17408 13670 17460 13676
rect 16856 13524 16908 13530
rect 16856 13466 16908 13472
rect 16580 13388 16632 13394
rect 16580 13330 16632 13336
rect 17052 13190 17080 13654
rect 17222 13560 17278 13569
rect 17222 13495 17278 13504
rect 17040 13184 17092 13190
rect 17236 13161 17264 13495
rect 17420 13394 17448 13670
rect 17592 13456 17644 13462
rect 17592 13398 17644 13404
rect 17408 13388 17460 13394
rect 17408 13330 17460 13336
rect 17316 13320 17368 13326
rect 17316 13262 17368 13268
rect 17040 13126 17092 13132
rect 17222 13152 17278 13161
rect 16948 12776 17000 12782
rect 17052 12730 17080 13126
rect 17222 13087 17278 13096
rect 17000 12724 17080 12730
rect 16948 12718 17080 12724
rect 16960 12702 17080 12718
rect 16948 12640 17000 12646
rect 16948 12582 17000 12588
rect 16304 12436 16356 12442
rect 16304 12378 16356 12384
rect 16212 12300 16264 12306
rect 16212 12242 16264 12248
rect 16120 11280 16172 11286
rect 16120 11222 16172 11228
rect 16212 11212 16264 11218
rect 16212 11154 16264 11160
rect 16224 11014 16252 11154
rect 16316 11014 16344 12378
rect 16854 12336 16910 12345
rect 16672 12300 16724 12306
rect 16854 12271 16856 12280
rect 16672 12242 16724 12248
rect 16908 12271 16910 12280
rect 16856 12242 16908 12248
rect 16396 11688 16448 11694
rect 16396 11630 16448 11636
rect 16408 11558 16436 11630
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 16212 11008 16264 11014
rect 16212 10950 16264 10956
rect 16304 11008 16356 11014
rect 16304 10950 16356 10956
rect 16224 10742 16252 10950
rect 16212 10736 16264 10742
rect 16212 10678 16264 10684
rect 16028 10124 16080 10130
rect 16028 10066 16080 10072
rect 15568 9988 15620 9994
rect 15568 9930 15620 9936
rect 16040 9722 16068 10066
rect 16316 9926 16344 10950
rect 16408 10266 16436 11494
rect 16684 11150 16712 12242
rect 16868 11898 16896 12242
rect 16856 11892 16908 11898
rect 16856 11834 16908 11840
rect 16868 11286 16896 11834
rect 16856 11280 16908 11286
rect 16856 11222 16908 11228
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 16396 10260 16448 10266
rect 16396 10202 16448 10208
rect 16304 9920 16356 9926
rect 16304 9862 16356 9868
rect 16672 9920 16724 9926
rect 16672 9862 16724 9868
rect 16028 9716 16080 9722
rect 16028 9658 16080 9664
rect 16316 9625 16344 9862
rect 16302 9616 16358 9625
rect 16302 9551 16358 9560
rect 16396 9580 16448 9586
rect 16396 9522 16448 9528
rect 16028 9512 16080 9518
rect 16028 9454 16080 9460
rect 16040 9042 16068 9454
rect 15936 9036 15988 9042
rect 15936 8978 15988 8984
rect 16028 9036 16080 9042
rect 16028 8978 16080 8984
rect 15476 8832 15528 8838
rect 15476 8774 15528 8780
rect 15948 8634 15976 8978
rect 16408 8974 16436 9522
rect 16684 9518 16712 9862
rect 16960 9586 16988 12582
rect 17052 11354 17080 12702
rect 17328 12374 17356 13262
rect 17420 12986 17448 13330
rect 17408 12980 17460 12986
rect 17408 12922 17460 12928
rect 17500 12776 17552 12782
rect 17500 12718 17552 12724
rect 17316 12368 17368 12374
rect 17316 12310 17368 12316
rect 17314 12200 17370 12209
rect 17314 12135 17370 12144
rect 17328 12102 17356 12135
rect 17512 12102 17540 12718
rect 17604 12458 17632 13398
rect 17696 13394 17724 13942
rect 18708 13870 18736 13942
rect 18236 13864 18288 13870
rect 18236 13806 18288 13812
rect 18604 13864 18656 13870
rect 18604 13806 18656 13812
rect 18696 13864 18748 13870
rect 18696 13806 18748 13812
rect 17868 13728 17920 13734
rect 17868 13670 17920 13676
rect 17880 13462 17908 13670
rect 18248 13530 18276 13806
rect 18236 13524 18288 13530
rect 18236 13466 18288 13472
rect 17868 13456 17920 13462
rect 17868 13398 17920 13404
rect 17684 13388 17736 13394
rect 17684 13330 17736 13336
rect 17696 12646 17724 13330
rect 18248 12782 18276 13466
rect 18616 13190 18644 13806
rect 18604 13184 18656 13190
rect 18604 13126 18656 13132
rect 18236 12776 18288 12782
rect 18236 12718 18288 12724
rect 18328 12776 18380 12782
rect 18328 12718 18380 12724
rect 17684 12640 17736 12646
rect 17684 12582 17736 12588
rect 17774 12472 17830 12481
rect 17604 12430 17774 12458
rect 17774 12407 17776 12416
rect 17828 12407 17830 12416
rect 17776 12378 17828 12384
rect 18340 12170 18368 12718
rect 18328 12164 18380 12170
rect 18328 12106 18380 12112
rect 18420 12164 18472 12170
rect 18420 12106 18472 12112
rect 17316 12096 17368 12102
rect 17316 12038 17368 12044
rect 17500 12096 17552 12102
rect 17500 12038 17552 12044
rect 17684 12096 17736 12102
rect 17684 12038 17736 12044
rect 17512 11898 17540 12038
rect 17500 11892 17552 11898
rect 17500 11834 17552 11840
rect 17592 11892 17644 11898
rect 17592 11834 17644 11840
rect 17040 11348 17092 11354
rect 17040 11290 17092 11296
rect 17604 11082 17632 11834
rect 17696 11218 17724 12038
rect 18340 11937 18368 12106
rect 18326 11928 18382 11937
rect 18326 11863 18382 11872
rect 17960 11688 18012 11694
rect 17960 11630 18012 11636
rect 18328 11688 18380 11694
rect 18328 11630 18380 11636
rect 17776 11552 17828 11558
rect 17776 11494 17828 11500
rect 17788 11218 17816 11494
rect 17684 11212 17736 11218
rect 17684 11154 17736 11160
rect 17776 11212 17828 11218
rect 17776 11154 17828 11160
rect 17592 11076 17644 11082
rect 17592 11018 17644 11024
rect 17788 10470 17816 11154
rect 17868 11144 17920 11150
rect 17868 11086 17920 11092
rect 17880 10742 17908 11086
rect 17972 11014 18000 11630
rect 18052 11620 18104 11626
rect 18236 11620 18288 11626
rect 18104 11580 18236 11608
rect 18052 11562 18104 11568
rect 18236 11562 18288 11568
rect 18340 11082 18368 11630
rect 18328 11076 18380 11082
rect 18328 11018 18380 11024
rect 17960 11008 18012 11014
rect 17960 10950 18012 10956
rect 18328 10804 18380 10810
rect 18328 10746 18380 10752
rect 17868 10736 17920 10742
rect 17868 10678 17920 10684
rect 18236 10532 18288 10538
rect 18236 10474 18288 10480
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17776 10464 17828 10470
rect 17776 10406 17828 10412
rect 17420 10130 17448 10406
rect 18248 10198 18276 10474
rect 18236 10192 18288 10198
rect 18236 10134 18288 10140
rect 18340 10130 18368 10746
rect 17408 10124 17460 10130
rect 17408 10066 17460 10072
rect 17776 10124 17828 10130
rect 17776 10066 17828 10072
rect 18328 10124 18380 10130
rect 18328 10066 18380 10072
rect 17592 9988 17644 9994
rect 17592 9930 17644 9936
rect 16948 9580 17000 9586
rect 16948 9522 17000 9528
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 17224 9444 17276 9450
rect 17224 9386 17276 9392
rect 17236 9178 17264 9386
rect 17604 9382 17632 9930
rect 17788 9926 17816 10066
rect 17960 10056 18012 10062
rect 17960 9998 18012 10004
rect 17776 9920 17828 9926
rect 17776 9862 17828 9868
rect 17592 9376 17644 9382
rect 17592 9318 17644 9324
rect 17224 9172 17276 9178
rect 17224 9114 17276 9120
rect 16764 9036 16816 9042
rect 16764 8978 16816 8984
rect 17316 9036 17368 9042
rect 17368 8996 17448 9024
rect 17316 8978 17368 8984
rect 16120 8968 16172 8974
rect 16120 8910 16172 8916
rect 16396 8968 16448 8974
rect 16396 8910 16448 8916
rect 16132 8838 16160 8910
rect 16776 8838 16804 8978
rect 17224 8968 17276 8974
rect 17224 8910 17276 8916
rect 16120 8832 16172 8838
rect 16120 8774 16172 8780
rect 16764 8832 16816 8838
rect 16764 8774 16816 8780
rect 16856 8832 16908 8838
rect 16856 8774 16908 8780
rect 15936 8628 15988 8634
rect 15936 8570 15988 8576
rect 15752 8424 15804 8430
rect 15752 8366 15804 8372
rect 15764 7818 15792 8366
rect 15948 8362 15976 8570
rect 16132 8498 16160 8774
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 16776 8430 16804 8774
rect 16764 8424 16816 8430
rect 16764 8366 16816 8372
rect 15936 8356 15988 8362
rect 15936 8298 15988 8304
rect 16580 8288 16632 8294
rect 16580 8230 16632 8236
rect 16592 7954 16620 8230
rect 16580 7948 16632 7954
rect 16580 7890 16632 7896
rect 16212 7880 16264 7886
rect 16212 7822 16264 7828
rect 15752 7812 15804 7818
rect 15752 7754 15804 7760
rect 15764 7410 15792 7754
rect 15752 7404 15804 7410
rect 15752 7346 15804 7352
rect 16224 7206 16252 7822
rect 16304 7336 16356 7342
rect 16304 7278 16356 7284
rect 16212 7200 16264 7206
rect 16212 7142 16264 7148
rect 16224 6866 16252 7142
rect 16316 6934 16344 7278
rect 16304 6928 16356 6934
rect 16304 6870 16356 6876
rect 15660 6860 15712 6866
rect 16212 6860 16264 6866
rect 15712 6820 15884 6848
rect 15660 6802 15712 6808
rect 15752 6248 15804 6254
rect 15752 6190 15804 6196
rect 15658 5400 15714 5409
rect 15658 5335 15714 5344
rect 15568 5160 15620 5166
rect 15568 5102 15620 5108
rect 15580 4826 15608 5102
rect 15568 4820 15620 4826
rect 15568 4762 15620 4768
rect 15474 4584 15530 4593
rect 15396 4542 15474 4570
rect 15474 4519 15530 4528
rect 15488 4486 15516 4519
rect 15476 4480 15528 4486
rect 15476 4422 15528 4428
rect 15672 4128 15700 5335
rect 15764 5030 15792 6190
rect 15856 5302 15884 6820
rect 16212 6802 16264 6808
rect 15936 6724 15988 6730
rect 15936 6666 15988 6672
rect 15948 6186 15976 6666
rect 16224 6662 16252 6802
rect 16120 6656 16172 6662
rect 16120 6598 16172 6604
rect 16212 6656 16264 6662
rect 16212 6598 16264 6604
rect 16028 6384 16080 6390
rect 16028 6326 16080 6332
rect 15936 6180 15988 6186
rect 15936 6122 15988 6128
rect 15936 5636 15988 5642
rect 15936 5578 15988 5584
rect 15844 5296 15896 5302
rect 15844 5238 15896 5244
rect 15948 5166 15976 5578
rect 16040 5166 16068 6326
rect 16132 6254 16160 6598
rect 16304 6384 16356 6390
rect 16304 6326 16356 6332
rect 16120 6248 16172 6254
rect 16120 6190 16172 6196
rect 16120 6112 16172 6118
rect 16120 6054 16172 6060
rect 16132 5778 16160 6054
rect 16316 5778 16344 6326
rect 16120 5772 16172 5778
rect 16120 5714 16172 5720
rect 16304 5772 16356 5778
rect 16304 5714 16356 5720
rect 15936 5160 15988 5166
rect 15936 5102 15988 5108
rect 16028 5160 16080 5166
rect 16028 5102 16080 5108
rect 15752 5024 15804 5030
rect 15752 4966 15804 4972
rect 16132 4486 16160 5714
rect 16210 5536 16266 5545
rect 16210 5471 16266 5480
rect 16224 4622 16252 5471
rect 16316 5370 16344 5714
rect 16592 5710 16620 7890
rect 16672 7744 16724 7750
rect 16672 7686 16724 7692
rect 16684 7342 16712 7686
rect 16776 7546 16804 8366
rect 16868 7721 16896 8774
rect 17236 8616 17264 8910
rect 17420 8838 17448 8996
rect 17500 8968 17552 8974
rect 17498 8936 17500 8945
rect 17552 8936 17554 8945
rect 17498 8871 17554 8880
rect 17408 8832 17460 8838
rect 17408 8774 17460 8780
rect 17236 8588 17356 8616
rect 17222 8528 17278 8537
rect 17222 8463 17278 8472
rect 17236 8430 17264 8463
rect 17224 8424 17276 8430
rect 17224 8366 17276 8372
rect 17328 8090 17356 8588
rect 17500 8492 17552 8498
rect 17500 8434 17552 8440
rect 17408 8356 17460 8362
rect 17408 8298 17460 8304
rect 17224 8084 17276 8090
rect 17224 8026 17276 8032
rect 17316 8084 17368 8090
rect 17316 8026 17368 8032
rect 16948 7948 17000 7954
rect 16948 7890 17000 7896
rect 16854 7712 16910 7721
rect 16854 7647 16910 7656
rect 16960 7585 16988 7890
rect 16946 7576 17002 7585
rect 16764 7540 16816 7546
rect 16946 7511 17002 7520
rect 16764 7482 16816 7488
rect 17236 7410 17264 8026
rect 17224 7404 17276 7410
rect 17224 7346 17276 7352
rect 16672 7336 16724 7342
rect 16672 7278 16724 7284
rect 17224 6860 17276 6866
rect 17224 6802 17276 6808
rect 17040 6792 17092 6798
rect 17040 6734 17092 6740
rect 17132 6792 17184 6798
rect 17132 6734 17184 6740
rect 16762 6488 16818 6497
rect 16762 6423 16818 6432
rect 16776 6254 16804 6423
rect 16764 6248 16816 6254
rect 16764 6190 16816 6196
rect 16776 5914 16804 6190
rect 17052 5914 17080 6734
rect 17144 6662 17172 6734
rect 17236 6662 17264 6802
rect 17132 6656 17184 6662
rect 17132 6598 17184 6604
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 17132 6112 17184 6118
rect 17132 6054 17184 6060
rect 16764 5908 16816 5914
rect 16764 5850 16816 5856
rect 17040 5908 17092 5914
rect 17040 5850 17092 5856
rect 16580 5704 16632 5710
rect 16580 5646 16632 5652
rect 16304 5364 16356 5370
rect 16304 5306 16356 5312
rect 16578 4856 16634 4865
rect 16578 4791 16634 4800
rect 16592 4690 16620 4791
rect 16580 4684 16632 4690
rect 16580 4626 16632 4632
rect 16672 4684 16724 4690
rect 16672 4626 16724 4632
rect 16212 4616 16264 4622
rect 16212 4558 16264 4564
rect 16120 4480 16172 4486
rect 16120 4422 16172 4428
rect 15488 4100 15700 4128
rect 15384 2916 15436 2922
rect 15384 2858 15436 2864
rect 15292 2508 15344 2514
rect 15292 2450 15344 2456
rect 15200 2100 15252 2106
rect 15200 2042 15252 2048
rect 15304 1970 15332 2450
rect 15396 2378 15424 2858
rect 15384 2372 15436 2378
rect 15384 2314 15436 2320
rect 15488 2258 15516 4100
rect 15660 4004 15712 4010
rect 15660 3946 15712 3952
rect 15936 4004 15988 4010
rect 15936 3946 15988 3952
rect 15672 3602 15700 3946
rect 15660 3596 15712 3602
rect 15660 3538 15712 3544
rect 15672 3194 15700 3538
rect 15948 3534 15976 3946
rect 16224 3602 16252 4558
rect 16592 4282 16620 4626
rect 16684 4554 16712 4626
rect 16672 4548 16724 4554
rect 16672 4490 16724 4496
rect 16684 4282 16712 4490
rect 16580 4276 16632 4282
rect 16580 4218 16632 4224
rect 16672 4276 16724 4282
rect 16672 4218 16724 4224
rect 16488 3936 16540 3942
rect 16486 3904 16488 3913
rect 16580 3936 16632 3942
rect 16540 3904 16542 3913
rect 16580 3878 16632 3884
rect 16486 3839 16542 3848
rect 16592 3738 16620 3878
rect 16580 3732 16632 3738
rect 16580 3674 16632 3680
rect 16212 3596 16264 3602
rect 16212 3538 16264 3544
rect 15936 3528 15988 3534
rect 15936 3470 15988 3476
rect 15948 3398 15976 3470
rect 15936 3392 15988 3398
rect 15936 3334 15988 3340
rect 16120 3392 16172 3398
rect 16120 3334 16172 3340
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 15948 2990 15976 3334
rect 16132 2990 16160 3334
rect 16224 3126 16252 3538
rect 16212 3120 16264 3126
rect 16212 3062 16264 3068
rect 15936 2984 15988 2990
rect 15934 2952 15936 2961
rect 16120 2984 16172 2990
rect 15988 2952 15990 2961
rect 16120 2926 16172 2932
rect 16396 2984 16448 2990
rect 16396 2926 16448 2932
rect 15934 2887 15990 2896
rect 16408 2650 16436 2926
rect 16396 2644 16448 2650
rect 16396 2586 16448 2592
rect 15752 2508 15804 2514
rect 15752 2450 15804 2456
rect 15396 2230 15516 2258
rect 15292 1964 15344 1970
rect 15292 1906 15344 1912
rect 15396 800 15424 2230
rect 15764 2106 15792 2450
rect 15752 2100 15804 2106
rect 15752 2042 15804 2048
rect 16304 1896 16356 1902
rect 16304 1838 16356 1844
rect 16316 800 16344 1838
rect 17144 800 17172 6054
rect 17236 4826 17264 6598
rect 17420 6118 17448 8298
rect 17512 8022 17540 8434
rect 17500 8016 17552 8022
rect 17500 7958 17552 7964
rect 17500 7880 17552 7886
rect 17500 7822 17552 7828
rect 17512 7721 17540 7822
rect 17498 7712 17554 7721
rect 17498 7647 17554 7656
rect 17500 7268 17552 7274
rect 17500 7210 17552 7216
rect 17512 6866 17540 7210
rect 17500 6860 17552 6866
rect 17500 6802 17552 6808
rect 17408 6112 17460 6118
rect 17408 6054 17460 6060
rect 17224 4820 17276 4826
rect 17224 4762 17276 4768
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 17420 4214 17448 4558
rect 17500 4480 17552 4486
rect 17500 4422 17552 4428
rect 17512 4282 17540 4422
rect 17500 4276 17552 4282
rect 17500 4218 17552 4224
rect 17408 4208 17460 4214
rect 17408 4150 17460 4156
rect 17408 3596 17460 3602
rect 17408 3538 17460 3544
rect 17420 2922 17448 3538
rect 17408 2916 17460 2922
rect 17408 2858 17460 2864
rect 17604 2514 17632 9318
rect 17788 8537 17816 9862
rect 17972 9722 18000 9998
rect 18052 9920 18104 9926
rect 18052 9862 18104 9868
rect 17960 9716 18012 9722
rect 17960 9658 18012 9664
rect 18064 9518 18092 9862
rect 18328 9648 18380 9654
rect 18328 9590 18380 9596
rect 18052 9512 18104 9518
rect 18236 9512 18288 9518
rect 18052 9454 18104 9460
rect 18156 9472 18236 9500
rect 18064 8566 18092 9454
rect 18156 9382 18184 9472
rect 18236 9454 18288 9460
rect 18144 9376 18196 9382
rect 18144 9318 18196 9324
rect 18156 8838 18184 9318
rect 18144 8832 18196 8838
rect 18144 8774 18196 8780
rect 18052 8560 18104 8566
rect 17774 8528 17830 8537
rect 18052 8502 18104 8508
rect 17774 8463 17830 8472
rect 17960 8084 18012 8090
rect 17960 8026 18012 8032
rect 17684 7336 17736 7342
rect 17684 7278 17736 7284
rect 17696 4570 17724 7278
rect 17972 6254 18000 8026
rect 18064 6866 18092 8502
rect 18156 8294 18184 8774
rect 18340 8566 18368 9590
rect 18432 9110 18460 12106
rect 18616 10674 18644 13126
rect 18708 12714 18736 13806
rect 18696 12708 18748 12714
rect 18696 12650 18748 12656
rect 18880 12640 18932 12646
rect 18880 12582 18932 12588
rect 18972 12640 19024 12646
rect 18972 12582 19024 12588
rect 18696 12300 18748 12306
rect 18696 12242 18748 12248
rect 18708 11218 18736 12242
rect 18892 12073 18920 12582
rect 18984 12170 19012 12582
rect 19352 12442 19380 15506
rect 19536 14822 19564 15506
rect 19800 15360 19852 15366
rect 19800 15302 19852 15308
rect 19524 14816 19576 14822
rect 19524 14758 19576 14764
rect 19524 13728 19576 13734
rect 19524 13670 19576 13676
rect 19536 13326 19564 13670
rect 19616 13456 19668 13462
rect 19616 13398 19668 13404
rect 19524 13320 19576 13326
rect 19524 13262 19576 13268
rect 19430 13016 19486 13025
rect 19536 12986 19564 13262
rect 19430 12951 19432 12960
rect 19484 12951 19486 12960
rect 19524 12980 19576 12986
rect 19432 12922 19484 12928
rect 19524 12922 19576 12928
rect 19628 12866 19656 13398
rect 19536 12850 19656 12866
rect 19524 12844 19656 12850
rect 19576 12838 19656 12844
rect 19524 12786 19576 12792
rect 19623 12776 19675 12782
rect 19812 12764 19840 15302
rect 20364 15026 20392 15982
rect 20456 15910 20484 16934
rect 20548 16250 20576 19162
rect 20720 16992 20772 16998
rect 20720 16934 20772 16940
rect 20732 16590 20760 16934
rect 21748 16892 22044 16912
rect 21804 16890 21828 16892
rect 21884 16890 21908 16892
rect 21964 16890 21988 16892
rect 21826 16838 21828 16890
rect 21890 16838 21902 16890
rect 21964 16838 21966 16890
rect 21804 16836 21828 16838
rect 21884 16836 21908 16838
rect 21964 16836 21988 16838
rect 21748 16816 22044 16836
rect 22480 16794 22508 19162
rect 24412 17338 24440 19162
rect 24400 17332 24452 17338
rect 24400 17274 24452 17280
rect 22744 17264 22796 17270
rect 22744 17206 22796 17212
rect 22756 17134 22784 17206
rect 22744 17128 22796 17134
rect 22744 17070 22796 17076
rect 23112 17128 23164 17134
rect 23112 17070 23164 17076
rect 22468 16788 22520 16794
rect 22468 16730 22520 16736
rect 22100 16652 22152 16658
rect 22100 16594 22152 16600
rect 20720 16584 20772 16590
rect 20720 16526 20772 16532
rect 21456 16584 21508 16590
rect 21456 16526 21508 16532
rect 20536 16244 20588 16250
rect 20536 16186 20588 16192
rect 20996 16244 21048 16250
rect 20996 16186 21048 16192
rect 20444 15904 20496 15910
rect 20444 15846 20496 15852
rect 20456 15570 20484 15846
rect 20444 15564 20496 15570
rect 20444 15506 20496 15512
rect 20352 15020 20404 15026
rect 20352 14962 20404 14968
rect 20456 14958 20484 15506
rect 21008 15094 21036 16186
rect 21088 16176 21140 16182
rect 21088 16118 21140 16124
rect 21100 15638 21128 16118
rect 21468 15638 21496 16526
rect 22112 15978 22140 16594
rect 22376 16176 22428 16182
rect 22376 16118 22428 16124
rect 22100 15972 22152 15978
rect 22100 15914 22152 15920
rect 21748 15804 22044 15824
rect 21804 15802 21828 15804
rect 21884 15802 21908 15804
rect 21964 15802 21988 15804
rect 21826 15750 21828 15802
rect 21890 15750 21902 15802
rect 21964 15750 21966 15802
rect 21804 15748 21828 15750
rect 21884 15748 21908 15750
rect 21964 15748 21988 15750
rect 21748 15728 22044 15748
rect 21088 15632 21140 15638
rect 21088 15574 21140 15580
rect 21456 15632 21508 15638
rect 21456 15574 21508 15580
rect 21640 15496 21692 15502
rect 21640 15438 21692 15444
rect 22008 15496 22060 15502
rect 22008 15438 22060 15444
rect 20812 15088 20864 15094
rect 20812 15030 20864 15036
rect 20996 15088 21048 15094
rect 20996 15030 21048 15036
rect 21088 15088 21140 15094
rect 21088 15030 21140 15036
rect 20536 15020 20588 15026
rect 20536 14962 20588 14968
rect 19984 14952 20036 14958
rect 19982 14920 19984 14929
rect 20444 14952 20496 14958
rect 20036 14920 20038 14929
rect 20444 14894 20496 14900
rect 19982 14855 20038 14864
rect 20168 14816 20220 14822
rect 20168 14758 20220 14764
rect 19892 14476 19944 14482
rect 19892 14418 19944 14424
rect 19904 13870 19932 14418
rect 19984 14272 20036 14278
rect 19984 14214 20036 14220
rect 19892 13864 19944 13870
rect 19892 13806 19944 13812
rect 19675 12736 19840 12764
rect 19623 12718 19675 12724
rect 19524 12708 19576 12714
rect 19524 12650 19576 12656
rect 19340 12436 19392 12442
rect 19340 12378 19392 12384
rect 19536 12306 19564 12650
rect 19524 12300 19576 12306
rect 19524 12242 19576 12248
rect 19156 12232 19208 12238
rect 19156 12174 19208 12180
rect 18972 12164 19024 12170
rect 18972 12106 19024 12112
rect 18878 12064 18934 12073
rect 18878 11999 18934 12008
rect 19168 11830 19196 12174
rect 19616 12164 19668 12170
rect 19616 12106 19668 12112
rect 19524 12096 19576 12102
rect 19524 12038 19576 12044
rect 19156 11824 19208 11830
rect 19156 11766 19208 11772
rect 18880 11620 18932 11626
rect 18880 11562 18932 11568
rect 18892 11354 18920 11562
rect 19168 11558 19196 11766
rect 19156 11552 19208 11558
rect 19156 11494 19208 11500
rect 18880 11348 18932 11354
rect 18880 11290 18932 11296
rect 18696 11212 18748 11218
rect 18696 11154 18748 11160
rect 18892 11150 18920 11290
rect 18880 11144 18932 11150
rect 18880 11086 18932 11092
rect 19064 11076 19116 11082
rect 19064 11018 19116 11024
rect 18696 11008 18748 11014
rect 18696 10950 18748 10956
rect 18604 10668 18656 10674
rect 18604 10610 18656 10616
rect 18512 9580 18564 9586
rect 18512 9522 18564 9528
rect 18420 9104 18472 9110
rect 18420 9046 18472 9052
rect 18524 8838 18552 9522
rect 18708 9450 18736 10950
rect 18788 10532 18840 10538
rect 18788 10474 18840 10480
rect 18972 10532 19024 10538
rect 18972 10474 19024 10480
rect 18800 9722 18828 10474
rect 18788 9716 18840 9722
rect 18788 9658 18840 9664
rect 18696 9444 18748 9450
rect 18696 9386 18748 9392
rect 18800 9330 18828 9658
rect 18616 9302 18828 9330
rect 18616 9110 18644 9302
rect 18604 9104 18656 9110
rect 18604 9046 18656 9052
rect 18696 9104 18748 9110
rect 18696 9046 18748 9052
rect 18512 8832 18564 8838
rect 18512 8774 18564 8780
rect 18708 8673 18736 9046
rect 18694 8664 18750 8673
rect 18694 8599 18750 8608
rect 18328 8560 18380 8566
rect 18328 8502 18380 8508
rect 18144 8288 18196 8294
rect 18144 8230 18196 8236
rect 18340 8090 18368 8502
rect 18880 8356 18932 8362
rect 18880 8298 18932 8304
rect 18328 8084 18380 8090
rect 18328 8026 18380 8032
rect 18236 7880 18288 7886
rect 18236 7822 18288 7828
rect 18248 7546 18276 7822
rect 18892 7818 18920 8298
rect 18880 7812 18932 7818
rect 18880 7754 18932 7760
rect 18236 7540 18288 7546
rect 18236 7482 18288 7488
rect 18144 7336 18196 7342
rect 18144 7278 18196 7284
rect 18052 6860 18104 6866
rect 18052 6802 18104 6808
rect 18064 6390 18092 6802
rect 18156 6730 18184 7278
rect 18248 6934 18276 7482
rect 18892 7342 18920 7754
rect 18880 7336 18932 7342
rect 18880 7278 18932 7284
rect 18604 7200 18656 7206
rect 18604 7142 18656 7148
rect 18788 7200 18840 7206
rect 18788 7142 18840 7148
rect 18880 7200 18932 7206
rect 18984 7188 19012 10474
rect 19076 9586 19104 11018
rect 19168 10810 19196 11494
rect 19536 11014 19564 12038
rect 19628 11694 19656 12106
rect 19800 12096 19852 12102
rect 19800 12038 19852 12044
rect 19812 11694 19840 12038
rect 19616 11688 19668 11694
rect 19616 11630 19668 11636
rect 19800 11688 19852 11694
rect 19800 11630 19852 11636
rect 19248 11008 19300 11014
rect 19248 10950 19300 10956
rect 19524 11008 19576 11014
rect 19524 10950 19576 10956
rect 19156 10804 19208 10810
rect 19156 10746 19208 10752
rect 19260 9908 19288 10950
rect 19628 10742 19656 11630
rect 19616 10736 19668 10742
rect 19616 10678 19668 10684
rect 19628 10606 19656 10678
rect 19616 10600 19668 10606
rect 19616 10542 19668 10548
rect 19340 9920 19392 9926
rect 19260 9880 19340 9908
rect 19340 9862 19392 9868
rect 19708 9920 19760 9926
rect 19708 9862 19760 9868
rect 19156 9648 19208 9654
rect 19156 9590 19208 9596
rect 19246 9616 19302 9625
rect 19064 9580 19116 9586
rect 19064 9522 19116 9528
rect 19168 9042 19196 9590
rect 19246 9551 19248 9560
rect 19300 9551 19302 9560
rect 19248 9522 19300 9528
rect 19248 9444 19300 9450
rect 19248 9386 19300 9392
rect 19260 9042 19288 9386
rect 19156 9036 19208 9042
rect 19156 8978 19208 8984
rect 19248 9036 19300 9042
rect 19248 8978 19300 8984
rect 19720 8974 19748 9862
rect 19812 9654 19840 11630
rect 19996 11286 20024 14214
rect 19984 11280 20036 11286
rect 19984 11222 20036 11228
rect 20074 10568 20130 10577
rect 20074 10503 20130 10512
rect 20088 10266 20116 10503
rect 20076 10260 20128 10266
rect 20076 10202 20128 10208
rect 19800 9648 19852 9654
rect 19800 9590 19852 9596
rect 19984 9512 20036 9518
rect 19984 9454 20036 9460
rect 19340 8968 19392 8974
rect 19340 8910 19392 8916
rect 19708 8968 19760 8974
rect 19708 8910 19760 8916
rect 19352 8566 19380 8910
rect 19892 8832 19944 8838
rect 19892 8774 19944 8780
rect 19340 8560 19392 8566
rect 19340 8502 19392 8508
rect 19708 8356 19760 8362
rect 19708 8298 19760 8304
rect 19524 8084 19576 8090
rect 19524 8026 19576 8032
rect 19536 7274 19564 8026
rect 19720 7886 19748 8298
rect 19800 8288 19852 8294
rect 19800 8230 19852 8236
rect 19708 7880 19760 7886
rect 19708 7822 19760 7828
rect 19720 7342 19748 7822
rect 19812 7585 19840 8230
rect 19798 7576 19854 7585
rect 19798 7511 19854 7520
rect 19708 7336 19760 7342
rect 19708 7278 19760 7284
rect 19524 7268 19576 7274
rect 19524 7210 19576 7216
rect 18932 7160 19012 7188
rect 18880 7142 18932 7148
rect 18616 7002 18644 7142
rect 18512 6996 18564 7002
rect 18512 6938 18564 6944
rect 18604 6996 18656 7002
rect 18604 6938 18656 6944
rect 18236 6928 18288 6934
rect 18236 6870 18288 6876
rect 18144 6724 18196 6730
rect 18144 6666 18196 6672
rect 18236 6656 18288 6662
rect 18236 6598 18288 6604
rect 18052 6384 18104 6390
rect 18104 6344 18184 6372
rect 18052 6326 18104 6332
rect 17960 6248 18012 6254
rect 17960 6190 18012 6196
rect 18052 6180 18104 6186
rect 18052 6122 18104 6128
rect 17776 5772 17828 5778
rect 17776 5714 17828 5720
rect 17788 5166 17816 5714
rect 18064 5710 18092 6122
rect 18156 5778 18184 6344
rect 18248 6322 18276 6598
rect 18236 6316 18288 6322
rect 18236 6258 18288 6264
rect 18236 6180 18288 6186
rect 18236 6122 18288 6128
rect 18144 5772 18196 5778
rect 18144 5714 18196 5720
rect 18052 5704 18104 5710
rect 18052 5646 18104 5652
rect 17776 5160 17828 5166
rect 17776 5102 17828 5108
rect 17788 4826 17816 5102
rect 18064 4826 18092 5646
rect 18144 5364 18196 5370
rect 18144 5306 18196 5312
rect 17776 4820 17828 4826
rect 17776 4762 17828 4768
rect 18052 4820 18104 4826
rect 18052 4762 18104 4768
rect 18156 4690 18184 5306
rect 18248 5098 18276 6122
rect 18524 5166 18552 6938
rect 18696 6248 18748 6254
rect 18696 6190 18748 6196
rect 18708 5778 18736 6190
rect 18800 5846 18828 7142
rect 18788 5840 18840 5846
rect 18788 5782 18840 5788
rect 18696 5772 18748 5778
rect 18696 5714 18748 5720
rect 18708 5574 18736 5714
rect 18696 5568 18748 5574
rect 18696 5510 18748 5516
rect 18604 5296 18656 5302
rect 18604 5238 18656 5244
rect 18512 5160 18564 5166
rect 18512 5102 18564 5108
rect 18236 5092 18288 5098
rect 18236 5034 18288 5040
rect 18328 5024 18380 5030
rect 18328 4966 18380 4972
rect 18144 4684 18196 4690
rect 18144 4626 18196 4632
rect 18340 4622 18368 4966
rect 18616 4690 18644 5238
rect 18604 4684 18656 4690
rect 18604 4626 18656 4632
rect 18328 4616 18380 4622
rect 17696 4542 18000 4570
rect 18328 4558 18380 4564
rect 17972 4486 18000 4542
rect 17960 4480 18012 4486
rect 17960 4422 18012 4428
rect 18236 4004 18288 4010
rect 18236 3946 18288 3952
rect 18052 3732 18104 3738
rect 18052 3674 18104 3680
rect 17684 3664 17736 3670
rect 17736 3612 17816 3618
rect 17684 3606 17816 3612
rect 17696 3590 17816 3606
rect 17788 3369 17816 3590
rect 17868 3596 17920 3602
rect 17868 3538 17920 3544
rect 17774 3360 17830 3369
rect 17774 3295 17830 3304
rect 17788 3194 17816 3295
rect 17776 3188 17828 3194
rect 17776 3130 17828 3136
rect 17774 2952 17830 2961
rect 17684 2916 17736 2922
rect 17880 2922 17908 3538
rect 18064 3194 18092 3674
rect 18248 3670 18276 3946
rect 18236 3664 18288 3670
rect 18236 3606 18288 3612
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 18052 3188 18104 3194
rect 18052 3130 18104 3136
rect 18144 3188 18196 3194
rect 18144 3130 18196 3136
rect 18064 2990 18092 3130
rect 18052 2984 18104 2990
rect 18052 2926 18104 2932
rect 17774 2887 17830 2896
rect 17868 2916 17920 2922
rect 17684 2858 17736 2864
rect 17592 2508 17644 2514
rect 17592 2450 17644 2456
rect 17604 1902 17632 2450
rect 17696 2310 17724 2858
rect 17788 2802 17816 2887
rect 17868 2858 17920 2864
rect 18156 2836 18184 3130
rect 18340 2990 18368 3470
rect 18616 3398 18644 4626
rect 18786 4176 18842 4185
rect 18786 4111 18842 4120
rect 18800 4078 18828 4111
rect 18788 4072 18840 4078
rect 18788 4014 18840 4020
rect 18696 3596 18748 3602
rect 18696 3538 18748 3544
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 18708 3126 18736 3538
rect 18696 3120 18748 3126
rect 18696 3062 18748 3068
rect 18328 2984 18380 2990
rect 18328 2926 18380 2932
rect 18708 2854 18736 3062
rect 17972 2808 18184 2836
rect 18696 2848 18748 2854
rect 17972 2802 18000 2808
rect 17788 2774 18000 2802
rect 18696 2790 18748 2796
rect 17880 2582 17908 2774
rect 17868 2576 17920 2582
rect 17868 2518 17920 2524
rect 18892 2378 18920 7142
rect 19536 6866 19564 7210
rect 19064 6860 19116 6866
rect 18984 6820 19064 6848
rect 18984 4622 19012 6820
rect 19064 6802 19116 6808
rect 19248 6860 19300 6866
rect 19248 6802 19300 6808
rect 19524 6860 19576 6866
rect 19524 6802 19576 6808
rect 19064 6248 19116 6254
rect 19260 6236 19288 6802
rect 19338 6760 19394 6769
rect 19338 6695 19340 6704
rect 19392 6695 19394 6704
rect 19340 6666 19392 6672
rect 19432 6316 19484 6322
rect 19432 6258 19484 6264
rect 19340 6248 19392 6254
rect 19260 6208 19340 6236
rect 19064 6190 19116 6196
rect 19340 6190 19392 6196
rect 19076 5370 19104 6190
rect 19246 6080 19302 6089
rect 19246 6015 19302 6024
rect 19064 5364 19116 5370
rect 19064 5306 19116 5312
rect 19156 5364 19208 5370
rect 19156 5306 19208 5312
rect 19168 5137 19196 5306
rect 19154 5128 19210 5137
rect 19154 5063 19210 5072
rect 18972 4616 19024 4622
rect 18972 4558 19024 4564
rect 19260 4214 19288 6015
rect 19352 5846 19380 6190
rect 19340 5840 19392 5846
rect 19340 5782 19392 5788
rect 19340 5568 19392 5574
rect 19340 5510 19392 5516
rect 19352 5234 19380 5510
rect 19340 5228 19392 5234
rect 19340 5170 19392 5176
rect 19340 4684 19392 4690
rect 19340 4626 19392 4632
rect 19248 4208 19300 4214
rect 18970 4176 19026 4185
rect 19248 4150 19300 4156
rect 18970 4111 19026 4120
rect 18984 3233 19012 4111
rect 19248 3392 19300 3398
rect 19248 3334 19300 3340
rect 19260 3233 19288 3334
rect 18970 3224 19026 3233
rect 18970 3159 19026 3168
rect 19246 3224 19302 3233
rect 19246 3159 19302 3168
rect 18972 3120 19024 3126
rect 18972 3062 19024 3068
rect 18052 2372 18104 2378
rect 18052 2314 18104 2320
rect 18880 2372 18932 2378
rect 18880 2314 18932 2320
rect 17684 2304 17736 2310
rect 17684 2246 17736 2252
rect 17592 1896 17644 1902
rect 17592 1838 17644 1844
rect 18064 800 18092 2314
rect 18984 800 19012 3062
rect 19064 3052 19116 3058
rect 19064 2994 19116 3000
rect 19076 2689 19104 2994
rect 19062 2680 19118 2689
rect 19062 2615 19118 2624
rect 19260 2446 19288 3159
rect 19352 2650 19380 4626
rect 19444 4457 19472 6258
rect 19536 5760 19564 6802
rect 19812 5930 19840 7511
rect 19904 6882 19932 8774
rect 19996 8634 20024 9454
rect 19984 8628 20036 8634
rect 19984 8570 20036 8576
rect 20180 7954 20208 14758
rect 20548 14618 20576 14962
rect 20536 14612 20588 14618
rect 20536 14554 20588 14560
rect 20720 14544 20772 14550
rect 20548 14492 20720 14498
rect 20824 14521 20852 15030
rect 21008 14890 21036 15030
rect 20996 14884 21048 14890
rect 20996 14826 21048 14832
rect 20548 14486 20772 14492
rect 20810 14512 20866 14521
rect 20548 14470 20760 14486
rect 20444 13796 20496 13802
rect 20444 13738 20496 13744
rect 20456 13025 20484 13738
rect 20258 13016 20314 13025
rect 20258 12951 20314 12960
rect 20442 13016 20498 13025
rect 20442 12951 20498 12960
rect 20272 12442 20300 12951
rect 20260 12436 20312 12442
rect 20260 12378 20312 12384
rect 20548 12170 20576 14470
rect 20810 14447 20866 14456
rect 20720 14272 20772 14278
rect 21100 14226 21128 15030
rect 21652 14550 21680 15438
rect 22020 15094 22048 15438
rect 22008 15088 22060 15094
rect 21914 15056 21970 15065
rect 22008 15030 22060 15036
rect 22388 15026 22416 16118
rect 22480 15162 22508 16730
rect 22756 16454 22784 17070
rect 22560 16448 22612 16454
rect 22560 16390 22612 16396
rect 22744 16448 22796 16454
rect 22744 16390 22796 16396
rect 22572 16182 22600 16390
rect 22560 16176 22612 16182
rect 22560 16118 22612 16124
rect 22560 15972 22612 15978
rect 22560 15914 22612 15920
rect 22468 15156 22520 15162
rect 22468 15098 22520 15104
rect 22480 15065 22508 15098
rect 22466 15056 22522 15065
rect 21914 14991 21970 15000
rect 22376 15020 22428 15026
rect 21928 14958 21956 14991
rect 22572 15026 22600 15914
rect 23124 15638 23152 17070
rect 23572 17060 23624 17066
rect 23572 17002 23624 17008
rect 23584 15978 23612 17002
rect 24412 16810 24440 17274
rect 24412 16794 24532 16810
rect 24412 16788 24544 16794
rect 24412 16782 24492 16788
rect 24492 16730 24544 16736
rect 25044 16652 25096 16658
rect 25044 16594 25096 16600
rect 23848 16584 23900 16590
rect 23848 16526 23900 16532
rect 23860 16114 23888 16526
rect 25056 16114 25084 16594
rect 26344 16522 26372 19162
rect 28368 17338 28396 19162
rect 28356 17332 28408 17338
rect 28356 17274 28408 17280
rect 28908 17332 28960 17338
rect 28908 17274 28960 17280
rect 27528 17196 27580 17202
rect 27528 17138 27580 17144
rect 26332 16516 26384 16522
rect 26332 16458 26384 16464
rect 25412 16448 25464 16454
rect 25412 16390 25464 16396
rect 26148 16448 26200 16454
rect 26148 16390 26200 16396
rect 25424 16182 25452 16390
rect 25412 16176 25464 16182
rect 25412 16118 25464 16124
rect 26160 16114 26188 16390
rect 23848 16108 23900 16114
rect 23848 16050 23900 16056
rect 25044 16108 25096 16114
rect 25044 16050 25096 16056
rect 26148 16108 26200 16114
rect 26148 16050 26200 16056
rect 23664 16040 23716 16046
rect 23664 15982 23716 15988
rect 24124 16040 24176 16046
rect 24124 15982 24176 15988
rect 23572 15972 23624 15978
rect 23572 15914 23624 15920
rect 23584 15706 23612 15914
rect 23676 15910 23704 15982
rect 23664 15904 23716 15910
rect 23664 15846 23716 15852
rect 23572 15700 23624 15706
rect 23572 15642 23624 15648
rect 23112 15632 23164 15638
rect 23112 15574 23164 15580
rect 23124 15094 23152 15574
rect 23676 15366 23704 15846
rect 24136 15570 24164 15982
rect 24124 15564 24176 15570
rect 24124 15506 24176 15512
rect 24676 15564 24728 15570
rect 24676 15506 24728 15512
rect 23296 15360 23348 15366
rect 23296 15302 23348 15308
rect 23664 15360 23716 15366
rect 23664 15302 23716 15308
rect 23308 15094 23336 15302
rect 23112 15088 23164 15094
rect 23112 15030 23164 15036
rect 23296 15088 23348 15094
rect 23296 15030 23348 15036
rect 22466 14991 22522 15000
rect 22560 15020 22612 15026
rect 22376 14962 22428 14968
rect 22560 14962 22612 14968
rect 23124 14958 23152 15030
rect 21916 14952 21968 14958
rect 21916 14894 21968 14900
rect 23112 14952 23164 14958
rect 23112 14894 23164 14900
rect 22376 14816 22428 14822
rect 22376 14758 22428 14764
rect 21748 14716 22044 14736
rect 21804 14714 21828 14716
rect 21884 14714 21908 14716
rect 21964 14714 21988 14716
rect 21826 14662 21828 14714
rect 21890 14662 21902 14714
rect 21964 14662 21966 14714
rect 21804 14660 21828 14662
rect 21884 14660 21908 14662
rect 21964 14660 21988 14662
rect 21748 14640 22044 14660
rect 21640 14544 21692 14550
rect 21640 14486 21692 14492
rect 21652 14414 21680 14486
rect 21548 14408 21600 14414
rect 21546 14376 21548 14385
rect 21640 14408 21692 14414
rect 21600 14376 21602 14385
rect 21640 14350 21692 14356
rect 21546 14311 21602 14320
rect 20720 14214 20772 14220
rect 20732 14090 20760 14214
rect 20640 14062 20760 14090
rect 21008 14198 21128 14226
rect 21364 14272 21416 14278
rect 21364 14214 21416 14220
rect 22098 14240 22154 14249
rect 20640 12481 20668 14062
rect 21008 13870 21036 14198
rect 21088 14068 21140 14074
rect 21088 14010 21140 14016
rect 21180 14068 21232 14074
rect 21180 14010 21232 14016
rect 20720 13864 20772 13870
rect 20720 13806 20772 13812
rect 20996 13864 21048 13870
rect 20996 13806 21048 13812
rect 20626 12472 20682 12481
rect 20626 12407 20682 12416
rect 20640 12306 20668 12407
rect 20628 12300 20680 12306
rect 20628 12242 20680 12248
rect 20536 12164 20588 12170
rect 20536 12106 20588 12112
rect 20352 11008 20404 11014
rect 20352 10950 20404 10956
rect 20444 11008 20496 11014
rect 20444 10950 20496 10956
rect 20364 10606 20392 10950
rect 20352 10600 20404 10606
rect 20352 10542 20404 10548
rect 20364 10198 20392 10542
rect 20456 10266 20484 10950
rect 20732 10742 20760 13806
rect 20996 13524 21048 13530
rect 20996 13466 21048 13472
rect 20812 13456 20864 13462
rect 20812 13398 20864 13404
rect 20824 12918 20852 13398
rect 20904 13252 20956 13258
rect 20904 13194 20956 13200
rect 20812 12912 20864 12918
rect 20812 12854 20864 12860
rect 20916 12782 20944 13194
rect 20904 12776 20956 12782
rect 20904 12718 20956 12724
rect 20916 12374 20944 12718
rect 20904 12368 20956 12374
rect 20904 12310 20956 12316
rect 21008 12322 21036 13466
rect 21100 12442 21128 14010
rect 21192 13977 21220 14010
rect 21178 13968 21234 13977
rect 21178 13903 21234 13912
rect 21180 12640 21232 12646
rect 21180 12582 21232 12588
rect 21088 12436 21140 12442
rect 21088 12378 21140 12384
rect 21192 12322 21220 12582
rect 21008 12294 21220 12322
rect 21088 11824 21140 11830
rect 21088 11766 21140 11772
rect 21100 11694 21128 11766
rect 21088 11688 21140 11694
rect 21192 11665 21220 12294
rect 21088 11630 21140 11636
rect 21178 11656 21234 11665
rect 20904 11620 20956 11626
rect 20904 11562 20956 11568
rect 20916 11286 20944 11562
rect 20904 11280 20956 11286
rect 20904 11222 20956 11228
rect 20720 10736 20772 10742
rect 20720 10678 20772 10684
rect 20444 10260 20496 10266
rect 20444 10202 20496 10208
rect 20352 10192 20404 10198
rect 20352 10134 20404 10140
rect 20994 10160 21050 10169
rect 20812 10124 20864 10130
rect 20994 10095 21050 10104
rect 20812 10066 20864 10072
rect 20720 9920 20772 9926
rect 20720 9862 20772 9868
rect 20732 9586 20760 9862
rect 20824 9722 20852 10066
rect 21008 10062 21036 10095
rect 20996 10056 21048 10062
rect 20996 9998 21048 10004
rect 21100 9761 21128 11630
rect 21178 11591 21234 11600
rect 21180 11348 21232 11354
rect 21180 11290 21232 11296
rect 21192 10266 21220 11290
rect 21272 11144 21324 11150
rect 21272 11086 21324 11092
rect 21284 10810 21312 11086
rect 21272 10804 21324 10810
rect 21272 10746 21324 10752
rect 21180 10260 21232 10266
rect 21180 10202 21232 10208
rect 21180 9988 21232 9994
rect 21180 9930 21232 9936
rect 21086 9752 21142 9761
rect 20812 9716 20864 9722
rect 21086 9687 21142 9696
rect 20812 9658 20864 9664
rect 20720 9580 20772 9586
rect 20720 9522 20772 9528
rect 20824 9450 20852 9658
rect 21100 9518 21128 9687
rect 21088 9512 21140 9518
rect 21088 9454 21140 9460
rect 20260 9444 20312 9450
rect 20260 9386 20312 9392
rect 20812 9444 20864 9450
rect 20812 9386 20864 9392
rect 20272 8838 20300 9386
rect 21088 9376 21140 9382
rect 21192 9364 21220 9930
rect 21376 9926 21404 14214
rect 22098 14175 22154 14184
rect 22112 14006 22140 14175
rect 22388 14074 22416 14758
rect 22560 14408 22612 14414
rect 22560 14350 22612 14356
rect 22572 14074 22600 14350
rect 22376 14068 22428 14074
rect 22376 14010 22428 14016
rect 22560 14068 22612 14074
rect 22560 14010 22612 14016
rect 21824 14000 21876 14006
rect 21824 13942 21876 13948
rect 22100 14000 22152 14006
rect 22100 13942 22152 13948
rect 21836 13870 21864 13942
rect 21640 13864 21692 13870
rect 21640 13806 21692 13812
rect 21824 13864 21876 13870
rect 21824 13806 21876 13812
rect 22100 13864 22152 13870
rect 22100 13806 22152 13812
rect 21548 13388 21600 13394
rect 21548 13330 21600 13336
rect 21456 12300 21508 12306
rect 21456 12242 21508 12248
rect 21468 12102 21496 12242
rect 21456 12096 21508 12102
rect 21456 12038 21508 12044
rect 21364 9920 21416 9926
rect 21364 9862 21416 9868
rect 21272 9376 21324 9382
rect 21192 9336 21272 9364
rect 21088 9318 21140 9324
rect 21272 9318 21324 9324
rect 20904 8968 20956 8974
rect 21100 8945 21128 9318
rect 21284 8974 21312 9318
rect 21468 9042 21496 12038
rect 21560 9042 21588 13330
rect 21652 10248 21680 13806
rect 21748 13628 22044 13648
rect 21804 13626 21828 13628
rect 21884 13626 21908 13628
rect 21964 13626 21988 13628
rect 21826 13574 21828 13626
rect 21890 13574 21902 13626
rect 21964 13574 21966 13626
rect 21804 13572 21828 13574
rect 21884 13572 21908 13574
rect 21964 13572 21988 13574
rect 21748 13552 22044 13572
rect 22112 13462 22140 13806
rect 22192 13796 22244 13802
rect 22192 13738 22244 13744
rect 22100 13456 22152 13462
rect 22100 13398 22152 13404
rect 21824 13388 21876 13394
rect 21824 13330 21876 13336
rect 21916 13388 21968 13394
rect 21916 13330 21968 13336
rect 21836 12714 21864 13330
rect 21928 13274 21956 13330
rect 22204 13274 22232 13738
rect 21928 13246 22232 13274
rect 22572 13258 22600 14010
rect 23308 13938 23336 15030
rect 23676 14958 23704 15302
rect 23664 14952 23716 14958
rect 23662 14920 23664 14929
rect 23940 14952 23992 14958
rect 23716 14920 23718 14929
rect 23940 14894 23992 14900
rect 23662 14855 23718 14864
rect 23848 14884 23900 14890
rect 23848 14826 23900 14832
rect 23860 14550 23888 14826
rect 23848 14544 23900 14550
rect 23848 14486 23900 14492
rect 23952 14278 23980 14894
rect 24688 14890 24716 15506
rect 25056 15366 25084 16050
rect 26976 16040 27028 16046
rect 26976 15982 27028 15988
rect 27068 16040 27120 16046
rect 27068 15982 27120 15988
rect 26988 15706 27016 15982
rect 26976 15700 27028 15706
rect 26976 15642 27028 15648
rect 26056 15632 26108 15638
rect 26056 15574 26108 15580
rect 25044 15360 25096 15366
rect 25044 15302 25096 15308
rect 25964 15360 26016 15366
rect 25964 15302 26016 15308
rect 25056 15026 25084 15302
rect 25044 15020 25096 15026
rect 25044 14962 25096 14968
rect 25228 15020 25280 15026
rect 25228 14962 25280 14968
rect 24676 14884 24728 14890
rect 24676 14826 24728 14832
rect 25136 14884 25188 14890
rect 25136 14826 25188 14832
rect 24688 14385 24716 14826
rect 25148 14482 25176 14826
rect 24860 14476 24912 14482
rect 24860 14418 24912 14424
rect 25136 14476 25188 14482
rect 25136 14418 25188 14424
rect 24674 14376 24730 14385
rect 24674 14311 24730 14320
rect 23388 14272 23440 14278
rect 23388 14214 23440 14220
rect 23572 14272 23624 14278
rect 23572 14214 23624 14220
rect 23940 14272 23992 14278
rect 23940 14214 23992 14220
rect 24122 14240 24178 14249
rect 23296 13932 23348 13938
rect 23296 13874 23348 13880
rect 22928 13796 22980 13802
rect 22928 13738 22980 13744
rect 23020 13796 23072 13802
rect 23020 13738 23072 13744
rect 22744 13728 22796 13734
rect 22744 13670 22796 13676
rect 22560 13252 22612 13258
rect 21824 12708 21876 12714
rect 21824 12650 21876 12656
rect 21748 12540 22044 12560
rect 21804 12538 21828 12540
rect 21884 12538 21908 12540
rect 21964 12538 21988 12540
rect 21826 12486 21828 12538
rect 21890 12486 21902 12538
rect 21964 12486 21966 12538
rect 21804 12484 21828 12486
rect 21884 12484 21908 12486
rect 21964 12484 21988 12486
rect 21748 12464 22044 12484
rect 22112 12306 22140 13246
rect 22560 13194 22612 13200
rect 22468 12912 22520 12918
rect 22468 12854 22520 12860
rect 22652 12912 22704 12918
rect 22652 12854 22704 12860
rect 22480 12714 22508 12854
rect 22192 12708 22244 12714
rect 22192 12650 22244 12656
rect 22468 12708 22520 12714
rect 22468 12650 22520 12656
rect 21732 12300 21784 12306
rect 21732 12242 21784 12248
rect 22100 12300 22152 12306
rect 22100 12242 22152 12248
rect 21744 11665 21772 12242
rect 22112 11898 22140 12242
rect 22204 12102 22232 12650
rect 22560 12640 22612 12646
rect 22560 12582 22612 12588
rect 22572 12238 22600 12582
rect 22560 12232 22612 12238
rect 22560 12174 22612 12180
rect 22192 12096 22244 12102
rect 22192 12038 22244 12044
rect 22100 11892 22152 11898
rect 22100 11834 22152 11840
rect 22204 11694 22232 12038
rect 22192 11688 22244 11694
rect 21730 11656 21786 11665
rect 22192 11630 22244 11636
rect 21730 11591 21786 11600
rect 21748 11452 22044 11472
rect 21804 11450 21828 11452
rect 21884 11450 21908 11452
rect 21964 11450 21988 11452
rect 21826 11398 21828 11450
rect 21890 11398 21902 11450
rect 21964 11398 21966 11450
rect 21804 11396 21828 11398
rect 21884 11396 21908 11398
rect 21964 11396 21988 11398
rect 21748 11376 22044 11396
rect 22468 11212 22520 11218
rect 22468 11154 22520 11160
rect 21732 11008 21784 11014
rect 21732 10950 21784 10956
rect 22100 11008 22152 11014
rect 22100 10950 22152 10956
rect 21744 10810 21772 10950
rect 21732 10804 21784 10810
rect 21732 10746 21784 10752
rect 22112 10538 22140 10950
rect 22284 10804 22336 10810
rect 22284 10746 22336 10752
rect 22296 10577 22324 10746
rect 22282 10568 22338 10577
rect 22100 10532 22152 10538
rect 22282 10503 22338 10512
rect 22100 10474 22152 10480
rect 21748 10364 22044 10384
rect 21804 10362 21828 10364
rect 21884 10362 21908 10364
rect 21964 10362 21988 10364
rect 21826 10310 21828 10362
rect 21890 10310 21902 10362
rect 21964 10310 21966 10362
rect 21804 10308 21828 10310
rect 21884 10308 21908 10310
rect 21964 10308 21988 10310
rect 21748 10288 22044 10308
rect 21652 10220 21864 10248
rect 21732 9920 21784 9926
rect 21732 9862 21784 9868
rect 21744 9625 21772 9862
rect 21730 9616 21786 9625
rect 21730 9551 21786 9560
rect 21836 9568 21864 10220
rect 22112 10130 22140 10474
rect 22100 10124 22152 10130
rect 22100 10066 22152 10072
rect 22192 10056 22244 10062
rect 22192 9998 22244 10004
rect 21916 9580 21968 9586
rect 21836 9540 21916 9568
rect 21916 9522 21968 9528
rect 21638 9480 21694 9489
rect 21638 9415 21694 9424
rect 21652 9110 21680 9415
rect 21748 9276 22044 9296
rect 21804 9274 21828 9276
rect 21884 9274 21908 9276
rect 21964 9274 21988 9276
rect 21826 9222 21828 9274
rect 21890 9222 21902 9274
rect 21964 9222 21966 9274
rect 21804 9220 21828 9222
rect 21884 9220 21908 9222
rect 21964 9220 21988 9222
rect 21748 9200 22044 9220
rect 21640 9104 21692 9110
rect 21640 9046 21692 9052
rect 21456 9036 21508 9042
rect 21456 8978 21508 8984
rect 21548 9036 21600 9042
rect 21548 8978 21600 8984
rect 21272 8968 21324 8974
rect 20904 8910 20956 8916
rect 21086 8936 21142 8945
rect 20260 8832 20312 8838
rect 20260 8774 20312 8780
rect 20352 8832 20404 8838
rect 20352 8774 20404 8780
rect 20272 8634 20300 8774
rect 20260 8628 20312 8634
rect 20260 8570 20312 8576
rect 20364 8566 20392 8774
rect 20916 8634 20944 8910
rect 21272 8910 21324 8916
rect 21086 8871 21142 8880
rect 21548 8832 21600 8838
rect 21824 8832 21876 8838
rect 21548 8774 21600 8780
rect 21744 8792 21824 8820
rect 20904 8628 20956 8634
rect 20904 8570 20956 8576
rect 20352 8560 20404 8566
rect 20352 8502 20404 8508
rect 20364 8430 20392 8502
rect 21560 8430 21588 8774
rect 21640 8628 21692 8634
rect 21640 8570 21692 8576
rect 20352 8424 20404 8430
rect 20352 8366 20404 8372
rect 20720 8424 20772 8430
rect 20720 8366 20772 8372
rect 21548 8424 21600 8430
rect 21548 8366 21600 8372
rect 20168 7948 20220 7954
rect 20168 7890 20220 7896
rect 20180 7721 20208 7890
rect 20166 7712 20222 7721
rect 20166 7647 20222 7656
rect 20076 7336 20128 7342
rect 20076 7278 20128 7284
rect 20088 7206 20116 7278
rect 20260 7268 20312 7274
rect 20260 7210 20312 7216
rect 20076 7200 20128 7206
rect 20076 7142 20128 7148
rect 19904 6866 20116 6882
rect 19904 6860 20128 6866
rect 19904 6854 20076 6860
rect 20076 6802 20128 6808
rect 19892 6656 19944 6662
rect 19892 6598 19944 6604
rect 19904 6361 19932 6598
rect 19984 6384 20036 6390
rect 19890 6352 19946 6361
rect 19984 6326 20036 6332
rect 19890 6287 19946 6296
rect 19720 5902 19840 5930
rect 19616 5772 19668 5778
rect 19536 5732 19616 5760
rect 19616 5714 19668 5720
rect 19524 5024 19576 5030
rect 19524 4966 19576 4972
rect 19430 4448 19486 4457
rect 19430 4383 19486 4392
rect 19536 3738 19564 4966
rect 19720 4865 19748 5902
rect 19800 5840 19852 5846
rect 19800 5782 19852 5788
rect 19706 4856 19762 4865
rect 19706 4791 19762 4800
rect 19812 4486 19840 5782
rect 19996 4690 20024 6326
rect 19984 4684 20036 4690
rect 19984 4626 20036 4632
rect 20088 4570 20116 6802
rect 20168 6656 20220 6662
rect 20168 6598 20220 6604
rect 20180 6458 20208 6598
rect 20168 6452 20220 6458
rect 20168 6394 20220 6400
rect 20180 6254 20208 6394
rect 20168 6248 20220 6254
rect 20168 6190 20220 6196
rect 20180 5681 20208 6190
rect 20166 5672 20222 5681
rect 20166 5607 20222 5616
rect 20272 5302 20300 7210
rect 20732 7002 20760 8366
rect 21088 8084 21140 8090
rect 21088 8026 21140 8032
rect 21100 7954 21128 8026
rect 20904 7948 20956 7954
rect 20904 7890 20956 7896
rect 21088 7948 21140 7954
rect 21088 7890 21140 7896
rect 20916 7546 20944 7890
rect 20904 7540 20956 7546
rect 20904 7482 20956 7488
rect 21560 7342 21588 8366
rect 21180 7336 21232 7342
rect 21180 7278 21232 7284
rect 21548 7336 21600 7342
rect 21548 7278 21600 7284
rect 20812 7200 20864 7206
rect 20812 7142 20864 7148
rect 20720 6996 20772 7002
rect 20720 6938 20772 6944
rect 20628 6860 20680 6866
rect 20628 6802 20680 6808
rect 20536 6656 20588 6662
rect 20536 6598 20588 6604
rect 20548 6390 20576 6598
rect 20536 6384 20588 6390
rect 20536 6326 20588 6332
rect 20548 6254 20576 6326
rect 20640 6254 20668 6802
rect 20720 6452 20772 6458
rect 20720 6394 20772 6400
rect 20536 6248 20588 6254
rect 20536 6190 20588 6196
rect 20628 6248 20680 6254
rect 20628 6190 20680 6196
rect 20732 5914 20760 6394
rect 20720 5908 20772 5914
rect 20720 5850 20772 5856
rect 20260 5296 20312 5302
rect 20260 5238 20312 5244
rect 20732 5166 20760 5850
rect 20824 5370 20852 7142
rect 20904 6112 20956 6118
rect 20904 6054 20956 6060
rect 20916 5846 20944 6054
rect 20904 5840 20956 5846
rect 20904 5782 20956 5788
rect 21192 5409 21220 7278
rect 21272 6996 21324 7002
rect 21272 6938 21324 6944
rect 21364 6996 21416 7002
rect 21364 6938 21416 6944
rect 21284 5846 21312 6938
rect 21272 5840 21324 5846
rect 21270 5808 21272 5817
rect 21324 5808 21326 5817
rect 21270 5743 21326 5752
rect 21178 5400 21234 5409
rect 20812 5364 20864 5370
rect 21178 5335 21234 5344
rect 20812 5306 20864 5312
rect 20352 5160 20404 5166
rect 20720 5160 20772 5166
rect 20352 5102 20404 5108
rect 20442 5128 20498 5137
rect 20364 5030 20392 5102
rect 20996 5160 21048 5166
rect 20772 5120 20852 5148
rect 20720 5102 20772 5108
rect 20442 5063 20498 5072
rect 20352 5024 20404 5030
rect 20352 4966 20404 4972
rect 19904 4542 20116 4570
rect 19800 4480 19852 4486
rect 19800 4422 19852 4428
rect 19524 3732 19576 3738
rect 19524 3674 19576 3680
rect 19616 3528 19668 3534
rect 19616 3470 19668 3476
rect 19628 2650 19656 3470
rect 19340 2644 19392 2650
rect 19340 2586 19392 2592
rect 19616 2644 19668 2650
rect 19616 2586 19668 2592
rect 19812 2582 19840 4422
rect 19800 2576 19852 2582
rect 19800 2518 19852 2524
rect 19248 2440 19300 2446
rect 19248 2382 19300 2388
rect 19904 1442 19932 4542
rect 20260 4480 20312 4486
rect 20260 4422 20312 4428
rect 20168 4004 20220 4010
rect 20168 3946 20220 3952
rect 20076 3528 20128 3534
rect 20076 3470 20128 3476
rect 20088 2990 20116 3470
rect 20180 2990 20208 3946
rect 20272 3466 20300 4422
rect 20260 3460 20312 3466
rect 20364 3448 20392 4966
rect 20456 3738 20484 5063
rect 20720 4616 20772 4622
rect 20720 4558 20772 4564
rect 20732 4486 20760 4558
rect 20536 4480 20588 4486
rect 20720 4480 20772 4486
rect 20588 4440 20668 4468
rect 20536 4422 20588 4428
rect 20640 4078 20668 4440
rect 20720 4422 20772 4428
rect 20536 4072 20588 4078
rect 20536 4014 20588 4020
rect 20628 4072 20680 4078
rect 20628 4014 20680 4020
rect 20548 3913 20576 4014
rect 20534 3904 20590 3913
rect 20534 3839 20590 3848
rect 20444 3732 20496 3738
rect 20444 3674 20496 3680
rect 20444 3460 20496 3466
rect 20364 3420 20444 3448
rect 20260 3402 20312 3408
rect 20444 3402 20496 3408
rect 20352 3052 20404 3058
rect 20352 2994 20404 3000
rect 20076 2984 20128 2990
rect 20076 2926 20128 2932
rect 20168 2984 20220 2990
rect 20364 2961 20392 2994
rect 20168 2926 20220 2932
rect 20350 2952 20406 2961
rect 20456 2922 20484 3402
rect 20732 3058 20760 4422
rect 20824 4282 20852 5120
rect 20996 5102 21048 5108
rect 20904 5024 20956 5030
rect 20904 4966 20956 4972
rect 20916 4690 20944 4966
rect 20904 4684 20956 4690
rect 20904 4626 20956 4632
rect 20812 4276 20864 4282
rect 20812 4218 20864 4224
rect 20916 4146 20944 4626
rect 20904 4140 20956 4146
rect 20904 4082 20956 4088
rect 20810 3904 20866 3913
rect 20810 3839 20866 3848
rect 20824 3738 20852 3839
rect 20812 3732 20864 3738
rect 20812 3674 20864 3680
rect 21008 3602 21036 5102
rect 21180 4684 21232 4690
rect 21180 4626 21232 4632
rect 21086 4176 21142 4185
rect 21192 4146 21220 4626
rect 21272 4616 21324 4622
rect 21272 4558 21324 4564
rect 21086 4111 21088 4120
rect 21140 4111 21142 4120
rect 21180 4140 21232 4146
rect 21088 4082 21140 4088
rect 21180 4082 21232 4088
rect 21284 3602 21312 4558
rect 20996 3596 21048 3602
rect 20996 3538 21048 3544
rect 21272 3596 21324 3602
rect 21272 3538 21324 3544
rect 21284 3194 21312 3538
rect 21376 3534 21404 6938
rect 21652 6254 21680 8570
rect 21744 8537 21772 8792
rect 21824 8774 21876 8780
rect 22006 8800 22062 8809
rect 22006 8735 22062 8744
rect 21730 8528 21786 8537
rect 22020 8498 22048 8735
rect 21730 8463 21786 8472
rect 22008 8492 22060 8498
rect 21744 8430 21772 8463
rect 22008 8434 22060 8440
rect 22100 8492 22152 8498
rect 22100 8434 22152 8440
rect 21732 8424 21784 8430
rect 22112 8378 22140 8434
rect 22204 8430 22232 9998
rect 22480 9994 22508 11154
rect 22664 10674 22692 12854
rect 22756 12481 22784 13670
rect 22836 13252 22888 13258
rect 22836 13194 22888 13200
rect 22848 13161 22876 13194
rect 22834 13152 22890 13161
rect 22834 13087 22890 13096
rect 22848 12782 22876 13087
rect 22940 12986 22968 13738
rect 22928 12980 22980 12986
rect 22928 12922 22980 12928
rect 22836 12776 22888 12782
rect 22836 12718 22888 12724
rect 22742 12472 22798 12481
rect 22742 12407 22798 12416
rect 22756 11354 22784 12407
rect 22928 12300 22980 12306
rect 22928 12242 22980 12248
rect 22940 11354 22968 12242
rect 23032 11694 23060 13738
rect 23400 13394 23428 14214
rect 23480 13864 23532 13870
rect 23480 13806 23532 13812
rect 23388 13388 23440 13394
rect 23388 13330 23440 13336
rect 23296 13320 23348 13326
rect 23296 13262 23348 13268
rect 23308 12918 23336 13262
rect 23400 12986 23428 13330
rect 23388 12980 23440 12986
rect 23388 12922 23440 12928
rect 23296 12912 23348 12918
rect 23296 12854 23348 12860
rect 23112 12368 23164 12374
rect 23112 12310 23164 12316
rect 23124 12170 23152 12310
rect 23296 12232 23348 12238
rect 23492 12209 23520 13806
rect 23296 12174 23348 12180
rect 23478 12200 23534 12209
rect 23112 12164 23164 12170
rect 23112 12106 23164 12112
rect 23308 11694 23336 12174
rect 23478 12135 23534 12144
rect 23020 11688 23072 11694
rect 23296 11688 23348 11694
rect 23020 11630 23072 11636
rect 23202 11656 23258 11665
rect 23032 11558 23060 11630
rect 23296 11630 23348 11636
rect 23202 11591 23258 11600
rect 23020 11552 23072 11558
rect 23020 11494 23072 11500
rect 22744 11348 22796 11354
rect 22744 11290 22796 11296
rect 22928 11348 22980 11354
rect 22928 11290 22980 11296
rect 22926 11248 22982 11257
rect 22926 11183 22982 11192
rect 22940 10742 22968 11183
rect 22928 10736 22980 10742
rect 22928 10678 22980 10684
rect 22652 10668 22704 10674
rect 22652 10610 22704 10616
rect 23032 10266 23060 11494
rect 23216 11354 23244 11591
rect 23492 11354 23520 12135
rect 23204 11348 23256 11354
rect 23204 11290 23256 11296
rect 23480 11348 23532 11354
rect 23480 11290 23532 11296
rect 23584 11286 23612 14214
rect 24122 14175 24178 14184
rect 24136 14074 24164 14175
rect 24124 14068 24176 14074
rect 24124 14010 24176 14016
rect 24492 14000 24544 14006
rect 24492 13942 24544 13948
rect 24216 13320 24268 13326
rect 24216 13262 24268 13268
rect 23664 13252 23716 13258
rect 23664 13194 23716 13200
rect 23676 12782 23704 13194
rect 24228 13190 24256 13262
rect 24216 13184 24268 13190
rect 24216 13126 24268 13132
rect 24228 12986 24256 13126
rect 24216 12980 24268 12986
rect 24216 12922 24268 12928
rect 23664 12776 23716 12782
rect 23664 12718 23716 12724
rect 24504 12442 24532 13942
rect 24872 13938 24900 14418
rect 25044 14408 25096 14414
rect 25044 14350 25096 14356
rect 24860 13932 24912 13938
rect 24860 13874 24912 13880
rect 25056 13530 25084 14350
rect 25148 13802 25176 14418
rect 25240 14006 25268 14962
rect 25780 14476 25832 14482
rect 25780 14418 25832 14424
rect 25792 14278 25820 14418
rect 25780 14272 25832 14278
rect 25780 14214 25832 14220
rect 25228 14000 25280 14006
rect 25228 13942 25280 13948
rect 25136 13796 25188 13802
rect 25136 13738 25188 13744
rect 25044 13524 25096 13530
rect 25044 13466 25096 13472
rect 24860 13184 24912 13190
rect 24860 13126 24912 13132
rect 24872 12782 24900 13126
rect 24860 12776 24912 12782
rect 24860 12718 24912 12724
rect 24768 12640 24820 12646
rect 24768 12582 24820 12588
rect 24492 12436 24544 12442
rect 24492 12378 24544 12384
rect 23940 12368 23992 12374
rect 23940 12310 23992 12316
rect 23848 12300 23900 12306
rect 23848 12242 23900 12248
rect 23662 12064 23718 12073
rect 23662 11999 23718 12008
rect 23572 11280 23624 11286
rect 23572 11222 23624 11228
rect 23676 11218 23704 11999
rect 23860 11898 23888 12242
rect 23848 11892 23900 11898
rect 23848 11834 23900 11840
rect 23952 11762 23980 12310
rect 24216 12164 24268 12170
rect 24216 12106 24268 12112
rect 24124 12096 24176 12102
rect 24124 12038 24176 12044
rect 23940 11756 23992 11762
rect 23940 11698 23992 11704
rect 24136 11626 24164 12038
rect 24124 11620 24176 11626
rect 24124 11562 24176 11568
rect 23480 11212 23532 11218
rect 23480 11154 23532 11160
rect 23664 11212 23716 11218
rect 23664 11154 23716 11160
rect 23492 10742 23520 11154
rect 24136 11121 24164 11562
rect 24122 11112 24178 11121
rect 24122 11047 24178 11056
rect 23480 10736 23532 10742
rect 23478 10704 23480 10713
rect 23532 10704 23534 10713
rect 23478 10639 23534 10648
rect 23204 10600 23256 10606
rect 23204 10542 23256 10548
rect 23020 10260 23072 10266
rect 23020 10202 23072 10208
rect 23216 10130 23244 10542
rect 23204 10124 23256 10130
rect 23204 10066 23256 10072
rect 22468 9988 22520 9994
rect 22468 9930 22520 9936
rect 23216 9722 23244 10066
rect 23940 9920 23992 9926
rect 23940 9862 23992 9868
rect 23386 9752 23442 9761
rect 23204 9716 23256 9722
rect 23386 9687 23442 9696
rect 23204 9658 23256 9664
rect 23400 9654 23428 9687
rect 23388 9648 23440 9654
rect 23294 9616 23350 9625
rect 23388 9590 23440 9596
rect 23294 9551 23350 9560
rect 23112 9512 23164 9518
rect 23112 9454 23164 9460
rect 23020 9376 23072 9382
rect 23020 9318 23072 9324
rect 22376 9036 22428 9042
rect 22376 8978 22428 8984
rect 22284 8968 22336 8974
rect 22284 8910 22336 8916
rect 21732 8366 21784 8372
rect 22020 8362 22140 8378
rect 22192 8424 22244 8430
rect 22192 8366 22244 8372
rect 22296 8362 22324 8910
rect 22388 8634 22416 8978
rect 22560 8968 22612 8974
rect 22560 8910 22612 8916
rect 22572 8809 22600 8910
rect 22558 8800 22614 8809
rect 22558 8735 22614 8744
rect 22376 8628 22428 8634
rect 22376 8570 22428 8576
rect 22008 8356 22140 8362
rect 22060 8350 22140 8356
rect 22284 8356 22336 8362
rect 22008 8298 22060 8304
rect 22284 8298 22336 8304
rect 21748 8188 22044 8208
rect 21804 8186 21828 8188
rect 21884 8186 21908 8188
rect 21964 8186 21988 8188
rect 21826 8134 21828 8186
rect 21890 8134 21902 8186
rect 21964 8134 21966 8186
rect 21804 8132 21828 8134
rect 21884 8132 21908 8134
rect 21964 8132 21988 8134
rect 21748 8112 22044 8132
rect 22284 7744 22336 7750
rect 22098 7712 22154 7721
rect 22388 7732 22416 8570
rect 22744 8356 22796 8362
rect 22744 8298 22796 8304
rect 22336 7704 22416 7732
rect 22468 7744 22520 7750
rect 22284 7686 22336 7692
rect 22468 7686 22520 7692
rect 22098 7647 22154 7656
rect 22112 7342 22140 7647
rect 22100 7336 22152 7342
rect 22100 7278 22152 7284
rect 22284 7268 22336 7274
rect 22284 7210 22336 7216
rect 21748 7100 22044 7120
rect 21804 7098 21828 7100
rect 21884 7098 21908 7100
rect 21964 7098 21988 7100
rect 21826 7046 21828 7098
rect 21890 7046 21902 7098
rect 21964 7046 21966 7098
rect 21804 7044 21828 7046
rect 21884 7044 21908 7046
rect 21964 7044 21988 7046
rect 21748 7024 22044 7044
rect 21824 6792 21876 6798
rect 21822 6760 21824 6769
rect 21876 6760 21878 6769
rect 21822 6695 21878 6704
rect 21640 6248 21692 6254
rect 21640 6190 21692 6196
rect 21548 5772 21600 5778
rect 21548 5714 21600 5720
rect 21560 5234 21588 5714
rect 21548 5228 21600 5234
rect 21548 5170 21600 5176
rect 21548 4820 21600 4826
rect 21548 4762 21600 4768
rect 21560 4554 21588 4762
rect 21548 4548 21600 4554
rect 21548 4490 21600 4496
rect 21364 3528 21416 3534
rect 21364 3470 21416 3476
rect 21272 3188 21324 3194
rect 21272 3130 21324 3136
rect 20720 3052 20772 3058
rect 20720 2994 20772 3000
rect 20350 2887 20406 2896
rect 20444 2916 20496 2922
rect 20444 2858 20496 2864
rect 20720 2848 20772 2854
rect 20720 2790 20772 2796
rect 19984 2508 20036 2514
rect 19984 2450 20036 2456
rect 19996 2038 20024 2450
rect 19984 2032 20036 2038
rect 19984 1974 20036 1980
rect 19812 1414 19932 1442
rect 19812 800 19840 1414
rect 20732 800 20760 2790
rect 21376 2428 21404 3470
rect 21548 3120 21600 3126
rect 21548 3062 21600 3068
rect 21560 2514 21588 3062
rect 21548 2508 21600 2514
rect 21548 2450 21600 2456
rect 21456 2440 21508 2446
rect 21376 2400 21456 2428
rect 21456 2382 21508 2388
rect 21468 1834 21496 2382
rect 21456 1828 21508 1834
rect 21456 1770 21508 1776
rect 21652 800 21680 6190
rect 21836 6186 21864 6695
rect 21824 6180 21876 6186
rect 21824 6122 21876 6128
rect 21748 6012 22044 6032
rect 21804 6010 21828 6012
rect 21884 6010 21908 6012
rect 21964 6010 21988 6012
rect 21826 5958 21828 6010
rect 21890 5958 21902 6010
rect 21964 5958 21966 6010
rect 21804 5956 21828 5958
rect 21884 5956 21908 5958
rect 21964 5956 21988 5958
rect 21748 5936 22044 5956
rect 22100 5908 22152 5914
rect 22100 5850 22152 5856
rect 21732 5568 21784 5574
rect 21784 5528 22048 5556
rect 21732 5510 21784 5516
rect 22020 5522 22048 5528
rect 22112 5522 22140 5850
rect 22020 5494 22140 5522
rect 21914 5400 21970 5409
rect 21914 5335 21970 5344
rect 22190 5400 22246 5409
rect 22190 5335 22192 5344
rect 21928 5302 21956 5335
rect 22244 5335 22246 5344
rect 22192 5306 22244 5312
rect 21916 5296 21968 5302
rect 21916 5238 21968 5244
rect 22296 5234 22324 7210
rect 22480 6662 22508 7686
rect 22558 6896 22614 6905
rect 22558 6831 22560 6840
rect 22612 6831 22614 6840
rect 22652 6860 22704 6866
rect 22560 6802 22612 6808
rect 22652 6802 22704 6808
rect 22468 6656 22520 6662
rect 22468 6598 22520 6604
rect 22664 6322 22692 6802
rect 22652 6316 22704 6322
rect 22652 6258 22704 6264
rect 22652 5772 22704 5778
rect 22652 5714 22704 5720
rect 22376 5636 22428 5642
rect 22376 5578 22428 5584
rect 22388 5409 22416 5578
rect 22374 5400 22430 5409
rect 22374 5335 22430 5344
rect 22284 5228 22336 5234
rect 22284 5170 22336 5176
rect 22664 5166 22692 5714
rect 22468 5160 22520 5166
rect 22468 5102 22520 5108
rect 22652 5160 22704 5166
rect 22652 5102 22704 5108
rect 22192 5092 22244 5098
rect 22192 5034 22244 5040
rect 21748 4924 22044 4944
rect 21804 4922 21828 4924
rect 21884 4922 21908 4924
rect 21964 4922 21988 4924
rect 21826 4870 21828 4922
rect 21890 4870 21902 4922
rect 21964 4870 21966 4922
rect 21804 4868 21828 4870
rect 21884 4868 21908 4870
rect 21964 4868 21988 4870
rect 21748 4848 22044 4868
rect 22204 4758 22232 5034
rect 22284 5024 22336 5030
rect 22284 4966 22336 4972
rect 22192 4752 22244 4758
rect 22192 4694 22244 4700
rect 22192 4480 22244 4486
rect 22192 4422 22244 4428
rect 22204 4282 22232 4422
rect 22192 4276 22244 4282
rect 22192 4218 22244 4224
rect 22006 4176 22062 4185
rect 22006 4111 22008 4120
rect 22060 4111 22062 4120
rect 22100 4140 22152 4146
rect 22008 4082 22060 4088
rect 22100 4082 22152 4088
rect 21748 3836 22044 3856
rect 21804 3834 21828 3836
rect 21884 3834 21908 3836
rect 21964 3834 21988 3836
rect 21826 3782 21828 3834
rect 21890 3782 21902 3834
rect 21964 3782 21966 3834
rect 21804 3780 21828 3782
rect 21884 3780 21908 3782
rect 21964 3780 21988 3782
rect 21748 3760 22044 3780
rect 21824 3392 21876 3398
rect 21824 3334 21876 3340
rect 21836 3126 21864 3334
rect 21824 3120 21876 3126
rect 21824 3062 21876 3068
rect 22112 3058 22140 4082
rect 22204 4010 22232 4218
rect 22192 4004 22244 4010
rect 22192 3946 22244 3952
rect 22190 3904 22246 3913
rect 22190 3839 22246 3848
rect 22100 3052 22152 3058
rect 22100 2994 22152 3000
rect 22204 2854 22232 3839
rect 22296 3040 22324 4966
rect 22480 4128 22508 5102
rect 22560 5024 22612 5030
rect 22560 4966 22612 4972
rect 22388 4100 22508 4128
rect 22388 3942 22416 4100
rect 22376 3936 22428 3942
rect 22376 3878 22428 3884
rect 22388 3738 22416 3878
rect 22376 3732 22428 3738
rect 22376 3674 22428 3680
rect 22468 3460 22520 3466
rect 22468 3402 22520 3408
rect 22376 3052 22428 3058
rect 22296 3012 22376 3040
rect 22376 2994 22428 3000
rect 22192 2848 22244 2854
rect 22192 2790 22244 2796
rect 21748 2748 22044 2768
rect 21804 2746 21828 2748
rect 21884 2746 21908 2748
rect 21964 2746 21988 2748
rect 21826 2694 21828 2746
rect 21890 2694 21902 2746
rect 21964 2694 21966 2746
rect 21804 2692 21828 2694
rect 21884 2692 21908 2694
rect 21964 2692 21988 2694
rect 21748 2672 22044 2692
rect 22388 2446 22416 2994
rect 22376 2440 22428 2446
rect 22376 2382 22428 2388
rect 22480 800 22508 3402
rect 22572 2990 22600 4966
rect 22664 4486 22692 5102
rect 22652 4480 22704 4486
rect 22652 4422 22704 4428
rect 22652 4072 22704 4078
rect 22756 4060 22784 8298
rect 22836 6656 22888 6662
rect 22836 6598 22888 6604
rect 22928 6656 22980 6662
rect 22928 6598 22980 6604
rect 22848 5914 22876 6598
rect 22940 6390 22968 6598
rect 22928 6384 22980 6390
rect 22928 6326 22980 6332
rect 22836 5908 22888 5914
rect 22836 5850 22888 5856
rect 22928 5772 22980 5778
rect 22928 5714 22980 5720
rect 22940 5234 22968 5714
rect 22836 5228 22888 5234
rect 22836 5170 22888 5176
rect 22928 5228 22980 5234
rect 22928 5170 22980 5176
rect 22704 4032 22784 4060
rect 22652 4014 22704 4020
rect 22664 3942 22692 4014
rect 22652 3936 22704 3942
rect 22652 3878 22704 3884
rect 22664 3194 22692 3878
rect 22744 3392 22796 3398
rect 22744 3334 22796 3340
rect 22652 3188 22704 3194
rect 22652 3130 22704 3136
rect 22756 2990 22784 3334
rect 22848 3233 22876 5170
rect 22928 4684 22980 4690
rect 23032 4672 23060 9318
rect 23124 9178 23152 9454
rect 23112 9172 23164 9178
rect 23112 9114 23164 9120
rect 23308 8294 23336 9551
rect 23952 8974 23980 9862
rect 24136 9489 24164 11047
rect 24228 10266 24256 12106
rect 24504 11694 24532 12378
rect 24492 11688 24544 11694
rect 24492 11630 24544 11636
rect 24780 11286 24808 12582
rect 24872 12442 24900 12718
rect 25318 12608 25374 12617
rect 25318 12543 25374 12552
rect 24860 12436 24912 12442
rect 24860 12378 24912 12384
rect 25332 12306 25360 12543
rect 25792 12442 25820 14214
rect 25976 12782 26004 15302
rect 26068 14958 26096 15574
rect 27080 15570 27108 15982
rect 27540 15638 27568 17138
rect 28356 17128 28408 17134
rect 28356 17070 28408 17076
rect 28724 17128 28776 17134
rect 28724 17070 28776 17076
rect 27620 16584 27672 16590
rect 27620 16526 27672 16532
rect 27632 16182 27660 16526
rect 27620 16176 27672 16182
rect 27620 16118 27672 16124
rect 27632 15638 27660 16118
rect 28368 16114 28396 17070
rect 28736 16454 28764 17070
rect 28724 16448 28776 16454
rect 28724 16390 28776 16396
rect 28356 16108 28408 16114
rect 28356 16050 28408 16056
rect 28264 16040 28316 16046
rect 28264 15982 28316 15988
rect 27712 15904 27764 15910
rect 27712 15846 27764 15852
rect 27160 15632 27212 15638
rect 27160 15574 27212 15580
rect 27528 15632 27580 15638
rect 27528 15574 27580 15580
rect 27620 15632 27672 15638
rect 27620 15574 27672 15580
rect 27068 15564 27120 15570
rect 27068 15506 27120 15512
rect 27080 15094 27108 15506
rect 27068 15088 27120 15094
rect 27068 15030 27120 15036
rect 26056 14952 26108 14958
rect 26056 14894 26108 14900
rect 26424 14884 26476 14890
rect 26424 14826 26476 14832
rect 26436 14550 26464 14826
rect 26424 14544 26476 14550
rect 26424 14486 26476 14492
rect 27172 14482 27200 15574
rect 27436 15496 27488 15502
rect 27436 15438 27488 15444
rect 27448 15094 27476 15438
rect 27436 15088 27488 15094
rect 27436 15030 27488 15036
rect 27344 14952 27396 14958
rect 27344 14894 27396 14900
rect 27160 14476 27212 14482
rect 27160 14418 27212 14424
rect 27356 14278 27384 14894
rect 26240 14272 26292 14278
rect 26240 14214 26292 14220
rect 26792 14272 26844 14278
rect 26792 14214 26844 14220
rect 27344 14272 27396 14278
rect 27344 14214 27396 14220
rect 26252 14113 26280 14214
rect 26238 14104 26294 14113
rect 26056 14068 26108 14074
rect 26238 14039 26294 14048
rect 26056 14010 26108 14016
rect 26068 13394 26096 14010
rect 26252 13938 26280 14039
rect 26240 13932 26292 13938
rect 26240 13874 26292 13880
rect 26240 13796 26292 13802
rect 26240 13738 26292 13744
rect 26252 13530 26280 13738
rect 26240 13524 26292 13530
rect 26240 13466 26292 13472
rect 26056 13388 26108 13394
rect 26056 13330 26108 13336
rect 26068 12918 26096 13330
rect 26332 13184 26384 13190
rect 26804 13161 26832 14214
rect 27356 13938 27384 14214
rect 27448 14006 27476 15030
rect 27528 14408 27580 14414
rect 27528 14350 27580 14356
rect 27436 14000 27488 14006
rect 27436 13942 27488 13948
rect 27344 13932 27396 13938
rect 27344 13874 27396 13880
rect 27160 13252 27212 13258
rect 27160 13194 27212 13200
rect 26332 13126 26384 13132
rect 26790 13152 26846 13161
rect 26238 13016 26294 13025
rect 26238 12951 26294 12960
rect 26056 12912 26108 12918
rect 26056 12854 26108 12860
rect 25964 12776 26016 12782
rect 25884 12736 25964 12764
rect 25780 12436 25832 12442
rect 25780 12378 25832 12384
rect 24952 12300 25004 12306
rect 24952 12242 25004 12248
rect 25320 12300 25372 12306
rect 25320 12242 25372 12248
rect 24964 11558 24992 12242
rect 25780 12096 25832 12102
rect 25780 12038 25832 12044
rect 25792 11762 25820 12038
rect 25780 11756 25832 11762
rect 25780 11698 25832 11704
rect 25136 11620 25188 11626
rect 25136 11562 25188 11568
rect 24952 11552 25004 11558
rect 24952 11494 25004 11500
rect 24768 11280 24820 11286
rect 24768 11222 24820 11228
rect 25148 11218 25176 11562
rect 25412 11552 25464 11558
rect 25464 11500 25544 11506
rect 25412 11494 25544 11500
rect 25424 11478 25544 11494
rect 24860 11212 24912 11218
rect 24860 11154 24912 11160
rect 25136 11212 25188 11218
rect 25136 11154 25188 11160
rect 24676 11008 24728 11014
rect 24676 10950 24728 10956
rect 24688 10606 24716 10950
rect 24676 10600 24728 10606
rect 24676 10542 24728 10548
rect 24872 10266 24900 11154
rect 25320 11144 25372 11150
rect 25320 11086 25372 11092
rect 24952 11076 25004 11082
rect 24952 11018 25004 11024
rect 24964 10606 24992 11018
rect 25044 10736 25096 10742
rect 25044 10678 25096 10684
rect 24952 10600 25004 10606
rect 24952 10542 25004 10548
rect 24216 10260 24268 10266
rect 24216 10202 24268 10208
rect 24860 10260 24912 10266
rect 24860 10202 24912 10208
rect 25056 9654 25084 10678
rect 25332 9926 25360 11086
rect 25320 9920 25372 9926
rect 25320 9862 25372 9868
rect 25044 9648 25096 9654
rect 24950 9616 25006 9625
rect 25044 9590 25096 9596
rect 24950 9551 25006 9560
rect 24964 9518 24992 9551
rect 24952 9512 25004 9518
rect 24122 9480 24178 9489
rect 24952 9454 25004 9460
rect 24122 9415 24178 9424
rect 24860 9376 24912 9382
rect 24860 9318 24912 9324
rect 24872 9110 24900 9318
rect 24860 9104 24912 9110
rect 24860 9046 24912 9052
rect 24400 9036 24452 9042
rect 24400 8978 24452 8984
rect 23940 8968 23992 8974
rect 23940 8910 23992 8916
rect 23480 8832 23532 8838
rect 23480 8774 23532 8780
rect 23492 8430 23520 8774
rect 23480 8424 23532 8430
rect 23480 8366 23532 8372
rect 23296 8288 23348 8294
rect 23296 8230 23348 8236
rect 23308 7750 23336 8230
rect 23296 7744 23348 7750
rect 23296 7686 23348 7692
rect 23112 7200 23164 7206
rect 23112 7142 23164 7148
rect 23124 6089 23152 7142
rect 23308 7002 23336 7686
rect 23492 7546 23520 8366
rect 23480 7540 23532 7546
rect 23480 7482 23532 7488
rect 23848 7336 23900 7342
rect 23848 7278 23900 7284
rect 23296 6996 23348 7002
rect 23296 6938 23348 6944
rect 23756 6724 23808 6730
rect 23756 6666 23808 6672
rect 23768 6254 23796 6666
rect 23756 6248 23808 6254
rect 23756 6190 23808 6196
rect 23664 6112 23716 6118
rect 23110 6080 23166 6089
rect 23664 6054 23716 6060
rect 23110 6015 23166 6024
rect 23676 5914 23704 6054
rect 23112 5908 23164 5914
rect 23112 5850 23164 5856
rect 23664 5908 23716 5914
rect 23664 5850 23716 5856
rect 22980 4644 23060 4672
rect 22928 4626 22980 4632
rect 22940 3913 22968 4626
rect 23020 4480 23072 4486
rect 23020 4422 23072 4428
rect 22926 3904 22982 3913
rect 22926 3839 22982 3848
rect 23032 3738 23060 4422
rect 23124 3738 23152 5850
rect 23204 5704 23256 5710
rect 23202 5672 23204 5681
rect 23256 5672 23258 5681
rect 23202 5607 23258 5616
rect 23860 4690 23888 7278
rect 23952 7206 23980 8910
rect 24412 8838 24440 8978
rect 24400 8832 24452 8838
rect 24400 8774 24452 8780
rect 24412 8022 24440 8774
rect 24964 8566 24992 9454
rect 25320 9376 25372 9382
rect 25240 9324 25320 9330
rect 25240 9318 25372 9324
rect 25240 9302 25360 9318
rect 25044 9036 25096 9042
rect 25044 8978 25096 8984
rect 24952 8560 25004 8566
rect 24766 8528 24822 8537
rect 24952 8502 25004 8508
rect 24766 8463 24822 8472
rect 24400 8016 24452 8022
rect 24400 7958 24452 7964
rect 24492 8016 24544 8022
rect 24492 7958 24544 7964
rect 24308 7948 24360 7954
rect 24308 7890 24360 7896
rect 24320 7342 24348 7890
rect 24504 7342 24532 7958
rect 24780 7478 24808 8463
rect 25056 8294 25084 8978
rect 25240 8430 25268 9302
rect 25412 9036 25464 9042
rect 25412 8978 25464 8984
rect 25424 8634 25452 8978
rect 25412 8628 25464 8634
rect 25412 8570 25464 8576
rect 25228 8424 25280 8430
rect 25228 8366 25280 8372
rect 24952 8288 25004 8294
rect 24950 8256 24952 8265
rect 25044 8288 25096 8294
rect 25004 8256 25006 8265
rect 25044 8230 25096 8236
rect 24950 8191 25006 8200
rect 24860 7812 24912 7818
rect 24860 7754 24912 7760
rect 24768 7472 24820 7478
rect 24768 7414 24820 7420
rect 24308 7336 24360 7342
rect 24308 7278 24360 7284
rect 24492 7336 24544 7342
rect 24492 7278 24544 7284
rect 23940 7200 23992 7206
rect 23940 7142 23992 7148
rect 24320 7002 24348 7278
rect 24124 6996 24176 7002
rect 24124 6938 24176 6944
rect 24308 6996 24360 7002
rect 24308 6938 24360 6944
rect 24032 6860 24084 6866
rect 24032 6802 24084 6808
rect 24044 6390 24072 6802
rect 24032 6384 24084 6390
rect 24032 6326 24084 6332
rect 24044 5914 24072 6326
rect 24032 5908 24084 5914
rect 24032 5850 24084 5856
rect 24032 5772 24084 5778
rect 24032 5714 24084 5720
rect 23938 5672 23994 5681
rect 23938 5607 23994 5616
rect 23952 5574 23980 5607
rect 24044 5574 24072 5714
rect 23940 5568 23992 5574
rect 23940 5510 23992 5516
rect 24032 5568 24084 5574
rect 24032 5510 24084 5516
rect 24136 5234 24164 6938
rect 24308 6860 24360 6866
rect 24308 6802 24360 6808
rect 24320 6662 24348 6802
rect 24872 6798 24900 7754
rect 25056 7721 25084 8230
rect 25240 7886 25268 8366
rect 25320 8288 25372 8294
rect 25320 8230 25372 8236
rect 25228 7880 25280 7886
rect 25228 7822 25280 7828
rect 25332 7750 25360 8230
rect 25320 7744 25372 7750
rect 25042 7712 25098 7721
rect 25320 7686 25372 7692
rect 25042 7647 25098 7656
rect 25056 7426 25084 7647
rect 25332 7546 25360 7686
rect 25320 7540 25372 7546
rect 25320 7482 25372 7488
rect 24964 7398 25084 7426
rect 24860 6792 24912 6798
rect 24860 6734 24912 6740
rect 24676 6724 24728 6730
rect 24676 6666 24728 6672
rect 24308 6656 24360 6662
rect 24308 6598 24360 6604
rect 24214 5944 24270 5953
rect 24214 5879 24270 5888
rect 24228 5370 24256 5879
rect 24216 5364 24268 5370
rect 24216 5306 24268 5312
rect 24124 5228 24176 5234
rect 24124 5170 24176 5176
rect 23940 4820 23992 4826
rect 23940 4762 23992 4768
rect 23848 4684 23900 4690
rect 23848 4626 23900 4632
rect 23664 4480 23716 4486
rect 23664 4422 23716 4428
rect 23754 4448 23810 4457
rect 23572 4276 23624 4282
rect 23572 4218 23624 4224
rect 23388 3936 23440 3942
rect 23386 3904 23388 3913
rect 23584 3913 23612 4218
rect 23440 3904 23442 3913
rect 23386 3839 23442 3848
rect 23570 3904 23626 3913
rect 23570 3839 23626 3848
rect 23020 3732 23072 3738
rect 23020 3674 23072 3680
rect 23112 3732 23164 3738
rect 23112 3674 23164 3680
rect 22834 3224 22890 3233
rect 22834 3159 22890 3168
rect 22560 2984 22612 2990
rect 22558 2952 22560 2961
rect 22744 2984 22796 2990
rect 22612 2952 22614 2961
rect 22744 2926 22796 2932
rect 22558 2887 22614 2896
rect 22572 2854 22600 2887
rect 22560 2848 22612 2854
rect 22560 2790 22612 2796
rect 22756 2310 22784 2926
rect 22836 2916 22888 2922
rect 22836 2858 22888 2864
rect 22848 2310 22876 2858
rect 23032 2582 23060 3674
rect 23124 3058 23152 3674
rect 23676 3670 23704 4422
rect 23754 4383 23810 4392
rect 23768 3670 23796 4383
rect 23860 4282 23888 4626
rect 23952 4282 23980 4762
rect 23848 4276 23900 4282
rect 23848 4218 23900 4224
rect 23940 4276 23992 4282
rect 23940 4218 23992 4224
rect 23860 3738 23888 4218
rect 23848 3732 23900 3738
rect 23848 3674 23900 3680
rect 23664 3664 23716 3670
rect 23664 3606 23716 3612
rect 23756 3664 23808 3670
rect 23756 3606 23808 3612
rect 23572 3596 23624 3602
rect 23572 3538 23624 3544
rect 23388 3528 23440 3534
rect 23386 3496 23388 3505
rect 23440 3496 23442 3505
rect 23442 3454 23520 3482
rect 23386 3431 23442 3440
rect 23492 3194 23520 3454
rect 23480 3188 23532 3194
rect 23480 3130 23532 3136
rect 23112 3052 23164 3058
rect 23112 2994 23164 3000
rect 23388 2848 23440 2854
rect 23388 2790 23440 2796
rect 23020 2576 23072 2582
rect 23020 2518 23072 2524
rect 22744 2304 22796 2310
rect 22744 2246 22796 2252
rect 22836 2304 22888 2310
rect 22836 2246 22888 2252
rect 23400 800 23428 2790
rect 23492 2582 23520 3130
rect 23584 3058 23612 3538
rect 23768 3534 23796 3606
rect 23756 3528 23808 3534
rect 23756 3470 23808 3476
rect 23572 3052 23624 3058
rect 23572 2994 23624 3000
rect 23480 2576 23532 2582
rect 23480 2518 23532 2524
rect 24136 2378 24164 5170
rect 24228 5166 24256 5306
rect 24216 5160 24268 5166
rect 24216 5102 24268 5108
rect 24228 4826 24256 5102
rect 24216 4820 24268 4826
rect 24216 4762 24268 4768
rect 24320 4078 24348 6598
rect 24584 6316 24636 6322
rect 24584 6258 24636 6264
rect 24596 6202 24624 6258
rect 24504 6174 24624 6202
rect 24504 6118 24532 6174
rect 24688 6168 24716 6666
rect 24860 6656 24912 6662
rect 24860 6598 24912 6604
rect 24872 6390 24900 6598
rect 24860 6384 24912 6390
rect 24860 6326 24912 6332
rect 24860 6180 24912 6186
rect 24688 6140 24808 6168
rect 24492 6112 24544 6118
rect 24398 6080 24454 6089
rect 24492 6054 24544 6060
rect 24398 6015 24454 6024
rect 24412 5778 24440 6015
rect 24400 5772 24452 5778
rect 24400 5714 24452 5720
rect 24676 5772 24728 5778
rect 24676 5714 24728 5720
rect 24400 5636 24452 5642
rect 24400 5578 24452 5584
rect 24412 4826 24440 5578
rect 24688 5302 24716 5714
rect 24676 5296 24728 5302
rect 24676 5238 24728 5244
rect 24490 5128 24546 5137
rect 24490 5063 24546 5072
rect 24674 5128 24730 5137
rect 24674 5063 24730 5072
rect 24400 4820 24452 4826
rect 24400 4762 24452 4768
rect 24504 4690 24532 5063
rect 24492 4684 24544 4690
rect 24492 4626 24544 4632
rect 24492 4480 24544 4486
rect 24492 4422 24544 4428
rect 24308 4072 24360 4078
rect 24308 4014 24360 4020
rect 24504 3398 24532 4422
rect 24688 4078 24716 5063
rect 24780 4078 24808 6140
rect 24860 6122 24912 6128
rect 24872 5846 24900 6122
rect 24860 5840 24912 5846
rect 24860 5782 24912 5788
rect 24872 4826 24900 5782
rect 24860 4820 24912 4826
rect 24860 4762 24912 4768
rect 24964 4729 24992 7398
rect 25320 7336 25372 7342
rect 25320 7278 25372 7284
rect 25332 7206 25360 7278
rect 25320 7200 25372 7206
rect 25320 7142 25372 7148
rect 25332 6866 25360 7142
rect 25320 6860 25372 6866
rect 25320 6802 25372 6808
rect 25412 6792 25464 6798
rect 25412 6734 25464 6740
rect 25136 6724 25188 6730
rect 25136 6666 25188 6672
rect 25148 6322 25176 6666
rect 25136 6316 25188 6322
rect 25136 6258 25188 6264
rect 25320 6248 25372 6254
rect 25320 6190 25372 6196
rect 25332 5846 25360 6190
rect 25320 5840 25372 5846
rect 25320 5782 25372 5788
rect 25044 5704 25096 5710
rect 25044 5646 25096 5652
rect 25056 5234 25084 5646
rect 25044 5228 25096 5234
rect 25044 5170 25096 5176
rect 25228 5228 25280 5234
rect 25228 5170 25280 5176
rect 24950 4720 25006 4729
rect 24950 4655 25006 4664
rect 25136 4684 25188 4690
rect 25136 4626 25188 4632
rect 24676 4072 24728 4078
rect 24676 4014 24728 4020
rect 24768 4072 24820 4078
rect 24768 4014 24820 4020
rect 25148 4010 25176 4626
rect 25136 4004 25188 4010
rect 25136 3946 25188 3952
rect 24952 3936 25004 3942
rect 24952 3878 25004 3884
rect 24860 3596 24912 3602
rect 24860 3538 24912 3544
rect 24584 3528 24636 3534
rect 24768 3528 24820 3534
rect 24584 3470 24636 3476
rect 24674 3496 24730 3505
rect 24596 3398 24624 3470
rect 24768 3470 24820 3476
rect 24674 3431 24730 3440
rect 24492 3392 24544 3398
rect 24492 3334 24544 3340
rect 24584 3392 24636 3398
rect 24584 3334 24636 3340
rect 24504 3126 24532 3334
rect 24492 3120 24544 3126
rect 24492 3062 24544 3068
rect 24596 2990 24624 3334
rect 24688 3097 24716 3431
rect 24674 3088 24730 3097
rect 24674 3023 24730 3032
rect 24584 2984 24636 2990
rect 24398 2952 24454 2961
rect 24308 2916 24360 2922
rect 24584 2926 24636 2932
rect 24398 2887 24454 2896
rect 24308 2858 24360 2864
rect 24320 2514 24348 2858
rect 24308 2508 24360 2514
rect 24308 2450 24360 2456
rect 24124 2372 24176 2378
rect 24124 2314 24176 2320
rect 24412 1578 24440 2887
rect 24780 2310 24808 3470
rect 24872 2990 24900 3538
rect 24860 2984 24912 2990
rect 24860 2926 24912 2932
rect 24872 2650 24900 2926
rect 24860 2644 24912 2650
rect 24860 2586 24912 2592
rect 24768 2304 24820 2310
rect 24768 2246 24820 2252
rect 24320 1550 24440 1578
rect 24320 800 24348 1550
rect 24964 1358 24992 3878
rect 25044 3732 25096 3738
rect 25044 3674 25096 3680
rect 25056 2514 25084 3674
rect 25240 3670 25268 5170
rect 25320 4684 25372 4690
rect 25320 4626 25372 4632
rect 25332 4146 25360 4626
rect 25424 4146 25452 6734
rect 25516 4865 25544 11478
rect 25792 11286 25820 11698
rect 25884 11558 25912 12736
rect 25964 12718 26016 12724
rect 25962 12608 26018 12617
rect 25962 12543 26018 12552
rect 25872 11552 25924 11558
rect 25872 11494 25924 11500
rect 25780 11280 25832 11286
rect 25780 11222 25832 11228
rect 25884 11150 25912 11494
rect 25872 11144 25924 11150
rect 25872 11086 25924 11092
rect 25976 11014 26004 12543
rect 26252 12442 26280 12951
rect 26344 12850 26372 13126
rect 26790 13087 26846 13096
rect 26804 12889 26832 13087
rect 27172 12918 27200 13194
rect 27448 13190 27476 13942
rect 27540 13870 27568 14350
rect 27528 13864 27580 13870
rect 27528 13806 27580 13812
rect 27724 13530 27752 15846
rect 28172 15632 28224 15638
rect 28172 15574 28224 15580
rect 28080 15564 28132 15570
rect 28080 15506 28132 15512
rect 27804 14952 27856 14958
rect 27856 14900 27936 14906
rect 27804 14894 27936 14900
rect 27816 14890 27936 14894
rect 27816 14884 27948 14890
rect 27816 14878 27896 14884
rect 27896 14826 27948 14832
rect 27712 13524 27764 13530
rect 27712 13466 27764 13472
rect 27436 13184 27488 13190
rect 27436 13126 27488 13132
rect 27712 12980 27764 12986
rect 27712 12922 27764 12928
rect 27160 12912 27212 12918
rect 26790 12880 26846 12889
rect 26332 12844 26384 12850
rect 27160 12854 27212 12860
rect 26790 12815 26846 12824
rect 26332 12786 26384 12792
rect 27724 12442 27752 12922
rect 26056 12436 26108 12442
rect 26056 12378 26108 12384
rect 26240 12436 26292 12442
rect 26240 12378 26292 12384
rect 27712 12436 27764 12442
rect 27712 12378 27764 12384
rect 26068 11014 26096 12378
rect 26252 12306 26280 12378
rect 26240 12300 26292 12306
rect 26240 12242 26292 12248
rect 26792 12300 26844 12306
rect 26792 12242 26844 12248
rect 27252 12300 27304 12306
rect 27252 12242 27304 12248
rect 27344 12300 27396 12306
rect 27344 12242 27396 12248
rect 26804 11558 26832 12242
rect 27160 12164 27212 12170
rect 27160 12106 27212 12112
rect 27172 11762 27200 12106
rect 27264 11898 27292 12242
rect 27356 12186 27384 12242
rect 27356 12170 27752 12186
rect 27356 12164 27764 12170
rect 27356 12158 27712 12164
rect 27252 11892 27304 11898
rect 27252 11834 27304 11840
rect 27160 11756 27212 11762
rect 27160 11698 27212 11704
rect 26792 11552 26844 11558
rect 26792 11494 26844 11500
rect 27172 11218 27200 11698
rect 26332 11212 26384 11218
rect 26332 11154 26384 11160
rect 27160 11212 27212 11218
rect 27160 11154 27212 11160
rect 25780 11008 25832 11014
rect 25780 10950 25832 10956
rect 25964 11008 26016 11014
rect 25964 10950 26016 10956
rect 26056 11008 26108 11014
rect 26056 10950 26108 10956
rect 25792 10606 25820 10950
rect 25596 10600 25648 10606
rect 25596 10542 25648 10548
rect 25780 10600 25832 10606
rect 25780 10542 25832 10548
rect 25608 9926 25636 10542
rect 26068 10198 26096 10950
rect 26148 10532 26200 10538
rect 26148 10474 26200 10480
rect 26056 10192 26108 10198
rect 26056 10134 26108 10140
rect 25596 9920 25648 9926
rect 25596 9862 25648 9868
rect 26160 9586 26188 10474
rect 26344 10266 26372 11154
rect 27158 11112 27214 11121
rect 27158 11047 27214 11056
rect 27172 11014 27200 11047
rect 27160 11008 27212 11014
rect 27160 10950 27212 10956
rect 27172 10606 27200 10950
rect 27250 10704 27306 10713
rect 27250 10639 27306 10648
rect 27264 10606 27292 10639
rect 27160 10600 27212 10606
rect 27160 10542 27212 10548
rect 27252 10600 27304 10606
rect 27252 10542 27304 10548
rect 27172 10470 27200 10542
rect 27068 10464 27120 10470
rect 27068 10406 27120 10412
rect 27160 10464 27212 10470
rect 27160 10406 27212 10412
rect 27080 10282 27108 10406
rect 26332 10260 26384 10266
rect 27080 10254 27200 10282
rect 26332 10202 26384 10208
rect 26344 9994 26372 10202
rect 26332 9988 26384 9994
rect 26332 9930 26384 9936
rect 26792 9648 26844 9654
rect 26792 9590 26844 9596
rect 26148 9580 26200 9586
rect 26148 9522 26200 9528
rect 26160 9042 26188 9522
rect 26148 9036 26200 9042
rect 26148 8978 26200 8984
rect 26608 8900 26660 8906
rect 26608 8842 26660 8848
rect 25872 8832 25924 8838
rect 25872 8774 25924 8780
rect 26240 8832 26292 8838
rect 26240 8774 26292 8780
rect 25884 8430 25912 8774
rect 26252 8430 26280 8774
rect 26516 8628 26568 8634
rect 26516 8570 26568 8576
rect 26528 8430 26556 8570
rect 25872 8424 25924 8430
rect 25872 8366 25924 8372
rect 26240 8424 26292 8430
rect 26240 8366 26292 8372
rect 26516 8424 26568 8430
rect 26516 8366 26568 8372
rect 25884 8022 25912 8366
rect 25872 8016 25924 8022
rect 25872 7958 25924 7964
rect 26516 8016 26568 8022
rect 26516 7958 26568 7964
rect 25884 7750 25912 7958
rect 26332 7948 26384 7954
rect 26332 7890 26384 7896
rect 26240 7812 26292 7818
rect 26240 7754 26292 7760
rect 25780 7744 25832 7750
rect 25780 7686 25832 7692
rect 25872 7744 25924 7750
rect 25872 7686 25924 7692
rect 25792 7041 25820 7686
rect 25964 7336 26016 7342
rect 25964 7278 26016 7284
rect 25976 7206 26004 7278
rect 26252 7274 26280 7754
rect 26240 7268 26292 7274
rect 26240 7210 26292 7216
rect 25964 7200 26016 7206
rect 26344 7177 26372 7890
rect 26528 7546 26556 7958
rect 26516 7540 26568 7546
rect 26516 7482 26568 7488
rect 25964 7142 26016 7148
rect 26330 7168 26386 7177
rect 25778 7032 25834 7041
rect 25778 6967 25834 6976
rect 25780 6792 25832 6798
rect 25780 6734 25832 6740
rect 25792 6458 25820 6734
rect 25780 6452 25832 6458
rect 25780 6394 25832 6400
rect 25594 6352 25650 6361
rect 25594 6287 25650 6296
rect 25608 6254 25636 6287
rect 25596 6248 25648 6254
rect 25872 6248 25924 6254
rect 25596 6190 25648 6196
rect 25700 6196 25872 6202
rect 25700 6190 25924 6196
rect 25608 5846 25636 6190
rect 25700 6174 25912 6190
rect 25596 5840 25648 5846
rect 25596 5782 25648 5788
rect 25502 4856 25558 4865
rect 25502 4791 25558 4800
rect 25596 4208 25648 4214
rect 25596 4150 25648 4156
rect 25320 4140 25372 4146
rect 25320 4082 25372 4088
rect 25412 4140 25464 4146
rect 25412 4082 25464 4088
rect 25608 3942 25636 4150
rect 25596 3936 25648 3942
rect 25596 3878 25648 3884
rect 25608 3738 25636 3878
rect 25596 3732 25648 3738
rect 25596 3674 25648 3680
rect 25228 3664 25280 3670
rect 25228 3606 25280 3612
rect 25318 3632 25374 3641
rect 25134 3088 25190 3097
rect 25240 3058 25268 3606
rect 25318 3567 25320 3576
rect 25372 3567 25374 3576
rect 25320 3538 25372 3544
rect 25332 3194 25360 3538
rect 25700 3369 25728 6174
rect 25976 5166 26004 7142
rect 26330 7103 26386 7112
rect 26422 7032 26478 7041
rect 26422 6967 26478 6976
rect 26332 6792 26384 6798
rect 26332 6734 26384 6740
rect 26240 6724 26292 6730
rect 26240 6666 26292 6672
rect 26252 5234 26280 6666
rect 26240 5228 26292 5234
rect 26240 5170 26292 5176
rect 25964 5160 26016 5166
rect 25964 5102 26016 5108
rect 25870 4856 25926 4865
rect 25870 4791 25926 4800
rect 25780 4616 25832 4622
rect 25780 4558 25832 4564
rect 25792 4486 25820 4558
rect 25780 4480 25832 4486
rect 25780 4422 25832 4428
rect 25792 4146 25820 4422
rect 25884 4185 25912 4791
rect 25870 4176 25926 4185
rect 25780 4140 25832 4146
rect 25976 4162 26004 5102
rect 26056 5024 26108 5030
rect 26056 4966 26108 4972
rect 26068 4826 26096 4966
rect 26056 4820 26108 4826
rect 26056 4762 26108 4768
rect 25976 4134 26188 4162
rect 25870 4111 25926 4120
rect 25780 4082 25832 4088
rect 25686 3360 25742 3369
rect 25686 3295 25742 3304
rect 25320 3188 25372 3194
rect 25320 3130 25372 3136
rect 25134 3023 25190 3032
rect 25228 3052 25280 3058
rect 25044 2508 25096 2514
rect 25044 2450 25096 2456
rect 24952 1352 25004 1358
rect 24952 1294 25004 1300
rect 25148 800 25176 3023
rect 25228 2994 25280 3000
rect 25884 2378 25912 4111
rect 26160 3482 26188 4134
rect 26344 4078 26372 6734
rect 26436 5846 26464 6967
rect 26516 6928 26568 6934
rect 26516 6870 26568 6876
rect 26528 6322 26556 6870
rect 26516 6316 26568 6322
rect 26516 6258 26568 6264
rect 26424 5840 26476 5846
rect 26424 5782 26476 5788
rect 26620 5574 26648 8842
rect 26700 8560 26752 8566
rect 26700 8502 26752 8508
rect 26712 7886 26740 8502
rect 26700 7880 26752 7886
rect 26700 7822 26752 7828
rect 26700 6860 26752 6866
rect 26804 6848 26832 9590
rect 27068 9580 27120 9586
rect 27068 9522 27120 9528
rect 26976 8288 27028 8294
rect 26976 8230 27028 8236
rect 26988 7886 27016 8230
rect 26976 7880 27028 7886
rect 26976 7822 27028 7828
rect 27080 7392 27108 9522
rect 27172 8974 27200 10254
rect 27252 10056 27304 10062
rect 27252 9998 27304 10004
rect 27264 9654 27292 9998
rect 27252 9648 27304 9654
rect 27252 9590 27304 9596
rect 27356 9194 27384 12158
rect 27712 12106 27764 12112
rect 27434 11928 27490 11937
rect 27434 11863 27490 11872
rect 27448 11762 27476 11863
rect 27436 11756 27488 11762
rect 27436 11698 27488 11704
rect 27804 11688 27856 11694
rect 27804 11630 27856 11636
rect 27528 11552 27580 11558
rect 27528 11494 27580 11500
rect 27540 10606 27568 11494
rect 27816 11257 27844 11630
rect 27802 11248 27858 11257
rect 27802 11183 27858 11192
rect 27804 11144 27856 11150
rect 27804 11086 27856 11092
rect 27816 10674 27844 11086
rect 27804 10668 27856 10674
rect 27804 10610 27856 10616
rect 27528 10600 27580 10606
rect 27528 10542 27580 10548
rect 27436 10124 27488 10130
rect 27436 10066 27488 10072
rect 27448 9722 27476 10066
rect 27540 9926 27568 10542
rect 27620 10532 27672 10538
rect 27620 10474 27672 10480
rect 27632 10266 27660 10474
rect 27620 10260 27672 10266
rect 27620 10202 27672 10208
rect 27712 10260 27764 10266
rect 27712 10202 27764 10208
rect 27724 10169 27752 10202
rect 27908 10198 27936 14826
rect 27988 14408 28040 14414
rect 27988 14350 28040 14356
rect 28000 14074 28028 14350
rect 28092 14074 28120 15506
rect 28184 15026 28212 15574
rect 28276 15162 28304 15982
rect 28540 15904 28592 15910
rect 28540 15846 28592 15852
rect 28552 15638 28580 15846
rect 28540 15632 28592 15638
rect 28540 15574 28592 15580
rect 28920 15570 28948 17274
rect 29368 16992 29420 16998
rect 29368 16934 29420 16940
rect 29276 16176 29328 16182
rect 29276 16118 29328 16124
rect 28908 15564 28960 15570
rect 29184 15564 29236 15570
rect 28960 15524 29040 15552
rect 28908 15506 28960 15512
rect 29012 15162 29040 15524
rect 29184 15506 29236 15512
rect 28264 15156 28316 15162
rect 28264 15098 28316 15104
rect 29000 15156 29052 15162
rect 29000 15098 29052 15104
rect 29196 15026 29224 15506
rect 29288 15502 29316 16118
rect 29380 16046 29408 16934
rect 30300 16658 30328 19162
rect 32232 17626 32260 19162
rect 32232 17598 32536 17626
rect 32144 17436 32440 17456
rect 32200 17434 32224 17436
rect 32280 17434 32304 17436
rect 32360 17434 32384 17436
rect 32222 17382 32224 17434
rect 32286 17382 32298 17434
rect 32360 17382 32362 17434
rect 32200 17380 32224 17382
rect 32280 17380 32304 17382
rect 32360 17380 32384 17382
rect 32144 17360 32440 17380
rect 30564 17128 30616 17134
rect 30748 17128 30800 17134
rect 30616 17088 30696 17116
rect 30564 17070 30616 17076
rect 30668 16658 30696 17088
rect 30748 17070 30800 17076
rect 30288 16652 30340 16658
rect 30288 16594 30340 16600
rect 30656 16652 30708 16658
rect 30656 16594 30708 16600
rect 30104 16516 30156 16522
rect 30104 16458 30156 16464
rect 29552 16448 29604 16454
rect 29552 16390 29604 16396
rect 29564 16046 29592 16390
rect 29368 16040 29420 16046
rect 29552 16040 29604 16046
rect 29420 15988 29500 15994
rect 29368 15982 29500 15988
rect 29552 15982 29604 15988
rect 29380 15966 29500 15982
rect 29368 15904 29420 15910
rect 29368 15846 29420 15852
rect 29380 15570 29408 15846
rect 29368 15564 29420 15570
rect 29368 15506 29420 15512
rect 29276 15496 29328 15502
rect 29276 15438 29328 15444
rect 29288 15162 29316 15438
rect 29276 15156 29328 15162
rect 29276 15098 29328 15104
rect 28172 15020 28224 15026
rect 28172 14962 28224 14968
rect 29184 15020 29236 15026
rect 29184 14962 29236 14968
rect 28184 14414 28212 14962
rect 29380 14550 29408 15506
rect 28264 14544 28316 14550
rect 29368 14544 29420 14550
rect 28264 14486 28316 14492
rect 28354 14512 28410 14521
rect 28172 14408 28224 14414
rect 28172 14350 28224 14356
rect 27988 14068 28040 14074
rect 27988 14010 28040 14016
rect 28080 14068 28132 14074
rect 28080 14010 28132 14016
rect 27896 10192 27948 10198
rect 27710 10160 27766 10169
rect 27896 10134 27948 10140
rect 27710 10095 27766 10104
rect 27528 9920 27580 9926
rect 27528 9862 27580 9868
rect 27436 9716 27488 9722
rect 27436 9658 27488 9664
rect 27436 9376 27488 9382
rect 27436 9318 27488 9324
rect 27264 9166 27384 9194
rect 27160 8968 27212 8974
rect 27160 8910 27212 8916
rect 27172 8430 27200 8910
rect 27160 8424 27212 8430
rect 27160 8366 27212 8372
rect 26988 7364 27108 7392
rect 26884 7336 26936 7342
rect 26884 7278 26936 7284
rect 26896 7177 26924 7278
rect 26882 7168 26938 7177
rect 26882 7103 26938 7112
rect 26752 6820 26832 6848
rect 26700 6802 26752 6808
rect 26804 6118 26832 6820
rect 26896 6730 26924 7103
rect 26884 6724 26936 6730
rect 26884 6666 26936 6672
rect 26792 6112 26844 6118
rect 26792 6054 26844 6060
rect 26700 5704 26752 5710
rect 26698 5672 26700 5681
rect 26752 5672 26754 5681
rect 26698 5607 26754 5616
rect 26608 5568 26660 5574
rect 26608 5510 26660 5516
rect 26712 5166 26740 5607
rect 26804 5574 26832 6054
rect 26988 5710 27016 7364
rect 27160 7336 27212 7342
rect 27160 7278 27212 7284
rect 27068 7268 27120 7274
rect 27068 7210 27120 7216
rect 27080 6866 27108 7210
rect 27172 6866 27200 7278
rect 27068 6860 27120 6866
rect 27068 6802 27120 6808
rect 27160 6860 27212 6866
rect 27160 6802 27212 6808
rect 27080 6254 27108 6802
rect 27172 6361 27200 6802
rect 27264 6497 27292 9166
rect 27448 9092 27476 9318
rect 27356 9064 27476 9092
rect 27356 8566 27384 9064
rect 27436 8900 27488 8906
rect 27436 8842 27488 8848
rect 27344 8560 27396 8566
rect 27344 8502 27396 8508
rect 27344 8424 27396 8430
rect 27344 8366 27396 8372
rect 27356 7834 27384 8366
rect 27448 7954 27476 8842
rect 27540 8294 27568 9862
rect 27620 9716 27672 9722
rect 27620 9658 27672 9664
rect 27632 9518 27660 9658
rect 28000 9586 28028 14010
rect 28184 13938 28212 14350
rect 28276 14074 28304 14486
rect 29368 14486 29420 14492
rect 28354 14447 28410 14456
rect 28368 14414 28396 14447
rect 28356 14408 28408 14414
rect 28356 14350 28408 14356
rect 29276 14340 29328 14346
rect 29276 14282 29328 14288
rect 28816 14272 28868 14278
rect 28816 14214 28868 14220
rect 28908 14272 28960 14278
rect 28908 14214 28960 14220
rect 28264 14068 28316 14074
rect 28264 14010 28316 14016
rect 28828 14006 28856 14214
rect 28816 14000 28868 14006
rect 28816 13942 28868 13948
rect 28172 13932 28224 13938
rect 28172 13874 28224 13880
rect 28184 13530 28212 13874
rect 28540 13864 28592 13870
rect 28540 13806 28592 13812
rect 28552 13530 28580 13806
rect 28828 13530 28856 13942
rect 28920 13938 28948 14214
rect 28908 13932 28960 13938
rect 28908 13874 28960 13880
rect 29090 13832 29146 13841
rect 29090 13767 29146 13776
rect 28172 13524 28224 13530
rect 28172 13466 28224 13472
rect 28540 13524 28592 13530
rect 28540 13466 28592 13472
rect 28816 13524 28868 13530
rect 28816 13466 28868 13472
rect 28184 13326 28212 13466
rect 28172 13320 28224 13326
rect 28172 13262 28224 13268
rect 28184 12986 28212 13262
rect 28264 13184 28316 13190
rect 28552 13172 28580 13466
rect 28724 13388 28776 13394
rect 28724 13330 28776 13336
rect 28552 13144 28672 13172
rect 28264 13126 28316 13132
rect 28172 12980 28224 12986
rect 28172 12922 28224 12928
rect 28276 11665 28304 13126
rect 28354 13016 28410 13025
rect 28354 12951 28410 12960
rect 28368 12918 28396 12951
rect 28356 12912 28408 12918
rect 28356 12854 28408 12860
rect 28540 12776 28592 12782
rect 28540 12718 28592 12724
rect 28552 12306 28580 12718
rect 28540 12300 28592 12306
rect 28540 12242 28592 12248
rect 28262 11656 28318 11665
rect 28262 11591 28318 11600
rect 28264 11552 28316 11558
rect 28264 11494 28316 11500
rect 28276 10538 28304 11494
rect 28264 10532 28316 10538
rect 28264 10474 28316 10480
rect 28356 9920 28408 9926
rect 28356 9862 28408 9868
rect 27988 9580 28040 9586
rect 27988 9522 28040 9528
rect 27620 9512 27672 9518
rect 27620 9454 27672 9460
rect 28368 8974 28396 9862
rect 28448 9512 28500 9518
rect 28448 9454 28500 9460
rect 28460 9042 28488 9454
rect 28448 9036 28500 9042
rect 28448 8978 28500 8984
rect 28356 8968 28408 8974
rect 28356 8910 28408 8916
rect 27620 8900 27672 8906
rect 27620 8842 27672 8848
rect 27632 8430 27660 8842
rect 27712 8832 27764 8838
rect 27712 8774 27764 8780
rect 27620 8424 27672 8430
rect 27620 8366 27672 8372
rect 27528 8288 27580 8294
rect 27528 8230 27580 8236
rect 27436 7948 27488 7954
rect 27436 7890 27488 7896
rect 27356 7806 27476 7834
rect 27448 6866 27476 7806
rect 27632 7154 27660 8366
rect 27724 8294 27752 8774
rect 28460 8634 28488 8978
rect 28538 8936 28594 8945
rect 28538 8871 28594 8880
rect 28552 8634 28580 8871
rect 28644 8838 28672 13144
rect 28736 12646 28764 13330
rect 28828 12986 28856 13466
rect 29104 13326 29132 13767
rect 29288 13530 29316 14282
rect 29276 13524 29328 13530
rect 29276 13466 29328 13472
rect 29092 13320 29144 13326
rect 29092 13262 29144 13268
rect 29184 13252 29236 13258
rect 29184 13194 29236 13200
rect 28816 12980 28868 12986
rect 28816 12922 28868 12928
rect 28724 12640 28776 12646
rect 28724 12582 28776 12588
rect 28736 12481 28764 12582
rect 28722 12472 28778 12481
rect 28722 12407 28778 12416
rect 28908 12232 28960 12238
rect 28908 12174 28960 12180
rect 28920 11694 28948 12174
rect 29196 12170 29224 13194
rect 29472 12170 29500 15966
rect 29564 15162 29592 15982
rect 30116 15162 30144 16458
rect 30300 16182 30328 16594
rect 30288 16176 30340 16182
rect 30288 16118 30340 16124
rect 30300 15706 30328 16118
rect 30668 15910 30696 16594
rect 30760 16590 30788 17070
rect 30748 16584 30800 16590
rect 30748 16526 30800 16532
rect 31944 16584 31996 16590
rect 31944 16526 31996 16532
rect 31116 16448 31168 16454
rect 31116 16390 31168 16396
rect 30748 16176 30800 16182
rect 30748 16118 30800 16124
rect 30656 15904 30708 15910
rect 30656 15846 30708 15852
rect 30288 15700 30340 15706
rect 30288 15642 30340 15648
rect 30760 15434 30788 16118
rect 31128 15706 31156 16390
rect 31956 15910 31984 16526
rect 32508 16454 32536 17598
rect 33784 17264 33836 17270
rect 33784 17206 33836 17212
rect 33324 16652 33376 16658
rect 33324 16594 33376 16600
rect 32588 16584 32640 16590
rect 32588 16526 32640 16532
rect 32496 16448 32548 16454
rect 32496 16390 32548 16396
rect 32144 16348 32440 16368
rect 32200 16346 32224 16348
rect 32280 16346 32304 16348
rect 32360 16346 32384 16348
rect 32222 16294 32224 16346
rect 32286 16294 32298 16346
rect 32360 16294 32362 16346
rect 32200 16292 32224 16294
rect 32280 16292 32304 16294
rect 32360 16292 32384 16294
rect 32144 16272 32440 16292
rect 32312 15972 32364 15978
rect 32312 15914 32364 15920
rect 31944 15904 31996 15910
rect 31944 15846 31996 15852
rect 31956 15706 31984 15846
rect 31116 15700 31168 15706
rect 31116 15642 31168 15648
rect 31944 15700 31996 15706
rect 31944 15642 31996 15648
rect 32324 15638 32352 15914
rect 32600 15910 32628 16526
rect 32864 16448 32916 16454
rect 32864 16390 32916 16396
rect 32680 16176 32732 16182
rect 32680 16118 32732 16124
rect 32588 15904 32640 15910
rect 32588 15846 32640 15852
rect 32312 15632 32364 15638
rect 32312 15574 32364 15580
rect 31300 15564 31352 15570
rect 31300 15506 31352 15512
rect 31760 15564 31812 15570
rect 31760 15506 31812 15512
rect 30748 15428 30800 15434
rect 30748 15370 30800 15376
rect 31312 15162 31340 15506
rect 31772 15162 31800 15506
rect 32036 15496 32088 15502
rect 32036 15438 32088 15444
rect 32048 15162 32076 15438
rect 32324 15348 32352 15574
rect 32600 15366 32628 15846
rect 32588 15360 32640 15366
rect 32324 15320 32536 15348
rect 32144 15260 32440 15280
rect 32200 15258 32224 15260
rect 32280 15258 32304 15260
rect 32360 15258 32384 15260
rect 32222 15206 32224 15258
rect 32286 15206 32298 15258
rect 32360 15206 32362 15258
rect 32200 15204 32224 15206
rect 32280 15204 32304 15206
rect 32360 15204 32384 15206
rect 32144 15184 32440 15204
rect 29552 15156 29604 15162
rect 29552 15098 29604 15104
rect 30104 15156 30156 15162
rect 30104 15098 30156 15104
rect 31300 15156 31352 15162
rect 31300 15098 31352 15104
rect 31760 15156 31812 15162
rect 31760 15098 31812 15104
rect 32036 15156 32088 15162
rect 32036 15098 32088 15104
rect 29552 14952 29604 14958
rect 29552 14894 29604 14900
rect 29828 14952 29880 14958
rect 29828 14894 29880 14900
rect 29564 14482 29592 14894
rect 29552 14476 29604 14482
rect 29552 14418 29604 14424
rect 29840 13938 29868 14894
rect 30116 14890 30144 15098
rect 30380 15020 30432 15026
rect 30380 14962 30432 14968
rect 30104 14884 30156 14890
rect 30104 14826 30156 14832
rect 30288 14816 30340 14822
rect 30288 14758 30340 14764
rect 30196 14476 30248 14482
rect 30196 14418 30248 14424
rect 30104 14408 30156 14414
rect 30104 14350 30156 14356
rect 29828 13932 29880 13938
rect 29828 13874 29880 13880
rect 30116 13870 30144 14350
rect 30208 13938 30236 14418
rect 30196 13932 30248 13938
rect 30196 13874 30248 13880
rect 29736 13864 29788 13870
rect 29736 13806 29788 13812
rect 30104 13864 30156 13870
rect 30104 13806 30156 13812
rect 29748 13530 29776 13806
rect 29828 13728 29880 13734
rect 29828 13670 29880 13676
rect 30012 13728 30064 13734
rect 30012 13670 30064 13676
rect 29736 13524 29788 13530
rect 29736 13466 29788 13472
rect 29748 13190 29776 13466
rect 29840 13394 29868 13670
rect 29828 13388 29880 13394
rect 29828 13330 29880 13336
rect 29736 13184 29788 13190
rect 29736 13126 29788 13132
rect 29840 12918 29868 13330
rect 30024 13190 30052 13670
rect 30012 13184 30064 13190
rect 30012 13126 30064 13132
rect 29828 12912 29880 12918
rect 29828 12854 29880 12860
rect 30024 12714 30052 13126
rect 30196 12776 30248 12782
rect 30196 12718 30248 12724
rect 30012 12708 30064 12714
rect 30012 12650 30064 12656
rect 30104 12300 30156 12306
rect 30104 12242 30156 12248
rect 29184 12164 29236 12170
rect 29184 12106 29236 12112
rect 29460 12164 29512 12170
rect 29460 12106 29512 12112
rect 29000 12096 29052 12102
rect 29000 12038 29052 12044
rect 29012 11898 29040 12038
rect 29000 11892 29052 11898
rect 29000 11834 29052 11840
rect 29012 11694 29040 11834
rect 28908 11688 28960 11694
rect 28908 11630 28960 11636
rect 29000 11688 29052 11694
rect 29000 11630 29052 11636
rect 29012 11354 29040 11630
rect 29092 11620 29144 11626
rect 29092 11562 29144 11568
rect 29000 11348 29052 11354
rect 29000 11290 29052 11296
rect 29104 10674 29132 11562
rect 29092 10668 29144 10674
rect 29092 10610 29144 10616
rect 28908 10464 28960 10470
rect 28908 10406 28960 10412
rect 28724 9988 28776 9994
rect 28724 9930 28776 9936
rect 28736 9518 28764 9930
rect 28920 9874 28948 10406
rect 29196 10198 29224 12106
rect 29368 11348 29420 11354
rect 29368 11290 29420 11296
rect 29380 10606 29408 11290
rect 29472 11218 29500 12106
rect 29460 11212 29512 11218
rect 29460 11154 29512 11160
rect 30116 11082 30144 12242
rect 30208 11898 30236 12718
rect 30300 12306 30328 14758
rect 30392 14618 30420 14962
rect 30380 14612 30432 14618
rect 30380 14554 30432 14560
rect 31772 14550 31800 15098
rect 32404 15088 32456 15094
rect 32402 15056 32404 15065
rect 32456 15056 32458 15065
rect 32402 14991 32458 15000
rect 32508 14618 32536 15320
rect 32588 15302 32640 15308
rect 32692 15094 32720 16118
rect 32876 16046 32904 16390
rect 33336 16114 33364 16594
rect 33692 16448 33744 16454
rect 33692 16390 33744 16396
rect 33704 16182 33732 16390
rect 33692 16176 33744 16182
rect 33692 16118 33744 16124
rect 33324 16108 33376 16114
rect 33324 16050 33376 16056
rect 32864 16040 32916 16046
rect 32864 15982 32916 15988
rect 33692 15972 33744 15978
rect 33692 15914 33744 15920
rect 32772 15904 32824 15910
rect 32772 15846 32824 15852
rect 32784 15706 32812 15846
rect 33704 15706 33732 15914
rect 32772 15700 32824 15706
rect 32772 15642 32824 15648
rect 33692 15700 33744 15706
rect 33692 15642 33744 15648
rect 32680 15088 32732 15094
rect 32680 15030 32732 15036
rect 32692 14958 32720 15030
rect 32680 14952 32732 14958
rect 32680 14894 32732 14900
rect 32312 14612 32364 14618
rect 32312 14554 32364 14560
rect 32496 14612 32548 14618
rect 32496 14554 32548 14560
rect 31760 14544 31812 14550
rect 31760 14486 31812 14492
rect 32324 14498 32352 14554
rect 32324 14482 32536 14498
rect 32324 14476 32548 14482
rect 32324 14470 32496 14476
rect 32496 14418 32548 14424
rect 32784 14414 32812 15642
rect 32864 15360 32916 15366
rect 32864 15302 32916 15308
rect 32876 15162 32904 15302
rect 32864 15156 32916 15162
rect 32864 15098 32916 15104
rect 33704 15026 33732 15642
rect 33796 15638 33824 17206
rect 34256 17202 34284 19162
rect 34244 17196 34296 17202
rect 34244 17138 34296 17144
rect 34152 17128 34204 17134
rect 34152 17070 34204 17076
rect 34164 16658 34192 17070
rect 34256 16794 34284 17138
rect 34336 17128 34388 17134
rect 34336 17070 34388 17076
rect 34244 16788 34296 16794
rect 34244 16730 34296 16736
rect 34152 16652 34204 16658
rect 34152 16594 34204 16600
rect 34348 16046 34376 17070
rect 34612 16584 34664 16590
rect 34612 16526 34664 16532
rect 35072 16584 35124 16590
rect 35072 16526 35124 16532
rect 34336 16040 34388 16046
rect 34336 15982 34388 15988
rect 33784 15632 33836 15638
rect 33784 15574 33836 15580
rect 34348 15366 34376 15982
rect 34624 15910 34652 16526
rect 35084 15910 35112 16526
rect 35716 16176 35768 16182
rect 35716 16118 35768 16124
rect 34612 15904 34664 15910
rect 34612 15846 34664 15852
rect 35072 15904 35124 15910
rect 35072 15846 35124 15852
rect 35624 15904 35676 15910
rect 35624 15846 35676 15852
rect 35084 15638 35112 15846
rect 35072 15632 35124 15638
rect 35072 15574 35124 15580
rect 34796 15564 34848 15570
rect 34796 15506 34848 15512
rect 34336 15360 34388 15366
rect 34336 15302 34388 15308
rect 34244 15156 34296 15162
rect 34244 15098 34296 15104
rect 33692 15020 33744 15026
rect 33692 14962 33744 14968
rect 33324 14476 33376 14482
rect 33324 14418 33376 14424
rect 31208 14408 31260 14414
rect 31208 14350 31260 14356
rect 32772 14408 32824 14414
rect 32772 14350 32824 14356
rect 33048 14408 33100 14414
rect 33048 14350 33100 14356
rect 30380 14272 30432 14278
rect 30380 14214 30432 14220
rect 30472 14272 30524 14278
rect 30472 14214 30524 14220
rect 30392 14074 30420 14214
rect 30380 14068 30432 14074
rect 30380 14010 30432 14016
rect 30288 12300 30340 12306
rect 30288 12242 30340 12248
rect 30196 11892 30248 11898
rect 30196 11834 30248 11840
rect 30196 11552 30248 11558
rect 30196 11494 30248 11500
rect 30104 11076 30156 11082
rect 30104 11018 30156 11024
rect 30208 10810 30236 11494
rect 30104 10804 30156 10810
rect 30104 10746 30156 10752
rect 30196 10804 30248 10810
rect 30196 10746 30248 10752
rect 30116 10713 30144 10746
rect 30102 10704 30158 10713
rect 30102 10639 30158 10648
rect 29368 10600 29420 10606
rect 29368 10542 29420 10548
rect 29184 10192 29236 10198
rect 29184 10134 29236 10140
rect 30288 10124 30340 10130
rect 30288 10066 30340 10072
rect 30300 9926 30328 10066
rect 29092 9920 29144 9926
rect 28920 9846 29040 9874
rect 29092 9862 29144 9868
rect 30104 9920 30156 9926
rect 30104 9862 30156 9868
rect 30288 9920 30340 9926
rect 30288 9862 30340 9868
rect 28920 9722 28948 9846
rect 28908 9716 28960 9722
rect 28908 9658 28960 9664
rect 28724 9512 28776 9518
rect 28724 9454 28776 9460
rect 28816 8968 28868 8974
rect 28868 8928 28948 8956
rect 28816 8910 28868 8916
rect 28632 8832 28684 8838
rect 28632 8774 28684 8780
rect 28448 8628 28500 8634
rect 28448 8570 28500 8576
rect 28540 8628 28592 8634
rect 28540 8570 28592 8576
rect 28920 8566 28948 8928
rect 28908 8560 28960 8566
rect 27894 8528 27950 8537
rect 28908 8502 28960 8508
rect 27894 8463 27950 8472
rect 28540 8492 28592 8498
rect 27908 8430 27936 8463
rect 28540 8434 28592 8440
rect 27896 8424 27948 8430
rect 27896 8366 27948 8372
rect 27712 8288 27764 8294
rect 27712 8230 27764 8236
rect 28172 8288 28224 8294
rect 28172 8230 28224 8236
rect 27896 8016 27948 8022
rect 27896 7958 27948 7964
rect 27908 7342 27936 7958
rect 27988 7744 28040 7750
rect 27988 7686 28040 7692
rect 27896 7336 27948 7342
rect 27896 7278 27948 7284
rect 27804 7268 27856 7274
rect 27804 7210 27856 7216
rect 27540 7126 27660 7154
rect 27436 6860 27488 6866
rect 27436 6802 27488 6808
rect 27250 6488 27306 6497
rect 27250 6423 27306 6432
rect 27158 6352 27214 6361
rect 27158 6287 27214 6296
rect 27068 6248 27120 6254
rect 27068 6190 27120 6196
rect 26976 5704 27028 5710
rect 26976 5646 27028 5652
rect 26792 5568 26844 5574
rect 26792 5510 26844 5516
rect 26804 5302 26832 5510
rect 26792 5296 26844 5302
rect 26792 5238 26844 5244
rect 26988 5234 27016 5646
rect 26976 5228 27028 5234
rect 26976 5170 27028 5176
rect 26700 5160 26752 5166
rect 26700 5102 26752 5108
rect 27172 5098 27200 6287
rect 27540 5545 27568 7126
rect 27816 7041 27844 7210
rect 27802 7032 27858 7041
rect 27802 6967 27858 6976
rect 27620 6316 27672 6322
rect 27620 6258 27672 6264
rect 27632 6100 27660 6258
rect 27804 6248 27856 6254
rect 27804 6190 27856 6196
rect 27712 6112 27764 6118
rect 27632 6072 27712 6100
rect 27712 6054 27764 6060
rect 27816 5953 27844 6190
rect 27802 5944 27858 5953
rect 27802 5879 27858 5888
rect 27804 5568 27856 5574
rect 27526 5536 27582 5545
rect 27804 5510 27856 5516
rect 27526 5471 27582 5480
rect 27252 5364 27304 5370
rect 27252 5306 27304 5312
rect 27264 5137 27292 5306
rect 27250 5128 27306 5137
rect 27160 5092 27212 5098
rect 27250 5063 27306 5072
rect 27160 5034 27212 5040
rect 27160 4684 27212 4690
rect 27160 4626 27212 4632
rect 26608 4548 26660 4554
rect 26660 4508 26832 4536
rect 26608 4490 26660 4496
rect 26332 4072 26384 4078
rect 26332 4014 26384 4020
rect 26344 3738 26372 4014
rect 26516 4004 26568 4010
rect 26516 3946 26568 3952
rect 26332 3732 26384 3738
rect 26332 3674 26384 3680
rect 26424 3732 26476 3738
rect 26424 3674 26476 3680
rect 26160 3454 26372 3482
rect 26344 3398 26372 3454
rect 26148 3392 26200 3398
rect 26146 3360 26148 3369
rect 26332 3392 26384 3398
rect 26200 3360 26202 3369
rect 26332 3334 26384 3340
rect 26146 3295 26202 3304
rect 26436 2904 26464 3674
rect 26528 3602 26556 3946
rect 26804 3602 26832 4508
rect 27172 3942 27200 4626
rect 27264 4078 27292 5063
rect 27436 4684 27488 4690
rect 27436 4626 27488 4632
rect 27448 4593 27476 4626
rect 27434 4584 27490 4593
rect 27434 4519 27490 4528
rect 27448 4282 27476 4519
rect 27436 4276 27488 4282
rect 27436 4218 27488 4224
rect 27252 4072 27304 4078
rect 27252 4014 27304 4020
rect 27620 4072 27672 4078
rect 27620 4014 27672 4020
rect 27160 3936 27212 3942
rect 27160 3878 27212 3884
rect 26882 3768 26938 3777
rect 26882 3703 26938 3712
rect 26516 3596 26568 3602
rect 26792 3596 26844 3602
rect 26568 3556 26740 3584
rect 26516 3538 26568 3544
rect 26516 3460 26568 3466
rect 26516 3402 26568 3408
rect 26068 2876 26464 2904
rect 25872 2372 25924 2378
rect 25872 2314 25924 2320
rect 26068 800 26096 2876
rect 26528 2854 26556 3402
rect 26608 2916 26660 2922
rect 26608 2858 26660 2864
rect 26516 2848 26568 2854
rect 26436 2808 26516 2836
rect 26436 2650 26464 2808
rect 26516 2790 26568 2796
rect 26620 2650 26648 2858
rect 26712 2650 26740 3556
rect 26792 3538 26844 3544
rect 26792 3460 26844 3466
rect 26792 3402 26844 3408
rect 26804 3369 26832 3402
rect 26790 3360 26846 3369
rect 26790 3295 26846 3304
rect 26424 2644 26476 2650
rect 26424 2586 26476 2592
rect 26608 2644 26660 2650
rect 26608 2586 26660 2592
rect 26700 2644 26752 2650
rect 26700 2586 26752 2592
rect 26896 800 26924 3703
rect 27264 3398 27292 4014
rect 27632 3534 27660 4014
rect 27816 4010 27844 5510
rect 27908 5166 27936 7278
rect 28000 7041 28028 7686
rect 28080 7336 28132 7342
rect 28080 7278 28132 7284
rect 27986 7032 28042 7041
rect 28092 7002 28120 7278
rect 27986 6967 28042 6976
rect 28080 6996 28132 7002
rect 28080 6938 28132 6944
rect 27988 5568 28040 5574
rect 27988 5510 28040 5516
rect 28000 5409 28028 5510
rect 27986 5400 28042 5409
rect 28184 5370 28212 8230
rect 28448 7744 28500 7750
rect 28448 7686 28500 7692
rect 28460 7410 28488 7686
rect 28448 7404 28500 7410
rect 28448 7346 28500 7352
rect 28264 7200 28316 7206
rect 28264 7142 28316 7148
rect 28276 6934 28304 7142
rect 28448 6996 28500 7002
rect 28448 6938 28500 6944
rect 28264 6928 28316 6934
rect 28264 6870 28316 6876
rect 28264 6792 28316 6798
rect 28264 6734 28316 6740
rect 28276 6186 28304 6734
rect 28356 6384 28408 6390
rect 28356 6326 28408 6332
rect 28264 6180 28316 6186
rect 28264 6122 28316 6128
rect 28264 5908 28316 5914
rect 28264 5850 28316 5856
rect 27986 5335 28042 5344
rect 28172 5364 28224 5370
rect 28172 5306 28224 5312
rect 27896 5160 27948 5166
rect 27896 5102 27948 5108
rect 28080 5160 28132 5166
rect 28184 5148 28212 5306
rect 28276 5166 28304 5850
rect 28368 5166 28396 6326
rect 28460 6322 28488 6938
rect 28552 6934 28580 8434
rect 28724 8424 28776 8430
rect 28724 8366 28776 8372
rect 28736 7546 28764 8366
rect 28920 8022 28948 8502
rect 28908 8016 28960 8022
rect 28908 7958 28960 7964
rect 28816 7948 28868 7954
rect 28816 7890 28868 7896
rect 28828 7546 28856 7890
rect 28724 7540 28776 7546
rect 28724 7482 28776 7488
rect 28816 7540 28868 7546
rect 28816 7482 28868 7488
rect 29012 7410 29040 9846
rect 29104 9450 29132 9862
rect 30116 9466 30144 9862
rect 30300 9654 30328 9862
rect 30288 9648 30340 9654
rect 30288 9590 30340 9596
rect 30300 9518 30328 9590
rect 29092 9444 29144 9450
rect 29092 9386 29144 9392
rect 29932 9438 30144 9466
rect 30288 9512 30340 9518
rect 30288 9454 30340 9460
rect 29104 7954 29132 9386
rect 29932 9382 29960 9438
rect 29920 9376 29972 9382
rect 29920 9318 29972 9324
rect 30012 9376 30064 9382
rect 30012 9318 30064 9324
rect 30024 9042 30052 9318
rect 30116 9042 30144 9438
rect 30392 9110 30420 14010
rect 30484 13530 30512 14214
rect 31220 13802 31248 14350
rect 31944 14272 31996 14278
rect 31944 14214 31996 14220
rect 31956 13938 31984 14214
rect 32144 14172 32440 14192
rect 32200 14170 32224 14172
rect 32280 14170 32304 14172
rect 32360 14170 32384 14172
rect 32222 14118 32224 14170
rect 32286 14118 32298 14170
rect 32360 14118 32362 14170
rect 32200 14116 32224 14118
rect 32280 14116 32304 14118
rect 32360 14116 32384 14118
rect 32144 14096 32440 14116
rect 31944 13932 31996 13938
rect 31944 13874 31996 13880
rect 31208 13796 31260 13802
rect 31208 13738 31260 13744
rect 32128 13796 32180 13802
rect 32128 13738 32180 13744
rect 30930 13560 30986 13569
rect 30472 13524 30524 13530
rect 31220 13530 31248 13738
rect 32140 13682 32168 13738
rect 32048 13654 32168 13682
rect 30930 13495 30986 13504
rect 31208 13524 31260 13530
rect 30472 13466 30524 13472
rect 30944 13394 30972 13495
rect 31208 13466 31260 13472
rect 30932 13388 30984 13394
rect 30932 13330 30984 13336
rect 30944 12986 30972 13330
rect 31668 13320 31720 13326
rect 31668 13262 31720 13268
rect 30932 12980 30984 12986
rect 30932 12922 30984 12928
rect 31680 12850 31708 13262
rect 32048 13190 32076 13654
rect 32496 13388 32548 13394
rect 32496 13330 32548 13336
rect 32036 13184 32088 13190
rect 32036 13126 32088 13132
rect 31668 12844 31720 12850
rect 31668 12786 31720 12792
rect 31392 12776 31444 12782
rect 31390 12744 31392 12753
rect 31576 12776 31628 12782
rect 31444 12744 31446 12753
rect 31208 12708 31260 12714
rect 31446 12702 31524 12730
rect 31576 12718 31628 12724
rect 31390 12679 31446 12688
rect 31208 12650 31260 12656
rect 30748 11824 30800 11830
rect 30748 11766 30800 11772
rect 30760 11354 30788 11766
rect 30748 11348 30800 11354
rect 30748 11290 30800 11296
rect 30472 11008 30524 11014
rect 30472 10950 30524 10956
rect 30932 11008 30984 11014
rect 30932 10950 30984 10956
rect 30484 10810 30512 10950
rect 30472 10804 30524 10810
rect 30472 10746 30524 10752
rect 30484 10577 30512 10746
rect 30944 10606 30972 10950
rect 31220 10810 31248 12650
rect 31392 12640 31444 12646
rect 31392 12582 31444 12588
rect 31404 12481 31432 12582
rect 31390 12472 31446 12481
rect 31390 12407 31446 12416
rect 31496 11558 31524 12702
rect 31588 12170 31616 12718
rect 32048 12646 32076 13126
rect 32144 13084 32440 13104
rect 32200 13082 32224 13084
rect 32280 13082 32304 13084
rect 32360 13082 32384 13084
rect 32222 13030 32224 13082
rect 32286 13030 32298 13082
rect 32360 13030 32362 13082
rect 32200 13028 32224 13030
rect 32280 13028 32304 13030
rect 32360 13028 32384 13030
rect 32144 13008 32440 13028
rect 32126 12744 32182 12753
rect 32126 12679 32128 12688
rect 32180 12679 32182 12688
rect 32128 12650 32180 12656
rect 32036 12640 32088 12646
rect 32036 12582 32088 12588
rect 31576 12164 31628 12170
rect 31576 12106 31628 12112
rect 31668 11756 31720 11762
rect 31760 11756 31812 11762
rect 31720 11716 31760 11744
rect 31668 11698 31720 11704
rect 31760 11698 31812 11704
rect 31760 11620 31812 11626
rect 31760 11562 31812 11568
rect 31484 11552 31536 11558
rect 31484 11494 31536 11500
rect 31576 11212 31628 11218
rect 31576 11154 31628 11160
rect 31208 10804 31260 10810
rect 31208 10746 31260 10752
rect 30932 10600 30984 10606
rect 30470 10568 30526 10577
rect 30932 10542 30984 10548
rect 30470 10503 30526 10512
rect 30840 10464 30892 10470
rect 30840 10406 30892 10412
rect 30852 10266 30880 10406
rect 30840 10260 30892 10266
rect 30840 10202 30892 10208
rect 30656 9444 30708 9450
rect 30656 9386 30708 9392
rect 30840 9444 30892 9450
rect 30840 9386 30892 9392
rect 30288 9104 30340 9110
rect 30286 9072 30288 9081
rect 30380 9104 30432 9110
rect 30340 9072 30342 9081
rect 30012 9036 30064 9042
rect 30012 8978 30064 8984
rect 30104 9036 30156 9042
rect 30380 9046 30432 9052
rect 30286 9007 30342 9016
rect 30104 8978 30156 8984
rect 29460 8968 29512 8974
rect 29460 8910 29512 8916
rect 29276 8832 29328 8838
rect 29276 8774 29328 8780
rect 29368 8832 29420 8838
rect 29368 8774 29420 8780
rect 29288 8498 29316 8774
rect 29276 8492 29328 8498
rect 29276 8434 29328 8440
rect 29380 8430 29408 8774
rect 29368 8424 29420 8430
rect 29368 8366 29420 8372
rect 29472 8276 29500 8910
rect 30024 8566 30052 8978
rect 30012 8560 30064 8566
rect 30012 8502 30064 8508
rect 29288 8248 29500 8276
rect 29550 8256 29606 8265
rect 29092 7948 29144 7954
rect 29092 7890 29144 7896
rect 29090 7848 29146 7857
rect 29090 7783 29092 7792
rect 29144 7783 29146 7792
rect 29092 7754 29144 7760
rect 29000 7404 29052 7410
rect 29000 7346 29052 7352
rect 29288 7274 29316 8248
rect 29550 8191 29606 8200
rect 29368 8016 29420 8022
rect 29368 7958 29420 7964
rect 29380 7750 29408 7958
rect 29460 7880 29512 7886
rect 29460 7822 29512 7828
rect 29368 7744 29420 7750
rect 29368 7686 29420 7692
rect 29276 7268 29328 7274
rect 29328 7228 29408 7256
rect 29276 7210 29328 7216
rect 28998 7168 29054 7177
rect 28998 7103 29054 7112
rect 29012 6934 29040 7103
rect 29090 7032 29146 7041
rect 29090 6967 29146 6976
rect 29104 6934 29132 6967
rect 28540 6928 28592 6934
rect 29000 6928 29052 6934
rect 28540 6870 28592 6876
rect 28736 6866 28948 6882
rect 29000 6870 29052 6876
rect 29092 6928 29144 6934
rect 29092 6870 29144 6876
rect 28724 6860 28948 6866
rect 28776 6854 28948 6860
rect 28724 6802 28776 6808
rect 28920 6780 28948 6854
rect 29092 6792 29144 6798
rect 28920 6752 29092 6780
rect 29092 6734 29144 6740
rect 28816 6724 28868 6730
rect 29380 6712 29408 7228
rect 29472 6866 29500 7822
rect 29564 7721 29592 8191
rect 29644 8084 29696 8090
rect 29644 8026 29696 8032
rect 29550 7712 29606 7721
rect 29550 7647 29606 7656
rect 29656 7290 29684 8026
rect 29920 7948 29972 7954
rect 29920 7890 29972 7896
rect 29828 7880 29880 7886
rect 29932 7857 29960 7890
rect 29828 7822 29880 7828
rect 29918 7848 29974 7857
rect 29840 7478 29868 7822
rect 29918 7783 29974 7792
rect 29920 7744 29972 7750
rect 29920 7686 29972 7692
rect 29828 7472 29880 7478
rect 29828 7414 29880 7420
rect 29564 7274 29684 7290
rect 29552 7268 29684 7274
rect 29604 7262 29684 7268
rect 29552 7210 29604 7216
rect 29932 7002 29960 7686
rect 30012 7268 30064 7274
rect 30012 7210 30064 7216
rect 29920 6996 29972 7002
rect 29920 6938 29972 6944
rect 30024 6866 30052 7210
rect 29460 6860 29512 6866
rect 29460 6802 29512 6808
rect 30012 6860 30064 6866
rect 30012 6802 30064 6808
rect 28816 6666 28868 6672
rect 29288 6684 29408 6712
rect 29552 6724 29604 6730
rect 28632 6656 28684 6662
rect 28632 6598 28684 6604
rect 28448 6316 28500 6322
rect 28448 6258 28500 6264
rect 28644 5710 28672 6598
rect 28722 6352 28778 6361
rect 28722 6287 28724 6296
rect 28776 6287 28778 6296
rect 28828 6304 28856 6666
rect 28828 6276 28948 6304
rect 28724 6258 28776 6264
rect 28816 6180 28868 6186
rect 28920 6168 28948 6276
rect 29092 6180 29144 6186
rect 28920 6140 29092 6168
rect 28816 6122 28868 6128
rect 29092 6122 29144 6128
rect 28632 5704 28684 5710
rect 28632 5646 28684 5652
rect 28132 5120 28212 5148
rect 28264 5160 28316 5166
rect 28080 5102 28132 5108
rect 28264 5102 28316 5108
rect 28356 5160 28408 5166
rect 28356 5102 28408 5108
rect 28632 4684 28684 4690
rect 28632 4626 28684 4632
rect 27896 4480 27948 4486
rect 27896 4422 27948 4428
rect 27908 4078 27936 4422
rect 27896 4072 27948 4078
rect 27896 4014 27948 4020
rect 28172 4072 28224 4078
rect 28172 4014 28224 4020
rect 27804 4004 27856 4010
rect 27804 3946 27856 3952
rect 27620 3528 27672 3534
rect 27620 3470 27672 3476
rect 26976 3392 27028 3398
rect 26976 3334 27028 3340
rect 27252 3392 27304 3398
rect 27252 3334 27304 3340
rect 27436 3392 27488 3398
rect 27436 3334 27488 3340
rect 26988 2990 27016 3334
rect 27448 3194 27476 3334
rect 27436 3188 27488 3194
rect 27488 3148 27752 3176
rect 27436 3130 27488 3136
rect 27724 2990 27752 3148
rect 27816 3126 27844 3946
rect 27908 3466 27936 4014
rect 28080 3596 28132 3602
rect 28080 3538 28132 3544
rect 27986 3496 28042 3505
rect 27896 3460 27948 3466
rect 27986 3431 28042 3440
rect 27896 3402 27948 3408
rect 27804 3120 27856 3126
rect 27804 3062 27856 3068
rect 26976 2984 27028 2990
rect 26976 2926 27028 2932
rect 27712 2984 27764 2990
rect 27712 2926 27764 2932
rect 28000 1816 28028 3431
rect 28092 2582 28120 3538
rect 28184 3194 28212 4014
rect 28356 4004 28408 4010
rect 28356 3946 28408 3952
rect 28264 3596 28316 3602
rect 28264 3538 28316 3544
rect 28276 3194 28304 3538
rect 28172 3188 28224 3194
rect 28172 3130 28224 3136
rect 28264 3188 28316 3194
rect 28264 3130 28316 3136
rect 28368 3058 28396 3946
rect 28644 3942 28672 4626
rect 28632 3936 28684 3942
rect 28446 3904 28502 3913
rect 28632 3878 28684 3884
rect 28446 3839 28502 3848
rect 28460 3058 28488 3839
rect 28828 3233 28856 6122
rect 29104 5953 29132 6122
rect 29090 5944 29146 5953
rect 29090 5879 29146 5888
rect 29092 5772 29144 5778
rect 29092 5714 29144 5720
rect 28998 5400 29054 5409
rect 28998 5335 29054 5344
rect 29012 5098 29040 5335
rect 29104 5302 29132 5714
rect 29288 5574 29316 6684
rect 29552 6666 29604 6672
rect 29564 6322 29592 6666
rect 29552 6316 29604 6322
rect 29552 6258 29604 6264
rect 30012 6248 30064 6254
rect 30116 6236 30144 8978
rect 30564 8492 30616 8498
rect 30564 8434 30616 8440
rect 30196 8016 30248 8022
rect 30196 7958 30248 7964
rect 30208 7546 30236 7958
rect 30196 7540 30248 7546
rect 30196 7482 30248 7488
rect 30576 6866 30604 8434
rect 30668 8430 30696 9386
rect 30748 8968 30800 8974
rect 30748 8910 30800 8916
rect 30656 8424 30708 8430
rect 30656 8366 30708 8372
rect 30656 8288 30708 8294
rect 30656 8230 30708 8236
rect 30668 7206 30696 8230
rect 30760 8090 30788 8910
rect 30748 8084 30800 8090
rect 30748 8026 30800 8032
rect 30748 7336 30800 7342
rect 30748 7278 30800 7284
rect 30656 7200 30708 7206
rect 30656 7142 30708 7148
rect 30564 6860 30616 6866
rect 30564 6802 30616 6808
rect 30380 6656 30432 6662
rect 30380 6598 30432 6604
rect 30064 6208 30144 6236
rect 30012 6190 30064 6196
rect 29460 5772 29512 5778
rect 29460 5714 29512 5720
rect 29552 5772 29604 5778
rect 29552 5714 29604 5720
rect 30012 5772 30064 5778
rect 30012 5714 30064 5720
rect 29472 5642 29500 5714
rect 29368 5636 29420 5642
rect 29368 5578 29420 5584
rect 29460 5636 29512 5642
rect 29460 5578 29512 5584
rect 29276 5568 29328 5574
rect 29276 5510 29328 5516
rect 29092 5296 29144 5302
rect 29092 5238 29144 5244
rect 29000 5092 29052 5098
rect 29000 5034 29052 5040
rect 28906 4720 28962 4729
rect 28906 4655 28908 4664
rect 28960 4655 28962 4664
rect 29000 4684 29052 4690
rect 28908 4626 28960 4632
rect 29000 4626 29052 4632
rect 29012 3618 29040 4626
rect 29104 3670 29132 5238
rect 29380 4214 29408 5578
rect 29472 4690 29500 5578
rect 29564 5574 29592 5714
rect 29828 5704 29880 5710
rect 29828 5646 29880 5652
rect 29552 5568 29604 5574
rect 29552 5510 29604 5516
rect 29564 5409 29592 5510
rect 29550 5400 29606 5409
rect 29550 5335 29606 5344
rect 29840 5166 29868 5646
rect 29828 5160 29880 5166
rect 29828 5102 29880 5108
rect 29920 5160 29972 5166
rect 29920 5102 29972 5108
rect 29932 5030 29960 5102
rect 29736 5024 29788 5030
rect 29734 4992 29736 5001
rect 29920 5024 29972 5030
rect 29788 4992 29790 5001
rect 29734 4927 29790 4936
rect 29840 4972 29920 4978
rect 29840 4966 29972 4972
rect 29840 4950 29960 4966
rect 29840 4758 29868 4950
rect 29932 4901 29960 4950
rect 29828 4752 29880 4758
rect 29828 4694 29880 4700
rect 29460 4684 29512 4690
rect 30024 4672 30052 5714
rect 30104 5636 30156 5642
rect 30104 5578 30156 5584
rect 30116 5166 30144 5578
rect 30288 5568 30340 5574
rect 30288 5510 30340 5516
rect 30300 5166 30328 5510
rect 30392 5273 30420 6598
rect 30378 5264 30434 5273
rect 30378 5199 30434 5208
rect 30104 5160 30156 5166
rect 30104 5102 30156 5108
rect 30288 5160 30340 5166
rect 30288 5102 30340 5108
rect 30196 5092 30248 5098
rect 30196 5034 30248 5040
rect 29460 4626 29512 4632
rect 29932 4644 30052 4672
rect 29644 4480 29696 4486
rect 29644 4422 29696 4428
rect 29460 4276 29512 4282
rect 29460 4218 29512 4224
rect 29368 4208 29420 4214
rect 29368 4150 29420 4156
rect 28920 3602 29040 3618
rect 29092 3664 29144 3670
rect 29092 3606 29144 3612
rect 28908 3596 29040 3602
rect 28960 3590 29040 3596
rect 28908 3538 28960 3544
rect 28814 3224 28870 3233
rect 28724 3188 28776 3194
rect 28814 3159 28870 3168
rect 28724 3130 28776 3136
rect 28356 3052 28408 3058
rect 28356 2994 28408 3000
rect 28448 3052 28500 3058
rect 28448 2994 28500 3000
rect 28080 2576 28132 2582
rect 28080 2518 28132 2524
rect 27816 1788 28028 1816
rect 27816 800 27844 1788
rect 28736 800 28764 3130
rect 29012 2650 29040 3590
rect 29274 3360 29330 3369
rect 29274 3295 29330 3304
rect 29288 2990 29316 3295
rect 29472 2990 29500 4218
rect 29656 4146 29684 4422
rect 29644 4140 29696 4146
rect 29644 4082 29696 4088
rect 29932 3602 29960 4644
rect 30208 4622 30236 5034
rect 30654 4992 30710 5001
rect 30654 4927 30710 4936
rect 30668 4758 30696 4927
rect 30472 4752 30524 4758
rect 30472 4694 30524 4700
rect 30656 4752 30708 4758
rect 30656 4694 30708 4700
rect 30196 4616 30248 4622
rect 30010 4584 30066 4593
rect 30196 4558 30248 4564
rect 30010 4519 30066 4528
rect 30288 4548 30340 4554
rect 30024 4078 30052 4519
rect 30288 4490 30340 4496
rect 30300 4214 30328 4490
rect 30484 4486 30512 4694
rect 30472 4480 30524 4486
rect 30472 4422 30524 4428
rect 30288 4208 30340 4214
rect 30288 4150 30340 4156
rect 30012 4072 30064 4078
rect 30012 4014 30064 4020
rect 30196 4004 30248 4010
rect 30196 3946 30248 3952
rect 29920 3596 29972 3602
rect 29920 3538 29972 3544
rect 30208 3058 30236 3946
rect 30300 3602 30328 4150
rect 30484 4078 30512 4422
rect 30760 4078 30788 7278
rect 30472 4072 30524 4078
rect 30472 4014 30524 4020
rect 30748 4072 30800 4078
rect 30748 4014 30800 4020
rect 30484 3670 30512 4014
rect 30656 3936 30708 3942
rect 30656 3878 30708 3884
rect 30472 3664 30524 3670
rect 30472 3606 30524 3612
rect 30668 3602 30696 3878
rect 30852 3641 30880 9386
rect 30944 6662 30972 10542
rect 31588 10470 31616 11154
rect 31772 11082 31800 11562
rect 31760 11076 31812 11082
rect 31760 11018 31812 11024
rect 31944 11076 31996 11082
rect 31944 11018 31996 11024
rect 31576 10464 31628 10470
rect 31576 10406 31628 10412
rect 31588 10062 31616 10406
rect 31576 10056 31628 10062
rect 31576 9998 31628 10004
rect 31208 9920 31260 9926
rect 31208 9862 31260 9868
rect 31116 9376 31168 9382
rect 31116 9318 31168 9324
rect 31022 9072 31078 9081
rect 31022 9007 31078 9016
rect 31036 7546 31064 9007
rect 31024 7540 31076 7546
rect 31024 7482 31076 7488
rect 30932 6656 30984 6662
rect 30932 6598 30984 6604
rect 31128 6474 31156 9318
rect 31220 8838 31248 9862
rect 31208 8832 31260 8838
rect 31208 8774 31260 8780
rect 31300 8424 31352 8430
rect 31300 8366 31352 8372
rect 31312 8294 31340 8366
rect 31300 8288 31352 8294
rect 31300 8230 31352 8236
rect 31208 7948 31260 7954
rect 31208 7890 31260 7896
rect 31220 7750 31248 7890
rect 31208 7744 31260 7750
rect 31208 7686 31260 7692
rect 31220 7002 31248 7686
rect 31312 7342 31340 8230
rect 31484 7744 31536 7750
rect 31484 7686 31536 7692
rect 31496 7410 31524 7686
rect 31484 7404 31536 7410
rect 31484 7346 31536 7352
rect 31300 7336 31352 7342
rect 31300 7278 31352 7284
rect 31390 7032 31446 7041
rect 31208 6996 31260 7002
rect 31390 6967 31446 6976
rect 31208 6938 31260 6944
rect 31300 6860 31352 6866
rect 31300 6802 31352 6808
rect 30944 6446 31156 6474
rect 30838 3632 30894 3641
rect 30288 3596 30340 3602
rect 30288 3538 30340 3544
rect 30564 3596 30616 3602
rect 30564 3538 30616 3544
rect 30656 3596 30708 3602
rect 30838 3567 30894 3576
rect 30656 3538 30708 3544
rect 30196 3052 30248 3058
rect 30196 2994 30248 3000
rect 29276 2984 29328 2990
rect 29276 2926 29328 2932
rect 29460 2984 29512 2990
rect 29460 2926 29512 2932
rect 29472 2854 29500 2926
rect 30576 2922 30604 3538
rect 30748 3120 30800 3126
rect 30748 3062 30800 3068
rect 30564 2916 30616 2922
rect 30564 2858 30616 2864
rect 29460 2848 29512 2854
rect 29460 2790 29512 2796
rect 29550 2816 29606 2825
rect 29550 2751 29606 2760
rect 29000 2644 29052 2650
rect 29000 2586 29052 2592
rect 29564 800 29592 2751
rect 30760 2514 30788 3062
rect 30944 2961 30972 6446
rect 31312 6254 31340 6802
rect 31300 6248 31352 6254
rect 31300 6190 31352 6196
rect 31312 5778 31340 6190
rect 31404 6118 31432 6967
rect 31484 6384 31536 6390
rect 31482 6352 31484 6361
rect 31536 6352 31538 6361
rect 31482 6287 31538 6296
rect 31392 6112 31444 6118
rect 31484 6112 31536 6118
rect 31392 6054 31444 6060
rect 31482 6080 31484 6089
rect 31536 6080 31538 6089
rect 31482 6015 31538 6024
rect 31588 6066 31616 9998
rect 31760 9920 31812 9926
rect 31760 9862 31812 9868
rect 31772 9450 31800 9862
rect 31956 9654 31984 11018
rect 32048 10538 32076 12582
rect 32508 12374 32536 13330
rect 32680 13320 32732 13326
rect 32586 13288 32642 13297
rect 32680 13262 32732 13268
rect 32586 13223 32642 13232
rect 32600 13190 32628 13223
rect 32588 13184 32640 13190
rect 32588 13126 32640 13132
rect 32586 13016 32642 13025
rect 32692 12986 32720 13262
rect 32586 12951 32588 12960
rect 32640 12951 32642 12960
rect 32680 12980 32732 12986
rect 32588 12922 32640 12928
rect 32680 12922 32732 12928
rect 32496 12368 32548 12374
rect 32496 12310 32548 12316
rect 32588 12300 32640 12306
rect 32588 12242 32640 12248
rect 32144 11996 32440 12016
rect 32200 11994 32224 11996
rect 32280 11994 32304 11996
rect 32360 11994 32384 11996
rect 32222 11942 32224 11994
rect 32286 11942 32298 11994
rect 32360 11942 32362 11994
rect 32200 11940 32224 11942
rect 32280 11940 32304 11942
rect 32360 11940 32384 11942
rect 32144 11920 32440 11940
rect 32404 11756 32456 11762
rect 32404 11698 32456 11704
rect 32416 11286 32444 11698
rect 32600 11558 32628 12242
rect 32496 11552 32548 11558
rect 32496 11494 32548 11500
rect 32588 11552 32640 11558
rect 32588 11494 32640 11500
rect 32404 11280 32456 11286
rect 32404 11222 32456 11228
rect 32508 11082 32536 11494
rect 32588 11212 32640 11218
rect 32588 11154 32640 11160
rect 32496 11076 32548 11082
rect 32496 11018 32548 11024
rect 32144 10908 32440 10928
rect 32200 10906 32224 10908
rect 32280 10906 32304 10908
rect 32360 10906 32384 10908
rect 32222 10854 32224 10906
rect 32286 10854 32298 10906
rect 32360 10854 32362 10906
rect 32200 10852 32224 10854
rect 32280 10852 32304 10854
rect 32360 10852 32384 10854
rect 32144 10832 32440 10852
rect 32312 10600 32364 10606
rect 32310 10568 32312 10577
rect 32364 10568 32366 10577
rect 32036 10532 32088 10538
rect 32310 10503 32366 10512
rect 32036 10474 32088 10480
rect 32324 10062 32352 10503
rect 32600 10266 32628 11154
rect 32784 11150 32812 14350
rect 32956 14272 33008 14278
rect 32956 14214 33008 14220
rect 32968 13954 32996 14214
rect 33060 14074 33088 14350
rect 33048 14068 33100 14074
rect 33048 14010 33100 14016
rect 32968 13926 33088 13954
rect 33060 13870 33088 13926
rect 33048 13864 33100 13870
rect 33048 13806 33100 13812
rect 33140 13864 33192 13870
rect 33140 13806 33192 13812
rect 33060 13462 33088 13806
rect 33048 13456 33100 13462
rect 33048 13398 33100 13404
rect 33048 13252 33100 13258
rect 33048 13194 33100 13200
rect 33060 12782 33088 13194
rect 33152 12850 33180 13806
rect 33232 13320 33284 13326
rect 33232 13262 33284 13268
rect 33140 12844 33192 12850
rect 33140 12786 33192 12792
rect 33048 12776 33100 12782
rect 33048 12718 33100 12724
rect 33140 12436 33192 12442
rect 33140 12378 33192 12384
rect 32864 11688 32916 11694
rect 32864 11630 32916 11636
rect 32876 11218 32904 11630
rect 33152 11558 33180 12378
rect 33048 11552 33100 11558
rect 33046 11520 33048 11529
rect 33140 11552 33192 11558
rect 33100 11520 33102 11529
rect 33140 11494 33192 11500
rect 33046 11455 33102 11464
rect 33244 11354 33272 13262
rect 33336 12442 33364 14418
rect 33508 13728 33560 13734
rect 33704 13705 33732 14962
rect 33784 14952 33836 14958
rect 33784 14894 33836 14900
rect 33508 13670 33560 13676
rect 33690 13696 33746 13705
rect 33520 13394 33548 13670
rect 33690 13631 33746 13640
rect 33796 13433 33824 14894
rect 34152 14884 34204 14890
rect 34152 14826 34204 14832
rect 34164 14618 34192 14826
rect 34152 14612 34204 14618
rect 34152 14554 34204 14560
rect 34152 14476 34204 14482
rect 34152 14418 34204 14424
rect 34164 13870 34192 14418
rect 33876 13864 33928 13870
rect 33876 13806 33928 13812
rect 34152 13864 34204 13870
rect 34152 13806 34204 13812
rect 33782 13424 33838 13433
rect 33508 13388 33560 13394
rect 33782 13359 33838 13368
rect 33508 13330 33560 13336
rect 33416 13184 33468 13190
rect 33416 13126 33468 13132
rect 33428 12850 33456 13126
rect 33508 12980 33560 12986
rect 33508 12922 33560 12928
rect 33416 12844 33468 12850
rect 33416 12786 33468 12792
rect 33520 12594 33548 12922
rect 33784 12844 33836 12850
rect 33784 12786 33836 12792
rect 33428 12566 33548 12594
rect 33324 12436 33376 12442
rect 33324 12378 33376 12384
rect 33336 11898 33364 12378
rect 33324 11892 33376 11898
rect 33324 11834 33376 11840
rect 33428 11694 33456 12566
rect 33508 12436 33560 12442
rect 33508 12378 33560 12384
rect 33416 11688 33468 11694
rect 33416 11630 33468 11636
rect 33520 11626 33548 12378
rect 33796 12345 33824 12786
rect 33782 12336 33838 12345
rect 33782 12271 33838 12280
rect 33692 12232 33744 12238
rect 33692 12174 33744 12180
rect 33704 11830 33732 12174
rect 33692 11824 33744 11830
rect 33692 11766 33744 11772
rect 33508 11620 33560 11626
rect 33508 11562 33560 11568
rect 33600 11620 33652 11626
rect 33600 11562 33652 11568
rect 33232 11348 33284 11354
rect 33232 11290 33284 11296
rect 32864 11212 32916 11218
rect 32864 11154 32916 11160
rect 32772 11144 32824 11150
rect 32772 11086 32824 11092
rect 33140 11144 33192 11150
rect 33140 11086 33192 11092
rect 32588 10260 32640 10266
rect 32588 10202 32640 10208
rect 33152 10062 33180 11086
rect 33612 11082 33640 11562
rect 33704 11354 33732 11766
rect 33888 11762 33916 13806
rect 33968 13728 34020 13734
rect 33968 13670 34020 13676
rect 33980 12782 34008 13670
rect 34256 13394 34284 15098
rect 34336 14816 34388 14822
rect 34336 14758 34388 14764
rect 34348 14618 34376 14758
rect 34336 14612 34388 14618
rect 34336 14554 34388 14560
rect 34704 14612 34756 14618
rect 34704 14554 34756 14560
rect 34244 13388 34296 13394
rect 34244 13330 34296 13336
rect 34612 13388 34664 13394
rect 34612 13330 34664 13336
rect 34152 13320 34204 13326
rect 34152 13262 34204 13268
rect 34060 13184 34112 13190
rect 34060 13126 34112 13132
rect 33968 12776 34020 12782
rect 33968 12718 34020 12724
rect 34072 12714 34100 13126
rect 34164 12866 34192 13262
rect 34336 13252 34388 13258
rect 34336 13194 34388 13200
rect 34164 12850 34284 12866
rect 34164 12844 34296 12850
rect 34164 12838 34244 12844
rect 34060 12708 34112 12714
rect 34060 12650 34112 12656
rect 33966 12472 34022 12481
rect 33966 12407 34022 12416
rect 33980 12306 34008 12407
rect 34164 12374 34192 12838
rect 34244 12786 34296 12792
rect 34152 12368 34204 12374
rect 34152 12310 34204 12316
rect 34348 12306 34376 13194
rect 34520 12776 34572 12782
rect 34520 12718 34572 12724
rect 34532 12306 34560 12718
rect 34624 12646 34652 13330
rect 34612 12640 34664 12646
rect 34610 12608 34612 12617
rect 34664 12608 34666 12617
rect 34610 12543 34666 12552
rect 33968 12300 34020 12306
rect 33968 12242 34020 12248
rect 34336 12300 34388 12306
rect 34336 12242 34388 12248
rect 34520 12300 34572 12306
rect 34520 12242 34572 12248
rect 34348 11898 34376 12242
rect 34532 11898 34560 12242
rect 34152 11892 34204 11898
rect 34152 11834 34204 11840
rect 34336 11892 34388 11898
rect 34336 11834 34388 11840
rect 34520 11892 34572 11898
rect 34520 11834 34572 11840
rect 33876 11756 33928 11762
rect 33876 11698 33928 11704
rect 33692 11348 33744 11354
rect 33692 11290 33744 11296
rect 33784 11144 33836 11150
rect 33784 11086 33836 11092
rect 33600 11076 33652 11082
rect 33600 11018 33652 11024
rect 33796 10742 33824 11086
rect 33784 10736 33836 10742
rect 33784 10678 33836 10684
rect 34164 10606 34192 11834
rect 34336 11212 34388 11218
rect 34336 11154 34388 11160
rect 33692 10600 33744 10606
rect 33692 10542 33744 10548
rect 34152 10600 34204 10606
rect 34152 10542 34204 10548
rect 33232 10124 33284 10130
rect 33232 10066 33284 10072
rect 32312 10056 32364 10062
rect 32312 9998 32364 10004
rect 33140 10056 33192 10062
rect 33140 9998 33192 10004
rect 32956 9988 33008 9994
rect 32956 9930 33008 9936
rect 32144 9820 32440 9840
rect 32200 9818 32224 9820
rect 32280 9818 32304 9820
rect 32360 9818 32384 9820
rect 32222 9766 32224 9818
rect 32286 9766 32298 9818
rect 32360 9766 32362 9818
rect 32200 9764 32224 9766
rect 32280 9764 32304 9766
rect 32360 9764 32384 9766
rect 32144 9744 32440 9764
rect 31944 9648 31996 9654
rect 31944 9590 31996 9596
rect 31760 9444 31812 9450
rect 31760 9386 31812 9392
rect 32402 9072 32458 9081
rect 32458 9016 32536 9024
rect 32402 9007 32404 9016
rect 32456 8996 32536 9016
rect 32404 8978 32456 8984
rect 32144 8732 32440 8752
rect 32200 8730 32224 8732
rect 32280 8730 32304 8732
rect 32360 8730 32384 8732
rect 32222 8678 32224 8730
rect 32286 8678 32298 8730
rect 32360 8678 32362 8730
rect 32200 8676 32224 8678
rect 32280 8676 32304 8678
rect 32360 8676 32384 8678
rect 32144 8656 32440 8676
rect 32508 8634 32536 8996
rect 32772 8968 32824 8974
rect 32772 8910 32824 8916
rect 32496 8628 32548 8634
rect 32496 8570 32548 8576
rect 31852 8424 31904 8430
rect 31852 8366 31904 8372
rect 32036 8424 32088 8430
rect 32036 8366 32088 8372
rect 31864 8294 31892 8366
rect 31852 8288 31904 8294
rect 31852 8230 31904 8236
rect 32048 7410 32076 8366
rect 32312 8356 32364 8362
rect 32312 8298 32364 8304
rect 32324 8090 32352 8298
rect 32312 8084 32364 8090
rect 32312 8026 32364 8032
rect 32784 8022 32812 8910
rect 32772 8016 32824 8022
rect 32772 7958 32824 7964
rect 32496 7948 32548 7954
rect 32496 7890 32548 7896
rect 32144 7644 32440 7664
rect 32200 7642 32224 7644
rect 32280 7642 32304 7644
rect 32360 7642 32384 7644
rect 32222 7590 32224 7642
rect 32286 7590 32298 7642
rect 32360 7590 32362 7642
rect 32200 7588 32224 7590
rect 32280 7588 32304 7590
rect 32360 7588 32384 7590
rect 32144 7568 32440 7588
rect 32036 7404 32088 7410
rect 32036 7346 32088 7352
rect 31760 7200 31812 7206
rect 32404 7200 32456 7206
rect 31760 7142 31812 7148
rect 32402 7168 32404 7177
rect 32508 7188 32536 7890
rect 32456 7168 32536 7188
rect 32458 7160 32536 7168
rect 31668 6724 31720 6730
rect 31668 6666 31720 6672
rect 31680 6322 31708 6666
rect 31668 6316 31720 6322
rect 31668 6258 31720 6264
rect 31668 6180 31720 6186
rect 31772 6168 31800 7142
rect 32402 7103 32458 7112
rect 32968 6866 32996 9930
rect 33048 8288 33100 8294
rect 33048 8230 33100 8236
rect 32956 6860 33008 6866
rect 32956 6802 33008 6808
rect 32496 6792 32548 6798
rect 32496 6734 32548 6740
rect 31944 6656 31996 6662
rect 31944 6598 31996 6604
rect 31956 6458 31984 6598
rect 32144 6556 32440 6576
rect 32200 6554 32224 6556
rect 32280 6554 32304 6556
rect 32360 6554 32384 6556
rect 32222 6502 32224 6554
rect 32286 6502 32298 6554
rect 32360 6502 32362 6554
rect 32200 6500 32224 6502
rect 32280 6500 32304 6502
rect 32360 6500 32384 6502
rect 32144 6480 32440 6500
rect 31944 6452 31996 6458
rect 31944 6394 31996 6400
rect 31956 6186 31984 6394
rect 32036 6248 32088 6254
rect 32036 6190 32088 6196
rect 31720 6140 31800 6168
rect 31668 6122 31720 6128
rect 31666 6080 31722 6089
rect 31588 6038 31666 6066
rect 31390 5944 31446 5953
rect 31390 5879 31392 5888
rect 31444 5879 31446 5888
rect 31392 5850 31444 5856
rect 31024 5772 31076 5778
rect 31024 5714 31076 5720
rect 31300 5772 31352 5778
rect 31300 5714 31352 5720
rect 31036 5030 31064 5714
rect 31484 5704 31536 5710
rect 31484 5646 31536 5652
rect 31208 5636 31260 5642
rect 31208 5578 31260 5584
rect 31116 5568 31168 5574
rect 31116 5510 31168 5516
rect 31024 5024 31076 5030
rect 31024 4966 31076 4972
rect 31036 4282 31064 4966
rect 31024 4276 31076 4282
rect 31024 4218 31076 4224
rect 31024 3460 31076 3466
rect 31024 3402 31076 3408
rect 31036 2990 31064 3402
rect 31024 2984 31076 2990
rect 30930 2952 30986 2961
rect 31024 2926 31076 2932
rect 30930 2887 30986 2896
rect 31128 2514 31156 5510
rect 31220 5001 31248 5578
rect 31392 5160 31444 5166
rect 31392 5102 31444 5108
rect 31206 4992 31262 5001
rect 31206 4927 31262 4936
rect 31300 4208 31352 4214
rect 31300 4150 31352 4156
rect 31312 3369 31340 4150
rect 31404 4078 31432 5102
rect 31392 4072 31444 4078
rect 31392 4014 31444 4020
rect 31496 3942 31524 5646
rect 31588 4729 31616 6038
rect 31666 6015 31722 6024
rect 31668 5296 31720 5302
rect 31668 5238 31720 5244
rect 31680 5098 31708 5238
rect 31668 5092 31720 5098
rect 31668 5034 31720 5040
rect 31772 4758 31800 6140
rect 31944 6180 31996 6186
rect 31944 6122 31996 6128
rect 31852 6112 31904 6118
rect 31852 6054 31904 6060
rect 31942 6080 31998 6089
rect 31864 5574 31892 6054
rect 31942 6015 31998 6024
rect 31852 5568 31904 5574
rect 31852 5510 31904 5516
rect 31864 5234 31892 5510
rect 31956 5302 31984 6015
rect 32048 5953 32076 6190
rect 32508 6118 32536 6734
rect 32588 6656 32640 6662
rect 32588 6598 32640 6604
rect 32496 6112 32548 6118
rect 32496 6054 32548 6060
rect 32034 5944 32090 5953
rect 32034 5879 32090 5888
rect 31944 5296 31996 5302
rect 32048 5273 32076 5879
rect 32508 5778 32536 6054
rect 32496 5772 32548 5778
rect 32496 5714 32548 5720
rect 32144 5468 32440 5488
rect 32200 5466 32224 5468
rect 32280 5466 32304 5468
rect 32360 5466 32384 5468
rect 32222 5414 32224 5466
rect 32286 5414 32298 5466
rect 32360 5414 32362 5466
rect 32200 5412 32224 5414
rect 32280 5412 32304 5414
rect 32360 5412 32384 5414
rect 32144 5392 32440 5412
rect 32508 5370 32536 5714
rect 32600 5574 32628 6598
rect 32968 5846 32996 6802
rect 32956 5840 33008 5846
rect 32956 5782 33008 5788
rect 32588 5568 32640 5574
rect 32588 5510 32640 5516
rect 32772 5568 32824 5574
rect 32772 5510 32824 5516
rect 32496 5364 32548 5370
rect 32496 5306 32548 5312
rect 31944 5238 31996 5244
rect 32034 5264 32090 5273
rect 31852 5228 31904 5234
rect 32034 5199 32090 5208
rect 32128 5228 32180 5234
rect 31852 5170 31904 5176
rect 32128 5170 32180 5176
rect 31942 4992 31998 5001
rect 31942 4927 31998 4936
rect 31760 4752 31812 4758
rect 31574 4720 31630 4729
rect 31760 4694 31812 4700
rect 31574 4655 31630 4664
rect 31852 4548 31904 4554
rect 31852 4490 31904 4496
rect 31484 3936 31536 3942
rect 31484 3878 31536 3884
rect 31864 3738 31892 4490
rect 31956 4010 31984 4927
rect 32140 4468 32168 5170
rect 32600 5166 32628 5510
rect 32588 5160 32640 5166
rect 32588 5102 32640 5108
rect 32680 5024 32732 5030
rect 32680 4966 32732 4972
rect 32310 4856 32366 4865
rect 32310 4791 32366 4800
rect 32324 4554 32352 4791
rect 32312 4548 32364 4554
rect 32312 4490 32364 4496
rect 32496 4548 32548 4554
rect 32496 4490 32548 4496
rect 32048 4440 32168 4468
rect 32048 4282 32076 4440
rect 32144 4380 32440 4400
rect 32200 4378 32224 4380
rect 32280 4378 32304 4380
rect 32360 4378 32384 4380
rect 32222 4326 32224 4378
rect 32286 4326 32298 4378
rect 32360 4326 32362 4378
rect 32200 4324 32224 4326
rect 32280 4324 32304 4326
rect 32360 4324 32384 4326
rect 32144 4304 32440 4324
rect 32036 4276 32088 4282
rect 32036 4218 32088 4224
rect 32034 4176 32090 4185
rect 32034 4111 32090 4120
rect 32220 4140 32272 4146
rect 31944 4004 31996 4010
rect 31944 3946 31996 3952
rect 32048 3738 32076 4111
rect 32220 4082 32272 4088
rect 32232 3913 32260 4082
rect 32218 3904 32274 3913
rect 32218 3839 32274 3848
rect 31852 3732 31904 3738
rect 31852 3674 31904 3680
rect 32036 3732 32088 3738
rect 32036 3674 32088 3680
rect 31390 3632 31446 3641
rect 31390 3567 31446 3576
rect 31496 3590 31800 3618
rect 31298 3360 31354 3369
rect 31298 3295 31354 3304
rect 31208 2984 31260 2990
rect 31208 2926 31260 2932
rect 30748 2508 30800 2514
rect 30748 2450 30800 2456
rect 31116 2508 31168 2514
rect 31116 2450 31168 2456
rect 31220 2446 31248 2926
rect 31208 2440 31260 2446
rect 31208 2382 31260 2388
rect 30472 1352 30524 1358
rect 30472 1294 30524 1300
rect 30484 800 30512 1294
rect 31404 800 31432 3567
rect 31496 3233 31524 3590
rect 31772 3534 31800 3590
rect 31760 3528 31812 3534
rect 31944 3528 31996 3534
rect 31760 3470 31812 3476
rect 31850 3496 31906 3505
rect 31944 3470 31996 3476
rect 32034 3496 32090 3505
rect 31850 3431 31906 3440
rect 31482 3224 31538 3233
rect 31482 3159 31538 3168
rect 31496 2990 31524 3159
rect 31864 3126 31892 3431
rect 31852 3120 31904 3126
rect 31852 3062 31904 3068
rect 31484 2984 31536 2990
rect 31484 2926 31536 2932
rect 31956 2650 31984 3470
rect 32034 3431 32090 3440
rect 32048 3194 32076 3431
rect 32144 3292 32440 3312
rect 32200 3290 32224 3292
rect 32280 3290 32304 3292
rect 32360 3290 32384 3292
rect 32222 3238 32224 3290
rect 32286 3238 32298 3290
rect 32360 3238 32362 3290
rect 32200 3236 32224 3238
rect 32280 3236 32304 3238
rect 32360 3236 32384 3238
rect 32144 3216 32440 3236
rect 32036 3188 32088 3194
rect 32036 3130 32088 3136
rect 32128 3120 32180 3126
rect 32126 3088 32128 3097
rect 32180 3088 32182 3097
rect 32508 3058 32536 4490
rect 32586 4448 32642 4457
rect 32586 4383 32642 4392
rect 32600 4078 32628 4383
rect 32588 4072 32640 4078
rect 32588 4014 32640 4020
rect 32692 3534 32720 4966
rect 32784 4690 32812 5510
rect 32864 5364 32916 5370
rect 32864 5306 32916 5312
rect 32772 4684 32824 4690
rect 32772 4626 32824 4632
rect 32772 3936 32824 3942
rect 32876 3913 32904 5306
rect 32968 4554 32996 5782
rect 33060 5409 33088 8230
rect 33046 5400 33102 5409
rect 33046 5335 33102 5344
rect 32956 4548 33008 4554
rect 32956 4490 33008 4496
rect 32772 3878 32824 3884
rect 32862 3904 32918 3913
rect 32784 3738 32812 3878
rect 32862 3839 32918 3848
rect 32772 3732 32824 3738
rect 32772 3674 32824 3680
rect 32680 3528 32732 3534
rect 32680 3470 32732 3476
rect 32692 3194 32720 3470
rect 33060 3398 33088 5335
rect 33244 5166 33272 10066
rect 33508 10056 33560 10062
rect 33508 9998 33560 10004
rect 33520 9586 33548 9998
rect 33508 9580 33560 9586
rect 33508 9522 33560 9528
rect 33324 9512 33376 9518
rect 33324 9454 33376 9460
rect 33336 9178 33364 9454
rect 33520 9178 33548 9522
rect 33324 9172 33376 9178
rect 33324 9114 33376 9120
rect 33508 9172 33560 9178
rect 33508 9114 33560 9120
rect 33704 9110 33732 10542
rect 33876 9920 33928 9926
rect 33928 9880 34008 9908
rect 33876 9862 33928 9868
rect 33980 9518 34008 9880
rect 34164 9518 34192 10542
rect 34348 10470 34376 11154
rect 34428 11008 34480 11014
rect 34428 10950 34480 10956
rect 34336 10464 34388 10470
rect 34336 10406 34388 10412
rect 34348 10198 34376 10406
rect 34336 10192 34388 10198
rect 34336 10134 34388 10140
rect 34336 9920 34388 9926
rect 34336 9862 34388 9868
rect 34348 9654 34376 9862
rect 34336 9648 34388 9654
rect 34336 9590 34388 9596
rect 34348 9518 34376 9590
rect 33968 9512 34020 9518
rect 33968 9454 34020 9460
rect 34152 9512 34204 9518
rect 34152 9454 34204 9460
rect 34336 9512 34388 9518
rect 34336 9454 34388 9460
rect 33692 9104 33744 9110
rect 33692 9046 33744 9052
rect 33416 8832 33468 8838
rect 33416 8774 33468 8780
rect 33876 8832 33928 8838
rect 33876 8774 33928 8780
rect 33428 7002 33456 8774
rect 33692 8424 33744 8430
rect 33888 8401 33916 8774
rect 33692 8366 33744 8372
rect 33874 8392 33930 8401
rect 33704 7886 33732 8366
rect 33874 8327 33930 8336
rect 33782 8120 33838 8129
rect 33782 8055 33838 8064
rect 33796 7886 33824 8055
rect 33692 7880 33744 7886
rect 33692 7822 33744 7828
rect 33784 7880 33836 7886
rect 33784 7822 33836 7828
rect 33796 7410 33824 7822
rect 33888 7546 33916 8327
rect 33980 7750 34008 9454
rect 34440 9194 34468 10950
rect 34520 10804 34572 10810
rect 34520 10746 34572 10752
rect 34348 9166 34468 9194
rect 34532 9178 34560 10746
rect 34716 10606 34744 14554
rect 34808 14346 34836 15506
rect 35164 15360 35216 15366
rect 35164 15302 35216 15308
rect 35176 14958 35204 15302
rect 35348 15088 35400 15094
rect 35348 15030 35400 15036
rect 35164 14952 35216 14958
rect 35084 14912 35164 14940
rect 34796 14340 34848 14346
rect 34796 14282 34848 14288
rect 34888 14272 34940 14278
rect 34888 14214 34940 14220
rect 34900 13802 34928 14214
rect 34888 13796 34940 13802
rect 34888 13738 34940 13744
rect 34900 13190 34928 13738
rect 34888 13184 34940 13190
rect 34888 13126 34940 13132
rect 34980 13184 35032 13190
rect 34980 13126 35032 13132
rect 34992 12918 35020 13126
rect 34980 12912 35032 12918
rect 34980 12854 35032 12860
rect 35084 12753 35112 14912
rect 35164 14894 35216 14900
rect 35360 14550 35388 15030
rect 35440 14952 35492 14958
rect 35440 14894 35492 14900
rect 35348 14544 35400 14550
rect 35348 14486 35400 14492
rect 35452 14006 35480 14894
rect 35636 14890 35664 15846
rect 35728 15502 35756 16118
rect 35900 15904 35952 15910
rect 35900 15846 35952 15852
rect 35716 15496 35768 15502
rect 35716 15438 35768 15444
rect 35728 15094 35756 15438
rect 35716 15088 35768 15094
rect 35716 15030 35768 15036
rect 35624 14884 35676 14890
rect 35624 14826 35676 14832
rect 35348 14000 35400 14006
rect 35348 13942 35400 13948
rect 35440 14000 35492 14006
rect 35440 13942 35492 13948
rect 35636 13954 35664 14826
rect 35716 14272 35768 14278
rect 35716 14214 35768 14220
rect 35728 14074 35756 14214
rect 35716 14068 35768 14074
rect 35716 14010 35768 14016
rect 35360 13870 35388 13942
rect 35348 13864 35400 13870
rect 35348 13806 35400 13812
rect 35256 13796 35308 13802
rect 35256 13738 35308 13744
rect 35268 13190 35296 13738
rect 35348 13728 35400 13734
rect 35348 13670 35400 13676
rect 35256 13184 35308 13190
rect 35256 13126 35308 13132
rect 35256 12912 35308 12918
rect 35256 12854 35308 12860
rect 35070 12744 35126 12753
rect 34796 12708 34848 12714
rect 35070 12679 35126 12688
rect 34796 12650 34848 12656
rect 34808 12238 34836 12650
rect 35268 12442 35296 12854
rect 35360 12714 35388 13670
rect 35452 13462 35480 13942
rect 35636 13938 35756 13954
rect 35636 13932 35768 13938
rect 35636 13926 35716 13932
rect 35532 13728 35584 13734
rect 35532 13670 35584 13676
rect 35544 13530 35572 13670
rect 35532 13524 35584 13530
rect 35532 13466 35584 13472
rect 35440 13456 35492 13462
rect 35440 13398 35492 13404
rect 35348 12708 35400 12714
rect 35348 12650 35400 12656
rect 35256 12436 35308 12442
rect 35256 12378 35308 12384
rect 35636 12288 35664 13926
rect 35716 13874 35768 13880
rect 35912 13394 35940 15846
rect 36188 15706 36216 19162
rect 38120 16674 38148 19162
rect 39488 17128 39540 17134
rect 39488 17070 39540 17076
rect 39856 17128 39908 17134
rect 39856 17070 39908 17076
rect 39028 17060 39080 17066
rect 39028 17002 39080 17008
rect 38120 16646 38240 16674
rect 38212 16590 38240 16646
rect 38108 16584 38160 16590
rect 38108 16526 38160 16532
rect 38200 16584 38252 16590
rect 38200 16526 38252 16532
rect 37372 16448 37424 16454
rect 37372 16390 37424 16396
rect 37384 16046 37412 16390
rect 37372 16040 37424 16046
rect 37372 15982 37424 15988
rect 38120 15910 38148 16526
rect 38476 16448 38528 16454
rect 38476 16390 38528 16396
rect 37924 15904 37976 15910
rect 37924 15846 37976 15852
rect 38108 15904 38160 15910
rect 38108 15846 38160 15852
rect 36176 15700 36228 15706
rect 36176 15642 36228 15648
rect 36544 15564 36596 15570
rect 36544 15506 36596 15512
rect 36176 15360 36228 15366
rect 36176 15302 36228 15308
rect 36084 15088 36136 15094
rect 36084 15030 36136 15036
rect 36096 14414 36124 15030
rect 36084 14408 36136 14414
rect 36084 14350 36136 14356
rect 36096 14074 36124 14350
rect 36084 14068 36136 14074
rect 36084 14010 36136 14016
rect 35900 13388 35952 13394
rect 35900 13330 35952 13336
rect 35808 12640 35860 12646
rect 35808 12582 35860 12588
rect 35452 12260 35664 12288
rect 35716 12300 35768 12306
rect 34796 12232 34848 12238
rect 34796 12174 34848 12180
rect 34808 12102 34836 12174
rect 34796 12096 34848 12102
rect 34796 12038 34848 12044
rect 35164 11620 35216 11626
rect 35164 11562 35216 11568
rect 34704 10600 34756 10606
rect 34704 10542 34756 10548
rect 35072 10532 35124 10538
rect 35072 10474 35124 10480
rect 35084 10266 35112 10474
rect 35072 10260 35124 10266
rect 35072 10202 35124 10208
rect 34520 9172 34572 9178
rect 34244 8016 34296 8022
rect 34244 7958 34296 7964
rect 34256 7886 34284 7958
rect 34244 7880 34296 7886
rect 34164 7840 34244 7868
rect 33968 7744 34020 7750
rect 33968 7686 34020 7692
rect 33876 7540 33928 7546
rect 33876 7482 33928 7488
rect 33784 7404 33836 7410
rect 33784 7346 33836 7352
rect 33508 7200 33560 7206
rect 33508 7142 33560 7148
rect 33416 6996 33468 7002
rect 33416 6938 33468 6944
rect 33428 6798 33456 6938
rect 33416 6792 33468 6798
rect 33416 6734 33468 6740
rect 33520 6118 33548 7142
rect 33692 6792 33744 6798
rect 33692 6734 33744 6740
rect 33508 6112 33560 6118
rect 33508 6054 33560 6060
rect 33520 5574 33548 6054
rect 33600 5772 33652 5778
rect 33600 5714 33652 5720
rect 33508 5568 33560 5574
rect 33508 5510 33560 5516
rect 33508 5228 33560 5234
rect 33508 5170 33560 5176
rect 33232 5160 33284 5166
rect 33232 5102 33284 5108
rect 33324 5024 33376 5030
rect 33324 4966 33376 4972
rect 33138 4720 33194 4729
rect 33138 4655 33194 4664
rect 33152 4554 33180 4655
rect 33336 4604 33364 4966
rect 33520 4622 33548 5170
rect 33612 5030 33640 5714
rect 33600 5024 33652 5030
rect 33600 4966 33652 4972
rect 33508 4616 33560 4622
rect 33336 4576 33456 4604
rect 33140 4548 33192 4554
rect 33140 4490 33192 4496
rect 33324 4480 33376 4486
rect 33324 4422 33376 4428
rect 33138 3904 33194 3913
rect 33138 3839 33194 3848
rect 33048 3392 33100 3398
rect 33048 3334 33100 3340
rect 32770 3224 32826 3233
rect 32680 3188 32732 3194
rect 32770 3159 32826 3168
rect 32680 3130 32732 3136
rect 32126 3023 32182 3032
rect 32496 3052 32548 3058
rect 32548 3012 32628 3040
rect 32496 2994 32548 3000
rect 31944 2644 31996 2650
rect 31944 2586 31996 2592
rect 32600 2310 32628 3012
rect 32680 2916 32732 2922
rect 32680 2858 32732 2864
rect 32692 2650 32720 2858
rect 32680 2644 32732 2650
rect 32680 2586 32732 2592
rect 32588 2304 32640 2310
rect 32588 2246 32640 2252
rect 32144 2204 32440 2224
rect 32200 2202 32224 2204
rect 32280 2202 32304 2204
rect 32360 2202 32384 2204
rect 32222 2150 32224 2202
rect 32286 2150 32298 2202
rect 32360 2150 32362 2202
rect 32200 2148 32224 2150
rect 32280 2148 32304 2150
rect 32360 2148 32384 2150
rect 32144 2128 32440 2148
rect 32220 1420 32272 1426
rect 32220 1362 32272 1368
rect 32232 800 32260 1362
rect 32784 1358 32812 3159
rect 32956 2848 33008 2854
rect 32956 2790 33008 2796
rect 32968 2446 32996 2790
rect 32956 2440 33008 2446
rect 32956 2382 33008 2388
rect 32772 1352 32824 1358
rect 32772 1294 32824 1300
rect 33152 800 33180 3839
rect 33232 3392 33284 3398
rect 33232 3334 33284 3340
rect 33244 2990 33272 3334
rect 33336 3126 33364 4422
rect 33324 3120 33376 3126
rect 33324 3062 33376 3068
rect 33232 2984 33284 2990
rect 33232 2926 33284 2932
rect 33428 2922 33456 4576
rect 33508 4558 33560 4564
rect 33520 4078 33548 4558
rect 33508 4072 33560 4078
rect 33508 4014 33560 4020
rect 33508 3664 33560 3670
rect 33508 3606 33560 3612
rect 33520 3398 33548 3606
rect 33508 3392 33560 3398
rect 33508 3334 33560 3340
rect 33520 2990 33548 3334
rect 33508 2984 33560 2990
rect 33508 2926 33560 2932
rect 33416 2916 33468 2922
rect 33416 2858 33468 2864
rect 33704 2514 33732 6734
rect 33876 6452 33928 6458
rect 33876 6394 33928 6400
rect 33888 6361 33916 6394
rect 33874 6352 33930 6361
rect 33874 6287 33930 6296
rect 34164 5846 34192 7840
rect 34244 7822 34296 7828
rect 34244 6792 34296 6798
rect 34244 6734 34296 6740
rect 34256 6254 34284 6734
rect 34244 6248 34296 6254
rect 34242 6216 34244 6225
rect 34296 6216 34298 6225
rect 34242 6151 34298 6160
rect 34152 5840 34204 5846
rect 34152 5782 34204 5788
rect 34244 5160 34296 5166
rect 34244 5102 34296 5108
rect 33968 4480 34020 4486
rect 33968 4422 34020 4428
rect 33782 4312 33838 4321
rect 33980 4282 34008 4422
rect 34256 4282 34284 5102
rect 33782 4247 33838 4256
rect 33968 4276 34020 4282
rect 33796 2961 33824 4247
rect 33968 4218 34020 4224
rect 34244 4276 34296 4282
rect 34244 4218 34296 4224
rect 34256 4078 34284 4218
rect 34244 4072 34296 4078
rect 34244 4014 34296 4020
rect 33968 3596 34020 3602
rect 33968 3538 34020 3544
rect 33980 3058 34008 3538
rect 34348 3466 34376 9166
rect 34520 9114 34572 9120
rect 34532 9042 34560 9114
rect 34612 9104 34664 9110
rect 34612 9046 34664 9052
rect 34888 9104 34940 9110
rect 34888 9046 34940 9052
rect 34520 9036 34572 9042
rect 34520 8978 34572 8984
rect 34624 8090 34652 9046
rect 34704 9036 34756 9042
rect 34704 8978 34756 8984
rect 34612 8084 34664 8090
rect 34612 8026 34664 8032
rect 34520 7744 34572 7750
rect 34520 7686 34572 7692
rect 34532 6934 34560 7686
rect 34624 7546 34652 8026
rect 34716 7954 34744 8978
rect 34796 8968 34848 8974
rect 34796 8910 34848 8916
rect 34808 8634 34836 8910
rect 34900 8838 34928 9046
rect 34888 8832 34940 8838
rect 34888 8774 34940 8780
rect 35072 8832 35124 8838
rect 35072 8774 35124 8780
rect 34796 8628 34848 8634
rect 34796 8570 34848 8576
rect 35084 8430 35112 8774
rect 35176 8430 35204 11562
rect 35348 11552 35400 11558
rect 35348 11494 35400 11500
rect 35360 11218 35388 11494
rect 35452 11286 35480 12260
rect 35716 12242 35768 12248
rect 35532 12164 35584 12170
rect 35532 12106 35584 12112
rect 35544 11898 35572 12106
rect 35624 12096 35676 12102
rect 35624 12038 35676 12044
rect 35532 11892 35584 11898
rect 35532 11834 35584 11840
rect 35636 11626 35664 12038
rect 35624 11620 35676 11626
rect 35624 11562 35676 11568
rect 35440 11280 35492 11286
rect 35440 11222 35492 11228
rect 35348 11212 35400 11218
rect 35348 11154 35400 11160
rect 35452 10062 35480 11222
rect 35728 11082 35756 12242
rect 35716 11076 35768 11082
rect 35716 11018 35768 11024
rect 35820 10538 35848 12582
rect 35912 11354 35940 13330
rect 36188 13190 36216 15302
rect 36556 15026 36584 15506
rect 37188 15360 37240 15366
rect 37188 15302 37240 15308
rect 37464 15360 37516 15366
rect 37464 15302 37516 15308
rect 36452 15020 36504 15026
rect 36452 14962 36504 14968
rect 36544 15020 36596 15026
rect 36544 14962 36596 14968
rect 36464 14822 36492 14962
rect 36452 14816 36504 14822
rect 36452 14758 36504 14764
rect 36360 14544 36412 14550
rect 36360 14486 36412 14492
rect 36268 14476 36320 14482
rect 36268 14418 36320 14424
rect 36280 14278 36308 14418
rect 36268 14272 36320 14278
rect 36268 14214 36320 14220
rect 36176 13184 36228 13190
rect 36176 13126 36228 13132
rect 36188 12986 36216 13126
rect 36176 12980 36228 12986
rect 36176 12922 36228 12928
rect 36176 12776 36228 12782
rect 36176 12718 36228 12724
rect 36188 12322 36216 12718
rect 36280 12442 36308 14214
rect 36372 14074 36400 14486
rect 36360 14068 36412 14074
rect 36360 14010 36412 14016
rect 36358 13560 36414 13569
rect 36358 13495 36414 13504
rect 36372 13326 36400 13495
rect 36360 13320 36412 13326
rect 36360 13262 36412 13268
rect 36452 13184 36504 13190
rect 36452 13126 36504 13132
rect 36360 12980 36412 12986
rect 36360 12922 36412 12928
rect 36268 12436 36320 12442
rect 36268 12378 36320 12384
rect 36372 12322 36400 12922
rect 36464 12646 36492 13126
rect 36452 12640 36504 12646
rect 36452 12582 36504 12588
rect 36004 12294 36216 12322
rect 36280 12294 36400 12322
rect 35900 11348 35952 11354
rect 35900 11290 35952 11296
rect 36004 10674 36032 12294
rect 36084 12232 36136 12238
rect 36084 12174 36136 12180
rect 36096 11354 36124 12174
rect 36084 11348 36136 11354
rect 36084 11290 36136 11296
rect 35992 10668 36044 10674
rect 35992 10610 36044 10616
rect 35808 10532 35860 10538
rect 35808 10474 35860 10480
rect 36084 10124 36136 10130
rect 36084 10066 36136 10072
rect 35440 10056 35492 10062
rect 35440 9998 35492 10004
rect 35532 9920 35584 9926
rect 35532 9862 35584 9868
rect 35544 9518 35572 9862
rect 35900 9716 35952 9722
rect 35900 9658 35952 9664
rect 35532 9512 35584 9518
rect 35584 9472 35756 9500
rect 35532 9454 35584 9460
rect 35728 8974 35756 9472
rect 35532 8968 35584 8974
rect 35532 8910 35584 8916
rect 35716 8968 35768 8974
rect 35716 8910 35768 8916
rect 35072 8424 35124 8430
rect 35072 8366 35124 8372
rect 35164 8424 35216 8430
rect 35164 8366 35216 8372
rect 35440 8424 35492 8430
rect 35440 8366 35492 8372
rect 35452 8129 35480 8366
rect 35544 8294 35572 8910
rect 35532 8288 35584 8294
rect 35532 8230 35584 8236
rect 35438 8120 35494 8129
rect 35256 8084 35308 8090
rect 35438 8055 35440 8064
rect 35256 8026 35308 8032
rect 35492 8055 35494 8064
rect 35440 8026 35492 8032
rect 35268 7993 35296 8026
rect 35452 7995 35480 8026
rect 35254 7984 35310 7993
rect 34704 7948 34756 7954
rect 35254 7919 35310 7928
rect 34704 7890 34756 7896
rect 34612 7540 34664 7546
rect 34612 7482 34664 7488
rect 34716 7410 34744 7890
rect 34980 7880 35032 7886
rect 34980 7822 35032 7828
rect 34704 7404 34756 7410
rect 34704 7346 34756 7352
rect 34992 7342 35020 7822
rect 34612 7336 34664 7342
rect 34612 7278 34664 7284
rect 34980 7336 35032 7342
rect 34980 7278 35032 7284
rect 34520 6928 34572 6934
rect 34520 6870 34572 6876
rect 34624 6118 34652 7278
rect 34888 6384 34940 6390
rect 34888 6326 34940 6332
rect 34612 6112 34664 6118
rect 34612 6054 34664 6060
rect 34520 5568 34572 5574
rect 34520 5510 34572 5516
rect 34532 5098 34560 5510
rect 34520 5092 34572 5098
rect 34520 5034 34572 5040
rect 34428 4684 34480 4690
rect 34428 4626 34480 4632
rect 34440 4214 34468 4626
rect 34532 4622 34560 5034
rect 34520 4616 34572 4622
rect 34624 4593 34652 6054
rect 34900 5778 34928 6326
rect 35544 6322 35572 8230
rect 35622 8120 35678 8129
rect 35622 8055 35678 8064
rect 35636 8022 35664 8055
rect 35624 8016 35676 8022
rect 35624 7958 35676 7964
rect 35728 7886 35756 8910
rect 35912 8634 35940 9658
rect 35990 9616 36046 9625
rect 35990 9551 36046 9560
rect 36004 9382 36032 9551
rect 35992 9376 36044 9382
rect 35992 9318 36044 9324
rect 35900 8628 35952 8634
rect 35900 8570 35952 8576
rect 36096 8498 36124 10066
rect 36176 9920 36228 9926
rect 36176 9862 36228 9868
rect 36188 9518 36216 9862
rect 36176 9512 36228 9518
rect 36176 9454 36228 9460
rect 36176 9376 36228 9382
rect 36176 9318 36228 9324
rect 36084 8492 36136 8498
rect 36084 8434 36136 8440
rect 35808 8084 35860 8090
rect 35808 8026 35860 8032
rect 35716 7880 35768 7886
rect 35716 7822 35768 7828
rect 35624 6656 35676 6662
rect 35624 6598 35676 6604
rect 35636 6361 35664 6598
rect 35622 6352 35678 6361
rect 35532 6316 35584 6322
rect 35622 6287 35678 6296
rect 35532 6258 35584 6264
rect 35544 6202 35572 6258
rect 35636 6254 35664 6287
rect 35256 6180 35308 6186
rect 35256 6122 35308 6128
rect 35360 6174 35572 6202
rect 35624 6248 35676 6254
rect 35624 6190 35676 6196
rect 35268 5914 35296 6122
rect 35256 5908 35308 5914
rect 35256 5850 35308 5856
rect 35360 5778 35388 6174
rect 34888 5772 34940 5778
rect 34888 5714 34940 5720
rect 34980 5772 35032 5778
rect 34980 5714 35032 5720
rect 35164 5772 35216 5778
rect 35164 5714 35216 5720
rect 35348 5772 35400 5778
rect 35348 5714 35400 5720
rect 35440 5772 35492 5778
rect 35440 5714 35492 5720
rect 34992 5574 35020 5714
rect 35176 5642 35204 5714
rect 35164 5636 35216 5642
rect 35164 5578 35216 5584
rect 34980 5568 35032 5574
rect 34980 5510 35032 5516
rect 35256 5568 35308 5574
rect 35256 5510 35308 5516
rect 35268 5302 35296 5510
rect 35360 5370 35388 5714
rect 35348 5364 35400 5370
rect 35348 5306 35400 5312
rect 35256 5296 35308 5302
rect 35256 5238 35308 5244
rect 35452 4690 35480 5714
rect 34980 4684 35032 4690
rect 34980 4626 35032 4632
rect 35440 4684 35492 4690
rect 35440 4626 35492 4632
rect 34520 4558 34572 4564
rect 34610 4584 34666 4593
rect 34532 4282 34560 4558
rect 34610 4519 34666 4528
rect 34520 4276 34572 4282
rect 34520 4218 34572 4224
rect 34428 4208 34480 4214
rect 34428 4150 34480 4156
rect 34532 4078 34560 4218
rect 34520 4072 34572 4078
rect 34520 4014 34572 4020
rect 34992 4010 35020 4626
rect 35452 4486 35480 4626
rect 35440 4480 35492 4486
rect 35440 4422 35492 4428
rect 35636 4185 35664 6190
rect 35716 6180 35768 6186
rect 35716 6122 35768 6128
rect 35728 5574 35756 6122
rect 35716 5568 35768 5574
rect 35716 5510 35768 5516
rect 35820 4622 35848 8026
rect 35900 7880 35952 7886
rect 35900 7822 35952 7828
rect 35912 7478 35940 7822
rect 35900 7472 35952 7478
rect 35900 7414 35952 7420
rect 35992 7200 36044 7206
rect 35992 7142 36044 7148
rect 35900 6792 35952 6798
rect 35900 6734 35952 6740
rect 35912 5574 35940 6734
rect 36004 6254 36032 7142
rect 35992 6248 36044 6254
rect 35992 6190 36044 6196
rect 36004 5642 36032 6190
rect 36188 5760 36216 9318
rect 36280 8906 36308 12294
rect 36464 12102 36492 12582
rect 36452 12096 36504 12102
rect 36452 12038 36504 12044
rect 36464 11830 36492 12038
rect 36452 11824 36504 11830
rect 36452 11766 36504 11772
rect 36360 11144 36412 11150
rect 36360 11086 36412 11092
rect 36372 10810 36400 11086
rect 36452 11076 36504 11082
rect 36452 11018 36504 11024
rect 36360 10804 36412 10810
rect 36360 10746 36412 10752
rect 36464 10674 36492 11018
rect 36452 10668 36504 10674
rect 36452 10610 36504 10616
rect 36556 10062 36584 14962
rect 37200 14890 37228 15302
rect 37188 14884 37240 14890
rect 37188 14826 37240 14832
rect 37200 14618 37228 14826
rect 37188 14612 37240 14618
rect 37188 14554 37240 14560
rect 36728 14272 36780 14278
rect 36728 14214 36780 14220
rect 37004 14272 37056 14278
rect 37004 14214 37056 14220
rect 36634 13832 36690 13841
rect 36634 13767 36690 13776
rect 36648 13258 36676 13767
rect 36636 13252 36688 13258
rect 36636 13194 36688 13200
rect 36740 12782 36768 14214
rect 36820 13320 36872 13326
rect 36820 13262 36872 13268
rect 36832 13190 36860 13262
rect 36820 13184 36872 13190
rect 36820 13126 36872 13132
rect 36728 12776 36780 12782
rect 36728 12718 36780 12724
rect 36832 12238 36860 13126
rect 37016 12782 37044 14214
rect 37476 13938 37504 15302
rect 37936 14958 37964 15846
rect 38016 15360 38068 15366
rect 38016 15302 38068 15308
rect 37832 14952 37884 14958
rect 37832 14894 37884 14900
rect 37924 14952 37976 14958
rect 37924 14894 37976 14900
rect 37740 14816 37792 14822
rect 37740 14758 37792 14764
rect 37464 13932 37516 13938
rect 37464 13874 37516 13880
rect 37186 13016 37242 13025
rect 37186 12951 37242 12960
rect 37200 12782 37228 12951
rect 37752 12782 37780 14758
rect 37004 12776 37056 12782
rect 37004 12718 37056 12724
rect 37188 12776 37240 12782
rect 37188 12718 37240 12724
rect 37740 12776 37792 12782
rect 37740 12718 37792 12724
rect 36820 12232 36872 12238
rect 36820 12174 36872 12180
rect 36820 12096 36872 12102
rect 36820 12038 36872 12044
rect 36832 11762 36860 12038
rect 37016 11898 37044 12718
rect 37200 12442 37228 12718
rect 37188 12436 37240 12442
rect 37188 12378 37240 12384
rect 37752 12374 37780 12718
rect 37844 12374 37872 14894
rect 37936 14482 37964 14894
rect 37924 14476 37976 14482
rect 37924 14418 37976 14424
rect 37936 14006 37964 14418
rect 37924 14000 37976 14006
rect 37924 13942 37976 13948
rect 37924 13320 37976 13326
rect 37924 13262 37976 13268
rect 37740 12368 37792 12374
rect 37740 12310 37792 12316
rect 37832 12368 37884 12374
rect 37832 12310 37884 12316
rect 37832 12164 37884 12170
rect 37832 12106 37884 12112
rect 37004 11892 37056 11898
rect 37004 11834 37056 11840
rect 37844 11762 37872 12106
rect 36820 11756 36872 11762
rect 36820 11698 36872 11704
rect 37832 11756 37884 11762
rect 37832 11698 37884 11704
rect 36832 11286 36860 11698
rect 37464 11688 37516 11694
rect 37464 11630 37516 11636
rect 37280 11620 37332 11626
rect 37280 11562 37332 11568
rect 36820 11280 36872 11286
rect 36820 11222 36872 11228
rect 37096 11008 37148 11014
rect 37096 10950 37148 10956
rect 36636 10804 36688 10810
rect 36636 10746 36688 10752
rect 36544 10056 36596 10062
rect 36544 9998 36596 10004
rect 36556 9722 36584 9998
rect 36544 9716 36596 9722
rect 36544 9658 36596 9664
rect 36544 9444 36596 9450
rect 36544 9386 36596 9392
rect 36556 9178 36584 9386
rect 36452 9172 36504 9178
rect 36452 9114 36504 9120
rect 36544 9172 36596 9178
rect 36544 9114 36596 9120
rect 36464 9058 36492 9114
rect 36648 9058 36676 10746
rect 37108 10674 37136 10950
rect 36728 10668 36780 10674
rect 36728 10610 36780 10616
rect 37096 10668 37148 10674
rect 37096 10610 37148 10616
rect 36740 9654 36768 10610
rect 36820 10464 36872 10470
rect 36820 10406 36872 10412
rect 36832 10062 36860 10406
rect 36820 10056 36872 10062
rect 36820 9998 36872 10004
rect 36912 9920 36964 9926
rect 36912 9862 36964 9868
rect 36728 9648 36780 9654
rect 36728 9590 36780 9596
rect 36924 9518 36952 9862
rect 37096 9716 37148 9722
rect 37096 9658 37148 9664
rect 37108 9518 37136 9658
rect 36912 9512 36964 9518
rect 36912 9454 36964 9460
rect 37096 9512 37148 9518
rect 37096 9454 37148 9460
rect 37292 9110 37320 11562
rect 37370 11520 37426 11529
rect 37370 11455 37426 11464
rect 37384 11286 37412 11455
rect 37476 11354 37504 11630
rect 37464 11348 37516 11354
rect 37464 11290 37516 11296
rect 37372 11280 37424 11286
rect 37372 11222 37424 11228
rect 37936 10810 37964 13262
rect 38028 11082 38056 15302
rect 38120 14278 38148 15846
rect 38488 15502 38516 16390
rect 38936 16040 38988 16046
rect 38934 16008 38936 16017
rect 38988 16008 38990 16017
rect 38660 15972 38712 15978
rect 38934 15943 38990 15952
rect 38660 15914 38712 15920
rect 38476 15496 38528 15502
rect 38476 15438 38528 15444
rect 38672 15162 38700 15914
rect 38936 15360 38988 15366
rect 38936 15302 38988 15308
rect 38660 15156 38712 15162
rect 38660 15098 38712 15104
rect 38672 15026 38700 15098
rect 38660 15020 38712 15026
rect 38660 14962 38712 14968
rect 38384 14884 38436 14890
rect 38384 14826 38436 14832
rect 38396 14482 38424 14826
rect 38200 14476 38252 14482
rect 38200 14418 38252 14424
rect 38384 14476 38436 14482
rect 38384 14418 38436 14424
rect 38108 14272 38160 14278
rect 38108 14214 38160 14220
rect 38212 14074 38240 14418
rect 38200 14068 38252 14074
rect 38200 14010 38252 14016
rect 38108 13864 38160 13870
rect 38108 13806 38160 13812
rect 38120 13394 38148 13806
rect 38212 13462 38240 14010
rect 38292 14000 38344 14006
rect 38292 13942 38344 13948
rect 38200 13456 38252 13462
rect 38200 13398 38252 13404
rect 38304 13394 38332 13942
rect 38844 13796 38896 13802
rect 38844 13738 38896 13744
rect 38108 13388 38160 13394
rect 38108 13330 38160 13336
rect 38292 13388 38344 13394
rect 38292 13330 38344 13336
rect 38120 12986 38148 13330
rect 38856 12986 38884 13738
rect 38108 12980 38160 12986
rect 38108 12922 38160 12928
rect 38844 12980 38896 12986
rect 38844 12922 38896 12928
rect 38120 12646 38148 12922
rect 38752 12844 38804 12850
rect 38752 12786 38804 12792
rect 38660 12776 38712 12782
rect 38660 12718 38712 12724
rect 38108 12640 38160 12646
rect 38108 12582 38160 12588
rect 38292 12232 38344 12238
rect 38292 12174 38344 12180
rect 38304 11558 38332 12174
rect 38672 11626 38700 12718
rect 38764 12458 38792 12786
rect 38842 12744 38898 12753
rect 38842 12679 38898 12688
rect 38856 12646 38884 12679
rect 38844 12640 38896 12646
rect 38844 12582 38896 12588
rect 38764 12430 38884 12458
rect 38660 11620 38712 11626
rect 38660 11562 38712 11568
rect 38292 11552 38344 11558
rect 38292 11494 38344 11500
rect 38476 11348 38528 11354
rect 38476 11290 38528 11296
rect 38292 11144 38344 11150
rect 38292 11086 38344 11092
rect 38016 11076 38068 11082
rect 38016 11018 38068 11024
rect 37924 10804 37976 10810
rect 37924 10746 37976 10752
rect 38304 10606 38332 11086
rect 38292 10600 38344 10606
rect 38292 10542 38344 10548
rect 37924 10464 37976 10470
rect 37924 10406 37976 10412
rect 37936 9926 37964 10406
rect 37924 9920 37976 9926
rect 37924 9862 37976 9868
rect 37832 9648 37884 9654
rect 37830 9616 37832 9625
rect 37884 9616 37886 9625
rect 37830 9551 37886 9560
rect 37936 9518 37964 9862
rect 37924 9512 37976 9518
rect 37924 9454 37976 9460
rect 38304 9110 38332 10542
rect 38488 9654 38516 11290
rect 38568 10804 38620 10810
rect 38568 10746 38620 10752
rect 38580 10713 38608 10746
rect 38566 10704 38622 10713
rect 38566 10639 38622 10648
rect 38672 10538 38700 11562
rect 38856 11218 38884 12430
rect 38844 11212 38896 11218
rect 38844 11154 38896 11160
rect 38752 11144 38804 11150
rect 38752 11086 38804 11092
rect 38660 10532 38712 10538
rect 38660 10474 38712 10480
rect 38764 10470 38792 11086
rect 38844 10600 38896 10606
rect 38842 10568 38844 10577
rect 38896 10568 38898 10577
rect 38842 10503 38898 10512
rect 38948 10470 38976 15302
rect 39040 14550 39068 17002
rect 39212 16992 39264 16998
rect 39212 16934 39264 16940
rect 39224 16046 39252 16934
rect 39500 16590 39528 17070
rect 39488 16584 39540 16590
rect 39488 16526 39540 16532
rect 39868 16454 39896 17070
rect 40144 16794 40172 19162
rect 42076 17338 42104 19162
rect 42064 17332 42116 17338
rect 42064 17274 42116 17280
rect 40224 17128 40276 17134
rect 40224 17070 40276 17076
rect 40132 16788 40184 16794
rect 40132 16730 40184 16736
rect 39856 16448 39908 16454
rect 39856 16390 39908 16396
rect 40144 16182 40172 16730
rect 40236 16590 40264 17070
rect 40224 16584 40276 16590
rect 40224 16526 40276 16532
rect 40960 16584 41012 16590
rect 41012 16532 41092 16538
rect 40960 16526 41092 16532
rect 40132 16176 40184 16182
rect 40132 16118 40184 16124
rect 39212 16040 39264 16046
rect 39212 15982 39264 15988
rect 39224 15162 39252 15982
rect 40236 15706 40264 16526
rect 40972 16510 41092 16526
rect 40684 16448 40736 16454
rect 40684 16390 40736 16396
rect 40696 15892 40724 16390
rect 41064 15910 41092 16510
rect 41604 16516 41656 16522
rect 41604 16458 41656 16464
rect 41616 16114 41644 16458
rect 41604 16108 41656 16114
rect 41604 16050 41656 16056
rect 41616 15910 41644 16050
rect 40776 15904 40828 15910
rect 40696 15864 40776 15892
rect 40776 15846 40828 15852
rect 41052 15904 41104 15910
rect 41052 15846 41104 15852
rect 41604 15904 41656 15910
rect 41604 15846 41656 15852
rect 40040 15700 40092 15706
rect 40040 15642 40092 15648
rect 40224 15700 40276 15706
rect 40224 15642 40276 15648
rect 39856 15428 39908 15434
rect 39856 15370 39908 15376
rect 39868 15162 39896 15370
rect 39212 15156 39264 15162
rect 39212 15098 39264 15104
rect 39856 15156 39908 15162
rect 39856 15098 39908 15104
rect 39868 14550 39896 15098
rect 39028 14544 39080 14550
rect 39028 14486 39080 14492
rect 39856 14544 39908 14550
rect 39856 14486 39908 14492
rect 40052 14482 40080 15642
rect 40132 15496 40184 15502
rect 40132 15438 40184 15444
rect 40144 14890 40172 15438
rect 40500 15360 40552 15366
rect 40500 15302 40552 15308
rect 40132 14884 40184 14890
rect 40132 14826 40184 14832
rect 40040 14476 40092 14482
rect 40040 14418 40092 14424
rect 39304 14408 39356 14414
rect 39304 14350 39356 14356
rect 39488 14408 39540 14414
rect 39488 14350 39540 14356
rect 39028 14340 39080 14346
rect 39028 14282 39080 14288
rect 39040 14113 39068 14282
rect 39316 14249 39344 14350
rect 39302 14240 39358 14249
rect 39302 14175 39358 14184
rect 39026 14104 39082 14113
rect 39026 14039 39082 14048
rect 39316 13938 39344 14175
rect 39304 13932 39356 13938
rect 39304 13874 39356 13880
rect 39028 13864 39080 13870
rect 39028 13806 39080 13812
rect 39040 12646 39068 13806
rect 39212 13728 39264 13734
rect 39212 13670 39264 13676
rect 39304 13728 39356 13734
rect 39304 13670 39356 13676
rect 39224 13433 39252 13670
rect 39316 13462 39344 13670
rect 39500 13462 39528 14350
rect 40052 13938 40080 14418
rect 40040 13932 40092 13938
rect 40040 13874 40092 13880
rect 40144 13462 40172 14826
rect 40316 14612 40368 14618
rect 40316 14554 40368 14560
rect 40328 13841 40356 14554
rect 40408 14408 40460 14414
rect 40408 14350 40460 14356
rect 40314 13832 40370 13841
rect 40314 13767 40370 13776
rect 39304 13456 39356 13462
rect 39210 13424 39266 13433
rect 39304 13398 39356 13404
rect 39488 13456 39540 13462
rect 40132 13456 40184 13462
rect 39540 13404 39620 13410
rect 39488 13398 39620 13404
rect 40132 13398 40184 13404
rect 39210 13359 39266 13368
rect 39396 13388 39448 13394
rect 39500 13382 39620 13398
rect 40420 13394 40448 14350
rect 40512 13938 40540 15302
rect 40592 14816 40644 14822
rect 40592 14758 40644 14764
rect 40684 14816 40736 14822
rect 40684 14758 40736 14764
rect 40604 14482 40632 14758
rect 40592 14476 40644 14482
rect 40592 14418 40644 14424
rect 40696 13988 40724 14758
rect 40788 14550 40816 15846
rect 40866 15056 40922 15065
rect 41064 15026 41092 15846
rect 41616 15706 41644 15846
rect 41604 15700 41656 15706
rect 41604 15642 41656 15648
rect 41696 15428 41748 15434
rect 41696 15370 41748 15376
rect 40866 14991 40922 15000
rect 41052 15020 41104 15026
rect 40776 14544 40828 14550
rect 40776 14486 40828 14492
rect 40604 13960 40724 13988
rect 40500 13932 40552 13938
rect 40500 13874 40552 13880
rect 39396 13330 39448 13336
rect 39212 13184 39264 13190
rect 39212 13126 39264 13132
rect 39224 12782 39252 13126
rect 39408 12986 39436 13330
rect 39396 12980 39448 12986
rect 39396 12922 39448 12928
rect 39212 12776 39264 12782
rect 39210 12744 39212 12753
rect 39264 12744 39266 12753
rect 39210 12679 39266 12688
rect 39028 12640 39080 12646
rect 39028 12582 39080 12588
rect 39488 12640 39540 12646
rect 39488 12582 39540 12588
rect 39396 11212 39448 11218
rect 39396 11154 39448 11160
rect 39028 10736 39080 10742
rect 39028 10678 39080 10684
rect 39040 10606 39068 10678
rect 39408 10674 39436 11154
rect 39396 10668 39448 10674
rect 39396 10610 39448 10616
rect 39028 10600 39080 10606
rect 39028 10542 39080 10548
rect 38752 10464 38804 10470
rect 38752 10406 38804 10412
rect 38936 10464 38988 10470
rect 38936 10406 38988 10412
rect 38660 10124 38712 10130
rect 38660 10066 38712 10072
rect 38476 9648 38528 9654
rect 38476 9590 38528 9596
rect 38672 9450 38700 10066
rect 38764 9994 38792 10406
rect 38948 10198 38976 10406
rect 38936 10192 38988 10198
rect 38936 10134 38988 10140
rect 38752 9988 38804 9994
rect 38752 9930 38804 9936
rect 38948 9654 38976 10134
rect 39040 10130 39068 10542
rect 39028 10124 39080 10130
rect 39028 10066 39080 10072
rect 39040 9722 39068 10066
rect 39028 9716 39080 9722
rect 39028 9658 39080 9664
rect 38844 9648 38896 9654
rect 38844 9590 38896 9596
rect 38936 9648 38988 9654
rect 38936 9590 38988 9596
rect 38856 9489 38884 9590
rect 38842 9480 38898 9489
rect 38660 9444 38712 9450
rect 38842 9415 38898 9424
rect 38660 9386 38712 9392
rect 36464 9030 36676 9058
rect 37280 9104 37332 9110
rect 37280 9046 37332 9052
rect 38292 9104 38344 9110
rect 38292 9046 38344 9052
rect 36268 8900 36320 8906
rect 36268 8842 36320 8848
rect 36464 8634 36492 9030
rect 38476 8968 38528 8974
rect 38476 8910 38528 8916
rect 36728 8832 36780 8838
rect 36728 8774 36780 8780
rect 37188 8832 37240 8838
rect 37188 8774 37240 8780
rect 36452 8628 36504 8634
rect 36452 8570 36504 8576
rect 36740 8498 36768 8774
rect 36728 8492 36780 8498
rect 36728 8434 36780 8440
rect 36820 8492 36872 8498
rect 36820 8434 36872 8440
rect 36268 8288 36320 8294
rect 36268 8230 36320 8236
rect 36280 8090 36308 8230
rect 36268 8084 36320 8090
rect 36268 8026 36320 8032
rect 36634 7304 36690 7313
rect 36634 7239 36690 7248
rect 36648 7206 36676 7239
rect 36636 7200 36688 7206
rect 36636 7142 36688 7148
rect 36542 7032 36598 7041
rect 36542 6967 36598 6976
rect 36556 6730 36584 6967
rect 36452 6724 36504 6730
rect 36452 6666 36504 6672
rect 36544 6724 36596 6730
rect 36544 6666 36596 6672
rect 36096 5732 36216 5760
rect 35992 5636 36044 5642
rect 35992 5578 36044 5584
rect 35900 5568 35952 5574
rect 35900 5510 35952 5516
rect 35808 4616 35860 4622
rect 35808 4558 35860 4564
rect 35820 4282 35848 4558
rect 35808 4276 35860 4282
rect 35808 4218 35860 4224
rect 35622 4176 35678 4185
rect 35912 4162 35940 5510
rect 36004 5370 36032 5578
rect 35992 5364 36044 5370
rect 35992 5306 36044 5312
rect 36096 5166 36124 5732
rect 36176 5636 36228 5642
rect 36176 5578 36228 5584
rect 36188 5166 36216 5578
rect 36360 5568 36412 5574
rect 36360 5510 36412 5516
rect 36372 5166 36400 5510
rect 36464 5370 36492 6666
rect 36728 5568 36780 5574
rect 36728 5510 36780 5516
rect 36452 5364 36504 5370
rect 36452 5306 36504 5312
rect 36084 5160 36136 5166
rect 36084 5102 36136 5108
rect 36176 5160 36228 5166
rect 36176 5102 36228 5108
rect 36360 5160 36412 5166
rect 36360 5102 36412 5108
rect 35992 4616 36044 4622
rect 35992 4558 36044 4564
rect 35622 4111 35678 4120
rect 35820 4134 35940 4162
rect 34980 4004 35032 4010
rect 34980 3946 35032 3952
rect 34428 3596 34480 3602
rect 34428 3538 34480 3544
rect 34704 3596 34756 3602
rect 34704 3538 34756 3544
rect 34336 3460 34388 3466
rect 34336 3402 34388 3408
rect 33968 3052 34020 3058
rect 33968 2994 34020 3000
rect 33782 2952 33838 2961
rect 33782 2887 33838 2896
rect 33966 2952 34022 2961
rect 33966 2887 34022 2896
rect 33692 2508 33744 2514
rect 33692 2450 33744 2456
rect 33980 800 34008 2887
rect 34440 2310 34468 3538
rect 34520 3392 34572 3398
rect 34520 3334 34572 3340
rect 34532 3194 34560 3334
rect 34716 3194 34744 3538
rect 34886 3496 34942 3505
rect 34886 3431 34942 3440
rect 34520 3188 34572 3194
rect 34520 3130 34572 3136
rect 34704 3188 34756 3194
rect 34704 3130 34756 3136
rect 34796 2984 34848 2990
rect 34796 2926 34848 2932
rect 34808 2650 34836 2926
rect 34796 2644 34848 2650
rect 34796 2586 34848 2592
rect 34428 2304 34480 2310
rect 34428 2246 34480 2252
rect 34900 800 34928 3431
rect 35820 800 35848 4134
rect 36004 4078 36032 4558
rect 36084 4140 36136 4146
rect 36084 4082 36136 4088
rect 35992 4072 36044 4078
rect 35992 4014 36044 4020
rect 36004 3942 36032 4014
rect 35992 3936 36044 3942
rect 35992 3878 36044 3884
rect 35900 3596 35952 3602
rect 35900 3538 35952 3544
rect 35912 2854 35940 3538
rect 35900 2848 35952 2854
rect 35900 2790 35952 2796
rect 35912 2650 35940 2790
rect 35900 2644 35952 2650
rect 35900 2586 35952 2592
rect 36096 2514 36124 4082
rect 36188 3942 36216 5102
rect 36358 4720 36414 4729
rect 36464 4690 36492 5306
rect 36544 5092 36596 5098
rect 36544 5034 36596 5040
rect 36358 4655 36414 4664
rect 36452 4684 36504 4690
rect 36268 4276 36320 4282
rect 36268 4218 36320 4224
rect 36280 4078 36308 4218
rect 36268 4072 36320 4078
rect 36268 4014 36320 4020
rect 36176 3936 36228 3942
rect 36176 3878 36228 3884
rect 36188 2922 36216 3878
rect 36268 3664 36320 3670
rect 36268 3606 36320 3612
rect 36280 2990 36308 3606
rect 36372 3602 36400 4655
rect 36452 4626 36504 4632
rect 36452 4480 36504 4486
rect 36452 4422 36504 4428
rect 36464 4078 36492 4422
rect 36452 4072 36504 4078
rect 36452 4014 36504 4020
rect 36360 3596 36412 3602
rect 36360 3538 36412 3544
rect 36452 3392 36504 3398
rect 36452 3334 36504 3340
rect 36268 2984 36320 2990
rect 36268 2926 36320 2932
rect 36360 2984 36412 2990
rect 36464 2972 36492 3334
rect 36556 2990 36584 5034
rect 36634 4448 36690 4457
rect 36634 4383 36690 4392
rect 36648 3466 36676 4383
rect 36740 3738 36768 5510
rect 36832 4321 36860 8434
rect 37200 8430 37228 8774
rect 37188 8424 37240 8430
rect 37188 8366 37240 8372
rect 38488 8378 38516 8910
rect 38672 8498 38700 9386
rect 39500 9110 39528 12582
rect 39592 12442 39620 13382
rect 39672 13388 39724 13394
rect 39672 13330 39724 13336
rect 40408 13388 40460 13394
rect 40408 13330 40460 13336
rect 39580 12436 39632 12442
rect 39580 12378 39632 12384
rect 39684 12170 39712 13330
rect 39948 13320 40000 13326
rect 39948 13262 40000 13268
rect 39764 12368 39816 12374
rect 39764 12310 39816 12316
rect 39672 12164 39724 12170
rect 39672 12106 39724 12112
rect 39776 11898 39804 12310
rect 39960 12306 39988 13262
rect 40420 12986 40448 13330
rect 40408 12980 40460 12986
rect 40408 12922 40460 12928
rect 39948 12300 40000 12306
rect 39948 12242 40000 12248
rect 39856 12232 39908 12238
rect 39856 12174 39908 12180
rect 39764 11892 39816 11898
rect 39764 11834 39816 11840
rect 39868 11354 39896 12174
rect 39960 11898 39988 12242
rect 39948 11892 40000 11898
rect 39948 11834 40000 11840
rect 40408 11620 40460 11626
rect 40408 11562 40460 11568
rect 39764 11348 39816 11354
rect 39764 11290 39816 11296
rect 39856 11348 39908 11354
rect 39856 11290 39908 11296
rect 39776 11257 39804 11290
rect 39762 11248 39818 11257
rect 39762 11183 39818 11192
rect 39868 10198 39896 11290
rect 40420 11218 40448 11562
rect 40512 11286 40540 13874
rect 40604 13870 40632 13960
rect 40592 13864 40644 13870
rect 40592 13806 40644 13812
rect 40684 13864 40736 13870
rect 40684 13806 40736 13812
rect 40604 13190 40632 13806
rect 40696 13394 40724 13806
rect 40684 13388 40736 13394
rect 40684 13330 40736 13336
rect 40592 13184 40644 13190
rect 40592 13126 40644 13132
rect 40604 11286 40632 13126
rect 40696 12442 40724 13330
rect 40880 12986 40908 14991
rect 41052 14962 41104 14968
rect 41604 14952 41656 14958
rect 41604 14894 41656 14900
rect 41144 14884 41196 14890
rect 41144 14826 41196 14832
rect 41236 14884 41288 14890
rect 41236 14826 41288 14832
rect 41156 13530 41184 14826
rect 41248 14346 41276 14826
rect 41616 14550 41644 14894
rect 41708 14550 41736 15370
rect 42076 15162 42104 17274
rect 43628 17128 43680 17134
rect 43628 17070 43680 17076
rect 43076 16992 43128 16998
rect 43076 16934 43128 16940
rect 42540 16892 42836 16912
rect 42596 16890 42620 16892
rect 42676 16890 42700 16892
rect 42756 16890 42780 16892
rect 42618 16838 42620 16890
rect 42682 16838 42694 16890
rect 42756 16838 42758 16890
rect 42596 16836 42620 16838
rect 42676 16836 42700 16838
rect 42756 16836 42780 16838
rect 42540 16816 42836 16836
rect 43088 16522 43116 16934
rect 43076 16516 43128 16522
rect 42996 16476 43076 16504
rect 42156 16448 42208 16454
rect 42156 16390 42208 16396
rect 42168 16046 42196 16390
rect 42156 16040 42208 16046
rect 42156 15982 42208 15988
rect 41788 15156 41840 15162
rect 41788 15098 41840 15104
rect 42064 15156 42116 15162
rect 42064 15098 42116 15104
rect 41800 14822 41828 15098
rect 41970 15056 42026 15065
rect 42076 15026 42104 15098
rect 41970 14991 42026 15000
rect 42064 15020 42116 15026
rect 41880 14952 41932 14958
rect 41878 14920 41880 14929
rect 41932 14920 41934 14929
rect 41878 14855 41934 14864
rect 41788 14816 41840 14822
rect 41788 14758 41840 14764
rect 41604 14544 41656 14550
rect 41604 14486 41656 14492
rect 41696 14544 41748 14550
rect 41696 14486 41748 14492
rect 41236 14340 41288 14346
rect 41236 14282 41288 14288
rect 41420 14272 41472 14278
rect 41418 14240 41420 14249
rect 41472 14240 41474 14249
rect 41418 14175 41474 14184
rect 41236 14000 41288 14006
rect 41236 13942 41288 13948
rect 41052 13524 41104 13530
rect 41052 13466 41104 13472
rect 41144 13524 41196 13530
rect 41144 13466 41196 13472
rect 41064 13394 41092 13466
rect 41052 13388 41104 13394
rect 41052 13330 41104 13336
rect 41144 13252 41196 13258
rect 41144 13194 41196 13200
rect 41156 13002 41184 13194
rect 41248 13190 41276 13942
rect 41432 13802 41460 14175
rect 41420 13796 41472 13802
rect 41420 13738 41472 13744
rect 41432 13326 41460 13738
rect 41708 13530 41736 14486
rect 41984 14482 42012 14991
rect 42064 14962 42116 14968
rect 42168 14550 42196 15982
rect 42540 15804 42836 15824
rect 42596 15802 42620 15804
rect 42676 15802 42700 15804
rect 42756 15802 42780 15804
rect 42618 15750 42620 15802
rect 42682 15750 42694 15802
rect 42756 15750 42758 15802
rect 42596 15748 42620 15750
rect 42676 15748 42700 15750
rect 42756 15748 42780 15750
rect 42540 15728 42836 15748
rect 42248 15564 42300 15570
rect 42248 15506 42300 15512
rect 42260 14929 42288 15506
rect 42340 15496 42392 15502
rect 42340 15438 42392 15444
rect 42352 15144 42380 15438
rect 42892 15360 42944 15366
rect 42892 15302 42944 15308
rect 42432 15156 42484 15162
rect 42352 15116 42432 15144
rect 42352 14958 42380 15116
rect 42432 15098 42484 15104
rect 42904 14958 42932 15302
rect 42340 14952 42392 14958
rect 42246 14920 42302 14929
rect 42340 14894 42392 14900
rect 42892 14952 42944 14958
rect 42892 14894 42944 14900
rect 42246 14855 42302 14864
rect 42260 14618 42288 14855
rect 42540 14716 42836 14736
rect 42596 14714 42620 14716
rect 42676 14714 42700 14716
rect 42756 14714 42780 14716
rect 42618 14662 42620 14714
rect 42682 14662 42694 14714
rect 42756 14662 42758 14714
rect 42596 14660 42620 14662
rect 42676 14660 42700 14662
rect 42756 14660 42780 14662
rect 42540 14640 42836 14660
rect 42248 14612 42300 14618
rect 42248 14554 42300 14560
rect 42064 14544 42116 14550
rect 42064 14486 42116 14492
rect 42156 14544 42208 14550
rect 42156 14486 42208 14492
rect 41972 14476 42024 14482
rect 41972 14418 42024 14424
rect 41788 14340 41840 14346
rect 41788 14282 41840 14288
rect 41800 14074 41828 14282
rect 42076 14074 42104 14486
rect 42904 14346 42932 14894
rect 42996 14414 43024 16476
rect 43076 16458 43128 16464
rect 43444 16176 43496 16182
rect 43444 16118 43496 16124
rect 43456 15638 43484 16118
rect 43444 15632 43496 15638
rect 43444 15574 43496 15580
rect 43076 15360 43128 15366
rect 43076 15302 43128 15308
rect 43088 15094 43116 15302
rect 43076 15088 43128 15094
rect 43076 15030 43128 15036
rect 43088 14958 43116 15030
rect 43456 15026 43484 15574
rect 43640 15026 43668 17070
rect 44008 16182 44036 19162
rect 45940 17338 45968 19162
rect 45928 17332 45980 17338
rect 45928 17274 45980 17280
rect 46940 17128 46992 17134
rect 46940 17070 46992 17076
rect 47124 17128 47176 17134
rect 47124 17070 47176 17076
rect 46952 16454 46980 17070
rect 47032 16584 47084 16590
rect 47032 16526 47084 16532
rect 46940 16448 46992 16454
rect 46940 16390 46992 16396
rect 47044 16182 47072 16526
rect 43996 16176 44048 16182
rect 43996 16118 44048 16124
rect 47032 16176 47084 16182
rect 47032 16118 47084 16124
rect 46204 16040 46256 16046
rect 46202 16008 46204 16017
rect 46756 16040 46808 16046
rect 46256 16008 46258 16017
rect 46756 15982 46808 15988
rect 46202 15943 46258 15952
rect 46204 15564 46256 15570
rect 46204 15506 46256 15512
rect 43904 15360 43956 15366
rect 43904 15302 43956 15308
rect 43444 15020 43496 15026
rect 43444 14962 43496 14968
rect 43628 15020 43680 15026
rect 43628 14962 43680 14968
rect 43916 14958 43944 15302
rect 43076 14952 43128 14958
rect 43076 14894 43128 14900
rect 43168 14952 43220 14958
rect 43168 14894 43220 14900
rect 43904 14952 43956 14958
rect 43904 14894 43956 14900
rect 42984 14408 43036 14414
rect 42984 14350 43036 14356
rect 42892 14340 42944 14346
rect 42892 14282 42944 14288
rect 41788 14068 41840 14074
rect 41788 14010 41840 14016
rect 42064 14068 42116 14074
rect 42064 14010 42116 14016
rect 42524 14068 42576 14074
rect 42524 14010 42576 14016
rect 42536 13938 42564 14010
rect 42524 13932 42576 13938
rect 42524 13874 42576 13880
rect 41972 13864 42024 13870
rect 41972 13806 42024 13812
rect 42156 13864 42208 13870
rect 42156 13806 42208 13812
rect 41696 13524 41748 13530
rect 41696 13466 41748 13472
rect 41984 13326 42012 13806
rect 41420 13320 41472 13326
rect 41972 13320 42024 13326
rect 41472 13280 41552 13308
rect 41420 13262 41472 13268
rect 41236 13184 41288 13190
rect 41236 13126 41288 13132
rect 41340 13144 41460 13172
rect 41340 13002 41368 13144
rect 40868 12980 40920 12986
rect 41156 12974 41368 13002
rect 40868 12922 40920 12928
rect 40880 12782 40908 12922
rect 41328 12912 41380 12918
rect 41328 12854 41380 12860
rect 40868 12776 40920 12782
rect 41340 12753 41368 12854
rect 41432 12782 41460 13144
rect 41524 12986 41552 13280
rect 41972 13262 42024 13268
rect 41788 13184 41840 13190
rect 41788 13126 41840 13132
rect 41972 13184 42024 13190
rect 41972 13126 42024 13132
rect 41512 12980 41564 12986
rect 41512 12922 41564 12928
rect 41420 12776 41472 12782
rect 40868 12718 40920 12724
rect 41326 12744 41382 12753
rect 41420 12718 41472 12724
rect 41326 12679 41382 12688
rect 40684 12436 40736 12442
rect 40684 12378 40736 12384
rect 40868 12096 40920 12102
rect 40868 12038 40920 12044
rect 40880 11898 40908 12038
rect 40868 11892 40920 11898
rect 40868 11834 40920 11840
rect 40500 11280 40552 11286
rect 40500 11222 40552 11228
rect 40592 11280 40644 11286
rect 40592 11222 40644 11228
rect 40408 11212 40460 11218
rect 40408 11154 40460 11160
rect 40512 10742 40540 11222
rect 40500 10736 40552 10742
rect 40500 10678 40552 10684
rect 40684 10600 40736 10606
rect 40684 10542 40736 10548
rect 39856 10192 39908 10198
rect 39856 10134 39908 10140
rect 40316 10056 40368 10062
rect 40316 9998 40368 10004
rect 40328 9500 40356 9998
rect 40408 9512 40460 9518
rect 40328 9472 40408 9500
rect 40408 9454 40460 9460
rect 40040 9376 40092 9382
rect 40040 9318 40092 9324
rect 39488 9104 39540 9110
rect 39488 9046 39540 9052
rect 40052 9042 40080 9318
rect 40040 9036 40092 9042
rect 40040 8978 40092 8984
rect 38752 8968 38804 8974
rect 38752 8910 38804 8916
rect 38844 8968 38896 8974
rect 38844 8910 38896 8916
rect 38764 8634 38792 8910
rect 38752 8628 38804 8634
rect 38752 8570 38804 8576
rect 38660 8492 38712 8498
rect 38660 8434 38712 8440
rect 38384 8356 38436 8362
rect 38488 8350 38700 8378
rect 38384 8298 38436 8304
rect 38396 8129 38424 8298
rect 38382 8120 38438 8129
rect 38382 8055 38438 8064
rect 38016 8016 38068 8022
rect 38016 7958 38068 7964
rect 38476 8016 38528 8022
rect 38476 7958 38528 7964
rect 36910 7440 36966 7449
rect 36910 7375 36966 7384
rect 36924 6866 36952 7375
rect 37280 7200 37332 7206
rect 37280 7142 37332 7148
rect 36912 6860 36964 6866
rect 36912 6802 36964 6808
rect 37292 6798 37320 7142
rect 37922 6896 37978 6905
rect 37922 6831 37978 6840
rect 37280 6792 37332 6798
rect 37280 6734 37332 6740
rect 37292 5778 37320 6734
rect 37936 6390 37964 6831
rect 37924 6384 37976 6390
rect 37924 6326 37976 6332
rect 37004 5772 37056 5778
rect 37004 5714 37056 5720
rect 37280 5772 37332 5778
rect 37280 5714 37332 5720
rect 37740 5772 37792 5778
rect 37740 5714 37792 5720
rect 37016 5030 37044 5714
rect 37752 5370 37780 5714
rect 37924 5568 37976 5574
rect 37924 5510 37976 5516
rect 37740 5364 37792 5370
rect 37740 5306 37792 5312
rect 37936 5234 37964 5510
rect 38028 5370 38056 7958
rect 38292 7812 38344 7818
rect 38292 7754 38344 7760
rect 38304 5692 38332 7754
rect 38384 7268 38436 7274
rect 38384 7210 38436 7216
rect 38396 6866 38424 7210
rect 38384 6860 38436 6866
rect 38384 6802 38436 6808
rect 38396 5846 38424 6802
rect 38488 6798 38516 7958
rect 38672 7698 38700 8350
rect 38764 7818 38792 8570
rect 38856 8566 38884 8910
rect 40316 8900 40368 8906
rect 40316 8842 40368 8848
rect 38844 8560 38896 8566
rect 38844 8502 38896 8508
rect 40328 8430 40356 8842
rect 39948 8424 40000 8430
rect 40316 8424 40368 8430
rect 39948 8366 40000 8372
rect 40314 8392 40316 8401
rect 40368 8392 40370 8401
rect 39120 8084 39172 8090
rect 39120 8026 39172 8032
rect 39132 7954 39160 8026
rect 39120 7948 39172 7954
rect 39120 7890 39172 7896
rect 38752 7812 38804 7818
rect 38752 7754 38804 7760
rect 38672 7670 38792 7698
rect 38660 7200 38712 7206
rect 38660 7142 38712 7148
rect 38672 6905 38700 7142
rect 38764 7002 38792 7670
rect 39132 7206 39160 7890
rect 39304 7880 39356 7886
rect 39304 7822 39356 7828
rect 39672 7880 39724 7886
rect 39672 7822 39724 7828
rect 39212 7812 39264 7818
rect 39212 7754 39264 7760
rect 39224 7342 39252 7754
rect 39212 7336 39264 7342
rect 39212 7278 39264 7284
rect 39120 7200 39172 7206
rect 39120 7142 39172 7148
rect 38752 6996 38804 7002
rect 38752 6938 38804 6944
rect 39028 6996 39080 7002
rect 39028 6938 39080 6944
rect 38658 6896 38714 6905
rect 38658 6831 38714 6840
rect 38752 6860 38804 6866
rect 38752 6802 38804 6808
rect 38476 6792 38528 6798
rect 38476 6734 38528 6740
rect 38764 6730 38792 6802
rect 38660 6724 38712 6730
rect 38660 6666 38712 6672
rect 38752 6724 38804 6730
rect 38752 6666 38804 6672
rect 38672 6254 38700 6666
rect 38660 6248 38712 6254
rect 38936 6248 38988 6254
rect 38660 6190 38712 6196
rect 38856 6196 38936 6202
rect 38856 6190 38988 6196
rect 38384 5840 38436 5846
rect 38384 5782 38436 5788
rect 38672 5692 38700 6190
rect 38304 5664 38424 5692
rect 38396 5574 38424 5664
rect 38580 5664 38700 5692
rect 38856 6174 38976 6190
rect 38384 5568 38436 5574
rect 38384 5510 38436 5516
rect 38016 5364 38068 5370
rect 38016 5306 38068 5312
rect 37924 5228 37976 5234
rect 37924 5170 37976 5176
rect 38028 5166 38056 5306
rect 38396 5166 38424 5510
rect 38016 5160 38068 5166
rect 38016 5102 38068 5108
rect 38384 5160 38436 5166
rect 38384 5102 38436 5108
rect 37556 5092 37608 5098
rect 37556 5034 37608 5040
rect 37004 5024 37056 5030
rect 37004 4966 37056 4972
rect 37372 5024 37424 5030
rect 37372 4966 37424 4972
rect 37464 5024 37516 5030
rect 37464 4966 37516 4972
rect 36818 4312 36874 4321
rect 36818 4247 36874 4256
rect 36728 3732 36780 3738
rect 36728 3674 36780 3680
rect 36636 3460 36688 3466
rect 36636 3402 36688 3408
rect 36740 3058 36768 3674
rect 36728 3052 36780 3058
rect 36728 2994 36780 3000
rect 36912 3052 36964 3058
rect 36912 2994 36964 3000
rect 36412 2944 36492 2972
rect 36544 2984 36596 2990
rect 36360 2926 36412 2932
rect 36544 2926 36596 2932
rect 36176 2916 36228 2922
rect 36176 2858 36228 2864
rect 36084 2508 36136 2514
rect 36084 2450 36136 2456
rect 36636 2508 36688 2514
rect 36636 2450 36688 2456
rect 36648 800 36676 2450
rect 36924 1426 36952 2994
rect 37016 2582 37044 4966
rect 37188 4616 37240 4622
rect 37188 4558 37240 4564
rect 37200 4146 37228 4558
rect 37384 4486 37412 4966
rect 37372 4480 37424 4486
rect 37372 4422 37424 4428
rect 37188 4140 37240 4146
rect 37188 4082 37240 4088
rect 37476 3126 37504 4966
rect 37568 4622 37596 5034
rect 37924 4684 37976 4690
rect 37924 4626 37976 4632
rect 37556 4616 37608 4622
rect 37556 4558 37608 4564
rect 37936 4554 37964 4626
rect 38580 4554 38608 5664
rect 38752 5568 38804 5574
rect 38752 5510 38804 5516
rect 38660 4752 38712 4758
rect 38764 4729 38792 5510
rect 38660 4694 38712 4700
rect 38750 4720 38806 4729
rect 37924 4548 37976 4554
rect 37924 4490 37976 4496
rect 38568 4548 38620 4554
rect 38568 4490 38620 4496
rect 37936 4078 37964 4490
rect 37924 4072 37976 4078
rect 37924 4014 37976 4020
rect 37740 4004 37792 4010
rect 37740 3946 37792 3952
rect 37752 3738 37780 3946
rect 37740 3732 37792 3738
rect 37740 3674 37792 3680
rect 38016 3732 38068 3738
rect 38016 3674 38068 3680
rect 37464 3120 37516 3126
rect 37464 3062 37516 3068
rect 37752 2990 37780 3674
rect 38028 3369 38056 3674
rect 38476 3596 38528 3602
rect 38476 3538 38528 3544
rect 38488 3398 38516 3538
rect 38476 3392 38528 3398
rect 38014 3360 38070 3369
rect 38476 3334 38528 3340
rect 38014 3295 38070 3304
rect 38016 3188 38068 3194
rect 38016 3130 38068 3136
rect 38028 2990 38056 3130
rect 37740 2984 37792 2990
rect 37740 2926 37792 2932
rect 38016 2984 38068 2990
rect 38016 2926 38068 2932
rect 38488 2922 38516 3334
rect 38476 2916 38528 2922
rect 38476 2858 38528 2864
rect 37280 2848 37332 2854
rect 37280 2790 37332 2796
rect 37004 2576 37056 2582
rect 37004 2518 37056 2524
rect 37016 1850 37044 2518
rect 37292 2514 37320 2790
rect 37280 2508 37332 2514
rect 37280 2450 37332 2456
rect 37292 2310 37320 2450
rect 38672 2446 38700 4694
rect 38750 4655 38806 4664
rect 38752 4548 38804 4554
rect 38752 4490 38804 4496
rect 38764 4010 38792 4490
rect 38752 4004 38804 4010
rect 38752 3946 38804 3952
rect 38856 3738 38884 6174
rect 39040 5710 39068 6938
rect 39316 6730 39344 7822
rect 39684 7478 39712 7822
rect 39764 7744 39816 7750
rect 39764 7686 39816 7692
rect 39672 7472 39724 7478
rect 39672 7414 39724 7420
rect 39396 7336 39448 7342
rect 39396 7278 39448 7284
rect 39408 6866 39436 7278
rect 39684 7002 39712 7414
rect 39776 7274 39804 7686
rect 39764 7268 39816 7274
rect 39764 7210 39816 7216
rect 39672 6996 39724 7002
rect 39672 6938 39724 6944
rect 39776 6934 39804 7210
rect 39856 6996 39908 7002
rect 39856 6938 39908 6944
rect 39764 6928 39816 6934
rect 39764 6870 39816 6876
rect 39396 6860 39448 6866
rect 39396 6802 39448 6808
rect 39212 6724 39264 6730
rect 39212 6666 39264 6672
rect 39304 6724 39356 6730
rect 39304 6666 39356 6672
rect 39028 5704 39080 5710
rect 39028 5646 39080 5652
rect 39120 5636 39172 5642
rect 39120 5578 39172 5584
rect 39026 5536 39082 5545
rect 39026 5471 39082 5480
rect 39040 5302 39068 5471
rect 39132 5302 39160 5578
rect 39028 5296 39080 5302
rect 39028 5238 39080 5244
rect 39120 5296 39172 5302
rect 39120 5238 39172 5244
rect 38936 5160 38988 5166
rect 38936 5102 38988 5108
rect 38948 4078 38976 5102
rect 39028 5092 39080 5098
rect 39028 5034 39080 5040
rect 39040 4690 39068 5034
rect 39224 5030 39252 6666
rect 39408 6322 39436 6802
rect 39764 6656 39816 6662
rect 39868 6644 39896 6938
rect 39816 6616 39896 6644
rect 39764 6598 39816 6604
rect 39396 6316 39448 6322
rect 39396 6258 39448 6264
rect 39488 6112 39540 6118
rect 39488 6054 39540 6060
rect 39304 5704 39356 5710
rect 39304 5646 39356 5652
rect 39316 5166 39344 5646
rect 39304 5160 39356 5166
rect 39304 5102 39356 5108
rect 39212 5024 39264 5030
rect 39212 4966 39264 4972
rect 39028 4684 39080 4690
rect 39028 4626 39080 4632
rect 39040 4282 39068 4626
rect 39028 4276 39080 4282
rect 39028 4218 39080 4224
rect 38936 4072 38988 4078
rect 38936 4014 38988 4020
rect 38948 3738 38976 4014
rect 38844 3732 38896 3738
rect 38844 3674 38896 3680
rect 38936 3732 38988 3738
rect 38936 3674 38988 3680
rect 38752 3596 38804 3602
rect 38752 3538 38804 3544
rect 38764 3369 38792 3538
rect 38750 3360 38806 3369
rect 38750 3295 38806 3304
rect 38764 2854 38792 3295
rect 38844 2984 38896 2990
rect 38844 2926 38896 2932
rect 38752 2848 38804 2854
rect 38750 2816 38752 2825
rect 38804 2816 38806 2825
rect 38750 2751 38806 2760
rect 38660 2440 38712 2446
rect 38660 2382 38712 2388
rect 37280 2304 37332 2310
rect 37280 2246 37332 2252
rect 38476 2304 38528 2310
rect 38476 2246 38528 2252
rect 37016 1822 37596 1850
rect 36912 1420 36964 1426
rect 36912 1362 36964 1368
rect 37568 800 37596 1822
rect 38488 800 38516 2246
rect 38856 1306 38884 2926
rect 39040 2650 39068 4218
rect 39212 3528 39264 3534
rect 39212 3470 39264 3476
rect 39028 2644 39080 2650
rect 39028 2586 39080 2592
rect 39224 2582 39252 3470
rect 39500 3398 39528 6054
rect 39580 5704 39632 5710
rect 39580 5646 39632 5652
rect 39592 5370 39620 5646
rect 39776 5370 39804 6598
rect 39580 5364 39632 5370
rect 39580 5306 39632 5312
rect 39764 5364 39816 5370
rect 39764 5306 39816 5312
rect 39592 4758 39620 5306
rect 39764 4820 39816 4826
rect 39764 4762 39816 4768
rect 39580 4752 39632 4758
rect 39580 4694 39632 4700
rect 39580 4616 39632 4622
rect 39580 4558 39632 4564
rect 39592 4146 39620 4558
rect 39776 4214 39804 4762
rect 39856 4684 39908 4690
rect 39856 4626 39908 4632
rect 39868 4214 39896 4626
rect 39764 4208 39816 4214
rect 39764 4150 39816 4156
rect 39856 4208 39908 4214
rect 39856 4150 39908 4156
rect 39580 4140 39632 4146
rect 39580 4082 39632 4088
rect 39488 3392 39540 3398
rect 39488 3334 39540 3340
rect 39302 3224 39358 3233
rect 39302 3159 39358 3168
rect 39316 2990 39344 3159
rect 39960 3126 39988 8366
rect 40314 8327 40370 8336
rect 40328 7954 40356 8327
rect 40316 7948 40368 7954
rect 40316 7890 40368 7896
rect 40420 7342 40448 9454
rect 40592 8832 40644 8838
rect 40592 8774 40644 8780
rect 40604 8430 40632 8774
rect 40500 8424 40552 8430
rect 40500 8366 40552 8372
rect 40592 8424 40644 8430
rect 40592 8366 40644 8372
rect 40408 7336 40460 7342
rect 40408 7278 40460 7284
rect 40224 5704 40276 5710
rect 40420 5658 40448 7278
rect 40512 6390 40540 8366
rect 40592 7200 40644 7206
rect 40592 7142 40644 7148
rect 40500 6384 40552 6390
rect 40500 6326 40552 6332
rect 40500 6180 40552 6186
rect 40500 6122 40552 6128
rect 40512 6089 40540 6122
rect 40498 6080 40554 6089
rect 40498 6015 40554 6024
rect 40604 5930 40632 7142
rect 40224 5646 40276 5652
rect 40236 5030 40264 5646
rect 40328 5630 40448 5658
rect 40512 5902 40632 5930
rect 40224 5024 40276 5030
rect 40224 4966 40276 4972
rect 40236 4690 40264 4966
rect 40328 4865 40356 5630
rect 40512 5166 40540 5902
rect 40592 5568 40644 5574
rect 40592 5510 40644 5516
rect 40500 5160 40552 5166
rect 40500 5102 40552 5108
rect 40314 4856 40370 4865
rect 40314 4791 40370 4800
rect 40224 4684 40276 4690
rect 40224 4626 40276 4632
rect 40316 4684 40368 4690
rect 40316 4626 40368 4632
rect 40040 4548 40092 4554
rect 40040 4490 40092 4496
rect 39764 3120 39816 3126
rect 39764 3062 39816 3068
rect 39948 3120 40000 3126
rect 39948 3062 40000 3068
rect 39304 2984 39356 2990
rect 39304 2926 39356 2932
rect 39212 2576 39264 2582
rect 39026 2544 39082 2553
rect 39212 2518 39264 2524
rect 39776 2514 39804 3062
rect 39960 2990 39988 3062
rect 40052 3058 40080 4490
rect 40328 4282 40356 4626
rect 40316 4276 40368 4282
rect 40316 4218 40368 4224
rect 40408 4276 40460 4282
rect 40408 4218 40460 4224
rect 40316 3596 40368 3602
rect 40316 3538 40368 3544
rect 40132 3392 40184 3398
rect 40132 3334 40184 3340
rect 40144 3058 40172 3334
rect 40328 3233 40356 3538
rect 40314 3224 40370 3233
rect 40314 3159 40370 3168
rect 40328 3126 40356 3159
rect 40316 3120 40368 3126
rect 40316 3062 40368 3068
rect 40040 3052 40092 3058
rect 40040 2994 40092 3000
rect 40132 3052 40184 3058
rect 40132 2994 40184 3000
rect 39948 2984 40000 2990
rect 39948 2926 40000 2932
rect 40316 2848 40368 2854
rect 40236 2796 40316 2802
rect 40236 2790 40368 2796
rect 40236 2774 40356 2790
rect 39026 2479 39082 2488
rect 39764 2508 39816 2514
rect 39040 2446 39068 2479
rect 39764 2450 39816 2456
rect 39028 2440 39080 2446
rect 39028 2382 39080 2388
rect 38856 1278 39344 1306
rect 39316 800 39344 1278
rect 40236 800 40264 2774
rect 40420 2514 40448 4218
rect 40512 2990 40540 5102
rect 40604 3534 40632 5510
rect 40696 5001 40724 10542
rect 40868 10464 40920 10470
rect 40868 10406 40920 10412
rect 40880 8265 40908 10406
rect 41052 10056 41104 10062
rect 41052 9998 41104 10004
rect 41064 9081 41092 9998
rect 41432 9994 41460 12718
rect 41524 12238 41552 12922
rect 41800 12442 41828 13126
rect 41984 12646 42012 13126
rect 41972 12640 42024 12646
rect 41972 12582 42024 12588
rect 41788 12436 41840 12442
rect 41788 12378 41840 12384
rect 41880 12300 41932 12306
rect 41880 12242 41932 12248
rect 41512 12232 41564 12238
rect 41512 12174 41564 12180
rect 41524 11898 41552 12174
rect 41788 12096 41840 12102
rect 41788 12038 41840 12044
rect 41512 11892 41564 11898
rect 41512 11834 41564 11840
rect 41696 11756 41748 11762
rect 41696 11698 41748 11704
rect 41708 11218 41736 11698
rect 41800 11694 41828 12038
rect 41788 11688 41840 11694
rect 41788 11630 41840 11636
rect 41512 11212 41564 11218
rect 41512 11154 41564 11160
rect 41696 11212 41748 11218
rect 41696 11154 41748 11160
rect 41420 9988 41472 9994
rect 41420 9930 41472 9936
rect 41524 9926 41552 11154
rect 41708 10674 41736 11154
rect 41892 11082 41920 12242
rect 41984 11830 42012 12582
rect 42168 12238 42196 13806
rect 42540 13628 42836 13648
rect 42596 13626 42620 13628
rect 42676 13626 42700 13628
rect 42756 13626 42780 13628
rect 42618 13574 42620 13626
rect 42682 13574 42694 13626
rect 42756 13574 42758 13626
rect 42596 13572 42620 13574
rect 42676 13572 42700 13574
rect 42756 13572 42780 13574
rect 42540 13552 42836 13572
rect 42996 13530 43024 14350
rect 43180 14074 43208 14894
rect 46216 14890 46244 15506
rect 46204 14884 46256 14890
rect 46204 14826 46256 14832
rect 45192 14816 45244 14822
rect 45192 14758 45244 14764
rect 43444 14476 43496 14482
rect 43444 14418 43496 14424
rect 43168 14068 43220 14074
rect 43168 14010 43220 14016
rect 43350 13832 43406 13841
rect 43350 13767 43406 13776
rect 42984 13524 43036 13530
rect 42984 13466 43036 13472
rect 42996 12850 43024 13466
rect 43364 13394 43392 13767
rect 43456 13734 43484 14418
rect 43628 14340 43680 14346
rect 43628 14282 43680 14288
rect 43536 14272 43588 14278
rect 43536 14214 43588 14220
rect 43548 14074 43576 14214
rect 43536 14068 43588 14074
rect 43536 14010 43588 14016
rect 43640 13870 43668 14282
rect 43812 14272 43864 14278
rect 43812 14214 43864 14220
rect 43824 14006 43852 14214
rect 43994 14104 44050 14113
rect 43994 14039 43996 14048
rect 44048 14039 44050 14048
rect 43996 14010 44048 14016
rect 43812 14000 43864 14006
rect 43812 13942 43864 13948
rect 43904 13932 43956 13938
rect 43904 13874 43956 13880
rect 43536 13864 43588 13870
rect 43536 13806 43588 13812
rect 43628 13864 43680 13870
rect 43628 13806 43680 13812
rect 43444 13728 43496 13734
rect 43444 13670 43496 13676
rect 43548 13530 43576 13806
rect 43536 13524 43588 13530
rect 43536 13466 43588 13472
rect 43352 13388 43404 13394
rect 43352 13330 43404 13336
rect 43536 13388 43588 13394
rect 43536 13330 43588 13336
rect 43076 13184 43128 13190
rect 43076 13126 43128 13132
rect 42984 12844 43036 12850
rect 42984 12786 43036 12792
rect 42540 12540 42836 12560
rect 42596 12538 42620 12540
rect 42676 12538 42700 12540
rect 42756 12538 42780 12540
rect 42618 12486 42620 12538
rect 42682 12486 42694 12538
rect 42756 12486 42758 12538
rect 42596 12484 42620 12486
rect 42676 12484 42700 12486
rect 42756 12484 42780 12486
rect 42540 12464 42836 12484
rect 42996 12306 43024 12786
rect 43088 12442 43116 13126
rect 43364 12850 43392 13330
rect 43548 12918 43576 13330
rect 43536 12912 43588 12918
rect 43536 12854 43588 12860
rect 43352 12844 43404 12850
rect 43352 12786 43404 12792
rect 43364 12714 43392 12786
rect 43352 12708 43404 12714
rect 43352 12650 43404 12656
rect 43076 12436 43128 12442
rect 43076 12378 43128 12384
rect 42984 12300 43036 12306
rect 42984 12242 43036 12248
rect 42156 12232 42208 12238
rect 42156 12174 42208 12180
rect 41972 11824 42024 11830
rect 41972 11766 42024 11772
rect 41972 11688 42024 11694
rect 41972 11630 42024 11636
rect 41880 11076 41932 11082
rect 41880 11018 41932 11024
rect 41696 10668 41748 10674
rect 41696 10610 41748 10616
rect 41604 10192 41656 10198
rect 41604 10134 41656 10140
rect 41512 9920 41564 9926
rect 41512 9862 41564 9868
rect 41420 9648 41472 9654
rect 41420 9590 41472 9596
rect 41432 9518 41460 9590
rect 41236 9512 41288 9518
rect 41236 9454 41288 9460
rect 41420 9512 41472 9518
rect 41420 9454 41472 9460
rect 41050 9072 41106 9081
rect 41050 9007 41106 9016
rect 41064 8838 41092 9007
rect 41248 8838 41276 9454
rect 41052 8832 41104 8838
rect 41052 8774 41104 8780
rect 41236 8832 41288 8838
rect 41236 8774 41288 8780
rect 41248 8498 41276 8774
rect 41432 8634 41460 9454
rect 41420 8628 41472 8634
rect 41420 8570 41472 8576
rect 41236 8492 41288 8498
rect 41236 8434 41288 8440
rect 41524 8430 41552 9862
rect 41616 9722 41644 10134
rect 41788 10124 41840 10130
rect 41708 10084 41788 10112
rect 41604 9716 41656 9722
rect 41604 9658 41656 9664
rect 41602 9616 41658 9625
rect 41602 9551 41658 9560
rect 41616 9518 41644 9551
rect 41604 9512 41656 9518
rect 41604 9454 41656 9460
rect 41616 9382 41644 9454
rect 41708 9382 41736 10084
rect 41788 10066 41840 10072
rect 41604 9376 41656 9382
rect 41604 9318 41656 9324
rect 41696 9376 41748 9382
rect 41696 9318 41748 9324
rect 41616 8974 41644 9318
rect 41708 9042 41736 9318
rect 41696 9036 41748 9042
rect 41696 8978 41748 8984
rect 41604 8968 41656 8974
rect 41604 8910 41656 8916
rect 41512 8424 41564 8430
rect 41512 8366 41564 8372
rect 41708 8294 41736 8978
rect 41892 8634 41920 11018
rect 41984 10198 42012 11630
rect 42540 11452 42836 11472
rect 42596 11450 42620 11452
rect 42676 11450 42700 11452
rect 42756 11450 42780 11452
rect 42618 11398 42620 11450
rect 42682 11398 42694 11450
rect 42756 11398 42758 11450
rect 42596 11396 42620 11398
rect 42676 11396 42700 11398
rect 42756 11396 42780 11398
rect 42540 11376 42836 11396
rect 42064 11008 42116 11014
rect 42064 10950 42116 10956
rect 42076 10674 42104 10950
rect 42064 10668 42116 10674
rect 42064 10610 42116 10616
rect 42996 10606 43024 12242
rect 43364 11898 43392 12650
rect 43444 12232 43496 12238
rect 43444 12174 43496 12180
rect 43456 11898 43484 12174
rect 43352 11892 43404 11898
rect 43352 11834 43404 11840
rect 43444 11892 43496 11898
rect 43444 11834 43496 11840
rect 43444 11620 43496 11626
rect 43444 11562 43496 11568
rect 43456 11354 43484 11562
rect 43444 11348 43496 11354
rect 43444 11290 43496 11296
rect 43350 11248 43406 11257
rect 43350 11183 43352 11192
rect 43404 11183 43406 11192
rect 43352 11154 43404 11160
rect 43168 11144 43220 11150
rect 43168 11086 43220 11092
rect 43180 10742 43208 11086
rect 43364 10742 43392 11154
rect 43168 10736 43220 10742
rect 43168 10678 43220 10684
rect 43352 10736 43404 10742
rect 43352 10678 43404 10684
rect 42984 10600 43036 10606
rect 42984 10542 43036 10548
rect 43536 10464 43588 10470
rect 43536 10406 43588 10412
rect 42540 10364 42836 10384
rect 42596 10362 42620 10364
rect 42676 10362 42700 10364
rect 42756 10362 42780 10364
rect 42618 10310 42620 10362
rect 42682 10310 42694 10362
rect 42756 10310 42758 10362
rect 42596 10308 42620 10310
rect 42676 10308 42700 10310
rect 42756 10308 42780 10310
rect 42540 10288 42836 10308
rect 41972 10192 42024 10198
rect 41972 10134 42024 10140
rect 43548 9926 43576 10406
rect 42892 9920 42944 9926
rect 42892 9862 42944 9868
rect 43076 9920 43128 9926
rect 43076 9862 43128 9868
rect 43536 9920 43588 9926
rect 43536 9862 43588 9868
rect 42904 9586 42932 9862
rect 42892 9580 42944 9586
rect 42892 9522 42944 9528
rect 42984 9580 43036 9586
rect 42984 9522 43036 9528
rect 42340 9512 42392 9518
rect 42340 9454 42392 9460
rect 41970 9072 42026 9081
rect 41970 9007 41972 9016
rect 42024 9007 42026 9016
rect 41972 8978 42024 8984
rect 42248 8968 42300 8974
rect 42248 8910 42300 8916
rect 41972 8832 42024 8838
rect 41972 8774 42024 8780
rect 41880 8628 41932 8634
rect 41880 8570 41932 8576
rect 41984 8498 42012 8774
rect 41972 8492 42024 8498
rect 41972 8434 42024 8440
rect 41604 8288 41656 8294
rect 40866 8256 40922 8265
rect 41604 8230 41656 8236
rect 41696 8288 41748 8294
rect 41696 8230 41748 8236
rect 41880 8288 41932 8294
rect 41880 8230 41932 8236
rect 40866 8191 40922 8200
rect 40880 7857 40908 8191
rect 40866 7848 40922 7857
rect 41616 7818 41644 8230
rect 41708 7954 41736 8230
rect 41696 7948 41748 7954
rect 41696 7890 41748 7896
rect 40866 7783 40922 7792
rect 41604 7812 41656 7818
rect 41604 7754 41656 7760
rect 40868 7744 40920 7750
rect 40868 7686 40920 7692
rect 40880 5710 40908 7686
rect 41708 7546 41736 7890
rect 41892 7750 41920 8230
rect 42260 7886 42288 8910
rect 42352 8906 42380 9454
rect 42996 9382 43024 9522
rect 42984 9376 43036 9382
rect 42984 9318 43036 9324
rect 42540 9276 42836 9296
rect 42596 9274 42620 9276
rect 42676 9274 42700 9276
rect 42756 9274 42780 9276
rect 42618 9222 42620 9274
rect 42682 9222 42694 9274
rect 42756 9222 42758 9274
rect 42596 9220 42620 9222
rect 42676 9220 42700 9222
rect 42756 9220 42780 9222
rect 42540 9200 42836 9220
rect 43088 8906 43116 9862
rect 43536 9036 43588 9042
rect 43536 8978 43588 8984
rect 43352 8968 43404 8974
rect 43352 8910 43404 8916
rect 42340 8900 42392 8906
rect 42340 8842 42392 8848
rect 43076 8900 43128 8906
rect 43076 8842 43128 8848
rect 41972 7880 42024 7886
rect 41972 7822 42024 7828
rect 42248 7880 42300 7886
rect 42248 7822 42300 7828
rect 41880 7744 41932 7750
rect 41880 7686 41932 7692
rect 41984 7546 42012 7822
rect 41696 7540 41748 7546
rect 41696 7482 41748 7488
rect 41972 7540 42024 7546
rect 41972 7482 42024 7488
rect 42352 7342 42380 8842
rect 43260 8424 43312 8430
rect 43364 8412 43392 8910
rect 43312 8384 43392 8412
rect 43260 8366 43312 8372
rect 42540 8188 42836 8208
rect 42596 8186 42620 8188
rect 42676 8186 42700 8188
rect 42756 8186 42780 8188
rect 42618 8134 42620 8186
rect 42682 8134 42694 8186
rect 42756 8134 42758 8186
rect 42596 8132 42620 8134
rect 42676 8132 42700 8134
rect 42756 8132 42780 8134
rect 42540 8112 42836 8132
rect 43272 7993 43300 8366
rect 43548 8090 43576 8978
rect 43536 8084 43588 8090
rect 43536 8026 43588 8032
rect 43640 8022 43668 13806
rect 43916 13802 43944 13874
rect 43904 13796 43956 13802
rect 43904 13738 43956 13744
rect 45100 13728 45152 13734
rect 45100 13670 45152 13676
rect 44546 13424 44602 13433
rect 44546 13359 44548 13368
rect 44600 13359 44602 13368
rect 44548 13330 44600 13336
rect 43720 13184 43772 13190
rect 43720 13126 43772 13132
rect 43732 12918 43760 13126
rect 43720 12912 43772 12918
rect 43720 12854 43772 12860
rect 44560 12782 44588 13330
rect 44548 12776 44600 12782
rect 44548 12718 44600 12724
rect 44272 12708 44324 12714
rect 44272 12650 44324 12656
rect 44284 12306 44312 12650
rect 44272 12300 44324 12306
rect 44272 12242 44324 12248
rect 44916 12300 44968 12306
rect 44916 12242 44968 12248
rect 44180 12232 44232 12238
rect 44180 12174 44232 12180
rect 44456 12232 44508 12238
rect 44456 12174 44508 12180
rect 43904 11552 43956 11558
rect 43904 11494 43956 11500
rect 43916 11014 43944 11494
rect 44192 11218 44220 12174
rect 44468 11830 44496 12174
rect 44456 11824 44508 11830
rect 44456 11766 44508 11772
rect 44928 11694 44956 12242
rect 44916 11688 44968 11694
rect 44916 11630 44968 11636
rect 44548 11620 44600 11626
rect 44548 11562 44600 11568
rect 44180 11212 44232 11218
rect 44180 11154 44232 11160
rect 43904 11008 43956 11014
rect 43904 10950 43956 10956
rect 44364 11008 44416 11014
rect 44364 10950 44416 10956
rect 43916 10470 43944 10950
rect 44376 10606 44404 10950
rect 44560 10810 44588 11562
rect 45112 10810 45140 13670
rect 45204 13190 45232 14758
rect 46768 14414 46796 15982
rect 47136 15162 47164 17070
rect 47964 16726 47992 19162
rect 48136 17332 48188 17338
rect 48136 17274 48188 17280
rect 47952 16720 48004 16726
rect 47952 16662 48004 16668
rect 47308 16652 47360 16658
rect 47308 16594 47360 16600
rect 47216 16516 47268 16522
rect 47216 16458 47268 16464
rect 47228 15706 47256 16458
rect 47320 16182 47348 16594
rect 47400 16448 47452 16454
rect 47400 16390 47452 16396
rect 47308 16176 47360 16182
rect 47308 16118 47360 16124
rect 47412 16046 47440 16390
rect 47400 16040 47452 16046
rect 47400 15982 47452 15988
rect 47216 15700 47268 15706
rect 47216 15642 47268 15648
rect 47308 15360 47360 15366
rect 47308 15302 47360 15308
rect 47124 15156 47176 15162
rect 47124 15098 47176 15104
rect 47320 15094 47348 15302
rect 47308 15088 47360 15094
rect 47308 15030 47360 15036
rect 46848 14884 46900 14890
rect 46848 14826 46900 14832
rect 45836 14408 45888 14414
rect 45836 14350 45888 14356
rect 46756 14408 46808 14414
rect 46756 14350 46808 14356
rect 45848 14074 45876 14350
rect 45836 14068 45888 14074
rect 45836 14010 45888 14016
rect 45652 13796 45704 13802
rect 45652 13738 45704 13744
rect 45560 13728 45612 13734
rect 45560 13670 45612 13676
rect 45192 13184 45244 13190
rect 45192 13126 45244 13132
rect 45204 12986 45232 13126
rect 45192 12980 45244 12986
rect 45192 12922 45244 12928
rect 45572 12782 45600 13670
rect 45664 13462 45692 13738
rect 45848 13462 45876 14010
rect 46768 13870 46796 14350
rect 46860 14006 46888 14826
rect 47412 14482 47440 15982
rect 47964 15910 47992 16662
rect 47952 15904 48004 15910
rect 47952 15846 48004 15852
rect 47584 15564 47636 15570
rect 47584 15506 47636 15512
rect 47492 14612 47544 14618
rect 47492 14554 47544 14560
rect 47400 14476 47452 14482
rect 47400 14418 47452 14424
rect 47412 14346 47440 14418
rect 47400 14340 47452 14346
rect 47400 14282 47452 14288
rect 47504 14074 47532 14554
rect 47492 14068 47544 14074
rect 47492 14010 47544 14016
rect 46848 14000 46900 14006
rect 46848 13942 46900 13948
rect 46860 13870 46888 13942
rect 46756 13864 46808 13870
rect 46756 13806 46808 13812
rect 46848 13864 46900 13870
rect 46848 13806 46900 13812
rect 46112 13796 46164 13802
rect 46112 13738 46164 13744
rect 47308 13796 47360 13802
rect 47308 13738 47360 13744
rect 45652 13456 45704 13462
rect 45652 13398 45704 13404
rect 45836 13456 45888 13462
rect 45836 13398 45888 13404
rect 45560 12776 45612 12782
rect 45560 12718 45612 12724
rect 45836 12776 45888 12782
rect 45928 12776 45980 12782
rect 45836 12718 45888 12724
rect 45926 12744 45928 12753
rect 45980 12744 45982 12753
rect 45284 11756 45336 11762
rect 45284 11698 45336 11704
rect 44548 10804 44600 10810
rect 44548 10746 44600 10752
rect 45100 10804 45152 10810
rect 45100 10746 45152 10752
rect 44916 10668 44968 10674
rect 44916 10610 44968 10616
rect 44364 10600 44416 10606
rect 44364 10542 44416 10548
rect 43904 10464 43956 10470
rect 43904 10406 43956 10412
rect 44088 10464 44140 10470
rect 44088 10406 44140 10412
rect 43904 10124 43956 10130
rect 43904 10066 43956 10072
rect 43916 9926 43944 10066
rect 43904 9920 43956 9926
rect 43904 9862 43956 9868
rect 43916 9518 43944 9862
rect 43904 9512 43956 9518
rect 43904 9454 43956 9460
rect 44100 9450 44128 10406
rect 44180 9648 44232 9654
rect 44178 9616 44180 9625
rect 44232 9616 44234 9625
rect 44178 9551 44234 9560
rect 44088 9444 44140 9450
rect 44088 9386 44140 9392
rect 44100 8974 44128 9386
rect 44376 9042 44404 10542
rect 44824 10124 44876 10130
rect 44824 10066 44876 10072
rect 44836 9382 44864 10066
rect 44824 9376 44876 9382
rect 44824 9318 44876 9324
rect 44836 9110 44864 9318
rect 44824 9104 44876 9110
rect 44824 9046 44876 9052
rect 44364 9036 44416 9042
rect 44364 8978 44416 8984
rect 44088 8968 44140 8974
rect 44088 8910 44140 8916
rect 44272 8832 44324 8838
rect 44272 8774 44324 8780
rect 44640 8832 44692 8838
rect 44640 8774 44692 8780
rect 44284 8498 44312 8774
rect 44272 8492 44324 8498
rect 44272 8434 44324 8440
rect 44284 8090 44312 8434
rect 44652 8430 44680 8774
rect 44456 8424 44508 8430
rect 44456 8366 44508 8372
rect 44640 8424 44692 8430
rect 44640 8366 44692 8372
rect 44468 8090 44496 8366
rect 44272 8084 44324 8090
rect 44272 8026 44324 8032
rect 44456 8084 44508 8090
rect 44456 8026 44508 8032
rect 43628 8016 43680 8022
rect 43258 7984 43314 7993
rect 43628 7958 43680 7964
rect 43258 7919 43314 7928
rect 42432 7744 42484 7750
rect 42432 7686 42484 7692
rect 43076 7744 43128 7750
rect 43076 7686 43128 7692
rect 42444 7342 42472 7686
rect 42800 7540 42852 7546
rect 42852 7500 42932 7528
rect 42800 7482 42852 7488
rect 42340 7336 42392 7342
rect 42340 7278 42392 7284
rect 42432 7336 42484 7342
rect 42432 7278 42484 7284
rect 41052 7268 41104 7274
rect 41052 7210 41104 7216
rect 41064 6905 41092 7210
rect 41328 7200 41380 7206
rect 41328 7142 41380 7148
rect 41050 6896 41106 6905
rect 41050 6831 41106 6840
rect 41340 5914 41368 7142
rect 41604 6860 41656 6866
rect 41604 6802 41656 6808
rect 41788 6860 41840 6866
rect 41788 6802 41840 6808
rect 41616 5914 41644 6802
rect 41694 6080 41750 6089
rect 41694 6015 41750 6024
rect 41328 5908 41380 5914
rect 41328 5850 41380 5856
rect 41604 5908 41656 5914
rect 41604 5850 41656 5856
rect 41708 5778 41736 6015
rect 41696 5772 41748 5778
rect 41696 5714 41748 5720
rect 40868 5704 40920 5710
rect 40868 5646 40920 5652
rect 41144 5704 41196 5710
rect 41144 5646 41196 5652
rect 40776 5636 40828 5642
rect 40776 5578 40828 5584
rect 40788 5302 40816 5578
rect 40880 5370 40908 5646
rect 40958 5400 41014 5409
rect 40868 5364 40920 5370
rect 40958 5335 41014 5344
rect 40868 5306 40920 5312
rect 40972 5302 41000 5335
rect 40776 5296 40828 5302
rect 40776 5238 40828 5244
rect 40960 5296 41012 5302
rect 40960 5238 41012 5244
rect 41156 5234 41184 5646
rect 41800 5574 41828 6802
rect 41880 6656 41932 6662
rect 41880 6598 41932 6604
rect 41892 6254 41920 6598
rect 42444 6458 42472 7278
rect 42540 7100 42836 7120
rect 42596 7098 42620 7100
rect 42676 7098 42700 7100
rect 42756 7098 42780 7100
rect 42618 7046 42620 7098
rect 42682 7046 42694 7098
rect 42756 7046 42758 7098
rect 42596 7044 42620 7046
rect 42676 7044 42700 7046
rect 42756 7044 42780 7046
rect 42540 7024 42836 7044
rect 42524 6656 42576 6662
rect 42524 6598 42576 6604
rect 42432 6452 42484 6458
rect 42432 6394 42484 6400
rect 42064 6316 42116 6322
rect 42064 6258 42116 6264
rect 41880 6248 41932 6254
rect 41878 6216 41880 6225
rect 41932 6216 41934 6225
rect 41878 6151 41934 6160
rect 41892 5846 41920 6151
rect 41880 5840 41932 5846
rect 41880 5782 41932 5788
rect 41972 5772 42024 5778
rect 41972 5714 42024 5720
rect 41788 5568 41840 5574
rect 41788 5510 41840 5516
rect 41800 5370 41828 5510
rect 41984 5370 42012 5714
rect 41788 5364 41840 5370
rect 41788 5306 41840 5312
rect 41972 5364 42024 5370
rect 41972 5306 42024 5312
rect 41144 5228 41196 5234
rect 41144 5170 41196 5176
rect 41972 5160 42024 5166
rect 41972 5102 42024 5108
rect 41984 5030 42012 5102
rect 40868 5024 40920 5030
rect 40682 4992 40738 5001
rect 40868 4966 40920 4972
rect 41972 5024 42024 5030
rect 41972 4966 42024 4972
rect 40682 4927 40738 4936
rect 40696 3602 40724 4927
rect 40880 4486 40908 4966
rect 41972 4616 42024 4622
rect 41972 4558 42024 4564
rect 40868 4480 40920 4486
rect 40920 4440 41000 4468
rect 40868 4422 40920 4428
rect 40972 4078 41000 4440
rect 41984 4282 42012 4558
rect 41972 4276 42024 4282
rect 41972 4218 42024 4224
rect 40960 4072 41012 4078
rect 40960 4014 41012 4020
rect 41604 3936 41656 3942
rect 41604 3878 41656 3884
rect 41236 3732 41288 3738
rect 41236 3674 41288 3680
rect 40684 3596 40736 3602
rect 40684 3538 40736 3544
rect 40592 3528 40644 3534
rect 40592 3470 40644 3476
rect 40500 2984 40552 2990
rect 40500 2926 40552 2932
rect 40408 2508 40460 2514
rect 40408 2450 40460 2456
rect 40512 1970 40540 2926
rect 40604 2582 40632 3470
rect 41248 3194 41276 3674
rect 41616 3670 41644 3878
rect 41984 3738 42012 4218
rect 42076 4078 42104 6258
rect 42432 6248 42484 6254
rect 42536 6236 42564 6598
rect 42904 6458 42932 7500
rect 43088 6934 43116 7686
rect 43076 6928 43128 6934
rect 43076 6870 43128 6876
rect 42984 6792 43036 6798
rect 42984 6734 43036 6740
rect 42892 6452 42944 6458
rect 42892 6394 42944 6400
rect 42904 6254 42932 6394
rect 42484 6208 42564 6236
rect 42892 6248 42944 6254
rect 42432 6190 42484 6196
rect 42892 6190 42944 6196
rect 42246 6080 42302 6089
rect 42246 6015 42302 6024
rect 42260 5914 42288 6015
rect 42248 5908 42300 5914
rect 42248 5850 42300 5856
rect 42154 4720 42210 4729
rect 42154 4655 42156 4664
rect 42208 4655 42210 4664
rect 42156 4626 42208 4632
rect 42064 4072 42116 4078
rect 42064 4014 42116 4020
rect 42168 3942 42196 4626
rect 42444 4554 42472 6190
rect 42540 6012 42836 6032
rect 42596 6010 42620 6012
rect 42676 6010 42700 6012
rect 42756 6010 42780 6012
rect 42618 5958 42620 6010
rect 42682 5958 42694 6010
rect 42756 5958 42758 6010
rect 42596 5956 42620 5958
rect 42676 5956 42700 5958
rect 42756 5956 42780 5958
rect 42540 5936 42836 5956
rect 42904 5642 42932 6190
rect 42996 6186 43024 6734
rect 42984 6180 43036 6186
rect 42984 6122 43036 6128
rect 42996 5914 43024 6122
rect 42984 5908 43036 5914
rect 42984 5850 43036 5856
rect 42892 5636 42944 5642
rect 42892 5578 42944 5584
rect 42904 5370 42932 5578
rect 42892 5364 42944 5370
rect 42892 5306 42944 5312
rect 42904 5166 42932 5306
rect 42892 5160 42944 5166
rect 42892 5102 42944 5108
rect 42540 4924 42836 4944
rect 42596 4922 42620 4924
rect 42676 4922 42700 4924
rect 42756 4922 42780 4924
rect 42618 4870 42620 4922
rect 42682 4870 42694 4922
rect 42756 4870 42758 4922
rect 42596 4868 42620 4870
rect 42676 4868 42700 4870
rect 42756 4868 42780 4870
rect 42540 4848 42836 4868
rect 42432 4548 42484 4554
rect 42432 4490 42484 4496
rect 42444 4214 42472 4490
rect 42432 4208 42484 4214
rect 42432 4150 42484 4156
rect 42156 3936 42208 3942
rect 42156 3878 42208 3884
rect 42540 3836 42836 3856
rect 42596 3834 42620 3836
rect 42676 3834 42700 3836
rect 42756 3834 42780 3836
rect 42618 3782 42620 3834
rect 42682 3782 42694 3834
rect 42756 3782 42758 3834
rect 42596 3780 42620 3782
rect 42676 3780 42700 3782
rect 42756 3780 42780 3782
rect 42246 3768 42302 3777
rect 41972 3732 42024 3738
rect 42540 3760 42836 3780
rect 42246 3703 42302 3712
rect 41972 3674 42024 3680
rect 41420 3664 41472 3670
rect 41420 3606 41472 3612
rect 41604 3664 41656 3670
rect 41604 3606 41656 3612
rect 41236 3188 41288 3194
rect 41236 3130 41288 3136
rect 40776 3052 40828 3058
rect 40776 2994 40828 3000
rect 40788 2650 40816 2994
rect 41432 2650 41460 3606
rect 42064 3596 42116 3602
rect 42064 3538 42116 3544
rect 41970 3224 42026 3233
rect 42076 3194 42104 3538
rect 42260 3233 42288 3703
rect 43088 3602 43116 6870
rect 43272 4570 43300 7919
rect 44284 7886 44312 8026
rect 44272 7880 44324 7886
rect 44272 7822 44324 7828
rect 43352 7268 43404 7274
rect 43352 7210 43404 7216
rect 43364 6866 43392 7210
rect 44468 7206 44496 8026
rect 44456 7200 44508 7206
rect 44456 7142 44508 7148
rect 44652 6866 44680 8366
rect 44732 8356 44784 8362
rect 44732 8298 44784 8304
rect 44744 7886 44772 8298
rect 44824 7948 44876 7954
rect 44824 7890 44876 7896
rect 44732 7880 44784 7886
rect 44732 7822 44784 7828
rect 44744 7546 44772 7822
rect 44836 7546 44864 7890
rect 44732 7540 44784 7546
rect 44732 7482 44784 7488
rect 44824 7540 44876 7546
rect 44824 7482 44876 7488
rect 44732 7200 44784 7206
rect 44732 7142 44784 7148
rect 43352 6860 43404 6866
rect 43352 6802 43404 6808
rect 44640 6860 44692 6866
rect 44640 6802 44692 6808
rect 43364 6254 43392 6802
rect 43442 6760 43498 6769
rect 43442 6695 43498 6704
rect 43352 6248 43404 6254
rect 43352 6190 43404 6196
rect 43456 5846 43484 6695
rect 44180 6656 44232 6662
rect 43902 6624 43958 6633
rect 44180 6598 44232 6604
rect 43902 6559 43958 6568
rect 43720 6180 43772 6186
rect 43720 6122 43772 6128
rect 43444 5840 43496 5846
rect 43444 5782 43496 5788
rect 43352 5364 43404 5370
rect 43456 5352 43484 5782
rect 43732 5710 43760 6122
rect 43916 5778 43944 6559
rect 44088 6316 44140 6322
rect 44088 6258 44140 6264
rect 44100 5778 44128 6258
rect 43904 5772 43956 5778
rect 43904 5714 43956 5720
rect 44088 5772 44140 5778
rect 44088 5714 44140 5720
rect 43720 5704 43772 5710
rect 43720 5646 43772 5652
rect 43404 5324 43484 5352
rect 43352 5306 43404 5312
rect 43916 5302 43944 5714
rect 43904 5296 43956 5302
rect 43904 5238 43956 5244
rect 43628 5160 43680 5166
rect 43628 5102 43680 5108
rect 43640 4690 43668 5102
rect 43812 5092 43864 5098
rect 43812 5034 43864 5040
rect 43824 4758 43852 5034
rect 43812 4752 43864 4758
rect 43812 4694 43864 4700
rect 43628 4684 43680 4690
rect 43628 4626 43680 4632
rect 43180 4542 43300 4570
rect 43076 3596 43128 3602
rect 43076 3538 43128 3544
rect 42800 3392 42852 3398
rect 42800 3334 42852 3340
rect 42984 3392 43036 3398
rect 42984 3334 43036 3340
rect 42246 3224 42302 3233
rect 41970 3159 42026 3168
rect 42064 3188 42116 3194
rect 41984 3126 42012 3159
rect 42246 3159 42302 3168
rect 42064 3130 42116 3136
rect 41972 3120 42024 3126
rect 42812 3108 42840 3334
rect 42892 3120 42944 3126
rect 42812 3080 42892 3108
rect 41972 3062 42024 3068
rect 42892 3062 42944 3068
rect 42996 2990 43024 3334
rect 43180 3097 43208 4542
rect 43640 4486 43668 4626
rect 43628 4480 43680 4486
rect 43628 4422 43680 4428
rect 43640 4214 43668 4422
rect 43628 4208 43680 4214
rect 43628 4150 43680 4156
rect 43720 3596 43772 3602
rect 43720 3538 43772 3544
rect 43442 3224 43498 3233
rect 43442 3159 43444 3168
rect 43496 3159 43498 3168
rect 43628 3188 43680 3194
rect 43444 3130 43496 3136
rect 43628 3130 43680 3136
rect 43166 3088 43222 3097
rect 43166 3023 43222 3032
rect 42984 2984 43036 2990
rect 42984 2926 43036 2932
rect 42892 2916 42944 2922
rect 42892 2858 42944 2864
rect 42540 2748 42836 2768
rect 42596 2746 42620 2748
rect 42676 2746 42700 2748
rect 42756 2746 42780 2748
rect 42618 2694 42620 2746
rect 42682 2694 42694 2746
rect 42756 2694 42758 2746
rect 42596 2692 42620 2694
rect 42676 2692 42700 2694
rect 42756 2692 42780 2694
rect 42540 2672 42836 2692
rect 40776 2644 40828 2650
rect 40776 2586 40828 2592
rect 41420 2644 41472 2650
rect 41420 2586 41472 2592
rect 40592 2576 40644 2582
rect 40592 2518 40644 2524
rect 41052 2576 41104 2582
rect 41052 2518 41104 2524
rect 40500 1964 40552 1970
rect 40500 1906 40552 1912
rect 41064 800 41092 2518
rect 41972 2440 42024 2446
rect 41972 2382 42024 2388
rect 41984 800 42012 2382
rect 42156 2304 42208 2310
rect 42156 2246 42208 2252
rect 42432 2304 42484 2310
rect 42432 2246 42484 2252
rect 42168 2106 42196 2246
rect 42156 2100 42208 2106
rect 42156 2042 42208 2048
rect 42444 2038 42472 2246
rect 42904 2122 42932 2858
rect 43076 2848 43128 2854
rect 43076 2790 43128 2796
rect 43088 2378 43116 2790
rect 43076 2372 43128 2378
rect 43076 2314 43128 2320
rect 42720 2106 42932 2122
rect 42708 2100 42932 2106
rect 42760 2094 42932 2100
rect 42708 2042 42760 2048
rect 42432 2032 42484 2038
rect 42432 1974 42484 1980
rect 42904 800 42932 2094
rect 43640 1442 43668 3130
rect 43732 2854 43760 3538
rect 43916 3505 43944 5238
rect 44088 5228 44140 5234
rect 44088 5170 44140 5176
rect 44100 4758 44128 5170
rect 44192 5148 44220 6598
rect 44652 6322 44680 6802
rect 44744 6798 44772 7142
rect 44732 6792 44784 6798
rect 44732 6734 44784 6740
rect 44640 6316 44692 6322
rect 44640 6258 44692 6264
rect 44744 6254 44772 6734
rect 44364 6248 44416 6254
rect 44364 6190 44416 6196
rect 44732 6248 44784 6254
rect 44732 6190 44784 6196
rect 44822 6216 44878 6225
rect 44376 5778 44404 6190
rect 44364 5772 44416 5778
rect 44364 5714 44416 5720
rect 44456 5704 44508 5710
rect 44456 5646 44508 5652
rect 44468 5370 44496 5646
rect 44744 5642 44772 6190
rect 44928 6186 44956 10610
rect 45296 10062 45324 11698
rect 45650 11248 45706 11257
rect 45650 11183 45706 11192
rect 45376 11144 45428 11150
rect 45376 11086 45428 11092
rect 45560 11144 45612 11150
rect 45560 11086 45612 11092
rect 45388 10452 45416 11086
rect 45468 10464 45520 10470
rect 45388 10424 45468 10452
rect 45468 10406 45520 10412
rect 45284 10056 45336 10062
rect 45284 9998 45336 10004
rect 45296 9654 45324 9998
rect 45480 9994 45508 10406
rect 45572 10130 45600 11086
rect 45560 10124 45612 10130
rect 45560 10066 45612 10072
rect 45468 9988 45520 9994
rect 45468 9930 45520 9936
rect 45572 9654 45600 10066
rect 45284 9648 45336 9654
rect 45284 9590 45336 9596
rect 45560 9648 45612 9654
rect 45560 9590 45612 9596
rect 45664 9586 45692 11183
rect 45848 10470 45876 12718
rect 45926 12679 45982 12688
rect 46124 12374 46152 13738
rect 46204 13728 46256 13734
rect 46204 13670 46256 13676
rect 46216 13326 46244 13670
rect 47320 13462 47348 13738
rect 47308 13456 47360 13462
rect 47030 13424 47086 13433
rect 46848 13388 46900 13394
rect 46848 13330 46900 13336
rect 46940 13388 46992 13394
rect 47308 13398 47360 13404
rect 47030 13359 47086 13368
rect 46940 13330 46992 13336
rect 46204 13320 46256 13326
rect 46204 13262 46256 13268
rect 46572 13320 46624 13326
rect 46572 13262 46624 13268
rect 46112 12368 46164 12374
rect 46112 12310 46164 12316
rect 46584 12238 46612 13262
rect 46860 12850 46888 13330
rect 46952 12986 46980 13330
rect 47044 13326 47072 13359
rect 47032 13320 47084 13326
rect 47032 13262 47084 13268
rect 47216 13184 47268 13190
rect 47216 13126 47268 13132
rect 47228 12986 47256 13126
rect 47596 12986 47624 15506
rect 48148 14958 48176 17274
rect 49896 17134 49924 19162
rect 49976 17264 50028 17270
rect 49976 17206 50028 17212
rect 49884 17128 49936 17134
rect 49884 17070 49936 17076
rect 48780 17060 48832 17066
rect 48780 17002 48832 17008
rect 48792 16794 48820 17002
rect 49896 16794 49924 17070
rect 48780 16788 48832 16794
rect 48780 16730 48832 16736
rect 49884 16788 49936 16794
rect 49884 16730 49936 16736
rect 48228 16584 48280 16590
rect 48228 16526 48280 16532
rect 48240 14958 48268 16526
rect 48320 16448 48372 16454
rect 48320 16390 48372 16396
rect 48332 16114 48360 16390
rect 48320 16108 48372 16114
rect 48320 16050 48372 16056
rect 48332 15638 48360 16050
rect 48792 15706 48820 16730
rect 49424 16584 49476 16590
rect 49424 16526 49476 16532
rect 49436 15910 49464 16526
rect 49700 16448 49752 16454
rect 49700 16390 49752 16396
rect 49712 16250 49740 16390
rect 49700 16244 49752 16250
rect 49700 16186 49752 16192
rect 49424 15904 49476 15910
rect 49424 15846 49476 15852
rect 48780 15700 48832 15706
rect 48780 15642 48832 15648
rect 48320 15632 48372 15638
rect 48320 15574 48372 15580
rect 48792 15434 48820 15642
rect 48780 15428 48832 15434
rect 48780 15370 48832 15376
rect 48792 14958 48820 15370
rect 49436 15366 49464 15846
rect 49988 15706 50016 17206
rect 50344 17128 50396 17134
rect 50344 17070 50396 17076
rect 50356 16454 50384 17070
rect 50620 16516 50672 16522
rect 50620 16458 50672 16464
rect 50344 16448 50396 16454
rect 50344 16390 50396 16396
rect 50632 15910 50660 16458
rect 51828 16454 51856 19162
rect 52936 17436 53232 17456
rect 52992 17434 53016 17436
rect 53072 17434 53096 17436
rect 53152 17434 53176 17436
rect 53014 17382 53016 17434
rect 53078 17382 53090 17434
rect 53152 17382 53154 17434
rect 52992 17380 53016 17382
rect 53072 17380 53096 17382
rect 53152 17380 53176 17382
rect 52936 17360 53232 17380
rect 53852 17338 53880 19162
rect 53840 17332 53892 17338
rect 53840 17274 53892 17280
rect 52828 17060 52880 17066
rect 52828 17002 52880 17008
rect 52092 16584 52144 16590
rect 52092 16526 52144 16532
rect 51816 16448 51868 16454
rect 51816 16390 51868 16396
rect 52104 16250 52132 16526
rect 52092 16244 52144 16250
rect 52092 16186 52144 16192
rect 51632 16176 51684 16182
rect 51092 16102 51580 16130
rect 51632 16118 51684 16124
rect 51092 15910 51120 16102
rect 51552 16046 51580 16102
rect 51448 16040 51500 16046
rect 51448 15982 51500 15988
rect 51540 16040 51592 16046
rect 51540 15982 51592 15988
rect 50620 15904 50672 15910
rect 50620 15846 50672 15852
rect 50988 15904 51040 15910
rect 50988 15846 51040 15852
rect 51080 15904 51132 15910
rect 51080 15846 51132 15852
rect 49976 15700 50028 15706
rect 49976 15642 50028 15648
rect 49608 15564 49660 15570
rect 49608 15506 49660 15512
rect 49148 15360 49200 15366
rect 49148 15302 49200 15308
rect 49424 15360 49476 15366
rect 49424 15302 49476 15308
rect 49160 15094 49188 15302
rect 49148 15088 49200 15094
rect 49148 15030 49200 15036
rect 48136 14952 48188 14958
rect 48136 14894 48188 14900
rect 48228 14952 48280 14958
rect 48228 14894 48280 14900
rect 48780 14952 48832 14958
rect 48780 14894 48832 14900
rect 48240 14482 48268 14894
rect 48964 14816 49016 14822
rect 48964 14758 49016 14764
rect 48976 14482 49004 14758
rect 49160 14550 49188 15030
rect 49148 14544 49200 14550
rect 49148 14486 49200 14492
rect 48228 14476 48280 14482
rect 48228 14418 48280 14424
rect 48964 14476 49016 14482
rect 48964 14418 49016 14424
rect 47768 14408 47820 14414
rect 47768 14350 47820 14356
rect 46940 12980 46992 12986
rect 46940 12922 46992 12928
rect 47216 12980 47268 12986
rect 47216 12922 47268 12928
rect 47584 12980 47636 12986
rect 47584 12922 47636 12928
rect 47124 12912 47176 12918
rect 47124 12854 47176 12860
rect 46848 12844 46900 12850
rect 46848 12786 46900 12792
rect 46860 12306 46888 12786
rect 46940 12708 46992 12714
rect 46940 12650 46992 12656
rect 46848 12300 46900 12306
rect 46848 12242 46900 12248
rect 46952 12238 46980 12650
rect 47032 12300 47084 12306
rect 47032 12242 47084 12248
rect 46572 12232 46624 12238
rect 46572 12174 46624 12180
rect 46664 12232 46716 12238
rect 46664 12174 46716 12180
rect 46940 12232 46992 12238
rect 46940 12174 46992 12180
rect 46676 11286 46704 12174
rect 47044 12170 47072 12242
rect 47032 12164 47084 12170
rect 47032 12106 47084 12112
rect 47044 11694 47072 12106
rect 46848 11688 46900 11694
rect 46848 11630 46900 11636
rect 47032 11688 47084 11694
rect 47032 11630 47084 11636
rect 46664 11280 46716 11286
rect 46664 11222 46716 11228
rect 46860 11150 46888 11630
rect 46848 11144 46900 11150
rect 46848 11086 46900 11092
rect 46664 10804 46716 10810
rect 46664 10746 46716 10752
rect 45836 10464 45888 10470
rect 45836 10406 45888 10412
rect 45848 10266 45876 10406
rect 45836 10260 45888 10266
rect 45836 10202 45888 10208
rect 46020 10192 46072 10198
rect 46020 10134 46072 10140
rect 45652 9580 45704 9586
rect 45652 9522 45704 9528
rect 46032 9518 46060 10134
rect 46676 10130 46704 10746
rect 46940 10668 46992 10674
rect 46940 10610 46992 10616
rect 46952 10577 46980 10610
rect 46938 10568 46994 10577
rect 46938 10503 46994 10512
rect 46664 10124 46716 10130
rect 46664 10066 46716 10072
rect 46480 9920 46532 9926
rect 46400 9880 46480 9908
rect 46020 9512 46072 9518
rect 46020 9454 46072 9460
rect 45100 8968 45152 8974
rect 45100 8910 45152 8916
rect 45112 8294 45140 8910
rect 46112 8900 46164 8906
rect 46112 8842 46164 8848
rect 45560 8628 45612 8634
rect 45560 8570 45612 8576
rect 45468 8356 45520 8362
rect 45468 8298 45520 8304
rect 45100 8288 45152 8294
rect 45100 8230 45152 8236
rect 45112 8022 45140 8230
rect 45480 8090 45508 8298
rect 45468 8084 45520 8090
rect 45468 8026 45520 8032
rect 45100 8016 45152 8022
rect 45100 7958 45152 7964
rect 45192 7948 45244 7954
rect 45192 7890 45244 7896
rect 45204 7274 45232 7890
rect 45572 7478 45600 8570
rect 45744 8356 45796 8362
rect 45744 8298 45796 8304
rect 45756 8090 45784 8298
rect 45744 8084 45796 8090
rect 45744 8026 45796 8032
rect 45652 8016 45704 8022
rect 45652 7958 45704 7964
rect 45560 7472 45612 7478
rect 45560 7414 45612 7420
rect 45192 7268 45244 7274
rect 45192 7210 45244 7216
rect 45204 7002 45232 7210
rect 45192 6996 45244 7002
rect 45192 6938 45244 6944
rect 45572 6934 45600 7414
rect 45664 6934 45692 7958
rect 46124 7410 46152 8842
rect 46296 8832 46348 8838
rect 46296 8774 46348 8780
rect 46308 8634 46336 8774
rect 46296 8628 46348 8634
rect 46296 8570 46348 8576
rect 46308 8498 46336 8570
rect 46296 8492 46348 8498
rect 46296 8434 46348 8440
rect 46204 7744 46256 7750
rect 46202 7712 46204 7721
rect 46256 7712 46258 7721
rect 46202 7647 46258 7656
rect 46112 7404 46164 7410
rect 46112 7346 46164 7352
rect 46124 7313 46152 7346
rect 46110 7304 46166 7313
rect 46216 7274 46244 7647
rect 46308 7274 46336 8434
rect 46110 7239 46166 7248
rect 46204 7268 46256 7274
rect 46204 7210 46256 7216
rect 46296 7268 46348 7274
rect 46296 7210 46348 7216
rect 45560 6928 45612 6934
rect 45560 6870 45612 6876
rect 45652 6928 45704 6934
rect 45652 6870 45704 6876
rect 45100 6724 45152 6730
rect 45100 6666 45152 6672
rect 44822 6151 44878 6160
rect 44916 6180 44968 6186
rect 44836 5642 44864 6151
rect 44916 6122 44968 6128
rect 44732 5636 44784 5642
rect 44732 5578 44784 5584
rect 44824 5636 44876 5642
rect 44824 5578 44876 5584
rect 44456 5364 44508 5370
rect 44456 5306 44508 5312
rect 44732 5364 44784 5370
rect 44732 5306 44784 5312
rect 44548 5160 44600 5166
rect 44192 5120 44548 5148
rect 44548 5102 44600 5108
rect 44088 4752 44140 4758
rect 44088 4694 44140 4700
rect 44180 4480 44232 4486
rect 44180 4422 44232 4428
rect 44192 4282 44220 4422
rect 44180 4276 44232 4282
rect 44180 4218 44232 4224
rect 44180 4004 44232 4010
rect 44180 3946 44232 3952
rect 44192 3505 44220 3946
rect 44744 3942 44772 5306
rect 44836 5234 44864 5578
rect 44824 5228 44876 5234
rect 44824 5170 44876 5176
rect 44732 3936 44784 3942
rect 44732 3878 44784 3884
rect 44824 3936 44876 3942
rect 44824 3878 44876 3884
rect 44640 3528 44692 3534
rect 43902 3496 43958 3505
rect 43902 3431 43958 3440
rect 44178 3496 44234 3505
rect 44640 3470 44692 3476
rect 44178 3431 44234 3440
rect 43996 3392 44048 3398
rect 43996 3334 44048 3340
rect 44272 3392 44324 3398
rect 44272 3334 44324 3340
rect 44008 3194 44036 3334
rect 43996 3188 44048 3194
rect 43996 3130 44048 3136
rect 43996 2916 44048 2922
rect 43996 2858 44048 2864
rect 43720 2848 43772 2854
rect 43720 2790 43772 2796
rect 44008 2650 44036 2858
rect 43996 2644 44048 2650
rect 43996 2586 44048 2592
rect 44284 2446 44312 3334
rect 44652 2666 44680 3470
rect 44744 2990 44772 3878
rect 44836 3670 44864 3878
rect 44824 3664 44876 3670
rect 44824 3606 44876 3612
rect 44824 3460 44876 3466
rect 44824 3402 44876 3408
rect 44732 2984 44784 2990
rect 44732 2926 44784 2932
rect 44836 2825 44864 3402
rect 44928 3097 44956 6122
rect 45112 5778 45140 6666
rect 45572 6458 45600 6870
rect 46204 6860 46256 6866
rect 46204 6802 46256 6808
rect 46112 6656 46164 6662
rect 46112 6598 46164 6604
rect 45560 6452 45612 6458
rect 45560 6394 45612 6400
rect 46124 6254 46152 6598
rect 46216 6458 46244 6802
rect 46400 6798 46428 9880
rect 46480 9862 46532 9868
rect 46676 9654 46704 10066
rect 47044 9654 47072 11630
rect 47136 9994 47164 12854
rect 47308 12844 47360 12850
rect 47308 12786 47360 12792
rect 47320 10266 47348 12786
rect 47492 11620 47544 11626
rect 47492 11562 47544 11568
rect 47400 10464 47452 10470
rect 47400 10406 47452 10412
rect 47308 10260 47360 10266
rect 47308 10202 47360 10208
rect 47412 10198 47440 10406
rect 47400 10192 47452 10198
rect 47400 10134 47452 10140
rect 47216 10056 47268 10062
rect 47216 9998 47268 10004
rect 47124 9988 47176 9994
rect 47124 9930 47176 9936
rect 47228 9926 47256 9998
rect 47216 9920 47268 9926
rect 47216 9862 47268 9868
rect 46664 9648 46716 9654
rect 46664 9590 46716 9596
rect 47032 9648 47084 9654
rect 47032 9590 47084 9596
rect 47228 9450 47256 9862
rect 47504 9625 47532 11562
rect 47584 11212 47636 11218
rect 47584 11154 47636 11160
rect 47596 10810 47624 11154
rect 47584 10804 47636 10810
rect 47584 10746 47636 10752
rect 47584 10464 47636 10470
rect 47584 10406 47636 10412
rect 47596 10130 47624 10406
rect 47780 10266 47808 14350
rect 48044 14340 48096 14346
rect 48044 14282 48096 14288
rect 48056 13274 48084 14282
rect 48320 14272 48372 14278
rect 48320 14214 48372 14220
rect 48332 14074 48360 14214
rect 48976 14074 49004 14418
rect 49620 14278 49648 15506
rect 50252 15496 50304 15502
rect 50252 15438 50304 15444
rect 49792 14952 49844 14958
rect 49792 14894 49844 14900
rect 49148 14272 49200 14278
rect 49148 14214 49200 14220
rect 49608 14272 49660 14278
rect 49608 14214 49660 14220
rect 49160 14074 49188 14214
rect 48320 14068 48372 14074
rect 48320 14010 48372 14016
rect 48964 14068 49016 14074
rect 48964 14010 49016 14016
rect 49148 14068 49200 14074
rect 49148 14010 49200 14016
rect 48228 13932 48280 13938
rect 48228 13874 48280 13880
rect 48240 13462 48268 13874
rect 48332 13530 48360 14010
rect 48412 13932 48464 13938
rect 48412 13874 48464 13880
rect 48320 13524 48372 13530
rect 48320 13466 48372 13472
rect 48228 13456 48280 13462
rect 48228 13398 48280 13404
rect 48056 13246 48176 13274
rect 48148 13190 48176 13246
rect 48044 13184 48096 13190
rect 48044 13126 48096 13132
rect 48136 13184 48188 13190
rect 48136 13126 48188 13132
rect 48056 12986 48084 13126
rect 48044 12980 48096 12986
rect 48044 12922 48096 12928
rect 48056 11286 48084 12922
rect 48044 11280 48096 11286
rect 48044 11222 48096 11228
rect 47860 11144 47912 11150
rect 47860 11086 47912 11092
rect 47872 10810 47900 11086
rect 48240 10810 48268 13398
rect 48424 13326 48452 13874
rect 48964 13388 49016 13394
rect 48964 13330 49016 13336
rect 48412 13320 48464 13326
rect 48412 13262 48464 13268
rect 48688 13320 48740 13326
rect 48688 13262 48740 13268
rect 48700 13190 48728 13262
rect 48688 13184 48740 13190
rect 48688 13126 48740 13132
rect 48780 13184 48832 13190
rect 48780 13126 48832 13132
rect 48410 12880 48466 12889
rect 48700 12850 48728 13126
rect 48410 12815 48466 12824
rect 48688 12844 48740 12850
rect 48320 12300 48372 12306
rect 48320 12242 48372 12248
rect 48332 11762 48360 12242
rect 48424 11898 48452 12815
rect 48688 12786 48740 12792
rect 48504 12708 48556 12714
rect 48504 12650 48556 12656
rect 48516 12102 48544 12650
rect 48504 12096 48556 12102
rect 48504 12038 48556 12044
rect 48792 11898 48820 13126
rect 48976 12322 49004 13330
rect 49424 13320 49476 13326
rect 49424 13262 49476 13268
rect 49240 13184 49292 13190
rect 49240 13126 49292 13132
rect 49252 12918 49280 13126
rect 49240 12912 49292 12918
rect 49240 12854 49292 12860
rect 49252 12374 49280 12854
rect 49436 12782 49464 13262
rect 49620 12986 49648 14214
rect 49804 13530 49832 14894
rect 50264 13870 50292 15438
rect 50344 15360 50396 15366
rect 50344 15302 50396 15308
rect 50356 14958 50384 15302
rect 50344 14952 50396 14958
rect 50344 14894 50396 14900
rect 50632 14414 50660 15846
rect 50712 15632 50764 15638
rect 50712 15574 50764 15580
rect 50528 14408 50580 14414
rect 50528 14350 50580 14356
rect 50620 14408 50672 14414
rect 50620 14350 50672 14356
rect 50540 13870 50568 14350
rect 50632 14278 50660 14350
rect 50620 14272 50672 14278
rect 50620 14214 50672 14220
rect 50252 13864 50304 13870
rect 50252 13806 50304 13812
rect 50528 13864 50580 13870
rect 50528 13806 50580 13812
rect 50264 13530 50292 13806
rect 49792 13524 49844 13530
rect 49792 13466 49844 13472
rect 50252 13524 50304 13530
rect 50252 13466 50304 13472
rect 50724 12986 50752 15574
rect 51000 15094 51028 15846
rect 51356 15428 51408 15434
rect 51356 15370 51408 15376
rect 51368 15162 51396 15370
rect 51356 15156 51408 15162
rect 51356 15098 51408 15104
rect 50988 15088 51040 15094
rect 50988 15030 51040 15036
rect 51368 14414 51396 15098
rect 51356 14408 51408 14414
rect 51356 14350 51408 14356
rect 51460 14074 51488 15982
rect 51644 15570 51672 16118
rect 52460 16040 52512 16046
rect 52460 15982 52512 15988
rect 52472 15706 52500 15982
rect 52644 15904 52696 15910
rect 52644 15846 52696 15852
rect 52460 15700 52512 15706
rect 52460 15642 52512 15648
rect 52656 15638 52684 15846
rect 52644 15632 52696 15638
rect 52644 15574 52696 15580
rect 51632 15564 51684 15570
rect 51632 15506 51684 15512
rect 51644 15026 51672 15506
rect 51724 15496 51776 15502
rect 51724 15438 51776 15444
rect 51736 15162 51764 15438
rect 52276 15360 52328 15366
rect 52276 15302 52328 15308
rect 51724 15156 51776 15162
rect 51724 15098 51776 15104
rect 51632 15020 51684 15026
rect 51632 14962 51684 14968
rect 52288 14958 52316 15302
rect 52368 15020 52420 15026
rect 52368 14962 52420 14968
rect 52276 14952 52328 14958
rect 52276 14894 52328 14900
rect 52288 14550 52316 14894
rect 52380 14550 52408 14962
rect 52840 14958 52868 17002
rect 53472 16992 53524 16998
rect 53472 16934 53524 16940
rect 53380 16652 53432 16658
rect 53380 16594 53432 16600
rect 53288 16448 53340 16454
rect 53288 16390 53340 16396
rect 52936 16348 53232 16368
rect 52992 16346 53016 16348
rect 53072 16346 53096 16348
rect 53152 16346 53176 16348
rect 53014 16294 53016 16346
rect 53078 16294 53090 16346
rect 53152 16294 53154 16346
rect 52992 16292 53016 16294
rect 53072 16292 53096 16294
rect 53152 16292 53176 16294
rect 52936 16272 53232 16292
rect 53300 15570 53328 16390
rect 53392 15910 53420 16594
rect 53380 15904 53432 15910
rect 53380 15846 53432 15852
rect 53288 15564 53340 15570
rect 53288 15506 53340 15512
rect 52936 15260 53232 15280
rect 52992 15258 53016 15260
rect 53072 15258 53096 15260
rect 53152 15258 53176 15260
rect 53014 15206 53016 15258
rect 53078 15206 53090 15258
rect 53152 15206 53154 15258
rect 52992 15204 53016 15206
rect 53072 15204 53096 15206
rect 53152 15204 53176 15206
rect 52936 15184 53232 15204
rect 53300 15162 53328 15506
rect 53288 15156 53340 15162
rect 53288 15098 53340 15104
rect 52828 14952 52880 14958
rect 52828 14894 52880 14900
rect 52736 14884 52788 14890
rect 52736 14826 52788 14832
rect 52748 14618 52776 14826
rect 52840 14618 52868 14894
rect 52736 14612 52788 14618
rect 52736 14554 52788 14560
rect 52828 14612 52880 14618
rect 52828 14554 52880 14560
rect 52276 14544 52328 14550
rect 52276 14486 52328 14492
rect 52368 14544 52420 14550
rect 52368 14486 52420 14492
rect 52288 14074 52316 14486
rect 52644 14476 52696 14482
rect 52644 14418 52696 14424
rect 51448 14068 51500 14074
rect 51448 14010 51500 14016
rect 52276 14068 52328 14074
rect 52276 14010 52328 14016
rect 52460 13932 52512 13938
rect 52460 13874 52512 13880
rect 52092 13864 52144 13870
rect 52092 13806 52144 13812
rect 52184 13864 52236 13870
rect 52184 13806 52236 13812
rect 52104 13734 52132 13806
rect 50988 13728 51040 13734
rect 50988 13670 51040 13676
rect 51080 13728 51132 13734
rect 51080 13670 51132 13676
rect 52092 13728 52144 13734
rect 52092 13670 52144 13676
rect 51000 13530 51028 13670
rect 50988 13524 51040 13530
rect 50988 13466 51040 13472
rect 51092 13394 51120 13670
rect 51080 13388 51132 13394
rect 51080 13330 51132 13336
rect 49608 12980 49660 12986
rect 49608 12922 49660 12928
rect 50712 12980 50764 12986
rect 50712 12922 50764 12928
rect 50252 12912 50304 12918
rect 50252 12854 50304 12860
rect 50526 12880 50582 12889
rect 49424 12776 49476 12782
rect 49424 12718 49476 12724
rect 50068 12708 50120 12714
rect 50068 12650 50120 12656
rect 48884 12306 49004 12322
rect 49240 12368 49292 12374
rect 49240 12310 49292 12316
rect 48872 12300 49004 12306
rect 48924 12294 49004 12300
rect 49056 12300 49108 12306
rect 48872 12242 48924 12248
rect 49056 12242 49108 12248
rect 48964 12232 49016 12238
rect 48964 12174 49016 12180
rect 48412 11892 48464 11898
rect 48412 11834 48464 11840
rect 48780 11892 48832 11898
rect 48780 11834 48832 11840
rect 48320 11756 48372 11762
rect 48320 11698 48372 11704
rect 48424 11694 48452 11834
rect 48412 11688 48464 11694
rect 48412 11630 48464 11636
rect 48792 11286 48820 11834
rect 48976 11626 49004 12174
rect 49068 12170 49096 12242
rect 49056 12164 49108 12170
rect 49056 12106 49108 12112
rect 49068 11898 49096 12106
rect 50080 12102 50108 12650
rect 50264 12646 50292 12854
rect 50526 12815 50528 12824
rect 50580 12815 50582 12824
rect 50528 12786 50580 12792
rect 50252 12640 50304 12646
rect 50252 12582 50304 12588
rect 50264 12374 50292 12582
rect 50252 12368 50304 12374
rect 50252 12310 50304 12316
rect 50710 12336 50766 12345
rect 50710 12271 50712 12280
rect 50764 12271 50766 12280
rect 50712 12242 50764 12248
rect 50252 12164 50304 12170
rect 50252 12106 50304 12112
rect 50068 12096 50120 12102
rect 50068 12038 50120 12044
rect 49056 11892 49108 11898
rect 49056 11834 49108 11840
rect 50264 11694 50292 12106
rect 51092 12102 51120 13330
rect 52104 13326 52132 13670
rect 52092 13320 52144 13326
rect 52092 13262 52144 13268
rect 51724 13184 51776 13190
rect 51724 13126 51776 13132
rect 51908 13184 51960 13190
rect 51908 13126 51960 13132
rect 51540 12708 51592 12714
rect 51540 12650 51592 12656
rect 51448 12300 51500 12306
rect 51448 12242 51500 12248
rect 51264 12232 51316 12238
rect 51264 12174 51316 12180
rect 50528 12096 50580 12102
rect 50528 12038 50580 12044
rect 50620 12096 50672 12102
rect 50620 12038 50672 12044
rect 51080 12096 51132 12102
rect 51080 12038 51132 12044
rect 50540 11898 50568 12038
rect 50528 11892 50580 11898
rect 50528 11834 50580 11840
rect 50632 11762 50660 12038
rect 50896 11824 50948 11830
rect 50896 11766 50948 11772
rect 50620 11756 50672 11762
rect 50620 11698 50672 11704
rect 50252 11688 50304 11694
rect 50252 11630 50304 11636
rect 48964 11620 49016 11626
rect 48964 11562 49016 11568
rect 49424 11620 49476 11626
rect 49424 11562 49476 11568
rect 48780 11280 48832 11286
rect 48780 11222 48832 11228
rect 49332 11212 49384 11218
rect 49332 11154 49384 11160
rect 48504 11144 48556 11150
rect 48504 11086 48556 11092
rect 47860 10804 47912 10810
rect 47860 10746 47912 10752
rect 48228 10804 48280 10810
rect 48228 10746 48280 10752
rect 47768 10260 47820 10266
rect 47872 10248 47900 10746
rect 47952 10736 48004 10742
rect 47952 10678 48004 10684
rect 48320 10736 48372 10742
rect 48320 10678 48372 10684
rect 47964 10470 47992 10678
rect 47952 10464 48004 10470
rect 47952 10406 48004 10412
rect 48332 10266 48360 10678
rect 48320 10260 48372 10266
rect 47872 10220 47992 10248
rect 47768 10202 47820 10208
rect 47584 10124 47636 10130
rect 47584 10066 47636 10072
rect 47768 10124 47820 10130
rect 47768 10066 47820 10072
rect 47860 10124 47912 10130
rect 47860 10066 47912 10072
rect 47490 9616 47546 9625
rect 47490 9551 47546 9560
rect 47490 9480 47546 9489
rect 47216 9444 47268 9450
rect 47490 9415 47546 9424
rect 47216 9386 47268 9392
rect 47032 8832 47084 8838
rect 47032 8774 47084 8780
rect 46848 8424 46900 8430
rect 46848 8366 46900 8372
rect 46860 8242 46888 8366
rect 46860 8214 46980 8242
rect 46952 7886 46980 8214
rect 47044 8090 47072 8774
rect 47228 8401 47256 9386
rect 47400 9036 47452 9042
rect 47320 8996 47400 9024
rect 47320 8566 47348 8996
rect 47400 8978 47452 8984
rect 47400 8832 47452 8838
rect 47400 8774 47452 8780
rect 47308 8560 47360 8566
rect 47308 8502 47360 8508
rect 47308 8424 47360 8430
rect 47214 8392 47270 8401
rect 47308 8366 47360 8372
rect 47214 8327 47270 8336
rect 47032 8084 47084 8090
rect 47032 8026 47084 8032
rect 46940 7880 46992 7886
rect 46940 7822 46992 7828
rect 46664 7744 46716 7750
rect 46664 7686 46716 7692
rect 46676 7562 46704 7686
rect 46492 7546 46704 7562
rect 46492 7540 46716 7546
rect 46492 7534 46664 7540
rect 46492 7478 46520 7534
rect 46664 7482 46716 7488
rect 46480 7472 46532 7478
rect 46480 7414 46532 7420
rect 46480 7336 46532 7342
rect 46664 7336 46716 7342
rect 46532 7296 46664 7324
rect 46480 7278 46532 7284
rect 46664 7278 46716 7284
rect 46952 7274 46980 7822
rect 46940 7268 46992 7274
rect 46940 7210 46992 7216
rect 46952 7002 46980 7210
rect 46940 6996 46992 7002
rect 46940 6938 46992 6944
rect 46938 6896 46994 6905
rect 46938 6831 46994 6840
rect 46388 6792 46440 6798
rect 46388 6734 46440 6740
rect 46664 6792 46716 6798
rect 46664 6734 46716 6740
rect 46204 6452 46256 6458
rect 46204 6394 46256 6400
rect 46112 6248 46164 6254
rect 46112 6190 46164 6196
rect 45008 5772 45060 5778
rect 45008 5714 45060 5720
rect 45100 5772 45152 5778
rect 45100 5714 45152 5720
rect 45020 5370 45048 5714
rect 46124 5574 46152 6190
rect 46112 5568 46164 5574
rect 46112 5510 46164 5516
rect 46216 5522 46244 6394
rect 46296 6248 46348 6254
rect 46296 6190 46348 6196
rect 46308 5846 46336 6190
rect 46296 5840 46348 5846
rect 46296 5782 46348 5788
rect 46294 5536 46350 5545
rect 45008 5364 45060 5370
rect 45008 5306 45060 5312
rect 46124 5302 46152 5510
rect 46216 5494 46294 5522
rect 46294 5471 46350 5480
rect 46308 5302 46336 5471
rect 46112 5296 46164 5302
rect 46112 5238 46164 5244
rect 46296 5296 46348 5302
rect 46296 5238 46348 5244
rect 45008 5160 45060 5166
rect 45008 5102 45060 5108
rect 45020 3126 45048 5102
rect 46124 4690 46152 5238
rect 46112 4684 46164 4690
rect 46112 4626 46164 4632
rect 46296 4684 46348 4690
rect 46296 4626 46348 4632
rect 45652 4616 45704 4622
rect 45652 4558 45704 4564
rect 45560 4480 45612 4486
rect 45560 4422 45612 4428
rect 45100 4004 45152 4010
rect 45100 3946 45152 3952
rect 45112 3466 45140 3946
rect 45572 3602 45600 4422
rect 45664 4185 45692 4558
rect 45650 4176 45706 4185
rect 45650 4111 45652 4120
rect 45704 4111 45706 4120
rect 45652 4082 45704 4088
rect 45664 4051 45692 4082
rect 46308 4010 46336 4626
rect 46296 4004 46348 4010
rect 46296 3946 46348 3952
rect 46020 3936 46072 3942
rect 46020 3878 46072 3884
rect 46204 3936 46256 3942
rect 46204 3878 46256 3884
rect 45192 3596 45244 3602
rect 45192 3538 45244 3544
rect 45560 3596 45612 3602
rect 45560 3538 45612 3544
rect 45100 3460 45152 3466
rect 45100 3402 45152 3408
rect 45008 3120 45060 3126
rect 44914 3088 44970 3097
rect 45112 3097 45140 3402
rect 45008 3062 45060 3068
rect 45098 3088 45154 3097
rect 44914 3023 44970 3032
rect 45098 3023 45154 3032
rect 45008 2984 45060 2990
rect 45112 2972 45140 3023
rect 45204 2990 45232 3538
rect 45468 3528 45520 3534
rect 45468 3470 45520 3476
rect 45060 2944 45140 2972
rect 45192 2984 45244 2990
rect 45008 2926 45060 2932
rect 45192 2926 45244 2932
rect 45376 2916 45428 2922
rect 45376 2858 45428 2864
rect 44822 2816 44878 2825
rect 44822 2751 44878 2760
rect 45388 2666 45416 2858
rect 44652 2638 45416 2666
rect 44272 2440 44324 2446
rect 44272 2382 44324 2388
rect 44284 1970 44312 2382
rect 44272 1964 44324 1970
rect 44272 1906 44324 1912
rect 43640 1414 43760 1442
rect 43732 800 43760 1414
rect 44652 800 44680 2638
rect 45480 2553 45508 3470
rect 46032 2922 46060 3878
rect 46216 3738 46244 3878
rect 46308 3738 46336 3946
rect 46204 3732 46256 3738
rect 46204 3674 46256 3680
rect 46296 3732 46348 3738
rect 46296 3674 46348 3680
rect 46204 3596 46256 3602
rect 46204 3538 46256 3544
rect 46110 3496 46166 3505
rect 46110 3431 46166 3440
rect 46124 3194 46152 3431
rect 46112 3188 46164 3194
rect 46112 3130 46164 3136
rect 46124 2990 46152 3130
rect 46112 2984 46164 2990
rect 46112 2926 46164 2932
rect 46020 2916 46072 2922
rect 46020 2858 46072 2864
rect 45560 2848 45612 2854
rect 45560 2790 45612 2796
rect 45466 2544 45522 2553
rect 45466 2479 45522 2488
rect 45572 800 45600 2790
rect 46216 2650 46244 3538
rect 46400 3466 46428 6734
rect 46676 6118 46704 6734
rect 46952 6730 46980 6831
rect 46940 6724 46992 6730
rect 46940 6666 46992 6672
rect 47044 6497 47072 8026
rect 47228 7206 47256 8327
rect 47320 8090 47348 8366
rect 47308 8084 47360 8090
rect 47308 8026 47360 8032
rect 47412 7954 47440 8774
rect 47504 8430 47532 9415
rect 47780 9382 47808 10066
rect 47872 9654 47900 10066
rect 47860 9648 47912 9654
rect 47860 9590 47912 9596
rect 47768 9376 47820 9382
rect 47768 9318 47820 9324
rect 47768 8968 47820 8974
rect 47768 8910 47820 8916
rect 47780 8430 47808 8910
rect 47492 8424 47544 8430
rect 47492 8366 47544 8372
rect 47768 8424 47820 8430
rect 47768 8366 47820 8372
rect 47674 8120 47730 8129
rect 47674 8055 47730 8064
rect 47688 7954 47716 8055
rect 47400 7948 47452 7954
rect 47400 7890 47452 7896
rect 47676 7948 47728 7954
rect 47676 7890 47728 7896
rect 47306 7712 47362 7721
rect 47306 7647 47362 7656
rect 47216 7200 47268 7206
rect 47216 7142 47268 7148
rect 47216 6792 47268 6798
rect 47216 6734 47268 6740
rect 47030 6488 47086 6497
rect 47030 6423 47086 6432
rect 46756 6180 46808 6186
rect 46756 6122 46808 6128
rect 46848 6180 46900 6186
rect 46848 6122 46900 6128
rect 46664 6112 46716 6118
rect 46664 6054 46716 6060
rect 46664 5772 46716 5778
rect 46664 5714 46716 5720
rect 46676 5574 46704 5714
rect 46768 5710 46796 6122
rect 46756 5704 46808 5710
rect 46756 5646 46808 5652
rect 46664 5568 46716 5574
rect 46664 5510 46716 5516
rect 46572 5024 46624 5030
rect 46572 4966 46624 4972
rect 46584 4826 46612 4966
rect 46572 4820 46624 4826
rect 46572 4762 46624 4768
rect 46676 4729 46704 5510
rect 46662 4720 46718 4729
rect 46662 4655 46718 4664
rect 46756 4276 46808 4282
rect 46756 4218 46808 4224
rect 46768 3602 46796 4218
rect 46756 3596 46808 3602
rect 46756 3538 46808 3544
rect 46860 3466 46888 6122
rect 47044 4282 47072 6423
rect 47124 5296 47176 5302
rect 47124 5238 47176 5244
rect 47136 4758 47164 5238
rect 47228 4826 47256 6734
rect 47320 6458 47348 7647
rect 47412 6934 47440 7890
rect 47492 7812 47544 7818
rect 47676 7812 47728 7818
rect 47544 7772 47676 7800
rect 47492 7754 47544 7760
rect 47676 7754 47728 7760
rect 47504 7546 47532 7754
rect 47492 7540 47544 7546
rect 47492 7482 47544 7488
rect 47676 7540 47728 7546
rect 47676 7482 47728 7488
rect 47688 7274 47716 7482
rect 47676 7268 47728 7274
rect 47676 7210 47728 7216
rect 47780 7154 47808 8366
rect 47964 7936 47992 10220
rect 48320 10202 48372 10208
rect 48332 9586 48360 10202
rect 48412 9920 48464 9926
rect 48516 9908 48544 11086
rect 48872 11076 48924 11082
rect 48872 11018 48924 11024
rect 48780 11008 48832 11014
rect 48780 10950 48832 10956
rect 48792 10606 48820 10950
rect 48884 10606 48912 11018
rect 49344 10674 49372 11154
rect 49332 10668 49384 10674
rect 49332 10610 49384 10616
rect 48596 10600 48648 10606
rect 48596 10542 48648 10548
rect 48780 10600 48832 10606
rect 48780 10542 48832 10548
rect 48872 10600 48924 10606
rect 48872 10542 48924 10548
rect 48464 9880 48544 9908
rect 48608 9908 48636 10542
rect 48686 10432 48742 10441
rect 48686 10367 48742 10376
rect 48700 10130 48728 10367
rect 48688 10124 48740 10130
rect 48688 10066 48740 10072
rect 48688 9920 48740 9926
rect 48608 9880 48688 9908
rect 48412 9862 48464 9868
rect 48688 9862 48740 9868
rect 48320 9580 48372 9586
rect 48320 9522 48372 9528
rect 48044 9376 48096 9382
rect 48044 9318 48096 9324
rect 48056 8362 48084 9318
rect 48044 8356 48096 8362
rect 48044 8298 48096 8304
rect 48226 8120 48282 8129
rect 48226 8055 48282 8064
rect 47964 7908 48084 7936
rect 47952 7812 48004 7818
rect 47952 7754 48004 7760
rect 47964 7274 47992 7754
rect 47952 7268 48004 7274
rect 47952 7210 48004 7216
rect 47688 7126 47808 7154
rect 47400 6928 47452 6934
rect 47400 6870 47452 6876
rect 47400 6792 47452 6798
rect 47400 6734 47452 6740
rect 47308 6452 47360 6458
rect 47308 6394 47360 6400
rect 47412 6254 47440 6734
rect 47492 6656 47544 6662
rect 47492 6598 47544 6604
rect 47400 6248 47452 6254
rect 47400 6190 47452 6196
rect 47216 4820 47268 4826
rect 47216 4762 47268 4768
rect 47124 4752 47176 4758
rect 47124 4694 47176 4700
rect 47032 4276 47084 4282
rect 47032 4218 47084 4224
rect 46940 4072 46992 4078
rect 46940 4014 46992 4020
rect 47032 4072 47084 4078
rect 47032 4014 47084 4020
rect 46952 3670 46980 4014
rect 46940 3664 46992 3670
rect 47044 3641 47072 4014
rect 47228 3670 47256 4762
rect 47504 4758 47532 6598
rect 47492 4752 47544 4758
rect 47492 4694 47544 4700
rect 47584 4684 47636 4690
rect 47584 4626 47636 4632
rect 47492 3936 47544 3942
rect 47320 3896 47492 3924
rect 47216 3664 47268 3670
rect 46940 3606 46992 3612
rect 47030 3632 47086 3641
rect 47216 3606 47268 3612
rect 47030 3567 47086 3576
rect 46388 3460 46440 3466
rect 46388 3402 46440 3408
rect 46848 3460 46900 3466
rect 46848 3402 46900 3408
rect 47320 3398 47348 3896
rect 47492 3878 47544 3884
rect 47400 3664 47452 3670
rect 47596 3652 47624 4626
rect 47452 3624 47624 3652
rect 47400 3606 47452 3612
rect 47308 3392 47360 3398
rect 47308 3334 47360 3340
rect 46296 3120 46348 3126
rect 47032 3120 47084 3126
rect 46296 3062 46348 3068
rect 47030 3088 47032 3097
rect 47084 3088 47086 3097
rect 46308 2990 46336 3062
rect 47030 3023 47086 3032
rect 47044 2990 47072 3023
rect 46296 2984 46348 2990
rect 46296 2926 46348 2932
rect 47032 2984 47084 2990
rect 47032 2926 47084 2932
rect 46940 2848 46992 2854
rect 46386 2816 46442 2825
rect 46940 2790 46992 2796
rect 46386 2751 46442 2760
rect 46204 2644 46256 2650
rect 46204 2586 46256 2592
rect 46400 800 46428 2751
rect 46952 2650 46980 2790
rect 46940 2644 46992 2650
rect 46940 2586 46992 2592
rect 47596 2582 47624 3624
rect 47688 3369 47716 7126
rect 47952 6656 48004 6662
rect 47952 6598 48004 6604
rect 47964 6458 47992 6598
rect 47952 6452 48004 6458
rect 47952 6394 48004 6400
rect 47964 6254 47992 6394
rect 47952 6248 48004 6254
rect 47952 6190 48004 6196
rect 48056 5896 48084 7908
rect 48136 7880 48188 7886
rect 48136 7822 48188 7828
rect 48148 7313 48176 7822
rect 48240 7750 48268 8055
rect 48424 7818 48452 9862
rect 48700 9110 48728 9862
rect 48792 9382 48820 10542
rect 49344 10130 49372 10610
rect 49436 10606 49464 11562
rect 50908 11286 50936 11766
rect 51276 11354 51304 12174
rect 51264 11348 51316 11354
rect 51264 11290 51316 11296
rect 50896 11280 50948 11286
rect 50896 11222 50948 11228
rect 51460 11150 51488 12242
rect 50344 11144 50396 11150
rect 50344 11086 50396 11092
rect 51448 11144 51500 11150
rect 51448 11086 51500 11092
rect 50356 10674 50384 11086
rect 51356 11076 51408 11082
rect 51356 11018 51408 11024
rect 51080 11008 51132 11014
rect 51080 10950 51132 10956
rect 50344 10668 50396 10674
rect 50344 10610 50396 10616
rect 49424 10600 49476 10606
rect 49424 10542 49476 10548
rect 49514 10568 49570 10577
rect 49332 10124 49384 10130
rect 49332 10066 49384 10072
rect 49240 9580 49292 9586
rect 49240 9522 49292 9528
rect 48780 9376 48832 9382
rect 48780 9318 48832 9324
rect 48688 9104 48740 9110
rect 48688 9046 48740 9052
rect 48504 8560 48556 8566
rect 48556 8520 48912 8548
rect 48504 8502 48556 8508
rect 48884 8430 48912 8520
rect 48504 8424 48556 8430
rect 48502 8392 48504 8401
rect 48872 8424 48924 8430
rect 48556 8392 48558 8401
rect 48872 8366 48924 8372
rect 49252 8362 49280 9522
rect 49344 9178 49372 10066
rect 49436 9908 49464 10542
rect 49514 10503 49570 10512
rect 49608 10532 49660 10538
rect 49528 10470 49556 10503
rect 49608 10474 49660 10480
rect 49516 10464 49568 10470
rect 49516 10406 49568 10412
rect 49620 10266 49648 10474
rect 49608 10260 49660 10266
rect 49608 10202 49660 10208
rect 49608 9920 49660 9926
rect 49436 9880 49608 9908
rect 49608 9862 49660 9868
rect 50252 9920 50304 9926
rect 50252 9862 50304 9868
rect 49620 9722 49648 9862
rect 49608 9716 49660 9722
rect 49608 9658 49660 9664
rect 50264 9518 50292 9862
rect 49700 9512 49752 9518
rect 50252 9512 50304 9518
rect 49700 9454 49752 9460
rect 50250 9480 50252 9489
rect 50304 9480 50306 9489
rect 49332 9172 49384 9178
rect 49332 9114 49384 9120
rect 49514 8392 49570 8401
rect 48502 8327 48558 8336
rect 49240 8356 49292 8362
rect 49514 8327 49570 8336
rect 49240 8298 49292 8304
rect 49146 7984 49202 7993
rect 48780 7948 48832 7954
rect 49146 7919 49148 7928
rect 48780 7890 48832 7896
rect 49200 7919 49202 7928
rect 49148 7890 49200 7896
rect 48412 7812 48464 7818
rect 48412 7754 48464 7760
rect 48596 7812 48648 7818
rect 48596 7754 48648 7760
rect 48228 7744 48280 7750
rect 48228 7686 48280 7692
rect 48134 7304 48190 7313
rect 48134 7239 48136 7248
rect 48188 7239 48190 7248
rect 48136 7210 48188 7216
rect 48148 7179 48176 7210
rect 48240 5914 48268 7686
rect 48504 7268 48556 7274
rect 48504 7210 48556 7216
rect 48410 6896 48466 6905
rect 48410 6831 48412 6840
rect 48464 6831 48466 6840
rect 48412 6802 48464 6808
rect 48516 6458 48544 7210
rect 48608 7206 48636 7754
rect 48688 7404 48740 7410
rect 48688 7346 48740 7352
rect 48596 7200 48648 7206
rect 48596 7142 48648 7148
rect 48608 7002 48636 7142
rect 48596 6996 48648 7002
rect 48596 6938 48648 6944
rect 48608 6866 48636 6938
rect 48596 6860 48648 6866
rect 48596 6802 48648 6808
rect 48504 6452 48556 6458
rect 48504 6394 48556 6400
rect 48516 6322 48544 6394
rect 48504 6316 48556 6322
rect 48504 6258 48556 6264
rect 48228 5908 48280 5914
rect 48056 5868 48176 5896
rect 48044 5772 48096 5778
rect 48044 5714 48096 5720
rect 47768 5568 47820 5574
rect 47768 5510 47820 5516
rect 47952 5568 48004 5574
rect 47952 5510 48004 5516
rect 47780 3584 47808 5510
rect 47860 5160 47912 5166
rect 47860 5102 47912 5108
rect 47872 4622 47900 5102
rect 47964 5098 47992 5510
rect 47952 5092 48004 5098
rect 47952 5034 48004 5040
rect 47860 4616 47912 4622
rect 47860 4558 47912 4564
rect 47964 4282 47992 5034
rect 48056 5030 48084 5714
rect 48148 5352 48176 5868
rect 48228 5850 48280 5856
rect 48240 5778 48268 5850
rect 48228 5772 48280 5778
rect 48228 5714 48280 5720
rect 48700 5642 48728 7346
rect 48792 7274 48820 7890
rect 49160 7274 49188 7890
rect 48780 7268 48832 7274
rect 48780 7210 48832 7216
rect 49148 7268 49200 7274
rect 49148 7210 49200 7216
rect 48792 6225 48820 7210
rect 49054 6624 49110 6633
rect 49054 6559 49110 6568
rect 48778 6216 48834 6225
rect 48778 6151 48834 6160
rect 48688 5636 48740 5642
rect 48688 5578 48740 5584
rect 48412 5568 48464 5574
rect 48412 5510 48464 5516
rect 48148 5324 48268 5352
rect 48136 5228 48188 5234
rect 48136 5170 48188 5176
rect 48044 5024 48096 5030
rect 48044 4966 48096 4972
rect 47952 4276 48004 4282
rect 47952 4218 48004 4224
rect 47950 4176 48006 4185
rect 47950 4111 47952 4120
rect 48004 4111 48006 4120
rect 47952 4082 48004 4088
rect 48056 3738 48084 4966
rect 48148 4826 48176 5170
rect 48136 4820 48188 4826
rect 48136 4762 48188 4768
rect 48136 4684 48188 4690
rect 48136 4626 48188 4632
rect 48148 4486 48176 4626
rect 48136 4480 48188 4486
rect 48136 4422 48188 4428
rect 48044 3732 48096 3738
rect 48044 3674 48096 3680
rect 47860 3596 47912 3602
rect 47780 3556 47860 3584
rect 47860 3538 47912 3544
rect 47674 3360 47730 3369
rect 47674 3295 47730 3304
rect 48240 2990 48268 5324
rect 48424 4078 48452 5510
rect 48688 4480 48740 4486
rect 48502 4448 48558 4457
rect 48688 4422 48740 4428
rect 48502 4383 48558 4392
rect 48516 4078 48544 4383
rect 48700 4078 48728 4422
rect 48412 4072 48464 4078
rect 48412 4014 48464 4020
rect 48504 4072 48556 4078
rect 48688 4072 48740 4078
rect 48504 4014 48556 4020
rect 48608 4032 48688 4060
rect 48320 3936 48372 3942
rect 48372 3896 48452 3924
rect 48320 3878 48372 3884
rect 48424 3890 48452 3896
rect 48516 3890 48544 4014
rect 48424 3862 48544 3890
rect 48608 3194 48636 4032
rect 48688 4014 48740 4020
rect 48688 3392 48740 3398
rect 48792 3380 48820 6151
rect 49068 6118 49096 6559
rect 49056 6112 49108 6118
rect 49056 6054 49108 6060
rect 48872 5364 48924 5370
rect 48872 5306 48924 5312
rect 48884 4622 48912 5306
rect 48964 4752 49016 4758
rect 48964 4694 49016 4700
rect 48872 4616 48924 4622
rect 48872 4558 48924 4564
rect 48884 3942 48912 4558
rect 48872 3936 48924 3942
rect 48872 3878 48924 3884
rect 48976 3738 49004 4694
rect 49068 3738 49096 6054
rect 49148 5908 49200 5914
rect 49148 5850 49200 5856
rect 49160 5817 49188 5850
rect 49146 5808 49202 5817
rect 49146 5743 49202 5752
rect 49160 5710 49188 5743
rect 49148 5704 49200 5710
rect 49148 5646 49200 5652
rect 49148 4480 49200 4486
rect 49148 4422 49200 4428
rect 49160 4214 49188 4422
rect 49148 4208 49200 4214
rect 49148 4150 49200 4156
rect 49252 4146 49280 8298
rect 49528 8294 49556 8327
rect 49516 8288 49568 8294
rect 49516 8230 49568 8236
rect 49332 5636 49384 5642
rect 49332 5578 49384 5584
rect 49344 5166 49372 5578
rect 49528 5234 49556 8230
rect 49608 7744 49660 7750
rect 49608 7686 49660 7692
rect 49620 7410 49648 7686
rect 49608 7404 49660 7410
rect 49608 7346 49660 7352
rect 49712 6866 49740 9454
rect 50068 9444 50120 9450
rect 50356 9450 50384 10610
rect 50986 10568 51042 10577
rect 50986 10503 51042 10512
rect 50436 10260 50488 10266
rect 50436 10202 50488 10208
rect 50448 9738 50476 10202
rect 50448 9710 50752 9738
rect 50448 9654 50476 9710
rect 50436 9648 50488 9654
rect 50436 9590 50488 9596
rect 50528 9512 50580 9518
rect 50528 9454 50580 9460
rect 50250 9415 50306 9424
rect 50344 9444 50396 9450
rect 50068 9386 50120 9392
rect 50344 9386 50396 9392
rect 49976 9172 50028 9178
rect 49976 9114 50028 9120
rect 49792 8968 49844 8974
rect 49792 8910 49844 8916
rect 49804 7993 49832 8910
rect 49988 8906 50016 9114
rect 50080 8922 50108 9386
rect 50540 9110 50568 9454
rect 50528 9104 50580 9110
rect 50528 9046 50580 9052
rect 49976 8900 50028 8906
rect 50080 8894 50292 8922
rect 49976 8842 50028 8848
rect 49988 8480 50016 8842
rect 50068 8832 50120 8838
rect 50120 8792 50200 8820
rect 50068 8774 50120 8780
rect 50172 8498 50200 8792
rect 50264 8566 50292 8894
rect 50252 8560 50304 8566
rect 50252 8502 50304 8508
rect 50068 8492 50120 8498
rect 49988 8452 50068 8480
rect 50068 8434 50120 8440
rect 50160 8492 50212 8498
rect 50160 8434 50212 8440
rect 50264 8362 50292 8502
rect 50620 8492 50672 8498
rect 50620 8434 50672 8440
rect 50632 8362 50660 8434
rect 50252 8356 50304 8362
rect 50252 8298 50304 8304
rect 50620 8356 50672 8362
rect 50620 8298 50672 8304
rect 49884 8288 49936 8294
rect 49884 8230 49936 8236
rect 49790 7984 49846 7993
rect 49790 7919 49846 7928
rect 49896 7886 49924 8230
rect 50344 8084 50396 8090
rect 50344 8026 50396 8032
rect 49792 7880 49844 7886
rect 49792 7822 49844 7828
rect 49884 7880 49936 7886
rect 49884 7822 49936 7828
rect 50252 7880 50304 7886
rect 50252 7822 50304 7828
rect 49700 6860 49752 6866
rect 49700 6802 49752 6808
rect 49608 6656 49660 6662
rect 49660 6604 49740 6610
rect 49608 6598 49740 6604
rect 49620 6582 49740 6598
rect 49712 6118 49740 6582
rect 49700 6112 49752 6118
rect 49700 6054 49752 6060
rect 49700 5772 49752 5778
rect 49700 5714 49752 5720
rect 49516 5228 49568 5234
rect 49516 5170 49568 5176
rect 49332 5160 49384 5166
rect 49332 5102 49384 5108
rect 49528 5030 49556 5170
rect 49712 5166 49740 5714
rect 49700 5160 49752 5166
rect 49700 5102 49752 5108
rect 49516 5024 49568 5030
rect 49516 4966 49568 4972
rect 49240 4140 49292 4146
rect 49240 4082 49292 4088
rect 48964 3732 49016 3738
rect 48964 3674 49016 3680
rect 49056 3732 49108 3738
rect 49056 3674 49108 3680
rect 48872 3596 48924 3602
rect 48872 3538 48924 3544
rect 48884 3505 48912 3538
rect 48870 3496 48926 3505
rect 48870 3431 48926 3440
rect 48740 3352 48820 3380
rect 48688 3334 48740 3340
rect 48596 3188 48648 3194
rect 48596 3130 48648 3136
rect 49068 3126 49096 3674
rect 49332 3392 49384 3398
rect 49332 3334 49384 3340
rect 49056 3120 49108 3126
rect 49056 3062 49108 3068
rect 49344 2990 49372 3334
rect 49528 3233 49556 4966
rect 49804 4826 49832 7822
rect 50160 7404 50212 7410
rect 50160 7346 50212 7352
rect 50068 7336 50120 7342
rect 50068 7278 50120 7284
rect 49884 7268 49936 7274
rect 49884 7210 49936 7216
rect 49896 6866 49924 7210
rect 49884 6860 49936 6866
rect 49884 6802 49936 6808
rect 49976 6248 50028 6254
rect 49976 6190 50028 6196
rect 49988 5914 50016 6190
rect 50080 6118 50108 7278
rect 50068 6112 50120 6118
rect 50068 6054 50120 6060
rect 49976 5908 50028 5914
rect 49976 5850 50028 5856
rect 50080 4826 50108 6054
rect 50172 5574 50200 7346
rect 50264 5778 50292 7822
rect 50356 7342 50384 8026
rect 50632 7750 50660 8298
rect 50724 8294 50752 9710
rect 50896 9376 50948 9382
rect 50896 9318 50948 9324
rect 50908 9042 50936 9318
rect 50896 9036 50948 9042
rect 50896 8978 50948 8984
rect 50908 8498 50936 8978
rect 50896 8492 50948 8498
rect 50896 8434 50948 8440
rect 50804 8356 50856 8362
rect 50804 8298 50856 8304
rect 50712 8288 50764 8294
rect 50712 8230 50764 8236
rect 50724 7886 50752 8230
rect 50712 7880 50764 7886
rect 50712 7822 50764 7828
rect 50620 7744 50672 7750
rect 50724 7721 50752 7822
rect 50620 7686 50672 7692
rect 50710 7712 50766 7721
rect 50344 7336 50396 7342
rect 50344 7278 50396 7284
rect 50344 6860 50396 6866
rect 50344 6802 50396 6808
rect 50356 6458 50384 6802
rect 50434 6488 50490 6497
rect 50344 6452 50396 6458
rect 50434 6423 50490 6432
rect 50344 6394 50396 6400
rect 50448 6254 50476 6423
rect 50632 6390 50660 7686
rect 50710 7647 50766 7656
rect 50712 7200 50764 7206
rect 50712 7142 50764 7148
rect 50724 6866 50752 7142
rect 50712 6860 50764 6866
rect 50712 6802 50764 6808
rect 50816 6497 50844 8298
rect 51000 7426 51028 10503
rect 51092 10266 51120 10950
rect 51368 10742 51396 11018
rect 51460 10810 51488 11086
rect 51448 10804 51500 10810
rect 51448 10746 51500 10752
rect 51356 10736 51408 10742
rect 51356 10678 51408 10684
rect 51172 10464 51224 10470
rect 51172 10406 51224 10412
rect 51080 10260 51132 10266
rect 51080 10202 51132 10208
rect 51184 9194 51212 10406
rect 51552 10198 51580 12650
rect 51632 12640 51684 12646
rect 51632 12582 51684 12588
rect 51644 12170 51672 12582
rect 51736 12238 51764 13126
rect 51920 12782 51948 13126
rect 51908 12776 51960 12782
rect 51908 12718 51960 12724
rect 51724 12232 51776 12238
rect 51724 12174 51776 12180
rect 51632 12164 51684 12170
rect 51632 12106 51684 12112
rect 51736 11898 51764 12174
rect 51908 12164 51960 12170
rect 51908 12106 51960 12112
rect 51920 11898 51948 12106
rect 51724 11892 51776 11898
rect 51724 11834 51776 11840
rect 51908 11892 51960 11898
rect 51908 11834 51960 11840
rect 51632 11280 51684 11286
rect 51632 11222 51684 11228
rect 51540 10192 51592 10198
rect 51540 10134 51592 10140
rect 51264 10124 51316 10130
rect 51264 10066 51316 10072
rect 51276 9654 51304 10066
rect 51644 10062 51672 11222
rect 51724 11008 51776 11014
rect 51724 10950 51776 10956
rect 51736 10606 51764 10950
rect 51920 10742 51948 11834
rect 52000 11824 52052 11830
rect 52000 11766 52052 11772
rect 52012 11694 52040 11766
rect 52000 11688 52052 11694
rect 52000 11630 52052 11636
rect 51908 10736 51960 10742
rect 51908 10678 51960 10684
rect 51816 10668 51868 10674
rect 51816 10610 51868 10616
rect 51724 10600 51776 10606
rect 51722 10568 51724 10577
rect 51776 10568 51778 10577
rect 51722 10503 51778 10512
rect 51828 10418 51856 10610
rect 51736 10390 51856 10418
rect 51540 10056 51592 10062
rect 51540 9998 51592 10004
rect 51632 10056 51684 10062
rect 51632 9998 51684 10004
rect 51264 9648 51316 9654
rect 51264 9590 51316 9596
rect 51448 9376 51500 9382
rect 51448 9318 51500 9324
rect 51184 9166 51304 9194
rect 51172 9104 51224 9110
rect 51172 9046 51224 9052
rect 51184 8430 51212 9046
rect 51276 8945 51304 9166
rect 51460 9042 51488 9318
rect 51356 9036 51408 9042
rect 51356 8978 51408 8984
rect 51448 9036 51500 9042
rect 51448 8978 51500 8984
rect 51262 8936 51318 8945
rect 51262 8871 51318 8880
rect 51276 8498 51304 8871
rect 51264 8492 51316 8498
rect 51264 8434 51316 8440
rect 51172 8424 51224 8430
rect 51172 8366 51224 8372
rect 51080 8356 51132 8362
rect 51080 8298 51132 8304
rect 51092 8090 51120 8298
rect 51080 8084 51132 8090
rect 51080 8026 51132 8032
rect 51184 7750 51212 8366
rect 51368 8090 51396 8978
rect 51552 8838 51580 9998
rect 51736 9518 51764 10390
rect 52000 10260 52052 10266
rect 52000 10202 52052 10208
rect 51816 9920 51868 9926
rect 51816 9862 51868 9868
rect 51828 9518 51856 9862
rect 51724 9512 51776 9518
rect 51722 9480 51724 9489
rect 51816 9512 51868 9518
rect 51776 9480 51778 9489
rect 51816 9454 51868 9460
rect 51722 9415 51778 9424
rect 51828 8906 51856 9454
rect 51816 8900 51868 8906
rect 51816 8842 51868 8848
rect 51540 8832 51592 8838
rect 51540 8774 51592 8780
rect 51724 8832 51776 8838
rect 51724 8774 51776 8780
rect 51356 8084 51408 8090
rect 51356 8026 51408 8032
rect 51172 7744 51224 7750
rect 51172 7686 51224 7692
rect 51000 7398 51120 7426
rect 50988 7336 51040 7342
rect 50988 7278 51040 7284
rect 51000 7018 51028 7278
rect 50908 7002 51028 7018
rect 50908 6996 51040 7002
rect 50908 6990 50988 6996
rect 50802 6488 50858 6497
rect 50802 6423 50858 6432
rect 50620 6384 50672 6390
rect 50620 6326 50672 6332
rect 50436 6248 50488 6254
rect 50908 6202 50936 6990
rect 50988 6938 51040 6944
rect 50988 6860 51040 6866
rect 50988 6802 51040 6808
rect 50436 6190 50488 6196
rect 50816 6174 50936 6202
rect 50816 6118 50844 6174
rect 50804 6112 50856 6118
rect 50804 6054 50856 6060
rect 50896 6112 50948 6118
rect 50896 6054 50948 6060
rect 50908 5778 50936 6054
rect 50252 5772 50304 5778
rect 50252 5714 50304 5720
rect 50436 5772 50488 5778
rect 50436 5714 50488 5720
rect 50896 5772 50948 5778
rect 50896 5714 50948 5720
rect 50252 5636 50304 5642
rect 50252 5578 50304 5584
rect 50160 5568 50212 5574
rect 50160 5510 50212 5516
rect 50264 5370 50292 5578
rect 50344 5568 50396 5574
rect 50344 5510 50396 5516
rect 50252 5364 50304 5370
rect 50252 5306 50304 5312
rect 49792 4820 49844 4826
rect 49792 4762 49844 4768
rect 50068 4820 50120 4826
rect 50068 4762 50120 4768
rect 49608 4752 49660 4758
rect 49606 4720 49608 4729
rect 49660 4720 49662 4729
rect 50080 4706 50108 4762
rect 50356 4758 50384 5510
rect 50448 5370 50476 5714
rect 50436 5364 50488 5370
rect 50436 5306 50488 5312
rect 50620 5228 50672 5234
rect 50620 5170 50672 5176
rect 49712 4690 50108 4706
rect 50344 4752 50396 4758
rect 50344 4694 50396 4700
rect 49606 4655 49662 4664
rect 49700 4684 50108 4690
rect 49752 4678 50108 4684
rect 49700 4626 49752 4632
rect 50632 4622 50660 5170
rect 50908 5166 50936 5714
rect 51000 5642 51028 6802
rect 50988 5636 51040 5642
rect 50988 5578 51040 5584
rect 50896 5160 50948 5166
rect 50894 5128 50896 5137
rect 50948 5128 50950 5137
rect 50894 5063 50950 5072
rect 50896 4820 50948 4826
rect 50896 4762 50948 4768
rect 50620 4616 50672 4622
rect 50620 4558 50672 4564
rect 50620 4140 50672 4146
rect 50620 4082 50672 4088
rect 49792 4072 49844 4078
rect 49792 4014 49844 4020
rect 49882 4040 49938 4049
rect 49514 3224 49570 3233
rect 49514 3159 49570 3168
rect 48228 2984 48280 2990
rect 48228 2926 48280 2932
rect 49332 2984 49384 2990
rect 49332 2926 49384 2932
rect 48136 2916 48188 2922
rect 48136 2858 48188 2864
rect 48148 2650 48176 2858
rect 48320 2848 48372 2854
rect 48320 2790 48372 2796
rect 48136 2644 48188 2650
rect 48136 2586 48188 2592
rect 47584 2576 47636 2582
rect 47584 2518 47636 2524
rect 48332 2446 48360 2790
rect 49056 2508 49108 2514
rect 49056 2450 49108 2456
rect 48320 2440 48372 2446
rect 48320 2382 48372 2388
rect 47308 2372 47360 2378
rect 47308 2314 47360 2320
rect 47320 800 47348 2314
rect 48228 2304 48280 2310
rect 48228 2246 48280 2252
rect 48240 2106 48268 2246
rect 48228 2100 48280 2106
rect 48228 2042 48280 2048
rect 48332 1714 48360 2382
rect 48240 1686 48360 1714
rect 48240 800 48268 1686
rect 49068 800 49096 2450
rect 49344 2446 49372 2926
rect 49804 2582 49832 4014
rect 49882 3975 49938 3984
rect 49896 3738 49924 3975
rect 50068 3936 50120 3942
rect 50068 3878 50120 3884
rect 50252 3936 50304 3942
rect 50252 3878 50304 3884
rect 50080 3738 50108 3878
rect 49884 3732 49936 3738
rect 49884 3674 49936 3680
rect 50068 3732 50120 3738
rect 50068 3674 50120 3680
rect 49896 2990 49924 3674
rect 50080 3602 50108 3674
rect 50068 3596 50120 3602
rect 50068 3538 50120 3544
rect 50080 3194 50108 3538
rect 50264 3466 50292 3878
rect 50434 3768 50490 3777
rect 50434 3703 50490 3712
rect 50252 3460 50304 3466
rect 50252 3402 50304 3408
rect 50068 3188 50120 3194
rect 50068 3130 50120 3136
rect 50448 3058 50476 3703
rect 50632 3466 50660 4082
rect 50908 4049 50936 4762
rect 50988 4480 51040 4486
rect 50988 4422 51040 4428
rect 50894 4040 50950 4049
rect 50894 3975 50950 3984
rect 51000 3754 51028 4422
rect 51092 4026 51120 7398
rect 51172 6724 51224 6730
rect 51172 6666 51224 6672
rect 51184 4554 51212 6666
rect 51552 6633 51580 8774
rect 51736 8650 51764 8774
rect 51644 8622 51764 8650
rect 51644 8362 51672 8622
rect 51632 8356 51684 8362
rect 51632 8298 51684 8304
rect 52012 8294 52040 10202
rect 52000 8288 52052 8294
rect 52000 8230 52052 8236
rect 51998 7984 52054 7993
rect 51998 7919 52000 7928
rect 52052 7919 52054 7928
rect 52000 7890 52052 7896
rect 51908 7880 51960 7886
rect 51814 7848 51870 7857
rect 51908 7822 51960 7828
rect 51814 7783 51870 7792
rect 51632 7540 51684 7546
rect 51632 7482 51684 7488
rect 51644 7206 51672 7482
rect 51632 7200 51684 7206
rect 51632 7142 51684 7148
rect 51644 7002 51672 7142
rect 51632 6996 51684 7002
rect 51632 6938 51684 6944
rect 51538 6624 51594 6633
rect 51538 6559 51594 6568
rect 51828 5778 51856 7783
rect 51920 7410 51948 7822
rect 52012 7546 52040 7890
rect 52000 7540 52052 7546
rect 52000 7482 52052 7488
rect 51908 7404 51960 7410
rect 51908 7346 51960 7352
rect 51908 6248 51960 6254
rect 51906 6216 51908 6225
rect 51960 6216 51962 6225
rect 51906 6151 51962 6160
rect 51816 5772 51868 5778
rect 51816 5714 51868 5720
rect 51448 5568 51500 5574
rect 51448 5510 51500 5516
rect 51460 4554 51488 5510
rect 51828 5370 51856 5714
rect 51816 5364 51868 5370
rect 51816 5306 51868 5312
rect 51540 5024 51592 5030
rect 51540 4966 51592 4972
rect 51552 4758 51580 4966
rect 51540 4752 51592 4758
rect 51538 4720 51540 4729
rect 51816 4752 51868 4758
rect 51592 4720 51594 4729
rect 51816 4694 51868 4700
rect 51538 4655 51594 4664
rect 51172 4548 51224 4554
rect 51172 4490 51224 4496
rect 51448 4548 51500 4554
rect 51448 4490 51500 4496
rect 51540 4480 51592 4486
rect 51828 4468 51856 4694
rect 51920 4672 51948 6151
rect 52000 4684 52052 4690
rect 51920 4644 52000 4672
rect 52000 4626 52052 4632
rect 51592 4440 51856 4468
rect 51908 4480 51960 4486
rect 51540 4422 51592 4428
rect 51828 4078 51856 4440
rect 51906 4448 51908 4457
rect 51960 4448 51962 4457
rect 51906 4383 51962 4392
rect 51724 4072 51776 4078
rect 51092 3998 51212 4026
rect 51724 4014 51776 4020
rect 51816 4072 51868 4078
rect 51816 4014 51868 4020
rect 51080 3936 51132 3942
rect 51080 3878 51132 3884
rect 50816 3726 51028 3754
rect 50816 3670 50844 3726
rect 50804 3664 50856 3670
rect 50804 3606 50856 3612
rect 51092 3602 51120 3878
rect 51080 3596 51132 3602
rect 51184 3584 51212 3998
rect 51736 3777 51764 4014
rect 52000 4004 52052 4010
rect 52000 3946 52052 3952
rect 51722 3768 51778 3777
rect 51722 3703 51778 3712
rect 52012 3602 52040 3946
rect 51724 3596 51776 3602
rect 51184 3556 51304 3584
rect 51080 3538 51132 3544
rect 50620 3460 50672 3466
rect 50620 3402 50672 3408
rect 51172 3460 51224 3466
rect 51172 3402 51224 3408
rect 51184 3058 51212 3402
rect 50436 3052 50488 3058
rect 50436 2994 50488 3000
rect 51172 3052 51224 3058
rect 51172 2994 51224 3000
rect 49884 2984 49936 2990
rect 49884 2926 49936 2932
rect 50528 2984 50580 2990
rect 50528 2926 50580 2932
rect 49896 2650 49924 2926
rect 49884 2644 49936 2650
rect 49884 2586 49936 2592
rect 49792 2576 49844 2582
rect 49792 2518 49844 2524
rect 49332 2440 49384 2446
rect 49332 2382 49384 2388
rect 49344 2038 49372 2382
rect 49896 2378 49924 2586
rect 50540 2582 50568 2926
rect 51080 2916 51132 2922
rect 51080 2858 51132 2864
rect 50528 2576 50580 2582
rect 50528 2518 50580 2524
rect 51092 2514 51120 2858
rect 51276 2582 51304 3556
rect 51724 3538 51776 3544
rect 52000 3596 52052 3602
rect 52000 3538 52052 3544
rect 51736 3482 51764 3538
rect 51736 3454 52040 3482
rect 52104 3466 52132 13262
rect 52196 11200 52224 13806
rect 52368 13796 52420 13802
rect 52368 13738 52420 13744
rect 52380 13394 52408 13738
rect 52368 13388 52420 13394
rect 52368 13330 52420 13336
rect 52380 12918 52408 13330
rect 52368 12912 52420 12918
rect 52368 12854 52420 12860
rect 52276 12164 52328 12170
rect 52276 12106 52328 12112
rect 52288 11694 52316 12106
rect 52368 12096 52420 12102
rect 52368 12038 52420 12044
rect 52380 11898 52408 12038
rect 52472 11898 52500 13874
rect 52656 13870 52684 14418
rect 53392 14414 53420 15846
rect 53484 15570 53512 16934
rect 53748 16448 53800 16454
rect 53748 16390 53800 16396
rect 53760 16114 53788 16390
rect 53852 16232 53880 17274
rect 53932 17128 53984 17134
rect 53932 17070 53984 17076
rect 53944 16794 53972 17070
rect 53932 16788 53984 16794
rect 53984 16748 54064 16776
rect 53932 16730 53984 16736
rect 53932 16244 53984 16250
rect 53852 16204 53932 16232
rect 53932 16186 53984 16192
rect 53748 16108 53800 16114
rect 53748 16050 53800 16056
rect 53472 15564 53524 15570
rect 53472 15506 53524 15512
rect 53484 15094 53512 15506
rect 53472 15088 53524 15094
rect 53472 15030 53524 15036
rect 53760 15026 53788 16050
rect 54036 15706 54064 16748
rect 54024 15700 54076 15706
rect 54024 15642 54076 15648
rect 55680 15360 55732 15366
rect 55680 15302 55732 15308
rect 53748 15020 53800 15026
rect 53748 14962 53800 14968
rect 55692 14958 55720 15302
rect 53840 14952 53892 14958
rect 53840 14894 53892 14900
rect 55680 14952 55732 14958
rect 55680 14894 55732 14900
rect 53380 14408 53432 14414
rect 53380 14350 53432 14356
rect 53748 14408 53800 14414
rect 53748 14350 53800 14356
rect 52828 14272 52880 14278
rect 52828 14214 52880 14220
rect 52644 13864 52696 13870
rect 52644 13806 52696 13812
rect 52736 13864 52788 13870
rect 52736 13806 52788 13812
rect 52748 13682 52776 13806
rect 52656 13654 52776 13682
rect 52552 13184 52604 13190
rect 52552 13126 52604 13132
rect 52564 12986 52592 13126
rect 52552 12980 52604 12986
rect 52552 12922 52604 12928
rect 52564 12442 52592 12922
rect 52552 12436 52604 12442
rect 52552 12378 52604 12384
rect 52368 11892 52420 11898
rect 52368 11834 52420 11840
rect 52460 11892 52512 11898
rect 52460 11834 52512 11840
rect 52276 11688 52328 11694
rect 52276 11630 52328 11636
rect 52380 11286 52408 11834
rect 52460 11756 52512 11762
rect 52460 11698 52512 11704
rect 52368 11280 52420 11286
rect 52368 11222 52420 11228
rect 52276 11212 52328 11218
rect 52196 11172 52276 11200
rect 52276 11154 52328 11160
rect 52288 10470 52316 11154
rect 52276 10464 52328 10470
rect 52274 10432 52276 10441
rect 52328 10432 52330 10441
rect 52274 10367 52330 10376
rect 52368 9580 52420 9586
rect 52368 9522 52420 9528
rect 52380 9110 52408 9522
rect 52472 9110 52500 11698
rect 52564 11354 52592 12378
rect 52552 11348 52604 11354
rect 52552 11290 52604 11296
rect 52656 9518 52684 13654
rect 52840 12306 52868 14214
rect 52936 14172 53232 14192
rect 52992 14170 53016 14172
rect 53072 14170 53096 14172
rect 53152 14170 53176 14172
rect 53014 14118 53016 14170
rect 53078 14118 53090 14170
rect 53152 14118 53154 14170
rect 52992 14116 53016 14118
rect 53072 14116 53096 14118
rect 53152 14116 53176 14118
rect 52936 14096 53232 14116
rect 53760 14006 53788 14350
rect 53852 14278 53880 14894
rect 55496 14816 55548 14822
rect 55496 14758 55548 14764
rect 55508 14414 55536 14758
rect 55220 14408 55272 14414
rect 55220 14350 55272 14356
rect 55496 14408 55548 14414
rect 55496 14350 55548 14356
rect 53840 14272 53892 14278
rect 53840 14214 53892 14220
rect 54576 14272 54628 14278
rect 54576 14214 54628 14220
rect 53288 14000 53340 14006
rect 53288 13942 53340 13948
rect 53748 14000 53800 14006
rect 53748 13942 53800 13948
rect 52936 13084 53232 13104
rect 52992 13082 53016 13084
rect 53072 13082 53096 13084
rect 53152 13082 53176 13084
rect 53014 13030 53016 13082
rect 53078 13030 53090 13082
rect 53152 13030 53154 13082
rect 52992 13028 53016 13030
rect 53072 13028 53096 13030
rect 53152 13028 53176 13030
rect 52936 13008 53232 13028
rect 53300 12782 53328 13942
rect 53472 13252 53524 13258
rect 53472 13194 53524 13200
rect 54208 13252 54260 13258
rect 54208 13194 54260 13200
rect 53484 12782 53512 13194
rect 53656 12912 53708 12918
rect 53656 12854 53708 12860
rect 53288 12776 53340 12782
rect 53472 12776 53524 12782
rect 53340 12724 53420 12730
rect 53288 12718 53420 12724
rect 53472 12718 53524 12724
rect 53300 12702 53420 12718
rect 53392 12646 53420 12702
rect 53288 12640 53340 12646
rect 53288 12582 53340 12588
rect 53380 12640 53432 12646
rect 53380 12582 53432 12588
rect 52828 12300 52880 12306
rect 52828 12242 52880 12248
rect 52840 11626 52868 12242
rect 53300 12238 53328 12582
rect 53472 12300 53524 12306
rect 53472 12242 53524 12248
rect 53288 12232 53340 12238
rect 53288 12174 53340 12180
rect 52936 11996 53232 12016
rect 52992 11994 53016 11996
rect 53072 11994 53096 11996
rect 53152 11994 53176 11996
rect 53014 11942 53016 11994
rect 53078 11942 53090 11994
rect 53152 11942 53154 11994
rect 52992 11940 53016 11942
rect 53072 11940 53096 11942
rect 53152 11940 53176 11942
rect 52936 11920 53232 11940
rect 52828 11620 52880 11626
rect 52828 11562 52880 11568
rect 53196 11144 53248 11150
rect 53300 11098 53328 12174
rect 53484 11898 53512 12242
rect 53472 11892 53524 11898
rect 53472 11834 53524 11840
rect 53484 11150 53512 11834
rect 53564 11824 53616 11830
rect 53564 11766 53616 11772
rect 53576 11354 53604 11766
rect 53564 11348 53616 11354
rect 53564 11290 53616 11296
rect 53248 11092 53328 11098
rect 53196 11086 53328 11092
rect 53472 11144 53524 11150
rect 53472 11086 53524 11092
rect 53208 11070 53328 11086
rect 52936 10908 53232 10928
rect 52992 10906 53016 10908
rect 53072 10906 53096 10908
rect 53152 10906 53176 10908
rect 53014 10854 53016 10906
rect 53078 10854 53090 10906
rect 53152 10854 53154 10906
rect 52992 10852 53016 10854
rect 53072 10852 53096 10854
rect 53152 10852 53176 10854
rect 52936 10832 53232 10852
rect 52828 10464 52880 10470
rect 52828 10406 52880 10412
rect 52736 10124 52788 10130
rect 52736 10066 52788 10072
rect 52748 9874 52776 10066
rect 52840 9994 52868 10406
rect 52828 9988 52880 9994
rect 52828 9930 52880 9936
rect 52748 9846 52868 9874
rect 52644 9512 52696 9518
rect 52644 9454 52696 9460
rect 52368 9104 52420 9110
rect 52368 9046 52420 9052
rect 52460 9104 52512 9110
rect 52460 9046 52512 9052
rect 52736 9036 52788 9042
rect 52736 8978 52788 8984
rect 52276 8832 52328 8838
rect 52276 8774 52328 8780
rect 52288 8498 52316 8774
rect 52748 8634 52776 8978
rect 52840 8838 52868 9846
rect 52936 9820 53232 9840
rect 52992 9818 53016 9820
rect 53072 9818 53096 9820
rect 53152 9818 53176 9820
rect 53014 9766 53016 9818
rect 53078 9766 53090 9818
rect 53152 9766 53154 9818
rect 52992 9764 53016 9766
rect 53072 9764 53096 9766
rect 53152 9764 53176 9766
rect 52936 9744 53232 9764
rect 53300 9586 53328 11070
rect 53564 10124 53616 10130
rect 53564 10066 53616 10072
rect 53576 9586 53604 10066
rect 53288 9580 53340 9586
rect 53288 9522 53340 9528
rect 53564 9580 53616 9586
rect 53564 9522 53616 9528
rect 53564 9036 53616 9042
rect 53564 8978 53616 8984
rect 53288 8968 53340 8974
rect 53288 8910 53340 8916
rect 52828 8832 52880 8838
rect 52828 8774 52880 8780
rect 52736 8628 52788 8634
rect 52736 8570 52788 8576
rect 52840 8566 52868 8774
rect 52936 8732 53232 8752
rect 52992 8730 53016 8732
rect 53072 8730 53096 8732
rect 53152 8730 53176 8732
rect 53014 8678 53016 8730
rect 53078 8678 53090 8730
rect 53152 8678 53154 8730
rect 52992 8676 53016 8678
rect 53072 8676 53096 8678
rect 53152 8676 53176 8678
rect 52936 8656 53232 8676
rect 52828 8560 52880 8566
rect 52828 8502 52880 8508
rect 52184 8492 52236 8498
rect 52184 8434 52236 8440
rect 52276 8492 52328 8498
rect 52276 8434 52328 8440
rect 52196 8294 52224 8434
rect 52460 8356 52512 8362
rect 52460 8298 52512 8304
rect 52184 8288 52236 8294
rect 52184 8230 52236 8236
rect 52196 8090 52224 8230
rect 52184 8084 52236 8090
rect 52184 8026 52236 8032
rect 52472 7954 52500 8298
rect 52550 7984 52606 7993
rect 52460 7948 52512 7954
rect 52550 7919 52606 7928
rect 52460 7890 52512 7896
rect 52182 7712 52238 7721
rect 52182 7647 52238 7656
rect 52196 7206 52224 7647
rect 52564 7478 52592 7919
rect 53300 7750 53328 8910
rect 53576 8634 53604 8978
rect 53564 8628 53616 8634
rect 53564 8570 53616 8576
rect 53380 8084 53432 8090
rect 53380 8026 53432 8032
rect 53288 7744 53340 7750
rect 53288 7686 53340 7692
rect 52936 7644 53232 7664
rect 52992 7642 53016 7644
rect 53072 7642 53096 7644
rect 53152 7642 53176 7644
rect 53014 7590 53016 7642
rect 53078 7590 53090 7642
rect 53152 7590 53154 7642
rect 52992 7588 53016 7590
rect 53072 7588 53096 7590
rect 53152 7588 53176 7590
rect 52936 7568 53232 7588
rect 52552 7472 52604 7478
rect 53012 7472 53064 7478
rect 52552 7414 52604 7420
rect 53010 7440 53012 7449
rect 53064 7440 53066 7449
rect 53010 7375 53066 7384
rect 52736 7268 52788 7274
rect 52736 7210 52788 7216
rect 52184 7200 52236 7206
rect 52184 7142 52236 7148
rect 52196 6798 52224 7142
rect 52460 6860 52512 6866
rect 52460 6802 52512 6808
rect 52184 6792 52236 6798
rect 52184 6734 52236 6740
rect 52184 6452 52236 6458
rect 52184 6394 52236 6400
rect 52196 5914 52224 6394
rect 52368 6112 52420 6118
rect 52472 6100 52500 6802
rect 52552 6112 52604 6118
rect 52472 6072 52552 6100
rect 52368 6054 52420 6060
rect 52552 6054 52604 6060
rect 52184 5908 52236 5914
rect 52184 5850 52236 5856
rect 52276 5908 52328 5914
rect 52276 5850 52328 5856
rect 52288 4758 52316 5850
rect 52380 4758 52408 6054
rect 52564 5148 52592 6054
rect 52748 5234 52776 7210
rect 53300 6866 53328 7686
rect 53288 6860 53340 6866
rect 53288 6802 53340 6808
rect 53288 6656 53340 6662
rect 53288 6598 53340 6604
rect 52936 6556 53232 6576
rect 52992 6554 53016 6556
rect 53072 6554 53096 6556
rect 53152 6554 53176 6556
rect 53014 6502 53016 6554
rect 53078 6502 53090 6554
rect 53152 6502 53154 6554
rect 52992 6500 53016 6502
rect 53072 6500 53096 6502
rect 53152 6500 53176 6502
rect 52936 6480 53232 6500
rect 53300 6322 53328 6598
rect 53392 6322 53420 8026
rect 53576 7206 53604 8570
rect 53564 7200 53616 7206
rect 53564 7142 53616 7148
rect 53288 6316 53340 6322
rect 53288 6258 53340 6264
rect 53380 6316 53432 6322
rect 53380 6258 53432 6264
rect 53012 6248 53064 6254
rect 53010 6216 53012 6225
rect 53064 6216 53066 6225
rect 53010 6151 53066 6160
rect 52828 5840 52880 5846
rect 52828 5782 52880 5788
rect 52736 5228 52788 5234
rect 52736 5170 52788 5176
rect 52840 5166 52868 5782
rect 53300 5642 53328 6258
rect 53380 5772 53432 5778
rect 53380 5714 53432 5720
rect 53288 5636 53340 5642
rect 53288 5578 53340 5584
rect 52936 5468 53232 5488
rect 52992 5466 53016 5468
rect 53072 5466 53096 5468
rect 53152 5466 53176 5468
rect 53014 5414 53016 5466
rect 53078 5414 53090 5466
rect 53152 5414 53154 5466
rect 52992 5412 53016 5414
rect 53072 5412 53096 5414
rect 53152 5412 53176 5414
rect 52936 5392 53232 5412
rect 53392 5302 53420 5714
rect 53380 5296 53432 5302
rect 53380 5238 53432 5244
rect 52644 5160 52696 5166
rect 52564 5120 52644 5148
rect 52644 5102 52696 5108
rect 52828 5160 52880 5166
rect 52828 5102 52880 5108
rect 52552 5024 52604 5030
rect 52552 4966 52604 4972
rect 52276 4752 52328 4758
rect 52276 4694 52328 4700
rect 52368 4752 52420 4758
rect 52368 4694 52420 4700
rect 52368 4548 52420 4554
rect 52368 4490 52420 4496
rect 52184 4480 52236 4486
rect 52184 4422 52236 4428
rect 52196 4185 52224 4422
rect 52182 4176 52238 4185
rect 52182 4111 52184 4120
rect 52236 4111 52238 4120
rect 52184 4082 52236 4088
rect 52196 4051 52224 4082
rect 52380 3738 52408 4490
rect 52564 4214 52592 4966
rect 52656 4468 52684 5102
rect 52736 4480 52788 4486
rect 52656 4440 52736 4468
rect 52736 4422 52788 4428
rect 52552 4208 52604 4214
rect 52552 4150 52604 4156
rect 52552 4072 52604 4078
rect 52550 4040 52552 4049
rect 52748 4049 52776 4422
rect 52840 4146 52868 5102
rect 53668 4842 53696 12854
rect 54116 12232 54168 12238
rect 54116 12174 54168 12180
rect 53932 12096 53984 12102
rect 53932 12038 53984 12044
rect 53944 10674 53972 12038
rect 54128 11694 54156 12174
rect 54220 12170 54248 13194
rect 54208 12164 54260 12170
rect 54208 12106 54260 12112
rect 54588 11898 54616 14214
rect 55128 14000 55180 14006
rect 55128 13942 55180 13948
rect 55140 13530 55168 13942
rect 55232 13870 55260 14350
rect 55508 13870 55536 14350
rect 55588 14272 55640 14278
rect 55588 14214 55640 14220
rect 55600 14006 55628 14214
rect 55692 14074 55720 14894
rect 55784 14618 55812 19162
rect 57152 16040 57204 16046
rect 57152 15982 57204 15988
rect 56968 15904 57020 15910
rect 56968 15846 57020 15852
rect 56980 15570 57008 15846
rect 56876 15564 56928 15570
rect 56876 15506 56928 15512
rect 56968 15564 57020 15570
rect 56968 15506 57020 15512
rect 55864 15496 55916 15502
rect 55864 15438 55916 15444
rect 56784 15496 56836 15502
rect 56784 15438 56836 15444
rect 55876 14958 55904 15438
rect 55864 14952 55916 14958
rect 55864 14894 55916 14900
rect 56232 14952 56284 14958
rect 56232 14894 56284 14900
rect 55772 14612 55824 14618
rect 55772 14554 55824 14560
rect 55784 14074 55812 14554
rect 55864 14476 55916 14482
rect 55864 14418 55916 14424
rect 55680 14068 55732 14074
rect 55680 14010 55732 14016
rect 55772 14068 55824 14074
rect 55772 14010 55824 14016
rect 55588 14000 55640 14006
rect 55588 13942 55640 13948
rect 55220 13864 55272 13870
rect 55220 13806 55272 13812
rect 55496 13864 55548 13870
rect 55496 13806 55548 13812
rect 55128 13524 55180 13530
rect 55128 13466 55180 13472
rect 55140 12714 55168 13466
rect 55232 12850 55260 13806
rect 55600 13326 55628 13942
rect 55692 13394 55720 14010
rect 55876 13870 55904 14418
rect 55864 13864 55916 13870
rect 55864 13806 55916 13812
rect 55680 13388 55732 13394
rect 55680 13330 55732 13336
rect 55588 13320 55640 13326
rect 55588 13262 55640 13268
rect 56048 13320 56100 13326
rect 56048 13262 56100 13268
rect 56060 12918 56088 13262
rect 56048 12912 56100 12918
rect 56048 12854 56100 12860
rect 55220 12844 55272 12850
rect 55220 12786 55272 12792
rect 55128 12708 55180 12714
rect 55128 12650 55180 12656
rect 55864 12708 55916 12714
rect 55864 12650 55916 12656
rect 55680 12640 55732 12646
rect 55732 12588 55812 12594
rect 55680 12582 55812 12588
rect 55692 12566 55812 12582
rect 55404 12368 55456 12374
rect 55404 12310 55456 12316
rect 55128 12300 55180 12306
rect 55128 12242 55180 12248
rect 54576 11892 54628 11898
rect 54576 11834 54628 11840
rect 54116 11688 54168 11694
rect 54116 11630 54168 11636
rect 54128 11354 54156 11630
rect 54852 11552 54904 11558
rect 54852 11494 54904 11500
rect 55036 11552 55088 11558
rect 55036 11494 55088 11500
rect 54116 11348 54168 11354
rect 54116 11290 54168 11296
rect 53932 10668 53984 10674
rect 53932 10610 53984 10616
rect 53944 10266 53972 10610
rect 54484 10600 54536 10606
rect 54484 10542 54536 10548
rect 54392 10464 54444 10470
rect 54392 10406 54444 10412
rect 53932 10260 53984 10266
rect 53932 10202 53984 10208
rect 53840 10056 53892 10062
rect 53840 9998 53892 10004
rect 53852 9722 53880 9998
rect 53840 9716 53892 9722
rect 53840 9658 53892 9664
rect 53840 8356 53892 8362
rect 53840 8298 53892 8304
rect 53852 8022 53880 8298
rect 53944 8090 53972 10202
rect 54404 9722 54432 10406
rect 54496 10266 54524 10542
rect 54484 10260 54536 10266
rect 54484 10202 54536 10208
rect 54760 10056 54812 10062
rect 54760 9998 54812 10004
rect 54392 9716 54444 9722
rect 54392 9658 54444 9664
rect 54208 9104 54260 9110
rect 54208 9046 54260 9052
rect 54220 8430 54248 9046
rect 54300 8968 54352 8974
rect 54300 8910 54352 8916
rect 54208 8424 54260 8430
rect 54208 8366 54260 8372
rect 53932 8084 53984 8090
rect 53932 8026 53984 8032
rect 53840 8016 53892 8022
rect 53840 7958 53892 7964
rect 53748 7948 53800 7954
rect 53748 7890 53800 7896
rect 53760 7546 53788 7890
rect 53748 7540 53800 7546
rect 53748 7482 53800 7488
rect 54116 7200 54168 7206
rect 54116 7142 54168 7148
rect 54128 6934 54156 7142
rect 54220 7002 54248 8366
rect 54312 7750 54340 8910
rect 54772 8906 54800 9998
rect 54760 8900 54812 8906
rect 54760 8842 54812 8848
rect 54300 7744 54352 7750
rect 54300 7686 54352 7692
rect 54208 6996 54260 7002
rect 54208 6938 54260 6944
rect 54116 6928 54168 6934
rect 54116 6870 54168 6876
rect 53840 6792 53892 6798
rect 53840 6734 53892 6740
rect 53852 5710 53880 6734
rect 54024 6656 54076 6662
rect 54024 6598 54076 6604
rect 53840 5704 53892 5710
rect 53840 5646 53892 5652
rect 53852 5370 53880 5646
rect 53840 5364 53892 5370
rect 53840 5306 53892 5312
rect 54036 5302 54064 6598
rect 54024 5296 54076 5302
rect 54024 5238 54076 5244
rect 53668 4814 53788 4842
rect 53656 4752 53708 4758
rect 53656 4694 53708 4700
rect 53196 4684 53248 4690
rect 53248 4644 53328 4672
rect 53196 4626 53248 4632
rect 52936 4380 53232 4400
rect 52992 4378 53016 4380
rect 53072 4378 53096 4380
rect 53152 4378 53176 4380
rect 53014 4326 53016 4378
rect 53078 4326 53090 4378
rect 53152 4326 53154 4378
rect 52992 4324 53016 4326
rect 53072 4324 53096 4326
rect 53152 4324 53176 4326
rect 52936 4304 53232 4324
rect 53300 4214 53328 4644
rect 53288 4208 53340 4214
rect 53288 4150 53340 4156
rect 52828 4140 52880 4146
rect 52828 4082 52880 4088
rect 53668 4078 53696 4694
rect 53380 4072 53432 4078
rect 52604 4040 52606 4049
rect 52550 3975 52606 3984
rect 52734 4040 52790 4049
rect 53380 4014 53432 4020
rect 53564 4072 53616 4078
rect 53564 4014 53616 4020
rect 53656 4072 53708 4078
rect 53656 4014 53708 4020
rect 52734 3975 52790 3984
rect 52748 3890 52776 3975
rect 53392 3942 53420 4014
rect 52472 3862 52776 3890
rect 53288 3936 53340 3942
rect 53288 3878 53340 3884
rect 53380 3936 53432 3942
rect 53380 3878 53432 3884
rect 52368 3732 52420 3738
rect 52368 3674 52420 3680
rect 52184 3596 52236 3602
rect 52184 3538 52236 3544
rect 52368 3596 52420 3602
rect 52368 3538 52420 3544
rect 51540 3392 51592 3398
rect 51540 3334 51592 3340
rect 51816 3392 51868 3398
rect 51816 3334 51868 3340
rect 51552 2990 51580 3334
rect 51724 3052 51776 3058
rect 51724 2994 51776 3000
rect 51540 2984 51592 2990
rect 51540 2926 51592 2932
rect 51264 2576 51316 2582
rect 51264 2518 51316 2524
rect 51080 2508 51132 2514
rect 51080 2450 51132 2456
rect 50804 2440 50856 2446
rect 50804 2382 50856 2388
rect 49884 2372 49936 2378
rect 49884 2314 49936 2320
rect 49976 2100 50028 2106
rect 49976 2042 50028 2048
rect 49332 2032 49384 2038
rect 49332 1974 49384 1980
rect 49988 800 50016 2042
rect 50816 800 50844 2382
rect 51552 2310 51580 2926
rect 51540 2304 51592 2310
rect 51540 2246 51592 2252
rect 51552 2106 51580 2246
rect 51540 2100 51592 2106
rect 51540 2042 51592 2048
rect 51736 800 51764 2994
rect 51828 2854 51856 3334
rect 51816 2848 51868 2854
rect 51816 2790 51868 2796
rect 51920 2650 51948 3454
rect 52012 3346 52040 3454
rect 52092 3460 52144 3466
rect 52092 3402 52144 3408
rect 52196 3346 52224 3538
rect 52012 3318 52224 3346
rect 52196 3126 52224 3318
rect 52380 3194 52408 3538
rect 52472 3398 52500 3862
rect 53300 3398 53328 3878
rect 53392 3602 53420 3878
rect 53380 3596 53432 3602
rect 53380 3538 53432 3544
rect 52460 3392 52512 3398
rect 52460 3334 52512 3340
rect 52644 3392 52696 3398
rect 52644 3334 52696 3340
rect 53288 3392 53340 3398
rect 53288 3334 53340 3340
rect 52656 3194 52684 3334
rect 52936 3292 53232 3312
rect 52992 3290 53016 3292
rect 53072 3290 53096 3292
rect 53152 3290 53176 3292
rect 53014 3238 53016 3290
rect 53078 3238 53090 3290
rect 53152 3238 53154 3290
rect 52992 3236 53016 3238
rect 53072 3236 53096 3238
rect 53152 3236 53176 3238
rect 52936 3216 53232 3236
rect 52368 3188 52420 3194
rect 52368 3130 52420 3136
rect 52644 3188 52696 3194
rect 52644 3130 52696 3136
rect 52184 3120 52236 3126
rect 52184 3062 52236 3068
rect 52380 2938 52408 3130
rect 52288 2922 52408 2938
rect 52000 2916 52052 2922
rect 52000 2858 52052 2864
rect 52276 2916 52408 2922
rect 52328 2910 52408 2916
rect 52276 2858 52328 2864
rect 52012 2650 52040 2858
rect 51908 2644 51960 2650
rect 51908 2586 51960 2592
rect 52000 2644 52052 2650
rect 52000 2586 52052 2592
rect 52656 800 52684 3130
rect 53472 3120 53524 3126
rect 53472 3062 53524 3068
rect 53484 2582 53512 3062
rect 53576 2922 53604 4014
rect 53760 3602 53788 4814
rect 54024 4616 54076 4622
rect 54312 4593 54340 7686
rect 54772 6458 54800 8842
rect 54864 8838 54892 11494
rect 55048 11286 55076 11494
rect 55036 11280 55088 11286
rect 55036 11222 55088 11228
rect 54944 11212 54996 11218
rect 54944 11154 54996 11160
rect 54956 10810 54984 11154
rect 54944 10804 54996 10810
rect 54944 10746 54996 10752
rect 54956 10266 54984 10746
rect 54944 10260 54996 10266
rect 54944 10202 54996 10208
rect 54956 9518 54984 10202
rect 55140 9586 55168 12242
rect 55416 12102 55444 12310
rect 55496 12232 55548 12238
rect 55496 12174 55548 12180
rect 55220 12096 55272 12102
rect 55220 12038 55272 12044
rect 55404 12096 55456 12102
rect 55404 12038 55456 12044
rect 55232 11354 55260 12038
rect 55416 11830 55444 12038
rect 55508 11898 55536 12174
rect 55496 11892 55548 11898
rect 55496 11834 55548 11840
rect 55404 11824 55456 11830
rect 55404 11766 55456 11772
rect 55508 11762 55536 11834
rect 55784 11830 55812 12566
rect 55876 12374 55904 12650
rect 55864 12368 55916 12374
rect 55864 12310 55916 12316
rect 55956 12096 56008 12102
rect 55956 12038 56008 12044
rect 55968 11830 55996 12038
rect 56244 11898 56272 14894
rect 56416 14884 56468 14890
rect 56416 14826 56468 14832
rect 56428 14482 56456 14826
rect 56796 14550 56824 15438
rect 56888 15162 56916 15506
rect 56876 15156 56928 15162
rect 56876 15098 56928 15104
rect 56784 14544 56836 14550
rect 56784 14486 56836 14492
rect 56416 14476 56468 14482
rect 56416 14418 56468 14424
rect 56428 14074 56456 14418
rect 56980 14414 57008 15506
rect 56968 14408 57020 14414
rect 56968 14350 57020 14356
rect 56980 14278 57008 14350
rect 56784 14272 56836 14278
rect 56784 14214 56836 14220
rect 56968 14272 57020 14278
rect 56968 14214 57020 14220
rect 56416 14068 56468 14074
rect 56416 14010 56468 14016
rect 56796 13462 56824 14214
rect 56980 13870 57008 14214
rect 56968 13864 57020 13870
rect 56968 13806 57020 13812
rect 57164 13530 57192 15982
rect 57716 15638 57744 19162
rect 57704 15632 57756 15638
rect 57704 15574 57756 15580
rect 57244 14952 57296 14958
rect 57244 14894 57296 14900
rect 57256 14414 57284 14894
rect 57716 14618 57744 15574
rect 58164 15496 58216 15502
rect 58164 15438 58216 15444
rect 57980 15360 58032 15366
rect 57980 15302 58032 15308
rect 57992 14958 58020 15302
rect 57980 14952 58032 14958
rect 57980 14894 58032 14900
rect 57704 14612 57756 14618
rect 57704 14554 57756 14560
rect 57244 14408 57296 14414
rect 57244 14350 57296 14356
rect 58176 13870 58204 15438
rect 59740 15434 59768 19162
rect 61672 15706 61700 19162
rect 61660 15700 61712 15706
rect 61660 15642 61712 15648
rect 58900 15428 58952 15434
rect 58900 15370 58952 15376
rect 59728 15428 59780 15434
rect 59728 15370 59780 15376
rect 58912 15162 58940 15370
rect 58900 15156 58952 15162
rect 58900 15098 58952 15104
rect 58716 14952 58768 14958
rect 58716 14894 58768 14900
rect 58440 14000 58492 14006
rect 58440 13942 58492 13948
rect 58164 13864 58216 13870
rect 58084 13812 58164 13818
rect 58084 13806 58216 13812
rect 57888 13796 57940 13802
rect 57888 13738 57940 13744
rect 58084 13790 58204 13806
rect 57152 13524 57204 13530
rect 57152 13466 57204 13472
rect 56784 13456 56836 13462
rect 56784 13398 56836 13404
rect 57796 13456 57848 13462
rect 57796 13398 57848 13404
rect 56796 12918 56824 13398
rect 57336 13252 57388 13258
rect 57336 13194 57388 13200
rect 56784 12912 56836 12918
rect 56784 12854 56836 12860
rect 56876 12300 56928 12306
rect 56876 12242 56928 12248
rect 56888 12102 56916 12242
rect 56692 12096 56744 12102
rect 56692 12038 56744 12044
rect 56876 12096 56928 12102
rect 56876 12038 56928 12044
rect 56232 11892 56284 11898
rect 56232 11834 56284 11840
rect 55772 11824 55824 11830
rect 55772 11766 55824 11772
rect 55956 11824 56008 11830
rect 55956 11766 56008 11772
rect 55496 11756 55548 11762
rect 55496 11698 55548 11704
rect 56140 11688 56192 11694
rect 56140 11630 56192 11636
rect 55220 11348 55272 11354
rect 55220 11290 55272 11296
rect 55232 9926 55260 11290
rect 55772 11076 55824 11082
rect 55772 11018 55824 11024
rect 55496 10600 55548 10606
rect 55496 10542 55548 10548
rect 55404 10532 55456 10538
rect 55404 10474 55456 10480
rect 55416 10198 55444 10474
rect 55404 10192 55456 10198
rect 55404 10134 55456 10140
rect 55220 9920 55272 9926
rect 55220 9862 55272 9868
rect 55416 9722 55444 10134
rect 55404 9716 55456 9722
rect 55404 9658 55456 9664
rect 55128 9580 55180 9586
rect 55128 9522 55180 9528
rect 54944 9512 54996 9518
rect 54944 9454 54996 9460
rect 55416 9042 55444 9658
rect 55220 9036 55272 9042
rect 55220 8978 55272 8984
rect 55404 9036 55456 9042
rect 55404 8978 55456 8984
rect 55128 8968 55180 8974
rect 55128 8910 55180 8916
rect 54852 8832 54904 8838
rect 54852 8774 54904 8780
rect 55140 8090 55168 8910
rect 55232 8430 55260 8978
rect 55220 8424 55272 8430
rect 55220 8366 55272 8372
rect 55312 8356 55364 8362
rect 55312 8298 55364 8304
rect 55404 8356 55456 8362
rect 55404 8298 55456 8304
rect 55324 8090 55352 8298
rect 55128 8084 55180 8090
rect 55128 8026 55180 8032
rect 55312 8084 55364 8090
rect 55312 8026 55364 8032
rect 55036 6928 55088 6934
rect 54942 6896 54998 6905
rect 55140 6916 55168 8026
rect 55416 7886 55444 8298
rect 55404 7880 55456 7886
rect 55404 7822 55456 7828
rect 55416 7546 55444 7822
rect 55404 7540 55456 7546
rect 55404 7482 55456 7488
rect 55088 6888 55168 6916
rect 55036 6870 55088 6876
rect 54942 6831 54944 6840
rect 54996 6831 54998 6840
rect 54944 6802 54996 6808
rect 54956 6458 54984 6802
rect 54760 6452 54812 6458
rect 54760 6394 54812 6400
rect 54944 6452 54996 6458
rect 54944 6394 54996 6400
rect 54772 5846 54800 6394
rect 54760 5840 54812 5846
rect 54760 5782 54812 5788
rect 54956 5710 54984 6394
rect 55048 6225 55076 6870
rect 55508 6458 55536 10542
rect 55784 10266 55812 11018
rect 55956 11008 56008 11014
rect 55956 10950 56008 10956
rect 55968 10606 55996 10950
rect 56152 10810 56180 11630
rect 56416 11212 56468 11218
rect 56416 11154 56468 11160
rect 56140 10804 56192 10810
rect 56140 10746 56192 10752
rect 55956 10600 56008 10606
rect 55956 10542 56008 10548
rect 56428 10266 56456 11154
rect 56704 11014 56732 12038
rect 56888 11801 56916 12038
rect 56874 11792 56930 11801
rect 56784 11756 56836 11762
rect 56874 11727 56930 11736
rect 56784 11698 56836 11704
rect 56796 11150 56824 11698
rect 57348 11150 57376 13194
rect 57808 12850 57836 13398
rect 57796 12844 57848 12850
rect 57796 12786 57848 12792
rect 57900 12238 57928 13738
rect 58084 12374 58112 13790
rect 58452 13462 58480 13942
rect 58440 13456 58492 13462
rect 58440 13398 58492 13404
rect 58256 13388 58308 13394
rect 58256 13330 58308 13336
rect 58268 12986 58296 13330
rect 58256 12980 58308 12986
rect 58256 12922 58308 12928
rect 58452 12442 58480 13398
rect 58728 13190 58756 14894
rect 58912 14074 58940 15098
rect 63604 15026 63632 19162
rect 63592 15020 63644 15026
rect 63592 14962 63644 14968
rect 58900 14068 58952 14074
rect 58900 14010 58952 14016
rect 59176 13388 59228 13394
rect 59176 13330 59228 13336
rect 58716 13184 58768 13190
rect 58716 13126 58768 13132
rect 58900 12844 58952 12850
rect 58900 12786 58952 12792
rect 58440 12436 58492 12442
rect 58440 12378 58492 12384
rect 58072 12368 58124 12374
rect 58072 12310 58124 12316
rect 57888 12232 57940 12238
rect 57888 12174 57940 12180
rect 57796 12164 57848 12170
rect 57796 12106 57848 12112
rect 57808 11694 57836 12106
rect 57428 11688 57480 11694
rect 57428 11630 57480 11636
rect 57796 11688 57848 11694
rect 57796 11630 57848 11636
rect 57440 11218 57468 11630
rect 57612 11620 57664 11626
rect 57612 11562 57664 11568
rect 57428 11212 57480 11218
rect 57428 11154 57480 11160
rect 56784 11144 56836 11150
rect 56784 11086 56836 11092
rect 57336 11144 57388 11150
rect 57336 11086 57388 11092
rect 56600 11008 56652 11014
rect 56600 10950 56652 10956
rect 56692 11008 56744 11014
rect 56692 10950 56744 10956
rect 56508 10532 56560 10538
rect 56508 10474 56560 10480
rect 55772 10260 55824 10266
rect 55772 10202 55824 10208
rect 56416 10260 56468 10266
rect 56416 10202 56468 10208
rect 56520 10130 56548 10474
rect 56612 10470 56640 10950
rect 56796 10810 56824 11086
rect 57244 11008 57296 11014
rect 57244 10950 57296 10956
rect 56784 10804 56836 10810
rect 56784 10746 56836 10752
rect 56600 10464 56652 10470
rect 56600 10406 56652 10412
rect 56508 10124 56560 10130
rect 56508 10066 56560 10072
rect 56416 10056 56468 10062
rect 56416 9998 56468 10004
rect 56428 9722 56456 9998
rect 56048 9716 56100 9722
rect 56048 9658 56100 9664
rect 56416 9716 56468 9722
rect 56416 9658 56468 9664
rect 55680 9376 55732 9382
rect 55680 9318 55732 9324
rect 55588 6656 55640 6662
rect 55588 6598 55640 6604
rect 55496 6452 55548 6458
rect 55496 6394 55548 6400
rect 55034 6216 55090 6225
rect 55600 6186 55628 6598
rect 55692 6361 55720 9318
rect 55864 8628 55916 8634
rect 55864 8570 55916 8576
rect 55876 8430 55904 8570
rect 55864 8424 55916 8430
rect 55864 8366 55916 8372
rect 55956 8356 56008 8362
rect 55956 8298 56008 8304
rect 55772 8288 55824 8294
rect 55772 8230 55824 8236
rect 55784 7342 55812 8230
rect 55968 7818 55996 8298
rect 55956 7812 56008 7818
rect 55956 7754 56008 7760
rect 55864 7744 55916 7750
rect 55864 7686 55916 7692
rect 55876 7342 55904 7686
rect 55772 7336 55824 7342
rect 55772 7278 55824 7284
rect 55864 7336 55916 7342
rect 55864 7278 55916 7284
rect 55876 6662 55904 7278
rect 55956 6792 56008 6798
rect 55956 6734 56008 6740
rect 55968 6662 55996 6734
rect 55864 6656 55916 6662
rect 55864 6598 55916 6604
rect 55956 6656 56008 6662
rect 55956 6598 56008 6604
rect 55772 6452 55824 6458
rect 55772 6394 55824 6400
rect 55678 6352 55734 6361
rect 55678 6287 55734 6296
rect 55034 6151 55090 6160
rect 55588 6180 55640 6186
rect 55588 6122 55640 6128
rect 55128 5840 55180 5846
rect 55128 5782 55180 5788
rect 54944 5704 54996 5710
rect 54944 5646 54996 5652
rect 54668 5568 54720 5574
rect 54668 5510 54720 5516
rect 54680 5166 54708 5510
rect 54668 5160 54720 5166
rect 54668 5102 54720 5108
rect 54576 5092 54628 5098
rect 54576 5034 54628 5040
rect 54484 4684 54536 4690
rect 54484 4626 54536 4632
rect 54024 4558 54076 4564
rect 54298 4584 54354 4593
rect 53932 4004 53984 4010
rect 53932 3946 53984 3952
rect 53748 3596 53800 3602
rect 53748 3538 53800 3544
rect 53944 3466 53972 3946
rect 54036 3738 54064 4558
rect 54298 4519 54300 4528
rect 54352 4519 54354 4528
rect 54300 4490 54352 4496
rect 54496 4214 54524 4626
rect 54484 4208 54536 4214
rect 54484 4150 54536 4156
rect 54116 4140 54168 4146
rect 54116 4082 54168 4088
rect 54128 3913 54156 4082
rect 54114 3904 54170 3913
rect 54114 3839 54170 3848
rect 54024 3732 54076 3738
rect 54024 3674 54076 3680
rect 53840 3460 53892 3466
rect 53840 3402 53892 3408
rect 53932 3460 53984 3466
rect 53932 3402 53984 3408
rect 53852 3194 53880 3402
rect 53840 3188 53892 3194
rect 53840 3130 53892 3136
rect 54036 2972 54064 3674
rect 54588 3602 54616 5034
rect 54760 4684 54812 4690
rect 54760 4626 54812 4632
rect 54668 4548 54720 4554
rect 54668 4490 54720 4496
rect 54680 4185 54708 4490
rect 54666 4176 54722 4185
rect 54772 4146 54800 4626
rect 55034 4584 55090 4593
rect 55034 4519 55090 4528
rect 55048 4214 55076 4519
rect 55140 4486 55168 5782
rect 55600 5642 55628 6122
rect 55784 5846 55812 6394
rect 55864 6316 55916 6322
rect 55864 6258 55916 6264
rect 55876 5914 55904 6258
rect 55864 5908 55916 5914
rect 55864 5850 55916 5856
rect 55772 5840 55824 5846
rect 55772 5782 55824 5788
rect 55784 5642 55812 5782
rect 55588 5636 55640 5642
rect 55588 5578 55640 5584
rect 55772 5636 55824 5642
rect 55772 5578 55824 5584
rect 55496 5568 55548 5574
rect 55496 5510 55548 5516
rect 55220 5364 55272 5370
rect 55220 5306 55272 5312
rect 55232 5166 55260 5306
rect 55310 5264 55366 5273
rect 55310 5199 55366 5208
rect 55220 5160 55272 5166
rect 55220 5102 55272 5108
rect 55128 4480 55180 4486
rect 55128 4422 55180 4428
rect 55036 4208 55088 4214
rect 55036 4150 55088 4156
rect 54666 4111 54722 4120
rect 54760 4140 54812 4146
rect 54760 4082 54812 4088
rect 55048 4010 55076 4150
rect 55140 4078 55168 4422
rect 55232 4146 55260 5102
rect 55220 4140 55272 4146
rect 55220 4082 55272 4088
rect 55128 4072 55180 4078
rect 55128 4014 55180 4020
rect 55218 4040 55274 4049
rect 54668 4004 54720 4010
rect 54668 3946 54720 3952
rect 55036 4004 55088 4010
rect 55036 3946 55088 3952
rect 54680 3670 54708 3946
rect 54852 3936 54904 3942
rect 54852 3878 54904 3884
rect 54864 3738 54892 3878
rect 54852 3732 54904 3738
rect 54852 3674 54904 3680
rect 54668 3664 54720 3670
rect 54668 3606 54720 3612
rect 54576 3596 54628 3602
rect 54576 3538 54628 3544
rect 54944 3596 54996 3602
rect 54944 3538 54996 3544
rect 55036 3596 55088 3602
rect 55036 3538 55088 3544
rect 54668 3188 54720 3194
rect 54668 3130 54720 3136
rect 54392 3052 54444 3058
rect 54392 2994 54444 3000
rect 54116 2984 54168 2990
rect 54036 2944 54116 2972
rect 54116 2926 54168 2932
rect 53564 2916 53616 2922
rect 53564 2858 53616 2864
rect 53748 2848 53800 2854
rect 53748 2790 53800 2796
rect 53472 2576 53524 2582
rect 53472 2518 53524 2524
rect 53760 2514 53788 2790
rect 53748 2508 53800 2514
rect 53748 2450 53800 2456
rect 53472 2304 53524 2310
rect 53472 2246 53524 2252
rect 52936 2204 53232 2224
rect 52992 2202 53016 2204
rect 53072 2202 53096 2204
rect 53152 2202 53176 2204
rect 53014 2150 53016 2202
rect 53078 2150 53090 2202
rect 53152 2150 53154 2202
rect 52992 2148 53016 2150
rect 53072 2148 53096 2150
rect 53152 2148 53176 2150
rect 52936 2128 53232 2148
rect 53484 800 53512 2246
rect 54404 800 54432 2994
rect 54680 2650 54708 3130
rect 54956 2650 54984 3538
rect 55048 3058 55076 3538
rect 55140 3194 55168 4014
rect 55218 3975 55220 3984
rect 55272 3975 55274 3984
rect 55220 3946 55272 3952
rect 55324 3602 55352 5199
rect 55508 5166 55536 5510
rect 55784 5370 55812 5578
rect 56060 5574 56088 9658
rect 56520 9654 56548 10066
rect 56612 9926 56640 10406
rect 57256 10266 57284 10950
rect 57348 10674 57376 11086
rect 57336 10668 57388 10674
rect 57336 10610 57388 10616
rect 57348 10266 57376 10610
rect 57244 10260 57296 10266
rect 57244 10202 57296 10208
rect 57336 10260 57388 10266
rect 57336 10202 57388 10208
rect 56600 9920 56652 9926
rect 56600 9862 56652 9868
rect 56508 9648 56560 9654
rect 56508 9590 56560 9596
rect 56140 9512 56192 9518
rect 56140 9454 56192 9460
rect 56152 8974 56180 9454
rect 57336 9376 57388 9382
rect 57336 9318 57388 9324
rect 56140 8968 56192 8974
rect 56140 8910 56192 8916
rect 56416 8968 56468 8974
rect 56508 8968 56560 8974
rect 56416 8910 56468 8916
rect 56506 8936 56508 8945
rect 57060 8968 57112 8974
rect 56560 8936 56562 8945
rect 56324 8832 56376 8838
rect 56324 8774 56376 8780
rect 56140 8628 56192 8634
rect 56140 8570 56192 8576
rect 56152 8430 56180 8570
rect 56336 8430 56364 8774
rect 56140 8424 56192 8430
rect 56140 8366 56192 8372
rect 56324 8424 56376 8430
rect 56324 8366 56376 8372
rect 56140 7948 56192 7954
rect 56140 7890 56192 7896
rect 56152 7857 56180 7890
rect 56138 7848 56194 7857
rect 56336 7818 56364 8366
rect 56428 8362 56456 8910
rect 57060 8910 57112 8916
rect 56506 8871 56562 8880
rect 56508 8832 56560 8838
rect 56508 8774 56560 8780
rect 56520 8498 56548 8774
rect 56600 8628 56652 8634
rect 56600 8570 56652 8576
rect 56508 8492 56560 8498
rect 56508 8434 56560 8440
rect 56416 8356 56468 8362
rect 56416 8298 56468 8304
rect 56138 7783 56194 7792
rect 56324 7812 56376 7818
rect 56152 7546 56180 7783
rect 56324 7754 56376 7760
rect 56140 7540 56192 7546
rect 56140 7482 56192 7488
rect 56336 7410 56364 7754
rect 56324 7404 56376 7410
rect 56324 7346 56376 7352
rect 56612 7206 56640 8570
rect 56690 7984 56746 7993
rect 56690 7919 56692 7928
rect 56744 7919 56746 7928
rect 56692 7890 56744 7896
rect 57072 7546 57100 8910
rect 57060 7540 57112 7546
rect 57060 7482 57112 7488
rect 57072 7342 57100 7482
rect 57060 7336 57112 7342
rect 57060 7278 57112 7284
rect 56600 7200 56652 7206
rect 56600 7142 56652 7148
rect 56612 7002 56640 7142
rect 56600 6996 56652 7002
rect 56600 6938 56652 6944
rect 56140 6656 56192 6662
rect 56140 6598 56192 6604
rect 56152 5710 56180 6598
rect 56612 6390 56640 6938
rect 57348 6866 57376 9318
rect 57440 7857 57468 11154
rect 57624 10810 57652 11562
rect 58084 11354 58112 12310
rect 58164 12096 58216 12102
rect 58164 12038 58216 12044
rect 58176 11694 58204 12038
rect 58912 11898 58940 12786
rect 59188 12102 59216 13330
rect 59268 13184 59320 13190
rect 59268 13126 59320 13132
rect 59280 12850 59308 13126
rect 59268 12844 59320 12850
rect 59268 12786 59320 12792
rect 60004 12640 60056 12646
rect 60004 12582 60056 12588
rect 60016 12374 60044 12582
rect 60004 12368 60056 12374
rect 60004 12310 60056 12316
rect 60556 12300 60608 12306
rect 60556 12242 60608 12248
rect 59176 12096 59228 12102
rect 59176 12038 59228 12044
rect 59728 12096 59780 12102
rect 59728 12038 59780 12044
rect 58900 11892 58952 11898
rect 58900 11834 58952 11840
rect 58164 11688 58216 11694
rect 58164 11630 58216 11636
rect 58072 11348 58124 11354
rect 58072 11290 58124 11296
rect 59188 11286 59216 12038
rect 59544 11824 59596 11830
rect 59544 11766 59596 11772
rect 59268 11620 59320 11626
rect 59268 11562 59320 11568
rect 59176 11280 59228 11286
rect 59176 11222 59228 11228
rect 58808 11212 58860 11218
rect 58808 11154 58860 11160
rect 57612 10804 57664 10810
rect 57612 10746 57664 10752
rect 58348 10600 58400 10606
rect 58348 10542 58400 10548
rect 57796 10056 57848 10062
rect 57796 9998 57848 10004
rect 57808 9382 57836 9998
rect 58164 9920 58216 9926
rect 58164 9862 58216 9868
rect 58176 9722 58204 9862
rect 58164 9716 58216 9722
rect 58164 9658 58216 9664
rect 58360 9518 58388 10542
rect 58820 10470 58848 11154
rect 59176 11144 59228 11150
rect 59280 11098 59308 11562
rect 59556 11354 59584 11766
rect 59740 11694 59768 12038
rect 59728 11688 59780 11694
rect 59728 11630 59780 11636
rect 59544 11348 59596 11354
rect 59544 11290 59596 11296
rect 59228 11092 59308 11098
rect 59176 11086 59308 11092
rect 59188 11070 59308 11086
rect 59188 10554 59216 11070
rect 59268 11008 59320 11014
rect 59268 10950 59320 10956
rect 59280 10606 59308 10950
rect 59556 10674 59584 11290
rect 59544 10668 59596 10674
rect 59544 10610 59596 10616
rect 59096 10526 59216 10554
rect 59268 10600 59320 10606
rect 59268 10542 59320 10548
rect 59096 10470 59124 10526
rect 58808 10464 58860 10470
rect 58808 10406 58860 10412
rect 59084 10464 59136 10470
rect 59084 10406 59136 10412
rect 58440 10124 58492 10130
rect 58440 10066 58492 10072
rect 58348 9512 58400 9518
rect 58348 9454 58400 9460
rect 57796 9376 57848 9382
rect 57796 9318 57848 9324
rect 58256 8900 58308 8906
rect 58256 8842 58308 8848
rect 57704 8628 57756 8634
rect 57704 8570 57756 8576
rect 57716 8294 57744 8570
rect 57612 8288 57664 8294
rect 57612 8230 57664 8236
rect 57704 8288 57756 8294
rect 57704 8230 57756 8236
rect 57624 8090 57652 8230
rect 57612 8084 57664 8090
rect 57612 8026 57664 8032
rect 58164 8084 58216 8090
rect 58164 8026 58216 8032
rect 57520 7880 57572 7886
rect 57426 7848 57482 7857
rect 57520 7822 57572 7828
rect 57426 7783 57482 7792
rect 57532 6866 57560 7822
rect 57624 7478 57652 8026
rect 58176 7954 58204 8026
rect 58268 7954 58296 8842
rect 58360 8430 58388 9454
rect 58452 8838 58480 10066
rect 58624 8968 58676 8974
rect 58624 8910 58676 8916
rect 58440 8832 58492 8838
rect 58440 8774 58492 8780
rect 58348 8424 58400 8430
rect 58348 8366 58400 8372
rect 58452 8090 58480 8774
rect 58636 8634 58664 8910
rect 58624 8628 58676 8634
rect 58624 8570 58676 8576
rect 58532 8424 58584 8430
rect 58532 8366 58584 8372
rect 58440 8084 58492 8090
rect 58440 8026 58492 8032
rect 58164 7948 58216 7954
rect 58164 7890 58216 7896
rect 58256 7948 58308 7954
rect 58256 7890 58308 7896
rect 57612 7472 57664 7478
rect 57612 7414 57664 7420
rect 57704 7472 57756 7478
rect 57704 7414 57756 7420
rect 57624 6934 57652 7414
rect 57716 7002 57744 7414
rect 57796 7336 57848 7342
rect 57796 7278 57848 7284
rect 58072 7336 58124 7342
rect 58072 7278 58124 7284
rect 57704 6996 57756 7002
rect 57704 6938 57756 6944
rect 57612 6928 57664 6934
rect 57612 6870 57664 6876
rect 57336 6860 57388 6866
rect 57336 6802 57388 6808
rect 57520 6860 57572 6866
rect 57520 6802 57572 6808
rect 56600 6384 56652 6390
rect 56600 6326 56652 6332
rect 57532 6322 57560 6802
rect 57612 6656 57664 6662
rect 57612 6598 57664 6604
rect 57520 6316 57572 6322
rect 57520 6258 57572 6264
rect 57624 5846 57652 6598
rect 57716 6458 57744 6938
rect 57808 6866 57836 7278
rect 57980 7268 58032 7274
rect 57980 7210 58032 7216
rect 57796 6860 57848 6866
rect 57796 6802 57848 6808
rect 57992 6798 58020 7210
rect 58084 7206 58112 7278
rect 58072 7200 58124 7206
rect 58072 7142 58124 7148
rect 57980 6792 58032 6798
rect 57980 6734 58032 6740
rect 57704 6452 57756 6458
rect 57704 6394 57756 6400
rect 57796 6452 57848 6458
rect 57796 6394 57848 6400
rect 57808 5914 57836 6394
rect 57992 6202 58020 6734
rect 58084 6372 58112 7142
rect 58256 6792 58308 6798
rect 58256 6734 58308 6740
rect 58084 6344 58204 6372
rect 57992 6174 58112 6202
rect 57980 6112 58032 6118
rect 57980 6054 58032 6060
rect 57992 5914 58020 6054
rect 57796 5908 57848 5914
rect 57796 5850 57848 5856
rect 57980 5908 58032 5914
rect 57980 5850 58032 5856
rect 57336 5840 57388 5846
rect 57336 5782 57388 5788
rect 57612 5840 57664 5846
rect 57612 5782 57664 5788
rect 56508 5772 56560 5778
rect 56508 5714 56560 5720
rect 56140 5704 56192 5710
rect 56140 5646 56192 5652
rect 56048 5568 56100 5574
rect 56048 5510 56100 5516
rect 56232 5568 56284 5574
rect 56232 5510 56284 5516
rect 56060 5370 56088 5510
rect 55772 5364 55824 5370
rect 55772 5306 55824 5312
rect 56048 5364 56100 5370
rect 56048 5306 56100 5312
rect 55404 5160 55456 5166
rect 55404 5102 55456 5108
rect 55496 5160 55548 5166
rect 55496 5102 55548 5108
rect 55416 4758 55444 5102
rect 55404 4752 55456 4758
rect 55404 4694 55456 4700
rect 56060 4706 56088 5306
rect 56060 4678 56180 4706
rect 56048 4616 56100 4622
rect 56048 4558 56100 4564
rect 56060 3942 56088 4558
rect 56152 4214 56180 4678
rect 56140 4208 56192 4214
rect 56140 4150 56192 4156
rect 55588 3936 55640 3942
rect 55588 3878 55640 3884
rect 55680 3936 55732 3942
rect 55680 3878 55732 3884
rect 56048 3936 56100 3942
rect 56048 3878 56100 3884
rect 55312 3596 55364 3602
rect 55312 3538 55364 3544
rect 55128 3188 55180 3194
rect 55128 3130 55180 3136
rect 55036 3052 55088 3058
rect 55036 2994 55088 3000
rect 55324 2990 55352 3538
rect 55312 2984 55364 2990
rect 55312 2926 55364 2932
rect 55600 2922 55628 3878
rect 55692 3670 55720 3878
rect 56244 3738 56272 5510
rect 56414 5264 56470 5273
rect 56414 5199 56416 5208
rect 56468 5199 56470 5208
rect 56416 5170 56468 5176
rect 56520 5030 56548 5714
rect 57152 5704 57204 5710
rect 56598 5638 56654 5647
rect 57152 5646 57204 5652
rect 56598 5573 56654 5582
rect 56600 5568 56652 5573
rect 56600 5510 56652 5516
rect 57164 5166 57192 5646
rect 57152 5160 57204 5166
rect 57152 5102 57204 5108
rect 56508 5024 56560 5030
rect 56508 4966 56560 4972
rect 57060 5024 57112 5030
rect 57060 4966 57112 4972
rect 56232 3732 56284 3738
rect 56232 3674 56284 3680
rect 55680 3664 55732 3670
rect 55680 3606 55732 3612
rect 56140 3120 56192 3126
rect 56140 3062 56192 3068
rect 55128 2916 55180 2922
rect 55128 2858 55180 2864
rect 55588 2916 55640 2922
rect 55588 2858 55640 2864
rect 55140 2666 55168 2858
rect 54668 2644 54720 2650
rect 54668 2586 54720 2592
rect 54944 2644 54996 2650
rect 55140 2638 55260 2666
rect 54944 2586 54996 2592
rect 55232 898 55260 2638
rect 55956 2304 56008 2310
rect 55956 2246 56008 2252
rect 55968 1970 55996 2246
rect 55956 1964 56008 1970
rect 55956 1906 56008 1912
rect 55232 870 55352 898
rect 55324 800 55352 870
rect 56152 800 56180 3062
rect 56244 2990 56272 3674
rect 56520 3602 56548 4966
rect 57072 4826 57100 4966
rect 57348 4826 57376 5782
rect 57808 5778 57836 5850
rect 57796 5772 57848 5778
rect 57796 5714 57848 5720
rect 57992 5234 58020 5850
rect 58084 5778 58112 6174
rect 58072 5772 58124 5778
rect 58072 5714 58124 5720
rect 57980 5228 58032 5234
rect 57980 5170 58032 5176
rect 58084 4826 58112 5714
rect 58176 5710 58204 6344
rect 58268 6322 58296 6734
rect 58544 6730 58572 8366
rect 58716 7948 58768 7954
rect 58716 7890 58768 7896
rect 58728 7274 58756 7890
rect 58716 7268 58768 7274
rect 58716 7210 58768 7216
rect 58532 6724 58584 6730
rect 58532 6666 58584 6672
rect 58256 6316 58308 6322
rect 58256 6258 58308 6264
rect 58268 5778 58296 6258
rect 58348 6248 58400 6254
rect 58348 6190 58400 6196
rect 58360 5914 58388 6190
rect 58440 6112 58492 6118
rect 58544 6100 58572 6666
rect 58492 6072 58572 6100
rect 58440 6054 58492 6060
rect 58348 5908 58400 5914
rect 58348 5850 58400 5856
rect 58256 5772 58308 5778
rect 58256 5714 58308 5720
rect 58164 5704 58216 5710
rect 58164 5646 58216 5652
rect 57060 4820 57112 4826
rect 57336 4820 57388 4826
rect 57060 4762 57112 4768
rect 57256 4780 57336 4808
rect 57256 3602 57284 4780
rect 57336 4762 57388 4768
rect 58072 4820 58124 4826
rect 58072 4762 58124 4768
rect 58348 4684 58400 4690
rect 58348 4626 58400 4632
rect 58072 4072 58124 4078
rect 58072 4014 58124 4020
rect 57612 4004 57664 4010
rect 57612 3946 57664 3952
rect 57336 3936 57388 3942
rect 57336 3878 57388 3884
rect 57348 3670 57376 3878
rect 57336 3664 57388 3670
rect 57336 3606 57388 3612
rect 56508 3596 56560 3602
rect 56508 3538 56560 3544
rect 57244 3596 57296 3602
rect 57244 3538 57296 3544
rect 56322 3496 56378 3505
rect 56322 3431 56378 3440
rect 56336 3194 56364 3431
rect 56520 3194 56548 3538
rect 57060 3528 57112 3534
rect 57060 3470 57112 3476
rect 56324 3188 56376 3194
rect 56324 3130 56376 3136
rect 56508 3188 56560 3194
rect 56508 3130 56560 3136
rect 56232 2984 56284 2990
rect 56232 2926 56284 2932
rect 57072 800 57100 3470
rect 57256 3194 57284 3538
rect 57624 3194 57652 3946
rect 57980 3528 58032 3534
rect 57980 3470 58032 3476
rect 57992 3194 58020 3470
rect 57244 3188 57296 3194
rect 57244 3130 57296 3136
rect 57612 3188 57664 3194
rect 57612 3130 57664 3136
rect 57980 3188 58032 3194
rect 57980 3130 58032 3136
rect 57256 2650 57284 3130
rect 57888 3120 57940 3126
rect 57888 3062 57940 3068
rect 57244 2644 57296 2650
rect 57244 2586 57296 2592
rect 57900 800 57928 3062
rect 58084 2446 58112 4014
rect 58360 3602 58388 4626
rect 58452 4486 58480 6054
rect 58728 5914 58756 7210
rect 58820 6662 58848 10406
rect 59096 9994 59124 10406
rect 59084 9988 59136 9994
rect 59084 9930 59136 9936
rect 59452 9920 59504 9926
rect 59452 9862 59504 9868
rect 59268 9036 59320 9042
rect 59268 8978 59320 8984
rect 59084 8832 59136 8838
rect 59084 8774 59136 8780
rect 59096 8430 59124 8774
rect 59084 8424 59136 8430
rect 59084 8366 59136 8372
rect 59096 8022 59124 8366
rect 59280 8090 59308 8978
rect 59268 8084 59320 8090
rect 59268 8026 59320 8032
rect 59084 8016 59136 8022
rect 59084 7958 59136 7964
rect 59464 7818 59492 9862
rect 59452 7812 59504 7818
rect 59452 7754 59504 7760
rect 59636 7744 59688 7750
rect 59636 7686 59688 7692
rect 59648 7342 59676 7686
rect 59636 7336 59688 7342
rect 59636 7278 59688 7284
rect 59648 6866 59676 7278
rect 59740 6934 59768 11630
rect 60568 11558 60596 12242
rect 61108 11756 61160 11762
rect 61108 11698 61160 11704
rect 60832 11620 60884 11626
rect 60832 11562 60884 11568
rect 60556 11552 60608 11558
rect 60556 11494 60608 11500
rect 60464 11212 60516 11218
rect 60464 11154 60516 11160
rect 60476 10810 60504 11154
rect 60464 10804 60516 10810
rect 60464 10746 60516 10752
rect 60464 10056 60516 10062
rect 60464 9998 60516 10004
rect 59820 9920 59872 9926
rect 59820 9862 59872 9868
rect 59832 9382 59860 9862
rect 60476 9382 60504 9998
rect 60568 9518 60596 11494
rect 60844 10742 60872 11562
rect 61120 11558 61148 11698
rect 61108 11552 61160 11558
rect 61108 11494 61160 11500
rect 60832 10736 60884 10742
rect 60832 10678 60884 10684
rect 60556 9512 60608 9518
rect 60556 9454 60608 9460
rect 59820 9376 59872 9382
rect 59820 9318 59872 9324
rect 60464 9376 60516 9382
rect 60464 9318 60516 9324
rect 59832 8838 59860 9318
rect 60476 8906 60504 9318
rect 60648 9172 60700 9178
rect 60648 9114 60700 9120
rect 60464 8900 60516 8906
rect 60464 8842 60516 8848
rect 59820 8832 59872 8838
rect 59820 8774 59872 8780
rect 59832 8498 59860 8774
rect 59820 8492 59872 8498
rect 59820 8434 59872 8440
rect 60660 8430 60688 9114
rect 61120 8974 61148 11494
rect 61292 10464 61344 10470
rect 61292 10406 61344 10412
rect 61304 10130 61332 10406
rect 61844 10260 61896 10266
rect 61844 10202 61896 10208
rect 61292 10124 61344 10130
rect 61292 10066 61344 10072
rect 61304 9382 61332 10066
rect 61856 9926 61884 10202
rect 61844 9920 61896 9926
rect 61844 9862 61896 9868
rect 61292 9376 61344 9382
rect 61292 9318 61344 9324
rect 61108 8968 61160 8974
rect 61108 8910 61160 8916
rect 61120 8566 61148 8910
rect 61304 8566 61332 9318
rect 61856 9042 61884 9862
rect 61844 9036 61896 9042
rect 61844 8978 61896 8984
rect 61384 8968 61436 8974
rect 61384 8910 61436 8916
rect 61108 8560 61160 8566
rect 61108 8502 61160 8508
rect 61292 8560 61344 8566
rect 61292 8502 61344 8508
rect 60648 8424 60700 8430
rect 60648 8366 60700 8372
rect 60924 8288 60976 8294
rect 60924 8230 60976 8236
rect 60936 7954 60964 8230
rect 60924 7948 60976 7954
rect 60924 7890 60976 7896
rect 60936 7546 60964 7890
rect 59912 7540 59964 7546
rect 59912 7482 59964 7488
rect 60924 7540 60976 7546
rect 60924 7482 60976 7488
rect 59820 7336 59872 7342
rect 59820 7278 59872 7284
rect 59728 6928 59780 6934
rect 59728 6870 59780 6876
rect 59636 6860 59688 6866
rect 59636 6802 59688 6808
rect 59832 6746 59860 7278
rect 59924 6866 59952 7482
rect 59912 6860 59964 6866
rect 59912 6802 59964 6808
rect 60648 6860 60700 6866
rect 60648 6802 60700 6808
rect 59648 6718 59860 6746
rect 60004 6792 60056 6798
rect 60004 6734 60056 6740
rect 58808 6656 58860 6662
rect 58808 6598 58860 6604
rect 58716 5908 58768 5914
rect 58716 5850 58768 5856
rect 58900 5772 58952 5778
rect 58900 5714 58952 5720
rect 58912 5370 58940 5714
rect 59648 5642 59676 6718
rect 60016 6118 60044 6734
rect 60660 6254 60688 6802
rect 61304 6798 61332 8502
rect 61292 6792 61344 6798
rect 61292 6734 61344 6740
rect 60648 6248 60700 6254
rect 60648 6190 60700 6196
rect 60004 6112 60056 6118
rect 60004 6054 60056 6060
rect 60280 6112 60332 6118
rect 60280 6054 60332 6060
rect 60016 5953 60044 6054
rect 60002 5944 60058 5953
rect 60002 5879 60058 5888
rect 59636 5636 59688 5642
rect 59636 5578 59688 5584
rect 59268 5568 59320 5574
rect 59268 5510 59320 5516
rect 58900 5364 58952 5370
rect 58900 5306 58952 5312
rect 58624 5160 58676 5166
rect 58624 5102 58676 5108
rect 58440 4480 58492 4486
rect 58440 4422 58492 4428
rect 58452 4078 58480 4422
rect 58440 4072 58492 4078
rect 58440 4014 58492 4020
rect 58636 3618 58664 5102
rect 58912 4622 58940 5306
rect 59280 5166 59308 5510
rect 59084 5160 59136 5166
rect 59084 5102 59136 5108
rect 59268 5160 59320 5166
rect 59268 5102 59320 5108
rect 59096 4690 59124 5102
rect 59084 4684 59136 4690
rect 59084 4626 59136 4632
rect 59280 4622 59308 5102
rect 58900 4616 58952 4622
rect 58900 4558 58952 4564
rect 59268 4616 59320 4622
rect 59268 4558 59320 4564
rect 59360 4616 59412 4622
rect 59360 4558 59412 4564
rect 59280 4282 59308 4558
rect 59268 4276 59320 4282
rect 59268 4218 59320 4224
rect 58636 3602 58756 3618
rect 58348 3596 58400 3602
rect 58348 3538 58400 3544
rect 58532 3596 58584 3602
rect 58532 3538 58584 3544
rect 58636 3596 58768 3602
rect 58636 3590 58716 3596
rect 58544 3398 58572 3538
rect 58532 3392 58584 3398
rect 58532 3334 58584 3340
rect 58544 2650 58572 3334
rect 58636 3194 58664 3590
rect 58716 3538 58768 3544
rect 59372 3534 59400 4558
rect 59452 4548 59504 4554
rect 59452 4490 59504 4496
rect 59464 3602 59492 4490
rect 59544 4480 59596 4486
rect 59544 4422 59596 4428
rect 59556 4146 59584 4422
rect 59544 4140 59596 4146
rect 59544 4082 59596 4088
rect 59452 3596 59504 3602
rect 59452 3538 59504 3544
rect 59360 3528 59412 3534
rect 59360 3470 59412 3476
rect 59556 3194 59584 4082
rect 59648 3602 59676 5578
rect 59728 5568 59780 5574
rect 59728 5510 59780 5516
rect 59740 5166 59768 5510
rect 59728 5160 59780 5166
rect 59728 5102 59780 5108
rect 59820 5160 59872 5166
rect 59820 5102 59872 5108
rect 59832 4758 59860 5102
rect 60004 5024 60056 5030
rect 60004 4966 60056 4972
rect 59820 4752 59872 4758
rect 59820 4694 59872 4700
rect 60016 3754 60044 4966
rect 59924 3738 60044 3754
rect 59912 3732 60044 3738
rect 59964 3726 60044 3732
rect 59912 3674 59964 3680
rect 59636 3596 59688 3602
rect 59636 3538 59688 3544
rect 59820 3528 59872 3534
rect 59820 3470 59872 3476
rect 59832 3398 59860 3470
rect 59820 3392 59872 3398
rect 59820 3334 59872 3340
rect 58624 3188 58676 3194
rect 58624 3130 58676 3136
rect 59544 3188 59596 3194
rect 59544 3130 59596 3136
rect 59832 2990 59860 3334
rect 60016 2990 60044 3726
rect 60292 3602 60320 6054
rect 61304 5778 61332 6734
rect 61396 6322 61424 8910
rect 61856 8634 61884 8978
rect 61844 8628 61896 8634
rect 61844 8570 61896 8576
rect 61568 6792 61620 6798
rect 61568 6734 61620 6740
rect 61384 6316 61436 6322
rect 61384 6258 61436 6264
rect 61580 6118 61608 6734
rect 61568 6112 61620 6118
rect 61568 6054 61620 6060
rect 61292 5772 61344 5778
rect 61292 5714 61344 5720
rect 60464 5704 60516 5710
rect 60464 5646 60516 5652
rect 60476 5030 60504 5646
rect 61304 5370 61332 5714
rect 61292 5364 61344 5370
rect 61292 5306 61344 5312
rect 61016 5160 61068 5166
rect 61016 5102 61068 5108
rect 61028 5030 61056 5102
rect 61200 5092 61252 5098
rect 61200 5034 61252 5040
rect 60464 5024 60516 5030
rect 60464 4966 60516 4972
rect 61016 5024 61068 5030
rect 61016 4966 61068 4972
rect 60476 3670 60504 4966
rect 61028 4690 61056 4966
rect 61212 4690 61240 5034
rect 61580 4826 61608 6054
rect 61752 5568 61804 5574
rect 61752 5510 61804 5516
rect 61568 4820 61620 4826
rect 61568 4762 61620 4768
rect 61016 4684 61068 4690
rect 61016 4626 61068 4632
rect 61200 4684 61252 4690
rect 61200 4626 61252 4632
rect 61028 4146 61056 4626
rect 61212 4282 61240 4626
rect 61764 4622 61792 5510
rect 61752 4616 61804 4622
rect 61752 4558 61804 4564
rect 61476 4480 61528 4486
rect 61476 4422 61528 4428
rect 61200 4276 61252 4282
rect 61200 4218 61252 4224
rect 61016 4140 61068 4146
rect 61016 4082 61068 4088
rect 61488 4078 61516 4422
rect 61764 4146 61792 4558
rect 61752 4140 61804 4146
rect 61752 4082 61804 4088
rect 61476 4072 61528 4078
rect 61476 4014 61528 4020
rect 60464 3664 60516 3670
rect 60464 3606 60516 3612
rect 60280 3596 60332 3602
rect 60280 3538 60332 3544
rect 59820 2984 59872 2990
rect 59820 2926 59872 2932
rect 60004 2984 60056 2990
rect 60292 2961 60320 3538
rect 62304 3528 62356 3534
rect 62304 3470 62356 3476
rect 61292 3460 61344 3466
rect 61292 3402 61344 3408
rect 60556 3392 60608 3398
rect 60556 3334 60608 3340
rect 60568 3194 60596 3334
rect 61304 3194 61332 3402
rect 62212 3392 62264 3398
rect 62212 3334 62264 3340
rect 60556 3188 60608 3194
rect 60556 3130 60608 3136
rect 61292 3188 61344 3194
rect 61292 3130 61344 3136
rect 60004 2926 60056 2932
rect 60278 2952 60334 2961
rect 60278 2887 60280 2896
rect 60332 2887 60334 2896
rect 60280 2858 60332 2864
rect 59452 2848 59504 2854
rect 59452 2790 59504 2796
rect 58532 2644 58584 2650
rect 58532 2586 58584 2592
rect 59464 2582 59492 2790
rect 59452 2576 59504 2582
rect 59452 2518 59504 2524
rect 58072 2440 58124 2446
rect 58072 2382 58124 2388
rect 58808 2440 58860 2446
rect 58808 2382 58860 2388
rect 58820 800 58848 2382
rect 59728 2304 59780 2310
rect 59728 2246 59780 2252
rect 59912 2304 59964 2310
rect 59912 2246 59964 2252
rect 59740 800 59768 2246
rect 59924 2106 59952 2246
rect 59912 2100 59964 2106
rect 59912 2042 59964 2048
rect 60568 800 60596 3130
rect 62224 3126 62252 3334
rect 62316 3194 62344 3470
rect 62304 3188 62356 3194
rect 62304 3130 62356 3136
rect 60832 3120 60884 3126
rect 62212 3120 62264 3126
rect 60884 3068 61240 3074
rect 60832 3062 61240 3068
rect 62212 3062 62264 3068
rect 60844 3058 61240 3062
rect 60844 3052 61252 3058
rect 60844 3046 61200 3052
rect 61200 2994 61252 3000
rect 61212 2854 61240 2994
rect 61200 2848 61252 2854
rect 61200 2790 61252 2796
rect 62224 2650 62252 3062
rect 64144 2984 64196 2990
rect 64144 2926 64196 2932
rect 63224 2916 63276 2922
rect 63224 2858 63276 2864
rect 62212 2644 62264 2650
rect 62212 2586 62264 2592
rect 61476 2508 61528 2514
rect 61476 2450 61528 2456
rect 62396 2508 62448 2514
rect 62396 2450 62448 2456
rect 61488 2310 61516 2450
rect 62408 2310 62436 2450
rect 61476 2304 61528 2310
rect 61476 2246 61528 2252
rect 62396 2304 62448 2310
rect 62396 2246 62448 2252
rect 61488 800 61516 2246
rect 62408 800 62436 2246
rect 63236 800 63264 2858
rect 64156 800 64184 2926
rect 386 0 442 800
rect 1214 0 1270 800
rect 2134 0 2190 800
rect 2962 0 3018 800
rect 3882 0 3938 800
rect 4802 0 4858 800
rect 5630 0 5686 800
rect 6550 0 6606 800
rect 7470 0 7526 800
rect 8298 0 8354 800
rect 9218 0 9274 800
rect 10046 0 10102 800
rect 10966 0 11022 800
rect 11886 0 11942 800
rect 12714 0 12770 800
rect 13634 0 13690 800
rect 14554 0 14610 800
rect 15382 0 15438 800
rect 16302 0 16358 800
rect 17130 0 17186 800
rect 18050 0 18106 800
rect 18970 0 19026 800
rect 19798 0 19854 800
rect 20718 0 20774 800
rect 21638 0 21694 800
rect 22466 0 22522 800
rect 23386 0 23442 800
rect 24306 0 24362 800
rect 25134 0 25190 800
rect 26054 0 26110 800
rect 26882 0 26938 800
rect 27802 0 27858 800
rect 28722 0 28778 800
rect 29550 0 29606 800
rect 30470 0 30526 800
rect 31390 0 31446 800
rect 32218 0 32274 800
rect 33138 0 33194 800
rect 33966 0 34022 800
rect 34886 0 34942 800
rect 35806 0 35862 800
rect 36634 0 36690 800
rect 37554 0 37610 800
rect 38474 0 38530 800
rect 39302 0 39358 800
rect 40222 0 40278 800
rect 41050 0 41106 800
rect 41970 0 42026 800
rect 42890 0 42946 800
rect 43718 0 43774 800
rect 44638 0 44694 800
rect 45558 0 45614 800
rect 46386 0 46442 800
rect 47306 0 47362 800
rect 48226 0 48282 800
rect 49054 0 49110 800
rect 49974 0 50030 800
rect 50802 0 50858 800
rect 51722 0 51778 800
rect 52642 0 52698 800
rect 53470 0 53526 800
rect 54390 0 54446 800
rect 55310 0 55366 800
rect 56138 0 56194 800
rect 57058 0 57114 800
rect 57886 0 57942 800
rect 58806 0 58862 800
rect 59726 0 59782 800
rect 60554 0 60610 800
rect 61474 0 61530 800
rect 62394 0 62450 800
rect 63222 0 63278 800
rect 64142 0 64198 800
<< via2 >>
rect 3974 18808 4030 18864
rect 3146 14456 3202 14512
rect 386 3032 442 3088
rect 2778 4936 2834 4992
rect 4066 16632 4122 16688
rect 3974 13232 4030 13288
rect 4066 12144 4122 12200
rect 3974 10648 4030 10704
rect 3882 9968 3938 10024
rect 3882 7792 3938 7848
rect 3422 3712 3478 3768
rect 3698 2760 3754 2816
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11378 17434
rect 11378 17382 11408 17434
rect 11432 17382 11442 17434
rect 11442 17382 11488 17434
rect 11512 17382 11558 17434
rect 11558 17382 11568 17434
rect 11592 17382 11622 17434
rect 11622 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11378 16346
rect 11378 16294 11408 16346
rect 11432 16294 11442 16346
rect 11442 16294 11488 16346
rect 11512 16294 11558 16346
rect 11558 16294 11568 16346
rect 11592 16294 11622 16346
rect 11622 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11378 15258
rect 11378 15206 11408 15258
rect 11432 15206 11442 15258
rect 11442 15206 11488 15258
rect 11512 15206 11558 15258
rect 11558 15206 11568 15258
rect 11592 15206 11622 15258
rect 11622 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 6642 8356 6698 8392
rect 6642 8336 6644 8356
rect 6644 8336 6696 8356
rect 6696 8336 6698 8356
rect 6274 7404 6330 7440
rect 6274 7384 6276 7404
rect 6276 7384 6328 7404
rect 6328 7384 6330 7404
rect 4066 5480 4122 5536
rect 4526 4684 4582 4720
rect 4526 4664 4528 4684
rect 4528 4664 4580 4684
rect 4580 4664 4582 4684
rect 4066 4020 4068 4040
rect 4068 4020 4120 4040
rect 4120 4020 4122 4040
rect 4066 3984 4122 4020
rect 4802 3576 4858 3632
rect 4066 1128 4122 1184
rect 5814 4972 5816 4992
rect 5816 4972 5868 4992
rect 5868 4972 5870 4992
rect 5814 4936 5870 4972
rect 9402 13504 9458 13560
rect 9310 12280 9366 12336
rect 9862 13504 9918 13560
rect 9586 12824 9642 12880
rect 9494 12588 9496 12608
rect 9496 12588 9548 12608
rect 9548 12588 9550 12608
rect 9494 12552 9550 12588
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11378 14170
rect 11378 14118 11408 14170
rect 11432 14118 11442 14170
rect 11442 14118 11488 14170
rect 11512 14118 11558 14170
rect 11558 14118 11568 14170
rect 11592 14118 11622 14170
rect 11622 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 8482 10648 8538 10704
rect 7562 7948 7618 7984
rect 7562 7928 7564 7948
rect 7564 7928 7616 7948
rect 7616 7928 7618 7948
rect 8298 5092 8354 5128
rect 8298 5072 8300 5092
rect 8300 5072 8352 5092
rect 8352 5072 8354 5092
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11378 13082
rect 11378 13030 11408 13082
rect 11432 13030 11442 13082
rect 11442 13030 11488 13082
rect 11512 13030 11558 13082
rect 11558 13030 11568 13082
rect 11592 13030 11622 13082
rect 11622 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 12622 13640 12678 13696
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11378 11994
rect 11378 11942 11408 11994
rect 11432 11942 11442 11994
rect 11442 11942 11488 11994
rect 11512 11942 11558 11994
rect 11558 11942 11568 11994
rect 11592 11942 11622 11994
rect 11622 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11378 10906
rect 11378 10854 11408 10906
rect 11432 10854 11442 10906
rect 11442 10854 11488 10906
rect 11512 10854 11558 10906
rect 11558 10854 11568 10906
rect 11592 10854 11622 10906
rect 11622 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11378 9818
rect 11378 9766 11408 9818
rect 11432 9766 11442 9818
rect 11442 9766 11488 9818
rect 11512 9766 11558 9818
rect 11558 9766 11568 9818
rect 11592 9766 11622 9818
rect 11622 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 8942 4936 8998 4992
rect 7838 2932 7840 2952
rect 7840 2932 7892 2952
rect 7892 2932 7894 2952
rect 7838 2896 7894 2932
rect 10138 4800 10194 4856
rect 11150 8900 11206 8936
rect 11150 8880 11152 8900
rect 11152 8880 11204 8900
rect 11204 8880 11206 8900
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11378 8730
rect 11378 8678 11408 8730
rect 11432 8678 11442 8730
rect 11442 8678 11488 8730
rect 11512 8678 11558 8730
rect 11558 8678 11568 8730
rect 11592 8678 11622 8730
rect 11622 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11886 8628 11942 8664
rect 11886 8608 11888 8628
rect 11888 8608 11940 8628
rect 11940 8608 11942 8628
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11378 7642
rect 11378 7590 11408 7642
rect 11432 7590 11442 7642
rect 11442 7590 11488 7642
rect 11512 7590 11558 7642
rect 11558 7590 11568 7642
rect 11592 7590 11622 7642
rect 11622 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11886 7520 11942 7576
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11378 6554
rect 11378 6502 11408 6554
rect 11432 6502 11442 6554
rect 11442 6502 11488 6554
rect 11512 6502 11558 6554
rect 11558 6502 11568 6554
rect 11592 6502 11622 6554
rect 11622 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 10966 6024 11022 6080
rect 13082 13388 13138 13424
rect 13082 13368 13084 13388
rect 13084 13368 13136 13388
rect 13136 13368 13138 13388
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11378 5466
rect 11378 5414 11408 5466
rect 11432 5414 11442 5466
rect 11442 5414 11488 5466
rect 11512 5414 11558 5466
rect 11558 5414 11568 5466
rect 11592 5414 11622 5466
rect 11622 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11886 5072 11942 5128
rect 10690 2624 10746 2680
rect 12162 5072 12218 5128
rect 11150 4120 11206 4176
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11378 4378
rect 11378 4326 11408 4378
rect 11432 4326 11442 4378
rect 11442 4326 11488 4378
rect 11512 4326 11558 4378
rect 11558 4326 11568 4378
rect 11592 4326 11622 4378
rect 11622 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 13726 11736 13782 11792
rect 11610 3460 11666 3496
rect 11610 3440 11612 3460
rect 11612 3440 11664 3460
rect 11664 3440 11666 3460
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11378 3290
rect 11378 3238 11408 3290
rect 11432 3238 11442 3290
rect 11442 3238 11488 3290
rect 11512 3238 11558 3290
rect 11558 3238 11568 3290
rect 11592 3238 11622 3290
rect 11622 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 11150 2932 11152 2952
rect 11152 2932 11204 2952
rect 11204 2932 11206 2952
rect 11150 2896 11206 2932
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11378 2202
rect 11378 2150 11408 2202
rect 11432 2150 11442 2202
rect 11442 2150 11488 2202
rect 11512 2150 11558 2202
rect 11558 2150 11568 2202
rect 11592 2150 11622 2202
rect 11622 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 12254 4276 12310 4312
rect 12254 4256 12256 4276
rect 12256 4256 12308 4276
rect 12308 4256 12310 4276
rect 12438 4120 12494 4176
rect 12898 3168 12954 3224
rect 12990 2760 13046 2816
rect 16026 12688 16082 12744
rect 13450 6160 13506 6216
rect 15290 7656 15346 7712
rect 13542 4120 13598 4176
rect 13358 3712 13414 3768
rect 13818 3340 13820 3360
rect 13820 3340 13872 3360
rect 13872 3340 13874 3360
rect 13818 3304 13874 3340
rect 14830 3848 14886 3904
rect 17038 13932 17094 13968
rect 17222 14048 17278 14104
rect 17038 13912 17040 13932
rect 17040 13912 17092 13932
rect 17092 13912 17094 13932
rect 17222 13504 17278 13560
rect 17222 13096 17278 13152
rect 16854 12300 16910 12336
rect 16854 12280 16856 12300
rect 16856 12280 16908 12300
rect 16908 12280 16910 12300
rect 16302 9560 16358 9616
rect 17314 12144 17370 12200
rect 17774 12436 17830 12472
rect 17774 12416 17776 12436
rect 17776 12416 17828 12436
rect 17828 12416 17830 12436
rect 18326 11872 18382 11928
rect 15658 5344 15714 5400
rect 15474 4528 15530 4584
rect 16210 5480 16266 5536
rect 17498 8916 17500 8936
rect 17500 8916 17552 8936
rect 17552 8916 17554 8936
rect 17498 8880 17554 8916
rect 17222 8472 17278 8528
rect 16854 7656 16910 7712
rect 16946 7520 17002 7576
rect 16762 6432 16818 6488
rect 16578 4800 16634 4856
rect 16486 3884 16488 3904
rect 16488 3884 16540 3904
rect 16540 3884 16542 3904
rect 16486 3848 16542 3884
rect 15934 2932 15936 2952
rect 15936 2932 15988 2952
rect 15988 2932 15990 2952
rect 15934 2896 15990 2932
rect 17498 7656 17554 7712
rect 17774 8472 17830 8528
rect 19430 12980 19486 13016
rect 19430 12960 19432 12980
rect 19432 12960 19484 12980
rect 19484 12960 19486 12980
rect 21748 16890 21804 16892
rect 21828 16890 21884 16892
rect 21908 16890 21964 16892
rect 21988 16890 22044 16892
rect 21748 16838 21774 16890
rect 21774 16838 21804 16890
rect 21828 16838 21838 16890
rect 21838 16838 21884 16890
rect 21908 16838 21954 16890
rect 21954 16838 21964 16890
rect 21988 16838 22018 16890
rect 22018 16838 22044 16890
rect 21748 16836 21804 16838
rect 21828 16836 21884 16838
rect 21908 16836 21964 16838
rect 21988 16836 22044 16838
rect 21748 15802 21804 15804
rect 21828 15802 21884 15804
rect 21908 15802 21964 15804
rect 21988 15802 22044 15804
rect 21748 15750 21774 15802
rect 21774 15750 21804 15802
rect 21828 15750 21838 15802
rect 21838 15750 21884 15802
rect 21908 15750 21954 15802
rect 21954 15750 21964 15802
rect 21988 15750 22018 15802
rect 22018 15750 22044 15802
rect 21748 15748 21804 15750
rect 21828 15748 21884 15750
rect 21908 15748 21964 15750
rect 21988 15748 22044 15750
rect 19982 14900 19984 14920
rect 19984 14900 20036 14920
rect 20036 14900 20038 14920
rect 19982 14864 20038 14900
rect 18878 12008 18934 12064
rect 18694 8608 18750 8664
rect 19246 9580 19302 9616
rect 19246 9560 19248 9580
rect 19248 9560 19300 9580
rect 19300 9560 19302 9580
rect 20074 10512 20130 10568
rect 19798 7520 19854 7576
rect 17774 3304 17830 3360
rect 17774 2896 17830 2952
rect 18786 4120 18842 4176
rect 19338 6724 19394 6760
rect 19338 6704 19340 6724
rect 19340 6704 19392 6724
rect 19392 6704 19394 6724
rect 19246 6024 19302 6080
rect 19154 5072 19210 5128
rect 18970 4120 19026 4176
rect 18970 3168 19026 3224
rect 19246 3168 19302 3224
rect 19062 2624 19118 2680
rect 20258 12960 20314 13016
rect 20442 12960 20498 13016
rect 20810 14456 20866 14512
rect 21914 15000 21970 15056
rect 22466 15000 22522 15056
rect 21748 14714 21804 14716
rect 21828 14714 21884 14716
rect 21908 14714 21964 14716
rect 21988 14714 22044 14716
rect 21748 14662 21774 14714
rect 21774 14662 21804 14714
rect 21828 14662 21838 14714
rect 21838 14662 21884 14714
rect 21908 14662 21954 14714
rect 21954 14662 21964 14714
rect 21988 14662 22018 14714
rect 22018 14662 22044 14714
rect 21748 14660 21804 14662
rect 21828 14660 21884 14662
rect 21908 14660 21964 14662
rect 21988 14660 22044 14662
rect 21546 14356 21548 14376
rect 21548 14356 21600 14376
rect 21600 14356 21602 14376
rect 21546 14320 21602 14356
rect 20626 12416 20682 12472
rect 21178 13912 21234 13968
rect 20994 10104 21050 10160
rect 21178 11600 21234 11656
rect 21086 9696 21142 9752
rect 22098 14184 22154 14240
rect 21748 13626 21804 13628
rect 21828 13626 21884 13628
rect 21908 13626 21964 13628
rect 21988 13626 22044 13628
rect 21748 13574 21774 13626
rect 21774 13574 21804 13626
rect 21828 13574 21838 13626
rect 21838 13574 21884 13626
rect 21908 13574 21954 13626
rect 21954 13574 21964 13626
rect 21988 13574 22018 13626
rect 22018 13574 22044 13626
rect 21748 13572 21804 13574
rect 21828 13572 21884 13574
rect 21908 13572 21964 13574
rect 21988 13572 22044 13574
rect 23662 14900 23664 14920
rect 23664 14900 23716 14920
rect 23716 14900 23718 14920
rect 23662 14864 23718 14900
rect 24674 14320 24730 14376
rect 21748 12538 21804 12540
rect 21828 12538 21884 12540
rect 21908 12538 21964 12540
rect 21988 12538 22044 12540
rect 21748 12486 21774 12538
rect 21774 12486 21804 12538
rect 21828 12486 21838 12538
rect 21838 12486 21884 12538
rect 21908 12486 21954 12538
rect 21954 12486 21964 12538
rect 21988 12486 22018 12538
rect 22018 12486 22044 12538
rect 21748 12484 21804 12486
rect 21828 12484 21884 12486
rect 21908 12484 21964 12486
rect 21988 12484 22044 12486
rect 21730 11600 21786 11656
rect 21748 11450 21804 11452
rect 21828 11450 21884 11452
rect 21908 11450 21964 11452
rect 21988 11450 22044 11452
rect 21748 11398 21774 11450
rect 21774 11398 21804 11450
rect 21828 11398 21838 11450
rect 21838 11398 21884 11450
rect 21908 11398 21954 11450
rect 21954 11398 21964 11450
rect 21988 11398 22018 11450
rect 22018 11398 22044 11450
rect 21748 11396 21804 11398
rect 21828 11396 21884 11398
rect 21908 11396 21964 11398
rect 21988 11396 22044 11398
rect 22282 10512 22338 10568
rect 21748 10362 21804 10364
rect 21828 10362 21884 10364
rect 21908 10362 21964 10364
rect 21988 10362 22044 10364
rect 21748 10310 21774 10362
rect 21774 10310 21804 10362
rect 21828 10310 21838 10362
rect 21838 10310 21884 10362
rect 21908 10310 21954 10362
rect 21954 10310 21964 10362
rect 21988 10310 22018 10362
rect 22018 10310 22044 10362
rect 21748 10308 21804 10310
rect 21828 10308 21884 10310
rect 21908 10308 21964 10310
rect 21988 10308 22044 10310
rect 21730 9560 21786 9616
rect 21638 9424 21694 9480
rect 21748 9274 21804 9276
rect 21828 9274 21884 9276
rect 21908 9274 21964 9276
rect 21988 9274 22044 9276
rect 21748 9222 21774 9274
rect 21774 9222 21804 9274
rect 21828 9222 21838 9274
rect 21838 9222 21884 9274
rect 21908 9222 21954 9274
rect 21954 9222 21964 9274
rect 21988 9222 22018 9274
rect 22018 9222 22044 9274
rect 21748 9220 21804 9222
rect 21828 9220 21884 9222
rect 21908 9220 21964 9222
rect 21988 9220 22044 9222
rect 21086 8880 21142 8936
rect 20166 7656 20222 7712
rect 19890 6296 19946 6352
rect 19430 4392 19486 4448
rect 19706 4800 19762 4856
rect 20166 5616 20222 5672
rect 21270 5788 21272 5808
rect 21272 5788 21324 5808
rect 21324 5788 21326 5808
rect 21270 5752 21326 5788
rect 21178 5344 21234 5400
rect 20442 5072 20498 5128
rect 20534 3848 20590 3904
rect 20350 2896 20406 2952
rect 20810 3848 20866 3904
rect 21086 4140 21142 4176
rect 21086 4120 21088 4140
rect 21088 4120 21140 4140
rect 21140 4120 21142 4140
rect 22006 8744 22062 8800
rect 21730 8472 21786 8528
rect 22834 13096 22890 13152
rect 22742 12416 22798 12472
rect 23478 12144 23534 12200
rect 23202 11600 23258 11656
rect 22926 11192 22982 11248
rect 24122 14184 24178 14240
rect 23662 12008 23718 12064
rect 24122 11056 24178 11112
rect 23478 10684 23480 10704
rect 23480 10684 23532 10704
rect 23532 10684 23534 10704
rect 23478 10648 23534 10684
rect 23386 9696 23442 9752
rect 23294 9560 23350 9616
rect 22558 8744 22614 8800
rect 21748 8186 21804 8188
rect 21828 8186 21884 8188
rect 21908 8186 21964 8188
rect 21988 8186 22044 8188
rect 21748 8134 21774 8186
rect 21774 8134 21804 8186
rect 21828 8134 21838 8186
rect 21838 8134 21884 8186
rect 21908 8134 21954 8186
rect 21954 8134 21964 8186
rect 21988 8134 22018 8186
rect 22018 8134 22044 8186
rect 21748 8132 21804 8134
rect 21828 8132 21884 8134
rect 21908 8132 21964 8134
rect 21988 8132 22044 8134
rect 22098 7656 22154 7712
rect 21748 7098 21804 7100
rect 21828 7098 21884 7100
rect 21908 7098 21964 7100
rect 21988 7098 22044 7100
rect 21748 7046 21774 7098
rect 21774 7046 21804 7098
rect 21828 7046 21838 7098
rect 21838 7046 21884 7098
rect 21908 7046 21954 7098
rect 21954 7046 21964 7098
rect 21988 7046 22018 7098
rect 22018 7046 22044 7098
rect 21748 7044 21804 7046
rect 21828 7044 21884 7046
rect 21908 7044 21964 7046
rect 21988 7044 22044 7046
rect 21822 6740 21824 6760
rect 21824 6740 21876 6760
rect 21876 6740 21878 6760
rect 21822 6704 21878 6740
rect 21748 6010 21804 6012
rect 21828 6010 21884 6012
rect 21908 6010 21964 6012
rect 21988 6010 22044 6012
rect 21748 5958 21774 6010
rect 21774 5958 21804 6010
rect 21828 5958 21838 6010
rect 21838 5958 21884 6010
rect 21908 5958 21954 6010
rect 21954 5958 21964 6010
rect 21988 5958 22018 6010
rect 22018 5958 22044 6010
rect 21748 5956 21804 5958
rect 21828 5956 21884 5958
rect 21908 5956 21964 5958
rect 21988 5956 22044 5958
rect 21914 5344 21970 5400
rect 22190 5364 22246 5400
rect 22190 5344 22192 5364
rect 22192 5344 22244 5364
rect 22244 5344 22246 5364
rect 22558 6860 22614 6896
rect 22558 6840 22560 6860
rect 22560 6840 22612 6860
rect 22612 6840 22614 6860
rect 22374 5344 22430 5400
rect 21748 4922 21804 4924
rect 21828 4922 21884 4924
rect 21908 4922 21964 4924
rect 21988 4922 22044 4924
rect 21748 4870 21774 4922
rect 21774 4870 21804 4922
rect 21828 4870 21838 4922
rect 21838 4870 21884 4922
rect 21908 4870 21954 4922
rect 21954 4870 21964 4922
rect 21988 4870 22018 4922
rect 22018 4870 22044 4922
rect 21748 4868 21804 4870
rect 21828 4868 21884 4870
rect 21908 4868 21964 4870
rect 21988 4868 22044 4870
rect 22006 4140 22062 4176
rect 22006 4120 22008 4140
rect 22008 4120 22060 4140
rect 22060 4120 22062 4140
rect 21748 3834 21804 3836
rect 21828 3834 21884 3836
rect 21908 3834 21964 3836
rect 21988 3834 22044 3836
rect 21748 3782 21774 3834
rect 21774 3782 21804 3834
rect 21828 3782 21838 3834
rect 21838 3782 21884 3834
rect 21908 3782 21954 3834
rect 21954 3782 21964 3834
rect 21988 3782 22018 3834
rect 22018 3782 22044 3834
rect 21748 3780 21804 3782
rect 21828 3780 21884 3782
rect 21908 3780 21964 3782
rect 21988 3780 22044 3782
rect 22190 3848 22246 3904
rect 21748 2746 21804 2748
rect 21828 2746 21884 2748
rect 21908 2746 21964 2748
rect 21988 2746 22044 2748
rect 21748 2694 21774 2746
rect 21774 2694 21804 2746
rect 21828 2694 21838 2746
rect 21838 2694 21884 2746
rect 21908 2694 21954 2746
rect 21954 2694 21964 2746
rect 21988 2694 22018 2746
rect 22018 2694 22044 2746
rect 21748 2692 21804 2694
rect 21828 2692 21884 2694
rect 21908 2692 21964 2694
rect 21988 2692 22044 2694
rect 25318 12552 25374 12608
rect 26238 14048 26294 14104
rect 26238 12960 26294 13016
rect 24950 9560 25006 9616
rect 24122 9424 24178 9480
rect 23110 6024 23166 6080
rect 22926 3848 22982 3904
rect 23202 5652 23204 5672
rect 23204 5652 23256 5672
rect 23256 5652 23258 5672
rect 23202 5616 23258 5652
rect 24766 8472 24822 8528
rect 24950 8236 24952 8256
rect 24952 8236 25004 8256
rect 25004 8236 25006 8256
rect 24950 8200 25006 8236
rect 23938 5616 23994 5672
rect 25042 7656 25098 7712
rect 24214 5888 24270 5944
rect 23386 3884 23388 3904
rect 23388 3884 23440 3904
rect 23440 3884 23442 3904
rect 23386 3848 23442 3884
rect 23570 3848 23626 3904
rect 22834 3168 22890 3224
rect 22558 2932 22560 2952
rect 22560 2932 22612 2952
rect 22612 2932 22614 2952
rect 22558 2896 22614 2932
rect 23754 4392 23810 4448
rect 23386 3476 23388 3496
rect 23388 3476 23440 3496
rect 23440 3476 23442 3496
rect 23386 3440 23442 3476
rect 24398 6024 24454 6080
rect 24490 5072 24546 5128
rect 24674 5072 24730 5128
rect 24950 4664 25006 4720
rect 24674 3440 24730 3496
rect 24674 3032 24730 3088
rect 24398 2896 24454 2952
rect 25962 12552 26018 12608
rect 26790 13096 26846 13152
rect 26790 12824 26846 12880
rect 27158 11056 27214 11112
rect 27250 10648 27306 10704
rect 25778 6976 25834 7032
rect 25594 6296 25650 6352
rect 25502 4800 25558 4856
rect 25134 3032 25190 3088
rect 25318 3596 25374 3632
rect 25318 3576 25320 3596
rect 25320 3576 25372 3596
rect 25372 3576 25374 3596
rect 26330 7112 26386 7168
rect 26422 6976 26478 7032
rect 25870 4800 25926 4856
rect 25870 4120 25926 4176
rect 25686 3304 25742 3360
rect 27434 11872 27490 11928
rect 27802 11192 27858 11248
rect 32144 17434 32200 17436
rect 32224 17434 32280 17436
rect 32304 17434 32360 17436
rect 32384 17434 32440 17436
rect 32144 17382 32170 17434
rect 32170 17382 32200 17434
rect 32224 17382 32234 17434
rect 32234 17382 32280 17434
rect 32304 17382 32350 17434
rect 32350 17382 32360 17434
rect 32384 17382 32414 17434
rect 32414 17382 32440 17434
rect 32144 17380 32200 17382
rect 32224 17380 32280 17382
rect 32304 17380 32360 17382
rect 32384 17380 32440 17382
rect 27710 10104 27766 10160
rect 26882 7112 26938 7168
rect 26698 5652 26700 5672
rect 26700 5652 26752 5672
rect 26752 5652 26754 5672
rect 26698 5616 26754 5652
rect 28354 14456 28410 14512
rect 29090 13776 29146 13832
rect 28354 12960 28410 13016
rect 28262 11600 28318 11656
rect 28538 8880 28594 8936
rect 28722 12416 28778 12472
rect 32144 16346 32200 16348
rect 32224 16346 32280 16348
rect 32304 16346 32360 16348
rect 32384 16346 32440 16348
rect 32144 16294 32170 16346
rect 32170 16294 32200 16346
rect 32224 16294 32234 16346
rect 32234 16294 32280 16346
rect 32304 16294 32350 16346
rect 32350 16294 32360 16346
rect 32384 16294 32414 16346
rect 32414 16294 32440 16346
rect 32144 16292 32200 16294
rect 32224 16292 32280 16294
rect 32304 16292 32360 16294
rect 32384 16292 32440 16294
rect 32144 15258 32200 15260
rect 32224 15258 32280 15260
rect 32304 15258 32360 15260
rect 32384 15258 32440 15260
rect 32144 15206 32170 15258
rect 32170 15206 32200 15258
rect 32224 15206 32234 15258
rect 32234 15206 32280 15258
rect 32304 15206 32350 15258
rect 32350 15206 32360 15258
rect 32384 15206 32414 15258
rect 32414 15206 32440 15258
rect 32144 15204 32200 15206
rect 32224 15204 32280 15206
rect 32304 15204 32360 15206
rect 32384 15204 32440 15206
rect 32402 15036 32404 15056
rect 32404 15036 32456 15056
rect 32456 15036 32458 15056
rect 32402 15000 32458 15036
rect 30102 10648 30158 10704
rect 27894 8472 27950 8528
rect 27250 6432 27306 6488
rect 27158 6296 27214 6352
rect 27802 6976 27858 7032
rect 27802 5888 27858 5944
rect 27526 5480 27582 5536
rect 27250 5072 27306 5128
rect 26146 3340 26148 3360
rect 26148 3340 26200 3360
rect 26200 3340 26202 3360
rect 26146 3304 26202 3340
rect 27434 4528 27490 4584
rect 26882 3712 26938 3768
rect 26790 3304 26846 3360
rect 27986 6976 28042 7032
rect 27986 5344 28042 5400
rect 32144 14170 32200 14172
rect 32224 14170 32280 14172
rect 32304 14170 32360 14172
rect 32384 14170 32440 14172
rect 32144 14118 32170 14170
rect 32170 14118 32200 14170
rect 32224 14118 32234 14170
rect 32234 14118 32280 14170
rect 32304 14118 32350 14170
rect 32350 14118 32360 14170
rect 32384 14118 32414 14170
rect 32414 14118 32440 14170
rect 32144 14116 32200 14118
rect 32224 14116 32280 14118
rect 32304 14116 32360 14118
rect 32384 14116 32440 14118
rect 30930 13504 30986 13560
rect 31390 12724 31392 12744
rect 31392 12724 31444 12744
rect 31444 12724 31446 12744
rect 31390 12688 31446 12724
rect 31390 12416 31446 12472
rect 32144 13082 32200 13084
rect 32224 13082 32280 13084
rect 32304 13082 32360 13084
rect 32384 13082 32440 13084
rect 32144 13030 32170 13082
rect 32170 13030 32200 13082
rect 32224 13030 32234 13082
rect 32234 13030 32280 13082
rect 32304 13030 32350 13082
rect 32350 13030 32360 13082
rect 32384 13030 32414 13082
rect 32414 13030 32440 13082
rect 32144 13028 32200 13030
rect 32224 13028 32280 13030
rect 32304 13028 32360 13030
rect 32384 13028 32440 13030
rect 32126 12708 32182 12744
rect 32126 12688 32128 12708
rect 32128 12688 32180 12708
rect 32180 12688 32182 12708
rect 30470 10512 30526 10568
rect 30286 9052 30288 9072
rect 30288 9052 30340 9072
rect 30340 9052 30342 9072
rect 30286 9016 30342 9052
rect 29090 7812 29146 7848
rect 29090 7792 29092 7812
rect 29092 7792 29144 7812
rect 29144 7792 29146 7812
rect 29550 8200 29606 8256
rect 28998 7112 29054 7168
rect 29090 6976 29146 7032
rect 29550 7656 29606 7712
rect 29918 7792 29974 7848
rect 28722 6316 28778 6352
rect 28722 6296 28724 6316
rect 28724 6296 28776 6316
rect 28776 6296 28778 6316
rect 27986 3440 28042 3496
rect 28446 3848 28502 3904
rect 29090 5888 29146 5944
rect 28998 5344 29054 5400
rect 28906 4684 28962 4720
rect 28906 4664 28908 4684
rect 28908 4664 28960 4684
rect 28960 4664 28962 4684
rect 29550 5344 29606 5400
rect 29734 4972 29736 4992
rect 29736 4972 29788 4992
rect 29788 4972 29790 4992
rect 29734 4936 29790 4972
rect 30378 5208 30434 5264
rect 28814 3168 28870 3224
rect 29274 3304 29330 3360
rect 30654 4936 30710 4992
rect 30010 4528 30066 4584
rect 31022 9016 31078 9072
rect 31390 6976 31446 7032
rect 30838 3576 30894 3632
rect 29550 2760 29606 2816
rect 31482 6332 31484 6352
rect 31484 6332 31536 6352
rect 31536 6332 31538 6352
rect 31482 6296 31538 6332
rect 31482 6060 31484 6080
rect 31484 6060 31536 6080
rect 31536 6060 31538 6080
rect 31482 6024 31538 6060
rect 32586 13232 32642 13288
rect 32586 12980 32642 13016
rect 32586 12960 32588 12980
rect 32588 12960 32640 12980
rect 32640 12960 32642 12980
rect 32144 11994 32200 11996
rect 32224 11994 32280 11996
rect 32304 11994 32360 11996
rect 32384 11994 32440 11996
rect 32144 11942 32170 11994
rect 32170 11942 32200 11994
rect 32224 11942 32234 11994
rect 32234 11942 32280 11994
rect 32304 11942 32350 11994
rect 32350 11942 32360 11994
rect 32384 11942 32414 11994
rect 32414 11942 32440 11994
rect 32144 11940 32200 11942
rect 32224 11940 32280 11942
rect 32304 11940 32360 11942
rect 32384 11940 32440 11942
rect 32144 10906 32200 10908
rect 32224 10906 32280 10908
rect 32304 10906 32360 10908
rect 32384 10906 32440 10908
rect 32144 10854 32170 10906
rect 32170 10854 32200 10906
rect 32224 10854 32234 10906
rect 32234 10854 32280 10906
rect 32304 10854 32350 10906
rect 32350 10854 32360 10906
rect 32384 10854 32414 10906
rect 32414 10854 32440 10906
rect 32144 10852 32200 10854
rect 32224 10852 32280 10854
rect 32304 10852 32360 10854
rect 32384 10852 32440 10854
rect 32310 10548 32312 10568
rect 32312 10548 32364 10568
rect 32364 10548 32366 10568
rect 32310 10512 32366 10548
rect 33046 11500 33048 11520
rect 33048 11500 33100 11520
rect 33100 11500 33102 11520
rect 33046 11464 33102 11500
rect 33690 13640 33746 13696
rect 33782 13368 33838 13424
rect 33782 12280 33838 12336
rect 33966 12416 34022 12472
rect 34610 12588 34612 12608
rect 34612 12588 34664 12608
rect 34664 12588 34666 12608
rect 34610 12552 34666 12588
rect 32144 9818 32200 9820
rect 32224 9818 32280 9820
rect 32304 9818 32360 9820
rect 32384 9818 32440 9820
rect 32144 9766 32170 9818
rect 32170 9766 32200 9818
rect 32224 9766 32234 9818
rect 32234 9766 32280 9818
rect 32304 9766 32350 9818
rect 32350 9766 32360 9818
rect 32384 9766 32414 9818
rect 32414 9766 32440 9818
rect 32144 9764 32200 9766
rect 32224 9764 32280 9766
rect 32304 9764 32360 9766
rect 32384 9764 32440 9766
rect 32402 9036 32458 9072
rect 32402 9016 32404 9036
rect 32404 9016 32456 9036
rect 32456 9016 32458 9036
rect 32144 8730 32200 8732
rect 32224 8730 32280 8732
rect 32304 8730 32360 8732
rect 32384 8730 32440 8732
rect 32144 8678 32170 8730
rect 32170 8678 32200 8730
rect 32224 8678 32234 8730
rect 32234 8678 32280 8730
rect 32304 8678 32350 8730
rect 32350 8678 32360 8730
rect 32384 8678 32414 8730
rect 32414 8678 32440 8730
rect 32144 8676 32200 8678
rect 32224 8676 32280 8678
rect 32304 8676 32360 8678
rect 32384 8676 32440 8678
rect 32144 7642 32200 7644
rect 32224 7642 32280 7644
rect 32304 7642 32360 7644
rect 32384 7642 32440 7644
rect 32144 7590 32170 7642
rect 32170 7590 32200 7642
rect 32224 7590 32234 7642
rect 32234 7590 32280 7642
rect 32304 7590 32350 7642
rect 32350 7590 32360 7642
rect 32384 7590 32414 7642
rect 32414 7590 32440 7642
rect 32144 7588 32200 7590
rect 32224 7588 32280 7590
rect 32304 7588 32360 7590
rect 32384 7588 32440 7590
rect 32402 7148 32404 7168
rect 32404 7148 32456 7168
rect 32456 7148 32458 7168
rect 32402 7112 32458 7148
rect 32144 6554 32200 6556
rect 32224 6554 32280 6556
rect 32304 6554 32360 6556
rect 32384 6554 32440 6556
rect 32144 6502 32170 6554
rect 32170 6502 32200 6554
rect 32224 6502 32234 6554
rect 32234 6502 32280 6554
rect 32304 6502 32350 6554
rect 32350 6502 32360 6554
rect 32384 6502 32414 6554
rect 32414 6502 32440 6554
rect 32144 6500 32200 6502
rect 32224 6500 32280 6502
rect 32304 6500 32360 6502
rect 32384 6500 32440 6502
rect 31390 5908 31446 5944
rect 31390 5888 31392 5908
rect 31392 5888 31444 5908
rect 31444 5888 31446 5908
rect 30930 2896 30986 2952
rect 31206 4936 31262 4992
rect 31666 6024 31722 6080
rect 31942 6024 31998 6080
rect 32034 5888 32090 5944
rect 32144 5466 32200 5468
rect 32224 5466 32280 5468
rect 32304 5466 32360 5468
rect 32384 5466 32440 5468
rect 32144 5414 32170 5466
rect 32170 5414 32200 5466
rect 32224 5414 32234 5466
rect 32234 5414 32280 5466
rect 32304 5414 32350 5466
rect 32350 5414 32360 5466
rect 32384 5414 32414 5466
rect 32414 5414 32440 5466
rect 32144 5412 32200 5414
rect 32224 5412 32280 5414
rect 32304 5412 32360 5414
rect 32384 5412 32440 5414
rect 32034 5208 32090 5264
rect 31942 4936 31998 4992
rect 31574 4664 31630 4720
rect 32310 4800 32366 4856
rect 32144 4378 32200 4380
rect 32224 4378 32280 4380
rect 32304 4378 32360 4380
rect 32384 4378 32440 4380
rect 32144 4326 32170 4378
rect 32170 4326 32200 4378
rect 32224 4326 32234 4378
rect 32234 4326 32280 4378
rect 32304 4326 32350 4378
rect 32350 4326 32360 4378
rect 32384 4326 32414 4378
rect 32414 4326 32440 4378
rect 32144 4324 32200 4326
rect 32224 4324 32280 4326
rect 32304 4324 32360 4326
rect 32384 4324 32440 4326
rect 32034 4120 32090 4176
rect 32218 3848 32274 3904
rect 31390 3576 31446 3632
rect 31298 3304 31354 3360
rect 31850 3440 31906 3496
rect 31482 3168 31538 3224
rect 32034 3440 32090 3496
rect 32144 3290 32200 3292
rect 32224 3290 32280 3292
rect 32304 3290 32360 3292
rect 32384 3290 32440 3292
rect 32144 3238 32170 3290
rect 32170 3238 32200 3290
rect 32224 3238 32234 3290
rect 32234 3238 32280 3290
rect 32304 3238 32350 3290
rect 32350 3238 32360 3290
rect 32384 3238 32414 3290
rect 32414 3238 32440 3290
rect 32144 3236 32200 3238
rect 32224 3236 32280 3238
rect 32304 3236 32360 3238
rect 32384 3236 32440 3238
rect 32126 3068 32128 3088
rect 32128 3068 32180 3088
rect 32180 3068 32182 3088
rect 32126 3032 32182 3068
rect 32586 4392 32642 4448
rect 33046 5344 33102 5400
rect 32862 3848 32918 3904
rect 33874 8336 33930 8392
rect 33782 8064 33838 8120
rect 35070 12688 35126 12744
rect 33138 4664 33194 4720
rect 33138 3848 33194 3904
rect 32770 3168 32826 3224
rect 32144 2202 32200 2204
rect 32224 2202 32280 2204
rect 32304 2202 32360 2204
rect 32384 2202 32440 2204
rect 32144 2150 32170 2202
rect 32170 2150 32200 2202
rect 32224 2150 32234 2202
rect 32234 2150 32280 2202
rect 32304 2150 32350 2202
rect 32350 2150 32360 2202
rect 32384 2150 32414 2202
rect 32414 2150 32440 2202
rect 32144 2148 32200 2150
rect 32224 2148 32280 2150
rect 32304 2148 32360 2150
rect 32384 2148 32440 2150
rect 33874 6296 33930 6352
rect 34242 6196 34244 6216
rect 34244 6196 34296 6216
rect 34296 6196 34298 6216
rect 34242 6160 34298 6196
rect 33782 4256 33838 4312
rect 36358 13504 36414 13560
rect 35438 8084 35494 8120
rect 35438 8064 35440 8084
rect 35440 8064 35492 8084
rect 35492 8064 35494 8084
rect 35254 7928 35310 7984
rect 35622 8064 35678 8120
rect 35990 9560 36046 9616
rect 35622 6296 35678 6352
rect 34610 4528 34666 4584
rect 36634 13776 36690 13832
rect 37186 12960 37242 13016
rect 37370 11464 37426 11520
rect 38934 15988 38936 16008
rect 38936 15988 38988 16008
rect 38988 15988 38990 16008
rect 38934 15952 38990 15988
rect 38842 12688 38898 12744
rect 37830 9596 37832 9616
rect 37832 9596 37884 9616
rect 37884 9596 37886 9616
rect 37830 9560 37886 9596
rect 38566 10648 38622 10704
rect 38842 10548 38844 10568
rect 38844 10548 38896 10568
rect 38896 10548 38898 10568
rect 38842 10512 38898 10548
rect 39302 14184 39358 14240
rect 39026 14048 39082 14104
rect 40314 13776 40370 13832
rect 39210 13368 39266 13424
rect 40866 15000 40922 15056
rect 39210 12724 39212 12744
rect 39212 12724 39264 12744
rect 39264 12724 39266 12744
rect 39210 12688 39266 12724
rect 38842 9424 38898 9480
rect 36634 7248 36690 7304
rect 36542 6976 36598 7032
rect 35622 4120 35678 4176
rect 33782 2896 33838 2952
rect 33966 2896 34022 2952
rect 34886 3440 34942 3496
rect 36358 4664 36414 4720
rect 36634 4392 36690 4448
rect 39762 11192 39818 11248
rect 42540 16890 42596 16892
rect 42620 16890 42676 16892
rect 42700 16890 42756 16892
rect 42780 16890 42836 16892
rect 42540 16838 42566 16890
rect 42566 16838 42596 16890
rect 42620 16838 42630 16890
rect 42630 16838 42676 16890
rect 42700 16838 42746 16890
rect 42746 16838 42756 16890
rect 42780 16838 42810 16890
rect 42810 16838 42836 16890
rect 42540 16836 42596 16838
rect 42620 16836 42676 16838
rect 42700 16836 42756 16838
rect 42780 16836 42836 16838
rect 41970 15000 42026 15056
rect 41878 14900 41880 14920
rect 41880 14900 41932 14920
rect 41932 14900 41934 14920
rect 41878 14864 41934 14900
rect 41418 14220 41420 14240
rect 41420 14220 41472 14240
rect 41472 14220 41474 14240
rect 41418 14184 41474 14220
rect 42540 15802 42596 15804
rect 42620 15802 42676 15804
rect 42700 15802 42756 15804
rect 42780 15802 42836 15804
rect 42540 15750 42566 15802
rect 42566 15750 42596 15802
rect 42620 15750 42630 15802
rect 42630 15750 42676 15802
rect 42700 15750 42746 15802
rect 42746 15750 42756 15802
rect 42780 15750 42810 15802
rect 42810 15750 42836 15802
rect 42540 15748 42596 15750
rect 42620 15748 42676 15750
rect 42700 15748 42756 15750
rect 42780 15748 42836 15750
rect 42246 14864 42302 14920
rect 42540 14714 42596 14716
rect 42620 14714 42676 14716
rect 42700 14714 42756 14716
rect 42780 14714 42836 14716
rect 42540 14662 42566 14714
rect 42566 14662 42596 14714
rect 42620 14662 42630 14714
rect 42630 14662 42676 14714
rect 42700 14662 42746 14714
rect 42746 14662 42756 14714
rect 42780 14662 42810 14714
rect 42810 14662 42836 14714
rect 42540 14660 42596 14662
rect 42620 14660 42676 14662
rect 42700 14660 42756 14662
rect 42780 14660 42836 14662
rect 46202 15988 46204 16008
rect 46204 15988 46256 16008
rect 46256 15988 46258 16008
rect 46202 15952 46258 15988
rect 41326 12688 41382 12744
rect 38382 8064 38438 8120
rect 36910 7384 36966 7440
rect 37922 6840 37978 6896
rect 40314 8372 40316 8392
rect 40316 8372 40368 8392
rect 40368 8372 40370 8392
rect 38658 6840 38714 6896
rect 36818 4256 36874 4312
rect 38014 3304 38070 3360
rect 38750 4664 38806 4720
rect 39026 5480 39082 5536
rect 38750 3304 38806 3360
rect 38750 2796 38752 2816
rect 38752 2796 38804 2816
rect 38804 2796 38806 2816
rect 38750 2760 38806 2796
rect 39302 3168 39358 3224
rect 40314 8336 40370 8372
rect 40498 6024 40554 6080
rect 40314 4800 40370 4856
rect 39026 2488 39082 2544
rect 40314 3168 40370 3224
rect 42540 13626 42596 13628
rect 42620 13626 42676 13628
rect 42700 13626 42756 13628
rect 42780 13626 42836 13628
rect 42540 13574 42566 13626
rect 42566 13574 42596 13626
rect 42620 13574 42630 13626
rect 42630 13574 42676 13626
rect 42700 13574 42746 13626
rect 42746 13574 42756 13626
rect 42780 13574 42810 13626
rect 42810 13574 42836 13626
rect 42540 13572 42596 13574
rect 42620 13572 42676 13574
rect 42700 13572 42756 13574
rect 42780 13572 42836 13574
rect 43350 13776 43406 13832
rect 43994 14068 44050 14104
rect 43994 14048 43996 14068
rect 43996 14048 44048 14068
rect 44048 14048 44050 14068
rect 42540 12538 42596 12540
rect 42620 12538 42676 12540
rect 42700 12538 42756 12540
rect 42780 12538 42836 12540
rect 42540 12486 42566 12538
rect 42566 12486 42596 12538
rect 42620 12486 42630 12538
rect 42630 12486 42676 12538
rect 42700 12486 42746 12538
rect 42746 12486 42756 12538
rect 42780 12486 42810 12538
rect 42810 12486 42836 12538
rect 42540 12484 42596 12486
rect 42620 12484 42676 12486
rect 42700 12484 42756 12486
rect 42780 12484 42836 12486
rect 41050 9016 41106 9072
rect 41602 9560 41658 9616
rect 42540 11450 42596 11452
rect 42620 11450 42676 11452
rect 42700 11450 42756 11452
rect 42780 11450 42836 11452
rect 42540 11398 42566 11450
rect 42566 11398 42596 11450
rect 42620 11398 42630 11450
rect 42630 11398 42676 11450
rect 42700 11398 42746 11450
rect 42746 11398 42756 11450
rect 42780 11398 42810 11450
rect 42810 11398 42836 11450
rect 42540 11396 42596 11398
rect 42620 11396 42676 11398
rect 42700 11396 42756 11398
rect 42780 11396 42836 11398
rect 43350 11212 43406 11248
rect 43350 11192 43352 11212
rect 43352 11192 43404 11212
rect 43404 11192 43406 11212
rect 42540 10362 42596 10364
rect 42620 10362 42676 10364
rect 42700 10362 42756 10364
rect 42780 10362 42836 10364
rect 42540 10310 42566 10362
rect 42566 10310 42596 10362
rect 42620 10310 42630 10362
rect 42630 10310 42676 10362
rect 42700 10310 42746 10362
rect 42746 10310 42756 10362
rect 42780 10310 42810 10362
rect 42810 10310 42836 10362
rect 42540 10308 42596 10310
rect 42620 10308 42676 10310
rect 42700 10308 42756 10310
rect 42780 10308 42836 10310
rect 41970 9036 42026 9072
rect 41970 9016 41972 9036
rect 41972 9016 42024 9036
rect 42024 9016 42026 9036
rect 40866 8200 40922 8256
rect 40866 7792 40922 7848
rect 42540 9274 42596 9276
rect 42620 9274 42676 9276
rect 42700 9274 42756 9276
rect 42780 9274 42836 9276
rect 42540 9222 42566 9274
rect 42566 9222 42596 9274
rect 42620 9222 42630 9274
rect 42630 9222 42676 9274
rect 42700 9222 42746 9274
rect 42746 9222 42756 9274
rect 42780 9222 42810 9274
rect 42810 9222 42836 9274
rect 42540 9220 42596 9222
rect 42620 9220 42676 9222
rect 42700 9220 42756 9222
rect 42780 9220 42836 9222
rect 42540 8186 42596 8188
rect 42620 8186 42676 8188
rect 42700 8186 42756 8188
rect 42780 8186 42836 8188
rect 42540 8134 42566 8186
rect 42566 8134 42596 8186
rect 42620 8134 42630 8186
rect 42630 8134 42676 8186
rect 42700 8134 42746 8186
rect 42746 8134 42756 8186
rect 42780 8134 42810 8186
rect 42810 8134 42836 8186
rect 42540 8132 42596 8134
rect 42620 8132 42676 8134
rect 42700 8132 42756 8134
rect 42780 8132 42836 8134
rect 44546 13388 44602 13424
rect 44546 13368 44548 13388
rect 44548 13368 44600 13388
rect 44600 13368 44602 13388
rect 45926 12724 45928 12744
rect 45928 12724 45980 12744
rect 45980 12724 45982 12744
rect 44178 9596 44180 9616
rect 44180 9596 44232 9616
rect 44232 9596 44234 9616
rect 44178 9560 44234 9596
rect 43258 7928 43314 7984
rect 41050 6840 41106 6896
rect 41694 6024 41750 6080
rect 40958 5344 41014 5400
rect 42540 7098 42596 7100
rect 42620 7098 42676 7100
rect 42700 7098 42756 7100
rect 42780 7098 42836 7100
rect 42540 7046 42566 7098
rect 42566 7046 42596 7098
rect 42620 7046 42630 7098
rect 42630 7046 42676 7098
rect 42700 7046 42746 7098
rect 42746 7046 42756 7098
rect 42780 7046 42810 7098
rect 42810 7046 42836 7098
rect 42540 7044 42596 7046
rect 42620 7044 42676 7046
rect 42700 7044 42756 7046
rect 42780 7044 42836 7046
rect 41878 6196 41880 6216
rect 41880 6196 41932 6216
rect 41932 6196 41934 6216
rect 41878 6160 41934 6196
rect 40682 4936 40738 4992
rect 42246 6024 42302 6080
rect 42154 4684 42210 4720
rect 42154 4664 42156 4684
rect 42156 4664 42208 4684
rect 42208 4664 42210 4684
rect 42540 6010 42596 6012
rect 42620 6010 42676 6012
rect 42700 6010 42756 6012
rect 42780 6010 42836 6012
rect 42540 5958 42566 6010
rect 42566 5958 42596 6010
rect 42620 5958 42630 6010
rect 42630 5958 42676 6010
rect 42700 5958 42746 6010
rect 42746 5958 42756 6010
rect 42780 5958 42810 6010
rect 42810 5958 42836 6010
rect 42540 5956 42596 5958
rect 42620 5956 42676 5958
rect 42700 5956 42756 5958
rect 42780 5956 42836 5958
rect 42540 4922 42596 4924
rect 42620 4922 42676 4924
rect 42700 4922 42756 4924
rect 42780 4922 42836 4924
rect 42540 4870 42566 4922
rect 42566 4870 42596 4922
rect 42620 4870 42630 4922
rect 42630 4870 42676 4922
rect 42700 4870 42746 4922
rect 42746 4870 42756 4922
rect 42780 4870 42810 4922
rect 42810 4870 42836 4922
rect 42540 4868 42596 4870
rect 42620 4868 42676 4870
rect 42700 4868 42756 4870
rect 42780 4868 42836 4870
rect 42540 3834 42596 3836
rect 42620 3834 42676 3836
rect 42700 3834 42756 3836
rect 42780 3834 42836 3836
rect 42540 3782 42566 3834
rect 42566 3782 42596 3834
rect 42620 3782 42630 3834
rect 42630 3782 42676 3834
rect 42700 3782 42746 3834
rect 42746 3782 42756 3834
rect 42780 3782 42810 3834
rect 42810 3782 42836 3834
rect 42540 3780 42596 3782
rect 42620 3780 42676 3782
rect 42700 3780 42756 3782
rect 42780 3780 42836 3782
rect 42246 3712 42302 3768
rect 41970 3168 42026 3224
rect 43442 6704 43498 6760
rect 43902 6568 43958 6624
rect 42246 3168 42302 3224
rect 43442 3188 43498 3224
rect 43442 3168 43444 3188
rect 43444 3168 43496 3188
rect 43496 3168 43498 3188
rect 43166 3032 43222 3088
rect 42540 2746 42596 2748
rect 42620 2746 42676 2748
rect 42700 2746 42756 2748
rect 42780 2746 42836 2748
rect 42540 2694 42566 2746
rect 42566 2694 42596 2746
rect 42620 2694 42630 2746
rect 42630 2694 42676 2746
rect 42700 2694 42746 2746
rect 42746 2694 42756 2746
rect 42780 2694 42810 2746
rect 42810 2694 42836 2746
rect 42540 2692 42596 2694
rect 42620 2692 42676 2694
rect 42700 2692 42756 2694
rect 42780 2692 42836 2694
rect 44822 6160 44878 6216
rect 45650 11192 45706 11248
rect 45926 12688 45982 12724
rect 47030 13368 47086 13424
rect 52936 17434 52992 17436
rect 53016 17434 53072 17436
rect 53096 17434 53152 17436
rect 53176 17434 53232 17436
rect 52936 17382 52962 17434
rect 52962 17382 52992 17434
rect 53016 17382 53026 17434
rect 53026 17382 53072 17434
rect 53096 17382 53142 17434
rect 53142 17382 53152 17434
rect 53176 17382 53206 17434
rect 53206 17382 53232 17434
rect 52936 17380 52992 17382
rect 53016 17380 53072 17382
rect 53096 17380 53152 17382
rect 53176 17380 53232 17382
rect 46938 10512 46994 10568
rect 46202 7692 46204 7712
rect 46204 7692 46256 7712
rect 46256 7692 46258 7712
rect 46202 7656 46258 7692
rect 46110 7248 46166 7304
rect 43902 3440 43958 3496
rect 44178 3440 44234 3496
rect 48410 12824 48466 12880
rect 52936 16346 52992 16348
rect 53016 16346 53072 16348
rect 53096 16346 53152 16348
rect 53176 16346 53232 16348
rect 52936 16294 52962 16346
rect 52962 16294 52992 16346
rect 53016 16294 53026 16346
rect 53026 16294 53072 16346
rect 53096 16294 53142 16346
rect 53142 16294 53152 16346
rect 53176 16294 53206 16346
rect 53206 16294 53232 16346
rect 52936 16292 52992 16294
rect 53016 16292 53072 16294
rect 53096 16292 53152 16294
rect 53176 16292 53232 16294
rect 52936 15258 52992 15260
rect 53016 15258 53072 15260
rect 53096 15258 53152 15260
rect 53176 15258 53232 15260
rect 52936 15206 52962 15258
rect 52962 15206 52992 15258
rect 53016 15206 53026 15258
rect 53026 15206 53072 15258
rect 53096 15206 53142 15258
rect 53142 15206 53152 15258
rect 53176 15206 53206 15258
rect 53206 15206 53232 15258
rect 52936 15204 52992 15206
rect 53016 15204 53072 15206
rect 53096 15204 53152 15206
rect 53176 15204 53232 15206
rect 50526 12844 50582 12880
rect 50526 12824 50528 12844
rect 50528 12824 50580 12844
rect 50580 12824 50582 12844
rect 50710 12300 50766 12336
rect 50710 12280 50712 12300
rect 50712 12280 50764 12300
rect 50764 12280 50766 12300
rect 47490 9560 47546 9616
rect 47490 9424 47546 9480
rect 47214 8336 47270 8392
rect 46938 6840 46994 6896
rect 46294 5480 46350 5536
rect 45650 4140 45706 4176
rect 45650 4120 45652 4140
rect 45652 4120 45704 4140
rect 45704 4120 45706 4140
rect 44914 3032 44970 3088
rect 45098 3032 45154 3088
rect 44822 2760 44878 2816
rect 46110 3440 46166 3496
rect 45466 2488 45522 2544
rect 47674 8064 47730 8120
rect 47306 7656 47362 7712
rect 47030 6432 47086 6488
rect 46662 4664 46718 4720
rect 48686 10376 48742 10432
rect 48226 8064 48282 8120
rect 47030 3576 47086 3632
rect 47030 3068 47032 3088
rect 47032 3068 47084 3088
rect 47084 3068 47086 3088
rect 47030 3032 47086 3068
rect 46386 2760 46442 2816
rect 48502 8372 48504 8392
rect 48504 8372 48556 8392
rect 48556 8372 48558 8392
rect 48502 8336 48558 8372
rect 49514 10512 49570 10568
rect 50250 9460 50252 9480
rect 50252 9460 50304 9480
rect 50304 9460 50306 9480
rect 49514 8336 49570 8392
rect 49146 7948 49202 7984
rect 49146 7928 49148 7948
rect 49148 7928 49200 7948
rect 49200 7928 49202 7948
rect 48134 7268 48190 7304
rect 48134 7248 48136 7268
rect 48136 7248 48188 7268
rect 48188 7248 48190 7268
rect 48410 6860 48466 6896
rect 48410 6840 48412 6860
rect 48412 6840 48464 6860
rect 48464 6840 48466 6860
rect 49054 6568 49110 6624
rect 48778 6160 48834 6216
rect 47950 4140 48006 4176
rect 47950 4120 47952 4140
rect 47952 4120 48004 4140
rect 48004 4120 48006 4140
rect 47674 3304 47730 3360
rect 48502 4392 48558 4448
rect 49146 5752 49202 5808
rect 50250 9424 50306 9460
rect 50986 10512 51042 10568
rect 49790 7928 49846 7984
rect 48870 3440 48926 3496
rect 50434 6432 50490 6488
rect 50710 7656 50766 7712
rect 51722 10548 51724 10568
rect 51724 10548 51776 10568
rect 51776 10548 51778 10568
rect 51722 10512 51778 10548
rect 51262 8880 51318 8936
rect 51722 9460 51724 9480
rect 51724 9460 51776 9480
rect 51776 9460 51778 9480
rect 51722 9424 51778 9460
rect 50802 6432 50858 6488
rect 49606 4700 49608 4720
rect 49608 4700 49660 4720
rect 49660 4700 49662 4720
rect 49606 4664 49662 4700
rect 50894 5108 50896 5128
rect 50896 5108 50948 5128
rect 50948 5108 50950 5128
rect 50894 5072 50950 5108
rect 49514 3168 49570 3224
rect 49882 3984 49938 4040
rect 50434 3712 50490 3768
rect 50894 3984 50950 4040
rect 51998 7948 52054 7984
rect 51998 7928 52000 7948
rect 52000 7928 52052 7948
rect 52052 7928 52054 7948
rect 51814 7792 51870 7848
rect 51538 6568 51594 6624
rect 51906 6196 51908 6216
rect 51908 6196 51960 6216
rect 51960 6196 51962 6216
rect 51906 6160 51962 6196
rect 51538 4700 51540 4720
rect 51540 4700 51592 4720
rect 51592 4700 51594 4720
rect 51538 4664 51594 4700
rect 51906 4428 51908 4448
rect 51908 4428 51960 4448
rect 51960 4428 51962 4448
rect 51906 4392 51962 4428
rect 51722 3712 51778 3768
rect 52274 10412 52276 10432
rect 52276 10412 52328 10432
rect 52328 10412 52330 10432
rect 52274 10376 52330 10412
rect 52936 14170 52992 14172
rect 53016 14170 53072 14172
rect 53096 14170 53152 14172
rect 53176 14170 53232 14172
rect 52936 14118 52962 14170
rect 52962 14118 52992 14170
rect 53016 14118 53026 14170
rect 53026 14118 53072 14170
rect 53096 14118 53142 14170
rect 53142 14118 53152 14170
rect 53176 14118 53206 14170
rect 53206 14118 53232 14170
rect 52936 14116 52992 14118
rect 53016 14116 53072 14118
rect 53096 14116 53152 14118
rect 53176 14116 53232 14118
rect 52936 13082 52992 13084
rect 53016 13082 53072 13084
rect 53096 13082 53152 13084
rect 53176 13082 53232 13084
rect 52936 13030 52962 13082
rect 52962 13030 52992 13082
rect 53016 13030 53026 13082
rect 53026 13030 53072 13082
rect 53096 13030 53142 13082
rect 53142 13030 53152 13082
rect 53176 13030 53206 13082
rect 53206 13030 53232 13082
rect 52936 13028 52992 13030
rect 53016 13028 53072 13030
rect 53096 13028 53152 13030
rect 53176 13028 53232 13030
rect 52936 11994 52992 11996
rect 53016 11994 53072 11996
rect 53096 11994 53152 11996
rect 53176 11994 53232 11996
rect 52936 11942 52962 11994
rect 52962 11942 52992 11994
rect 53016 11942 53026 11994
rect 53026 11942 53072 11994
rect 53096 11942 53142 11994
rect 53142 11942 53152 11994
rect 53176 11942 53206 11994
rect 53206 11942 53232 11994
rect 52936 11940 52992 11942
rect 53016 11940 53072 11942
rect 53096 11940 53152 11942
rect 53176 11940 53232 11942
rect 52936 10906 52992 10908
rect 53016 10906 53072 10908
rect 53096 10906 53152 10908
rect 53176 10906 53232 10908
rect 52936 10854 52962 10906
rect 52962 10854 52992 10906
rect 53016 10854 53026 10906
rect 53026 10854 53072 10906
rect 53096 10854 53142 10906
rect 53142 10854 53152 10906
rect 53176 10854 53206 10906
rect 53206 10854 53232 10906
rect 52936 10852 52992 10854
rect 53016 10852 53072 10854
rect 53096 10852 53152 10854
rect 53176 10852 53232 10854
rect 52936 9818 52992 9820
rect 53016 9818 53072 9820
rect 53096 9818 53152 9820
rect 53176 9818 53232 9820
rect 52936 9766 52962 9818
rect 52962 9766 52992 9818
rect 53016 9766 53026 9818
rect 53026 9766 53072 9818
rect 53096 9766 53142 9818
rect 53142 9766 53152 9818
rect 53176 9766 53206 9818
rect 53206 9766 53232 9818
rect 52936 9764 52992 9766
rect 53016 9764 53072 9766
rect 53096 9764 53152 9766
rect 53176 9764 53232 9766
rect 52936 8730 52992 8732
rect 53016 8730 53072 8732
rect 53096 8730 53152 8732
rect 53176 8730 53232 8732
rect 52936 8678 52962 8730
rect 52962 8678 52992 8730
rect 53016 8678 53026 8730
rect 53026 8678 53072 8730
rect 53096 8678 53142 8730
rect 53142 8678 53152 8730
rect 53176 8678 53206 8730
rect 53206 8678 53232 8730
rect 52936 8676 52992 8678
rect 53016 8676 53072 8678
rect 53096 8676 53152 8678
rect 53176 8676 53232 8678
rect 52550 7928 52606 7984
rect 52182 7656 52238 7712
rect 52936 7642 52992 7644
rect 53016 7642 53072 7644
rect 53096 7642 53152 7644
rect 53176 7642 53232 7644
rect 52936 7590 52962 7642
rect 52962 7590 52992 7642
rect 53016 7590 53026 7642
rect 53026 7590 53072 7642
rect 53096 7590 53142 7642
rect 53142 7590 53152 7642
rect 53176 7590 53206 7642
rect 53206 7590 53232 7642
rect 52936 7588 52992 7590
rect 53016 7588 53072 7590
rect 53096 7588 53152 7590
rect 53176 7588 53232 7590
rect 53010 7420 53012 7440
rect 53012 7420 53064 7440
rect 53064 7420 53066 7440
rect 53010 7384 53066 7420
rect 52936 6554 52992 6556
rect 53016 6554 53072 6556
rect 53096 6554 53152 6556
rect 53176 6554 53232 6556
rect 52936 6502 52962 6554
rect 52962 6502 52992 6554
rect 53016 6502 53026 6554
rect 53026 6502 53072 6554
rect 53096 6502 53142 6554
rect 53142 6502 53152 6554
rect 53176 6502 53206 6554
rect 53206 6502 53232 6554
rect 52936 6500 52992 6502
rect 53016 6500 53072 6502
rect 53096 6500 53152 6502
rect 53176 6500 53232 6502
rect 53010 6196 53012 6216
rect 53012 6196 53064 6216
rect 53064 6196 53066 6216
rect 53010 6160 53066 6196
rect 52936 5466 52992 5468
rect 53016 5466 53072 5468
rect 53096 5466 53152 5468
rect 53176 5466 53232 5468
rect 52936 5414 52962 5466
rect 52962 5414 52992 5466
rect 53016 5414 53026 5466
rect 53026 5414 53072 5466
rect 53096 5414 53142 5466
rect 53142 5414 53152 5466
rect 53176 5414 53206 5466
rect 53206 5414 53232 5466
rect 52936 5412 52992 5414
rect 53016 5412 53072 5414
rect 53096 5412 53152 5414
rect 53176 5412 53232 5414
rect 52182 4140 52238 4176
rect 52182 4120 52184 4140
rect 52184 4120 52236 4140
rect 52236 4120 52238 4140
rect 52936 4378 52992 4380
rect 53016 4378 53072 4380
rect 53096 4378 53152 4380
rect 53176 4378 53232 4380
rect 52936 4326 52962 4378
rect 52962 4326 52992 4378
rect 53016 4326 53026 4378
rect 53026 4326 53072 4378
rect 53096 4326 53142 4378
rect 53142 4326 53152 4378
rect 53176 4326 53206 4378
rect 53206 4326 53232 4378
rect 52936 4324 52992 4326
rect 53016 4324 53072 4326
rect 53096 4324 53152 4326
rect 53176 4324 53232 4326
rect 52550 4020 52552 4040
rect 52552 4020 52604 4040
rect 52604 4020 52606 4040
rect 52550 3984 52606 4020
rect 52734 3984 52790 4040
rect 52936 3290 52992 3292
rect 53016 3290 53072 3292
rect 53096 3290 53152 3292
rect 53176 3290 53232 3292
rect 52936 3238 52962 3290
rect 52962 3238 52992 3290
rect 53016 3238 53026 3290
rect 53026 3238 53072 3290
rect 53096 3238 53142 3290
rect 53142 3238 53152 3290
rect 53176 3238 53206 3290
rect 53206 3238 53232 3290
rect 52936 3236 52992 3238
rect 53016 3236 53072 3238
rect 53096 3236 53152 3238
rect 53176 3236 53232 3238
rect 54942 6860 54998 6896
rect 54942 6840 54944 6860
rect 54944 6840 54996 6860
rect 54996 6840 54998 6860
rect 56874 11736 56930 11792
rect 55034 6160 55090 6216
rect 55678 6296 55734 6352
rect 54298 4548 54354 4584
rect 54298 4528 54300 4548
rect 54300 4528 54352 4548
rect 54352 4528 54354 4548
rect 54114 3848 54170 3904
rect 54666 4120 54722 4176
rect 55034 4528 55090 4584
rect 55310 5208 55366 5264
rect 52936 2202 52992 2204
rect 53016 2202 53072 2204
rect 53096 2202 53152 2204
rect 53176 2202 53232 2204
rect 52936 2150 52962 2202
rect 52962 2150 52992 2202
rect 53016 2150 53026 2202
rect 53026 2150 53072 2202
rect 53096 2150 53142 2202
rect 53142 2150 53152 2202
rect 53176 2150 53206 2202
rect 53206 2150 53232 2202
rect 52936 2148 52992 2150
rect 53016 2148 53072 2150
rect 53096 2148 53152 2150
rect 53176 2148 53232 2150
rect 55218 4004 55274 4040
rect 55218 3984 55220 4004
rect 55220 3984 55272 4004
rect 55272 3984 55274 4004
rect 56506 8916 56508 8936
rect 56508 8916 56560 8936
rect 56560 8916 56562 8936
rect 56138 7792 56194 7848
rect 56506 8880 56562 8916
rect 56690 7948 56746 7984
rect 56690 7928 56692 7948
rect 56692 7928 56744 7948
rect 56744 7928 56746 7948
rect 57426 7792 57482 7848
rect 56414 5228 56470 5264
rect 56414 5208 56416 5228
rect 56416 5208 56468 5228
rect 56468 5208 56470 5228
rect 56598 5582 56654 5638
rect 56322 3440 56378 3496
rect 60002 5888 60058 5944
rect 60278 2916 60334 2952
rect 60278 2896 60280 2916
rect 60280 2896 60332 2916
rect 60332 2896 60334 2916
<< metal3 >>
rect 0 18866 800 18896
rect 3969 18866 4035 18869
rect 0 18864 4035 18866
rect 0 18808 3974 18864
rect 4030 18808 4035 18864
rect 0 18806 4035 18808
rect 0 18776 800 18806
rect 3969 18803 4035 18806
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 32132 17440 32452 17441
rect 32132 17376 32140 17440
rect 32204 17376 32220 17440
rect 32284 17376 32300 17440
rect 32364 17376 32380 17440
rect 32444 17376 32452 17440
rect 32132 17375 32452 17376
rect 52924 17440 53244 17441
rect 52924 17376 52932 17440
rect 52996 17376 53012 17440
rect 53076 17376 53092 17440
rect 53156 17376 53172 17440
rect 53236 17376 53244 17440
rect 52924 17375 53244 17376
rect 21736 16896 22056 16897
rect 21736 16832 21744 16896
rect 21808 16832 21824 16896
rect 21888 16832 21904 16896
rect 21968 16832 21984 16896
rect 22048 16832 22056 16896
rect 21736 16831 22056 16832
rect 42528 16896 42848 16897
rect 42528 16832 42536 16896
rect 42600 16832 42616 16896
rect 42680 16832 42696 16896
rect 42760 16832 42776 16896
rect 42840 16832 42848 16896
rect 42528 16831 42848 16832
rect 0 16690 800 16720
rect 4061 16690 4127 16693
rect 0 16688 4127 16690
rect 0 16632 4066 16688
rect 4122 16632 4127 16688
rect 0 16630 4127 16632
rect 0 16600 800 16630
rect 4061 16627 4127 16630
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 32132 16352 32452 16353
rect 32132 16288 32140 16352
rect 32204 16288 32220 16352
rect 32284 16288 32300 16352
rect 32364 16288 32380 16352
rect 32444 16288 32452 16352
rect 32132 16287 32452 16288
rect 52924 16352 53244 16353
rect 52924 16288 52932 16352
rect 52996 16288 53012 16352
rect 53076 16288 53092 16352
rect 53156 16288 53172 16352
rect 53236 16288 53244 16352
rect 52924 16287 53244 16288
rect 38929 16010 38995 16013
rect 46197 16010 46263 16013
rect 38929 16008 46263 16010
rect 38929 15952 38934 16008
rect 38990 15952 46202 16008
rect 46258 15952 46263 16008
rect 38929 15950 46263 15952
rect 38929 15947 38995 15950
rect 46197 15947 46263 15950
rect 21736 15808 22056 15809
rect 21736 15744 21744 15808
rect 21808 15744 21824 15808
rect 21888 15744 21904 15808
rect 21968 15744 21984 15808
rect 22048 15744 22056 15808
rect 21736 15743 22056 15744
rect 42528 15808 42848 15809
rect 42528 15744 42536 15808
rect 42600 15744 42616 15808
rect 42680 15744 42696 15808
rect 42760 15744 42776 15808
rect 42840 15744 42848 15808
rect 42528 15743 42848 15744
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 32132 15264 32452 15265
rect 32132 15200 32140 15264
rect 32204 15200 32220 15264
rect 32284 15200 32300 15264
rect 32364 15200 32380 15264
rect 32444 15200 32452 15264
rect 32132 15199 32452 15200
rect 52924 15264 53244 15265
rect 52924 15200 52932 15264
rect 52996 15200 53012 15264
rect 53076 15200 53092 15264
rect 53156 15200 53172 15264
rect 53236 15200 53244 15264
rect 52924 15199 53244 15200
rect 21909 15058 21975 15061
rect 22461 15058 22527 15061
rect 21909 15056 22527 15058
rect 21909 15000 21914 15056
rect 21970 15000 22466 15056
rect 22522 15000 22527 15056
rect 21909 14998 22527 15000
rect 21909 14995 21975 14998
rect 22461 14995 22527 14998
rect 32397 15058 32463 15061
rect 40861 15058 40927 15061
rect 41965 15058 42031 15061
rect 32397 15056 42031 15058
rect 32397 15000 32402 15056
rect 32458 15000 40866 15056
rect 40922 15000 41970 15056
rect 42026 15000 42031 15056
rect 32397 14998 42031 15000
rect 32397 14995 32463 14998
rect 40861 14995 40927 14998
rect 41965 14995 42031 14998
rect 19977 14922 20043 14925
rect 23657 14922 23723 14925
rect 19977 14920 23723 14922
rect 19977 14864 19982 14920
rect 20038 14864 23662 14920
rect 23718 14864 23723 14920
rect 19977 14862 23723 14864
rect 19977 14859 20043 14862
rect 23657 14859 23723 14862
rect 41873 14922 41939 14925
rect 42241 14922 42307 14925
rect 41873 14920 42307 14922
rect 41873 14864 41878 14920
rect 41934 14864 42246 14920
rect 42302 14864 42307 14920
rect 41873 14862 42307 14864
rect 41873 14859 41939 14862
rect 42241 14859 42307 14862
rect 21736 14720 22056 14721
rect 21736 14656 21744 14720
rect 21808 14656 21824 14720
rect 21888 14656 21904 14720
rect 21968 14656 21984 14720
rect 22048 14656 22056 14720
rect 21736 14655 22056 14656
rect 42528 14720 42848 14721
rect 42528 14656 42536 14720
rect 42600 14656 42616 14720
rect 42680 14656 42696 14720
rect 42760 14656 42776 14720
rect 42840 14656 42848 14720
rect 42528 14655 42848 14656
rect 0 14514 800 14544
rect 3141 14514 3207 14517
rect 0 14512 3207 14514
rect 0 14456 3146 14512
rect 3202 14456 3207 14512
rect 0 14454 3207 14456
rect 0 14424 800 14454
rect 3141 14451 3207 14454
rect 20805 14514 20871 14517
rect 28349 14514 28415 14517
rect 20805 14512 28415 14514
rect 20805 14456 20810 14512
rect 20866 14456 28354 14512
rect 28410 14456 28415 14512
rect 20805 14454 28415 14456
rect 20805 14451 20871 14454
rect 28349 14451 28415 14454
rect 21541 14378 21607 14381
rect 24669 14378 24735 14381
rect 21541 14376 24735 14378
rect 21541 14320 21546 14376
rect 21602 14320 24674 14376
rect 24730 14320 24735 14376
rect 21541 14318 24735 14320
rect 21541 14315 21607 14318
rect 24669 14315 24735 14318
rect 22093 14242 22159 14245
rect 24117 14242 24183 14245
rect 22093 14240 24183 14242
rect 22093 14184 22098 14240
rect 22154 14184 24122 14240
rect 24178 14184 24183 14240
rect 22093 14182 24183 14184
rect 22093 14179 22159 14182
rect 24117 14179 24183 14182
rect 39297 14242 39363 14245
rect 41413 14242 41479 14245
rect 39297 14240 41479 14242
rect 39297 14184 39302 14240
rect 39358 14184 41418 14240
rect 41474 14184 41479 14240
rect 39297 14182 41479 14184
rect 39297 14179 39363 14182
rect 41413 14179 41479 14182
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 32132 14176 32452 14177
rect 32132 14112 32140 14176
rect 32204 14112 32220 14176
rect 32284 14112 32300 14176
rect 32364 14112 32380 14176
rect 32444 14112 32452 14176
rect 32132 14111 32452 14112
rect 52924 14176 53244 14177
rect 52924 14112 52932 14176
rect 52996 14112 53012 14176
rect 53076 14112 53092 14176
rect 53156 14112 53172 14176
rect 53236 14112 53244 14176
rect 52924 14111 53244 14112
rect 17217 14106 17283 14109
rect 26233 14106 26299 14109
rect 17217 14104 26299 14106
rect 17217 14048 17222 14104
rect 17278 14048 26238 14104
rect 26294 14048 26299 14104
rect 17217 14046 26299 14048
rect 17217 14043 17283 14046
rect 26233 14043 26299 14046
rect 39021 14106 39087 14109
rect 43989 14106 44055 14109
rect 39021 14104 44055 14106
rect 39021 14048 39026 14104
rect 39082 14048 43994 14104
rect 44050 14048 44055 14104
rect 39021 14046 44055 14048
rect 39021 14043 39087 14046
rect 43989 14043 44055 14046
rect 17033 13970 17099 13973
rect 21173 13970 21239 13973
rect 17033 13968 21239 13970
rect 17033 13912 17038 13968
rect 17094 13912 21178 13968
rect 21234 13912 21239 13968
rect 17033 13910 21239 13912
rect 17033 13907 17099 13910
rect 21173 13907 21239 13910
rect 29085 13834 29151 13837
rect 36629 13834 36695 13837
rect 21590 13774 22202 13834
rect 12617 13698 12683 13701
rect 21590 13698 21650 13774
rect 12617 13696 21650 13698
rect 12617 13640 12622 13696
rect 12678 13640 21650 13696
rect 12617 13638 21650 13640
rect 22142 13698 22202 13774
rect 29085 13832 36695 13834
rect 29085 13776 29090 13832
rect 29146 13776 36634 13832
rect 36690 13776 36695 13832
rect 29085 13774 36695 13776
rect 29085 13771 29151 13774
rect 36629 13771 36695 13774
rect 40309 13834 40375 13837
rect 43345 13834 43411 13837
rect 40309 13832 43411 13834
rect 40309 13776 40314 13832
rect 40370 13776 43350 13832
rect 43406 13776 43411 13832
rect 40309 13774 43411 13776
rect 40309 13771 40375 13774
rect 43345 13771 43411 13774
rect 33685 13698 33751 13701
rect 22142 13696 33751 13698
rect 22142 13640 33690 13696
rect 33746 13640 33751 13696
rect 22142 13638 33751 13640
rect 12617 13635 12683 13638
rect 33685 13635 33751 13638
rect 21736 13632 22056 13633
rect 21736 13568 21744 13632
rect 21808 13568 21824 13632
rect 21888 13568 21904 13632
rect 21968 13568 21984 13632
rect 22048 13568 22056 13632
rect 21736 13567 22056 13568
rect 42528 13632 42848 13633
rect 42528 13568 42536 13632
rect 42600 13568 42616 13632
rect 42680 13568 42696 13632
rect 42760 13568 42776 13632
rect 42840 13568 42848 13632
rect 42528 13567 42848 13568
rect 9397 13562 9463 13565
rect 9857 13562 9923 13565
rect 17217 13562 17283 13565
rect 9397 13560 17283 13562
rect 9397 13504 9402 13560
rect 9458 13504 9862 13560
rect 9918 13504 17222 13560
rect 17278 13504 17283 13560
rect 9397 13502 17283 13504
rect 9397 13499 9463 13502
rect 9857 13499 9923 13502
rect 17217 13499 17283 13502
rect 30925 13562 30991 13565
rect 36353 13562 36419 13565
rect 30925 13560 36419 13562
rect 30925 13504 30930 13560
rect 30986 13504 36358 13560
rect 36414 13504 36419 13560
rect 30925 13502 36419 13504
rect 30925 13499 30991 13502
rect 36353 13499 36419 13502
rect 13077 13426 13143 13429
rect 33777 13426 33843 13429
rect 13077 13424 33843 13426
rect 13077 13368 13082 13424
rect 13138 13368 33782 13424
rect 33838 13368 33843 13424
rect 13077 13366 33843 13368
rect 13077 13363 13143 13366
rect 33777 13363 33843 13366
rect 39205 13426 39271 13429
rect 44541 13426 44607 13429
rect 47025 13426 47091 13429
rect 39205 13424 47091 13426
rect 39205 13368 39210 13424
rect 39266 13368 44546 13424
rect 44602 13368 47030 13424
rect 47086 13368 47091 13424
rect 39205 13366 47091 13368
rect 39205 13363 39271 13366
rect 44541 13363 44607 13366
rect 47025 13363 47091 13366
rect 3969 13290 4035 13293
rect 32581 13290 32647 13293
rect 3969 13288 32647 13290
rect 3969 13232 3974 13288
rect 4030 13232 32586 13288
rect 32642 13232 32647 13288
rect 3969 13230 32647 13232
rect 3969 13227 4035 13230
rect 32581 13227 32647 13230
rect 17217 13154 17283 13157
rect 22829 13154 22895 13157
rect 26785 13154 26851 13157
rect 17217 13152 26851 13154
rect 17217 13096 17222 13152
rect 17278 13096 22834 13152
rect 22890 13096 26790 13152
rect 26846 13096 26851 13152
rect 17217 13094 26851 13096
rect 17217 13091 17283 13094
rect 22829 13091 22895 13094
rect 26785 13091 26851 13094
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 32132 13088 32452 13089
rect 32132 13024 32140 13088
rect 32204 13024 32220 13088
rect 32284 13024 32300 13088
rect 32364 13024 32380 13088
rect 32444 13024 32452 13088
rect 32132 13023 32452 13024
rect 52924 13088 53244 13089
rect 52924 13024 52932 13088
rect 52996 13024 53012 13088
rect 53076 13024 53092 13088
rect 53156 13024 53172 13088
rect 53236 13024 53244 13088
rect 52924 13023 53244 13024
rect 19425 13018 19491 13021
rect 20253 13018 20319 13021
rect 19425 13016 20319 13018
rect 19425 12960 19430 13016
rect 19486 12960 20258 13016
rect 20314 12960 20319 13016
rect 19425 12958 20319 12960
rect 19425 12955 19491 12958
rect 20253 12955 20319 12958
rect 20437 13018 20503 13021
rect 26233 13018 26299 13021
rect 28349 13018 28415 13021
rect 20437 13016 28415 13018
rect 20437 12960 20442 13016
rect 20498 12960 26238 13016
rect 26294 12960 28354 13016
rect 28410 12960 28415 13016
rect 20437 12958 28415 12960
rect 20437 12955 20503 12958
rect 26233 12955 26299 12958
rect 28349 12955 28415 12958
rect 32581 13018 32647 13021
rect 37181 13018 37247 13021
rect 32581 13016 37247 13018
rect 32581 12960 32586 13016
rect 32642 12960 37186 13016
rect 37242 12960 37247 13016
rect 32581 12958 37247 12960
rect 32581 12955 32647 12958
rect 37181 12955 37247 12958
rect 9581 12882 9647 12885
rect 26785 12882 26851 12885
rect 48405 12882 48471 12885
rect 50521 12882 50587 12885
rect 9581 12880 23674 12882
rect 9581 12824 9586 12880
rect 9642 12824 23674 12880
rect 9581 12822 23674 12824
rect 9581 12819 9647 12822
rect 16021 12746 16087 12749
rect 16021 12744 23536 12746
rect 16021 12688 16026 12744
rect 16082 12688 23536 12744
rect 16021 12686 23536 12688
rect 16021 12683 16087 12686
rect 9489 12610 9555 12613
rect 9489 12608 21650 12610
rect 9489 12552 9494 12608
rect 9550 12552 21650 12608
rect 9489 12550 21650 12552
rect 9489 12547 9555 12550
rect 17769 12474 17835 12477
rect 20621 12474 20687 12477
rect 17769 12472 20687 12474
rect 17769 12416 17774 12472
rect 17830 12416 20626 12472
rect 20682 12416 20687 12472
rect 17769 12414 20687 12416
rect 17769 12411 17835 12414
rect 20621 12411 20687 12414
rect 9305 12338 9371 12341
rect 16849 12338 16915 12341
rect 9305 12336 16915 12338
rect 9305 12280 9310 12336
rect 9366 12280 16854 12336
rect 16910 12280 16915 12336
rect 9305 12278 16915 12280
rect 21590 12338 21650 12550
rect 21736 12544 22056 12545
rect 21736 12480 21744 12544
rect 21808 12480 21824 12544
rect 21888 12480 21904 12544
rect 21968 12480 21984 12544
rect 22048 12480 22056 12544
rect 21736 12479 22056 12480
rect 22737 12474 22803 12477
rect 22142 12472 22803 12474
rect 22142 12416 22742 12472
rect 22798 12416 22803 12472
rect 22142 12414 22803 12416
rect 23476 12474 23536 12686
rect 23614 12610 23674 12822
rect 26785 12880 50587 12882
rect 26785 12824 26790 12880
rect 26846 12824 48410 12880
rect 48466 12824 50526 12880
rect 50582 12824 50587 12880
rect 26785 12822 50587 12824
rect 26785 12819 26851 12822
rect 48405 12819 48471 12822
rect 50521 12819 50587 12822
rect 31385 12746 31451 12749
rect 32121 12746 32187 12749
rect 35065 12746 35131 12749
rect 31385 12744 35131 12746
rect 31385 12688 31390 12744
rect 31446 12688 32126 12744
rect 32182 12688 35070 12744
rect 35126 12688 35131 12744
rect 31385 12686 35131 12688
rect 31385 12683 31451 12686
rect 32121 12683 32187 12686
rect 35065 12683 35131 12686
rect 38837 12746 38903 12749
rect 39205 12746 39271 12749
rect 38837 12744 39271 12746
rect 38837 12688 38842 12744
rect 38898 12688 39210 12744
rect 39266 12688 39271 12744
rect 38837 12686 39271 12688
rect 38837 12683 38903 12686
rect 39205 12683 39271 12686
rect 41321 12746 41387 12749
rect 45921 12746 45987 12749
rect 41321 12744 45987 12746
rect 41321 12688 41326 12744
rect 41382 12688 45926 12744
rect 45982 12688 45987 12744
rect 41321 12686 45987 12688
rect 41321 12683 41387 12686
rect 45921 12683 45987 12686
rect 25313 12610 25379 12613
rect 25957 12610 26023 12613
rect 34605 12610 34671 12613
rect 23614 12608 34671 12610
rect 23614 12552 25318 12608
rect 25374 12552 25962 12608
rect 26018 12552 34610 12608
rect 34666 12552 34671 12608
rect 23614 12550 34671 12552
rect 25313 12547 25379 12550
rect 25957 12547 26023 12550
rect 34605 12547 34671 12550
rect 42528 12544 42848 12545
rect 42528 12480 42536 12544
rect 42600 12480 42616 12544
rect 42680 12480 42696 12544
rect 42760 12480 42776 12544
rect 42840 12480 42848 12544
rect 42528 12479 42848 12480
rect 28717 12474 28783 12477
rect 23476 12472 28783 12474
rect 23476 12416 28722 12472
rect 28778 12416 28783 12472
rect 23476 12414 28783 12416
rect 22142 12338 22202 12414
rect 22737 12411 22803 12414
rect 28717 12411 28783 12414
rect 31385 12474 31451 12477
rect 33961 12474 34027 12477
rect 31385 12472 34027 12474
rect 31385 12416 31390 12472
rect 31446 12416 33966 12472
rect 34022 12416 34027 12472
rect 31385 12414 34027 12416
rect 31385 12411 31451 12414
rect 33961 12411 34027 12414
rect 21590 12278 22202 12338
rect 33777 12338 33843 12341
rect 50705 12338 50771 12341
rect 33777 12336 50771 12338
rect 33777 12280 33782 12336
rect 33838 12280 50710 12336
rect 50766 12280 50771 12336
rect 33777 12278 50771 12280
rect 9305 12275 9371 12278
rect 16849 12275 16915 12278
rect 33777 12275 33843 12278
rect 50705 12275 50771 12278
rect 0 12202 800 12232
rect 4061 12202 4127 12205
rect 0 12200 4127 12202
rect 0 12144 4066 12200
rect 4122 12144 4127 12200
rect 0 12142 4127 12144
rect 0 12112 800 12142
rect 4061 12139 4127 12142
rect 17309 12202 17375 12205
rect 23473 12202 23539 12205
rect 17309 12200 23539 12202
rect 17309 12144 17314 12200
rect 17370 12144 23478 12200
rect 23534 12144 23539 12200
rect 17309 12142 23539 12144
rect 17309 12139 17375 12142
rect 23473 12139 23539 12142
rect 18873 12066 18939 12069
rect 23657 12066 23723 12069
rect 18873 12064 23723 12066
rect 18873 12008 18878 12064
rect 18934 12008 23662 12064
rect 23718 12008 23723 12064
rect 18873 12006 23723 12008
rect 18873 12003 18939 12006
rect 23657 12003 23723 12006
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 32132 12000 32452 12001
rect 32132 11936 32140 12000
rect 32204 11936 32220 12000
rect 32284 11936 32300 12000
rect 32364 11936 32380 12000
rect 32444 11936 32452 12000
rect 32132 11935 32452 11936
rect 52924 12000 53244 12001
rect 52924 11936 52932 12000
rect 52996 11936 53012 12000
rect 53076 11936 53092 12000
rect 53156 11936 53172 12000
rect 53236 11936 53244 12000
rect 52924 11935 53244 11936
rect 18321 11930 18387 11933
rect 27429 11930 27495 11933
rect 18321 11928 27495 11930
rect 18321 11872 18326 11928
rect 18382 11872 27434 11928
rect 27490 11872 27495 11928
rect 18321 11870 27495 11872
rect 18321 11867 18387 11870
rect 27429 11867 27495 11870
rect 13721 11794 13787 11797
rect 56869 11794 56935 11797
rect 13721 11792 56935 11794
rect 13721 11736 13726 11792
rect 13782 11736 56874 11792
rect 56930 11736 56935 11792
rect 13721 11734 56935 11736
rect 13721 11731 13787 11734
rect 56869 11731 56935 11734
rect 21173 11658 21239 11661
rect 21725 11658 21791 11661
rect 23197 11658 23263 11661
rect 28257 11658 28323 11661
rect 21173 11656 28323 11658
rect 21173 11600 21178 11656
rect 21234 11600 21730 11656
rect 21786 11600 23202 11656
rect 23258 11600 28262 11656
rect 28318 11600 28323 11656
rect 21173 11598 28323 11600
rect 21173 11595 21239 11598
rect 21725 11595 21791 11598
rect 23197 11595 23263 11598
rect 28257 11595 28323 11598
rect 33041 11522 33107 11525
rect 37365 11522 37431 11525
rect 33041 11520 37431 11522
rect 33041 11464 33046 11520
rect 33102 11464 37370 11520
rect 37426 11464 37431 11520
rect 33041 11462 37431 11464
rect 33041 11459 33107 11462
rect 37365 11459 37431 11462
rect 21736 11456 22056 11457
rect 21736 11392 21744 11456
rect 21808 11392 21824 11456
rect 21888 11392 21904 11456
rect 21968 11392 21984 11456
rect 22048 11392 22056 11456
rect 21736 11391 22056 11392
rect 42528 11456 42848 11457
rect 42528 11392 42536 11456
rect 42600 11392 42616 11456
rect 42680 11392 42696 11456
rect 42760 11392 42776 11456
rect 42840 11392 42848 11456
rect 42528 11391 42848 11392
rect 22921 11250 22987 11253
rect 27797 11250 27863 11253
rect 22921 11248 27863 11250
rect 22921 11192 22926 11248
rect 22982 11192 27802 11248
rect 27858 11192 27863 11248
rect 22921 11190 27863 11192
rect 22921 11187 22987 11190
rect 27797 11187 27863 11190
rect 39757 11250 39823 11253
rect 43345 11250 43411 11253
rect 45645 11250 45711 11253
rect 39757 11248 45711 11250
rect 39757 11192 39762 11248
rect 39818 11192 43350 11248
rect 43406 11192 45650 11248
rect 45706 11192 45711 11248
rect 39757 11190 45711 11192
rect 39757 11187 39823 11190
rect 43345 11187 43411 11190
rect 45645 11187 45711 11190
rect 24117 11114 24183 11117
rect 27153 11114 27219 11117
rect 24117 11112 27219 11114
rect 24117 11056 24122 11112
rect 24178 11056 27158 11112
rect 27214 11056 27219 11112
rect 24117 11054 27219 11056
rect 24117 11051 24183 11054
rect 27153 11051 27219 11054
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 32132 10912 32452 10913
rect 32132 10848 32140 10912
rect 32204 10848 32220 10912
rect 32284 10848 32300 10912
rect 32364 10848 32380 10912
rect 32444 10848 32452 10912
rect 32132 10847 32452 10848
rect 52924 10912 53244 10913
rect 52924 10848 52932 10912
rect 52996 10848 53012 10912
rect 53076 10848 53092 10912
rect 53156 10848 53172 10912
rect 53236 10848 53244 10912
rect 52924 10847 53244 10848
rect 3969 10706 4035 10709
rect 8477 10706 8543 10709
rect 3969 10704 8543 10706
rect 3969 10648 3974 10704
rect 4030 10648 8482 10704
rect 8538 10648 8543 10704
rect 3969 10646 8543 10648
rect 3969 10643 4035 10646
rect 8477 10643 8543 10646
rect 23473 10706 23539 10709
rect 27245 10706 27311 10709
rect 23473 10704 27311 10706
rect 23473 10648 23478 10704
rect 23534 10648 27250 10704
rect 27306 10648 27311 10704
rect 23473 10646 27311 10648
rect 23473 10643 23539 10646
rect 27245 10643 27311 10646
rect 30097 10706 30163 10709
rect 38561 10706 38627 10709
rect 30097 10704 38627 10706
rect 30097 10648 30102 10704
rect 30158 10648 38566 10704
rect 38622 10648 38627 10704
rect 30097 10646 38627 10648
rect 30097 10643 30163 10646
rect 38561 10643 38627 10646
rect 20069 10570 20135 10573
rect 22277 10570 22343 10573
rect 20069 10568 22343 10570
rect 20069 10512 20074 10568
rect 20130 10512 22282 10568
rect 22338 10512 22343 10568
rect 20069 10510 22343 10512
rect 20069 10507 20135 10510
rect 22277 10507 22343 10510
rect 30465 10570 30531 10573
rect 32305 10570 32371 10573
rect 30465 10568 32371 10570
rect 30465 10512 30470 10568
rect 30526 10512 32310 10568
rect 32366 10512 32371 10568
rect 30465 10510 32371 10512
rect 30465 10507 30531 10510
rect 32305 10507 32371 10510
rect 38837 10570 38903 10573
rect 46933 10570 46999 10573
rect 38837 10568 46999 10570
rect 38837 10512 38842 10568
rect 38898 10512 46938 10568
rect 46994 10512 46999 10568
rect 38837 10510 46999 10512
rect 38837 10507 38903 10510
rect 46933 10507 46999 10510
rect 49509 10570 49575 10573
rect 50981 10570 51047 10573
rect 51717 10570 51783 10573
rect 49509 10568 51783 10570
rect 49509 10512 49514 10568
rect 49570 10512 50986 10568
rect 51042 10512 51722 10568
rect 51778 10512 51783 10568
rect 49509 10510 51783 10512
rect 49509 10507 49575 10510
rect 50981 10507 51047 10510
rect 51717 10507 51783 10510
rect 48681 10434 48747 10437
rect 52269 10434 52335 10437
rect 48681 10432 52335 10434
rect 48681 10376 48686 10432
rect 48742 10376 52274 10432
rect 52330 10376 52335 10432
rect 48681 10374 52335 10376
rect 48681 10371 48747 10374
rect 52269 10371 52335 10374
rect 21736 10368 22056 10369
rect 21736 10304 21744 10368
rect 21808 10304 21824 10368
rect 21888 10304 21904 10368
rect 21968 10304 21984 10368
rect 22048 10304 22056 10368
rect 21736 10303 22056 10304
rect 42528 10368 42848 10369
rect 42528 10304 42536 10368
rect 42600 10304 42616 10368
rect 42680 10304 42696 10368
rect 42760 10304 42776 10368
rect 42840 10304 42848 10368
rect 42528 10303 42848 10304
rect 20989 10162 21055 10165
rect 27705 10162 27771 10165
rect 20989 10160 27771 10162
rect 20989 10104 20994 10160
rect 21050 10104 27710 10160
rect 27766 10104 27771 10160
rect 20989 10102 27771 10104
rect 20989 10099 21055 10102
rect 27705 10099 27771 10102
rect 0 10026 800 10056
rect 3877 10026 3943 10029
rect 0 10024 3943 10026
rect 0 9968 3882 10024
rect 3938 9968 3943 10024
rect 0 9966 3943 9968
rect 0 9936 800 9966
rect 3877 9963 3943 9966
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 32132 9824 32452 9825
rect 32132 9760 32140 9824
rect 32204 9760 32220 9824
rect 32284 9760 32300 9824
rect 32364 9760 32380 9824
rect 32444 9760 32452 9824
rect 32132 9759 32452 9760
rect 52924 9824 53244 9825
rect 52924 9760 52932 9824
rect 52996 9760 53012 9824
rect 53076 9760 53092 9824
rect 53156 9760 53172 9824
rect 53236 9760 53244 9824
rect 52924 9759 53244 9760
rect 21081 9754 21147 9757
rect 23381 9754 23447 9757
rect 21081 9752 23447 9754
rect 21081 9696 21086 9752
rect 21142 9696 23386 9752
rect 23442 9696 23447 9752
rect 21081 9694 23447 9696
rect 21081 9691 21147 9694
rect 23381 9691 23447 9694
rect 16297 9618 16363 9621
rect 19241 9618 19307 9621
rect 16297 9616 19307 9618
rect 16297 9560 16302 9616
rect 16358 9560 19246 9616
rect 19302 9560 19307 9616
rect 16297 9558 19307 9560
rect 16297 9555 16363 9558
rect 19241 9555 19307 9558
rect 21725 9618 21791 9621
rect 23289 9618 23355 9621
rect 24945 9618 25011 9621
rect 21725 9616 25011 9618
rect 21725 9560 21730 9616
rect 21786 9560 23294 9616
rect 23350 9560 24950 9616
rect 25006 9560 25011 9616
rect 21725 9558 25011 9560
rect 21725 9555 21791 9558
rect 23289 9555 23355 9558
rect 24945 9555 25011 9558
rect 35985 9618 36051 9621
rect 37825 9618 37891 9621
rect 35985 9616 37891 9618
rect 35985 9560 35990 9616
rect 36046 9560 37830 9616
rect 37886 9560 37891 9616
rect 35985 9558 37891 9560
rect 35985 9555 36051 9558
rect 37825 9555 37891 9558
rect 41597 9618 41663 9621
rect 44173 9618 44239 9621
rect 47485 9618 47551 9621
rect 41597 9616 47551 9618
rect 41597 9560 41602 9616
rect 41658 9560 44178 9616
rect 44234 9560 47490 9616
rect 47546 9560 47551 9616
rect 41597 9558 47551 9560
rect 41597 9555 41663 9558
rect 44173 9555 44239 9558
rect 47485 9555 47551 9558
rect 21633 9482 21699 9485
rect 24117 9482 24183 9485
rect 21633 9480 24183 9482
rect 21633 9424 21638 9480
rect 21694 9424 24122 9480
rect 24178 9424 24183 9480
rect 21633 9422 24183 9424
rect 21633 9419 21699 9422
rect 24117 9419 24183 9422
rect 38837 9482 38903 9485
rect 47485 9482 47551 9485
rect 38837 9480 47551 9482
rect 38837 9424 38842 9480
rect 38898 9424 47490 9480
rect 47546 9424 47551 9480
rect 38837 9422 47551 9424
rect 38837 9419 38903 9422
rect 47485 9419 47551 9422
rect 50245 9482 50311 9485
rect 51717 9482 51783 9485
rect 50245 9480 51783 9482
rect 50245 9424 50250 9480
rect 50306 9424 51722 9480
rect 51778 9424 51783 9480
rect 50245 9422 51783 9424
rect 50245 9419 50311 9422
rect 51717 9419 51783 9422
rect 21736 9280 22056 9281
rect 21736 9216 21744 9280
rect 21808 9216 21824 9280
rect 21888 9216 21904 9280
rect 21968 9216 21984 9280
rect 22048 9216 22056 9280
rect 21736 9215 22056 9216
rect 42528 9280 42848 9281
rect 42528 9216 42536 9280
rect 42600 9216 42616 9280
rect 42680 9216 42696 9280
rect 42760 9216 42776 9280
rect 42840 9216 42848 9280
rect 42528 9215 42848 9216
rect 30281 9074 30347 9077
rect 31017 9074 31083 9077
rect 32397 9074 32463 9077
rect 30281 9072 32463 9074
rect 30281 9016 30286 9072
rect 30342 9016 31022 9072
rect 31078 9016 32402 9072
rect 32458 9016 32463 9072
rect 30281 9014 32463 9016
rect 30281 9011 30347 9014
rect 31017 9011 31083 9014
rect 32397 9011 32463 9014
rect 41045 9074 41111 9077
rect 41965 9074 42031 9077
rect 41045 9072 42031 9074
rect 41045 9016 41050 9072
rect 41106 9016 41970 9072
rect 42026 9016 42031 9072
rect 41045 9014 42031 9016
rect 41045 9011 41111 9014
rect 41965 9011 42031 9014
rect 11145 8938 11211 8941
rect 17493 8938 17559 8941
rect 11145 8936 17559 8938
rect 11145 8880 11150 8936
rect 11206 8880 17498 8936
rect 17554 8880 17559 8936
rect 11145 8878 17559 8880
rect 11145 8875 11211 8878
rect 17493 8875 17559 8878
rect 21081 8938 21147 8941
rect 28533 8938 28599 8941
rect 21081 8936 28599 8938
rect 21081 8880 21086 8936
rect 21142 8880 28538 8936
rect 28594 8880 28599 8936
rect 21081 8878 28599 8880
rect 21081 8875 21147 8878
rect 28533 8875 28599 8878
rect 51257 8938 51323 8941
rect 56501 8938 56567 8941
rect 51257 8936 56567 8938
rect 51257 8880 51262 8936
rect 51318 8880 56506 8936
rect 56562 8880 56567 8936
rect 51257 8878 56567 8880
rect 51257 8875 51323 8878
rect 56501 8875 56567 8878
rect 22001 8802 22067 8805
rect 22553 8802 22619 8805
rect 22001 8800 22619 8802
rect 22001 8744 22006 8800
rect 22062 8744 22558 8800
rect 22614 8744 22619 8800
rect 22001 8742 22619 8744
rect 22001 8739 22067 8742
rect 22553 8739 22619 8742
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 32132 8736 32452 8737
rect 32132 8672 32140 8736
rect 32204 8672 32220 8736
rect 32284 8672 32300 8736
rect 32364 8672 32380 8736
rect 32444 8672 32452 8736
rect 32132 8671 32452 8672
rect 52924 8736 53244 8737
rect 52924 8672 52932 8736
rect 52996 8672 53012 8736
rect 53076 8672 53092 8736
rect 53156 8672 53172 8736
rect 53236 8672 53244 8736
rect 52924 8671 53244 8672
rect 11881 8666 11947 8669
rect 18689 8666 18755 8669
rect 11881 8664 18755 8666
rect 11881 8608 11886 8664
rect 11942 8608 18694 8664
rect 18750 8608 18755 8664
rect 11881 8606 18755 8608
rect 11881 8603 11947 8606
rect 18689 8603 18755 8606
rect 17217 8530 17283 8533
rect 17769 8530 17835 8533
rect 21725 8530 21791 8533
rect 17217 8528 21791 8530
rect 17217 8472 17222 8528
rect 17278 8472 17774 8528
rect 17830 8472 21730 8528
rect 21786 8472 21791 8528
rect 17217 8470 21791 8472
rect 17217 8467 17283 8470
rect 17769 8467 17835 8470
rect 21725 8467 21791 8470
rect 24761 8530 24827 8533
rect 27889 8530 27955 8533
rect 24761 8528 27955 8530
rect 24761 8472 24766 8528
rect 24822 8472 27894 8528
rect 27950 8472 27955 8528
rect 24761 8470 27955 8472
rect 24761 8467 24827 8470
rect 27889 8467 27955 8470
rect 6637 8394 6703 8397
rect 33869 8394 33935 8397
rect 6637 8392 33935 8394
rect 6637 8336 6642 8392
rect 6698 8336 33874 8392
rect 33930 8336 33935 8392
rect 6637 8334 33935 8336
rect 6637 8331 6703 8334
rect 33869 8331 33935 8334
rect 40309 8394 40375 8397
rect 47209 8394 47275 8397
rect 40309 8392 47275 8394
rect 40309 8336 40314 8392
rect 40370 8336 47214 8392
rect 47270 8336 47275 8392
rect 40309 8334 47275 8336
rect 40309 8331 40375 8334
rect 47209 8331 47275 8334
rect 48497 8394 48563 8397
rect 49509 8394 49575 8397
rect 48497 8392 49575 8394
rect 48497 8336 48502 8392
rect 48558 8336 49514 8392
rect 49570 8336 49575 8392
rect 48497 8334 49575 8336
rect 48497 8331 48563 8334
rect 49509 8331 49575 8334
rect 24945 8258 25011 8261
rect 28942 8258 28948 8260
rect 24945 8256 28948 8258
rect 24945 8200 24950 8256
rect 25006 8200 28948 8256
rect 24945 8198 28948 8200
rect 24945 8195 25011 8198
rect 28942 8196 28948 8198
rect 29012 8196 29018 8260
rect 29545 8258 29611 8261
rect 40861 8258 40927 8261
rect 29545 8256 40927 8258
rect 29545 8200 29550 8256
rect 29606 8200 40866 8256
rect 40922 8200 40927 8256
rect 29545 8198 40927 8200
rect 29545 8195 29611 8198
rect 40861 8195 40927 8198
rect 21736 8192 22056 8193
rect 21736 8128 21744 8192
rect 21808 8128 21824 8192
rect 21888 8128 21904 8192
rect 21968 8128 21984 8192
rect 22048 8128 22056 8192
rect 21736 8127 22056 8128
rect 42528 8192 42848 8193
rect 42528 8128 42536 8192
rect 42600 8128 42616 8192
rect 42680 8128 42696 8192
rect 42760 8128 42776 8192
rect 42840 8128 42848 8192
rect 42528 8127 42848 8128
rect 33777 8122 33843 8125
rect 35433 8122 35499 8125
rect 26926 8120 35499 8122
rect 26926 8064 33782 8120
rect 33838 8064 35438 8120
rect 35494 8064 35499 8120
rect 26926 8062 35499 8064
rect 7557 7986 7623 7989
rect 26926 7986 26986 8062
rect 33777 8059 33843 8062
rect 35433 8059 35499 8062
rect 35617 8122 35683 8125
rect 38377 8122 38443 8125
rect 35617 8120 38443 8122
rect 35617 8064 35622 8120
rect 35678 8064 38382 8120
rect 38438 8064 38443 8120
rect 35617 8062 38443 8064
rect 35617 8059 35683 8062
rect 38377 8059 38443 8062
rect 47669 8122 47735 8125
rect 48221 8122 48287 8125
rect 47669 8120 48287 8122
rect 47669 8064 47674 8120
rect 47730 8064 48226 8120
rect 48282 8064 48287 8120
rect 47669 8062 48287 8064
rect 47669 8059 47735 8062
rect 48221 8059 48287 8062
rect 35249 7986 35315 7989
rect 7557 7984 26986 7986
rect 7557 7928 7562 7984
rect 7618 7928 26986 7984
rect 7557 7926 26986 7928
rect 27110 7984 35315 7986
rect 27110 7928 35254 7984
rect 35310 7928 35315 7984
rect 27110 7926 35315 7928
rect 7557 7923 7623 7926
rect 0 7850 800 7880
rect 3877 7850 3943 7853
rect 27110 7850 27170 7926
rect 35249 7923 35315 7926
rect 43253 7986 43319 7989
rect 49141 7986 49207 7989
rect 43253 7984 49207 7986
rect 43253 7928 43258 7984
rect 43314 7928 49146 7984
rect 49202 7928 49207 7984
rect 43253 7926 49207 7928
rect 43253 7923 43319 7926
rect 49141 7923 49207 7926
rect 49785 7986 49851 7989
rect 51993 7986 52059 7989
rect 49785 7984 52059 7986
rect 49785 7928 49790 7984
rect 49846 7928 51998 7984
rect 52054 7928 52059 7984
rect 49785 7926 52059 7928
rect 49785 7923 49851 7926
rect 51993 7923 52059 7926
rect 52545 7986 52611 7989
rect 56685 7986 56751 7989
rect 52545 7984 56751 7986
rect 52545 7928 52550 7984
rect 52606 7928 56690 7984
rect 56746 7928 56751 7984
rect 52545 7926 56751 7928
rect 52545 7923 52611 7926
rect 56685 7923 56751 7926
rect 0 7790 3802 7850
rect 0 7760 800 7790
rect 3742 7306 3802 7790
rect 3877 7848 27170 7850
rect 3877 7792 3882 7848
rect 3938 7792 27170 7848
rect 3877 7790 27170 7792
rect 29085 7850 29151 7853
rect 29913 7850 29979 7853
rect 40861 7850 40927 7853
rect 51809 7850 51875 7853
rect 56133 7850 56199 7853
rect 57421 7850 57487 7853
rect 29085 7848 29979 7850
rect 29085 7792 29090 7848
rect 29146 7792 29918 7848
rect 29974 7792 29979 7848
rect 29085 7790 29979 7792
rect 3877 7787 3943 7790
rect 29085 7787 29151 7790
rect 29913 7787 29979 7790
rect 31940 7790 32644 7850
rect 15285 7714 15351 7717
rect 16849 7714 16915 7717
rect 17493 7714 17559 7717
rect 15285 7712 17559 7714
rect 15285 7656 15290 7712
rect 15346 7656 16854 7712
rect 16910 7656 17498 7712
rect 17554 7656 17559 7712
rect 15285 7654 17559 7656
rect 15285 7651 15351 7654
rect 16849 7651 16915 7654
rect 17493 7651 17559 7654
rect 20161 7714 20227 7717
rect 22093 7714 22159 7717
rect 20161 7712 22159 7714
rect 20161 7656 20166 7712
rect 20222 7656 22098 7712
rect 22154 7656 22159 7712
rect 20161 7654 22159 7656
rect 20161 7651 20227 7654
rect 22093 7651 22159 7654
rect 25037 7714 25103 7717
rect 29545 7714 29611 7717
rect 25037 7712 29611 7714
rect 25037 7656 25042 7712
rect 25098 7656 29550 7712
rect 29606 7656 29611 7712
rect 25037 7654 29611 7656
rect 25037 7651 25103 7654
rect 29545 7651 29611 7654
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 11881 7578 11947 7581
rect 16941 7578 17007 7581
rect 11881 7576 17007 7578
rect 11881 7520 11886 7576
rect 11942 7520 16946 7576
rect 17002 7520 17007 7576
rect 11881 7518 17007 7520
rect 11881 7515 11947 7518
rect 16941 7515 17007 7518
rect 19793 7578 19859 7581
rect 31940 7578 32000 7790
rect 32584 7714 32644 7790
rect 40861 7848 57487 7850
rect 40861 7792 40866 7848
rect 40922 7792 51814 7848
rect 51870 7792 56138 7848
rect 56194 7792 57426 7848
rect 57482 7792 57487 7848
rect 40861 7790 57487 7792
rect 40861 7787 40927 7790
rect 51809 7787 51875 7790
rect 56133 7787 56199 7790
rect 57421 7787 57487 7790
rect 46197 7714 46263 7717
rect 47301 7714 47367 7717
rect 32584 7712 47367 7714
rect 32584 7656 46202 7712
rect 46258 7656 47306 7712
rect 47362 7656 47367 7712
rect 32584 7654 47367 7656
rect 46197 7651 46263 7654
rect 47301 7651 47367 7654
rect 50705 7714 50771 7717
rect 52177 7714 52243 7717
rect 50705 7712 52243 7714
rect 50705 7656 50710 7712
rect 50766 7656 52182 7712
rect 52238 7656 52243 7712
rect 50705 7654 52243 7656
rect 50705 7651 50771 7654
rect 52177 7651 52243 7654
rect 32132 7648 32452 7649
rect 32132 7584 32140 7648
rect 32204 7584 32220 7648
rect 32284 7584 32300 7648
rect 32364 7584 32380 7648
rect 32444 7584 32452 7648
rect 32132 7583 32452 7584
rect 52924 7648 53244 7649
rect 52924 7584 52932 7648
rect 52996 7584 53012 7648
rect 53076 7584 53092 7648
rect 53156 7584 53172 7648
rect 53236 7584 53244 7648
rect 52924 7583 53244 7584
rect 19793 7576 32000 7578
rect 19793 7520 19798 7576
rect 19854 7520 32000 7576
rect 19793 7518 32000 7520
rect 19793 7515 19859 7518
rect 6269 7442 6335 7445
rect 36905 7442 36971 7445
rect 53005 7442 53071 7445
rect 6269 7440 53071 7442
rect 6269 7384 6274 7440
rect 6330 7384 36910 7440
rect 36966 7384 53010 7440
rect 53066 7384 53071 7440
rect 6269 7382 53071 7384
rect 6269 7379 6335 7382
rect 36905 7379 36971 7382
rect 53005 7379 53071 7382
rect 36629 7306 36695 7309
rect 3742 7304 36695 7306
rect 3742 7248 36634 7304
rect 36690 7248 36695 7304
rect 3742 7246 36695 7248
rect 36629 7243 36695 7246
rect 46105 7306 46171 7309
rect 48129 7306 48195 7309
rect 46105 7304 48195 7306
rect 46105 7248 46110 7304
rect 46166 7248 48134 7304
rect 48190 7248 48195 7304
rect 46105 7246 48195 7248
rect 46105 7243 46171 7246
rect 48129 7243 48195 7246
rect 26325 7170 26391 7173
rect 26877 7170 26943 7173
rect 26325 7168 26943 7170
rect 26325 7112 26330 7168
rect 26386 7112 26882 7168
rect 26938 7112 26943 7168
rect 26325 7110 26943 7112
rect 26325 7107 26391 7110
rect 26877 7107 26943 7110
rect 28993 7170 29059 7173
rect 32397 7170 32463 7173
rect 28993 7168 32463 7170
rect 28993 7112 28998 7168
rect 29054 7112 32402 7168
rect 32458 7112 32463 7168
rect 28993 7110 32463 7112
rect 28993 7107 29059 7110
rect 32397 7107 32463 7110
rect 21736 7104 22056 7105
rect 21736 7040 21744 7104
rect 21808 7040 21824 7104
rect 21888 7040 21904 7104
rect 21968 7040 21984 7104
rect 22048 7040 22056 7104
rect 21736 7039 22056 7040
rect 42528 7104 42848 7105
rect 42528 7040 42536 7104
rect 42600 7040 42616 7104
rect 42680 7040 42696 7104
rect 42760 7040 42776 7104
rect 42840 7040 42848 7104
rect 42528 7039 42848 7040
rect 25773 7034 25839 7037
rect 26417 7034 26483 7037
rect 27797 7034 27863 7037
rect 25773 7032 27863 7034
rect 25773 6976 25778 7032
rect 25834 6976 26422 7032
rect 26478 6976 27802 7032
rect 27858 6976 27863 7032
rect 25773 6974 27863 6976
rect 25773 6971 25839 6974
rect 26417 6971 26483 6974
rect 27797 6971 27863 6974
rect 27981 7034 28047 7037
rect 29085 7034 29151 7037
rect 27981 7032 29151 7034
rect 27981 6976 27986 7032
rect 28042 6976 29090 7032
rect 29146 6976 29151 7032
rect 27981 6974 29151 6976
rect 27981 6971 28047 6974
rect 29085 6971 29151 6974
rect 31385 7034 31451 7037
rect 36537 7034 36603 7037
rect 31385 7032 36603 7034
rect 31385 6976 31390 7032
rect 31446 6976 36542 7032
rect 36598 6976 36603 7032
rect 31385 6974 36603 6976
rect 31385 6971 31451 6974
rect 36537 6971 36603 6974
rect 22553 6898 22619 6901
rect 37917 6898 37983 6901
rect 38653 6898 38719 6901
rect 19382 6896 38719 6898
rect 19382 6840 22558 6896
rect 22614 6840 37922 6896
rect 37978 6840 38658 6896
rect 38714 6840 38719 6896
rect 19382 6838 38719 6840
rect 19382 6765 19442 6838
rect 22553 6835 22619 6838
rect 37917 6835 37983 6838
rect 38653 6835 38719 6838
rect 41045 6898 41111 6901
rect 46933 6898 46999 6901
rect 41045 6896 46999 6898
rect 41045 6840 41050 6896
rect 41106 6840 46938 6896
rect 46994 6840 46999 6896
rect 41045 6838 46999 6840
rect 41045 6835 41111 6838
rect 46933 6835 46999 6838
rect 48405 6898 48471 6901
rect 54937 6898 55003 6901
rect 48405 6896 55003 6898
rect 48405 6840 48410 6896
rect 48466 6840 54942 6896
rect 54998 6840 55003 6896
rect 48405 6838 55003 6840
rect 48405 6835 48471 6838
rect 54937 6835 55003 6838
rect 19333 6760 19442 6765
rect 19333 6704 19338 6760
rect 19394 6704 19442 6760
rect 19333 6702 19442 6704
rect 21817 6762 21883 6765
rect 43437 6762 43503 6765
rect 21817 6760 43503 6762
rect 21817 6704 21822 6760
rect 21878 6704 43442 6760
rect 43498 6704 43503 6760
rect 21817 6702 43503 6704
rect 19333 6699 19399 6702
rect 21817 6699 21883 6702
rect 43437 6699 43503 6702
rect 43897 6626 43963 6629
rect 46790 6626 46796 6628
rect 43897 6624 46796 6626
rect 43897 6568 43902 6624
rect 43958 6568 46796 6624
rect 43897 6566 46796 6568
rect 43897 6563 43963 6566
rect 46790 6564 46796 6566
rect 46860 6564 46866 6628
rect 49049 6626 49115 6629
rect 51533 6626 51599 6629
rect 49049 6624 51599 6626
rect 49049 6568 49054 6624
rect 49110 6568 51538 6624
rect 51594 6568 51599 6624
rect 49049 6566 51599 6568
rect 49049 6563 49115 6566
rect 51533 6563 51599 6566
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 32132 6560 32452 6561
rect 32132 6496 32140 6560
rect 32204 6496 32220 6560
rect 32284 6496 32300 6560
rect 32364 6496 32380 6560
rect 32444 6496 32452 6560
rect 32132 6495 32452 6496
rect 52924 6560 53244 6561
rect 52924 6496 52932 6560
rect 52996 6496 53012 6560
rect 53076 6496 53092 6560
rect 53156 6496 53172 6560
rect 53236 6496 53244 6560
rect 52924 6495 53244 6496
rect 16757 6490 16823 6493
rect 27245 6490 27311 6493
rect 47025 6490 47091 6493
rect 16757 6488 32000 6490
rect 16757 6432 16762 6488
rect 16818 6432 27250 6488
rect 27306 6432 32000 6488
rect 16757 6430 32000 6432
rect 16757 6427 16823 6430
rect 27245 6427 27311 6430
rect 19885 6354 19951 6357
rect 25589 6354 25655 6357
rect 27153 6354 27219 6357
rect 19885 6352 27219 6354
rect 19885 6296 19890 6352
rect 19946 6296 25594 6352
rect 25650 6296 27158 6352
rect 27214 6296 27219 6352
rect 19885 6294 27219 6296
rect 19885 6291 19951 6294
rect 25589 6291 25655 6294
rect 27153 6291 27219 6294
rect 28717 6354 28783 6357
rect 31477 6354 31543 6357
rect 28717 6352 31543 6354
rect 28717 6296 28722 6352
rect 28778 6296 31482 6352
rect 31538 6296 31543 6352
rect 28717 6294 31543 6296
rect 31940 6354 32000 6430
rect 33872 6488 47091 6490
rect 33872 6432 47030 6488
rect 47086 6432 47091 6488
rect 33872 6430 47091 6432
rect 33872 6357 33932 6430
rect 47025 6427 47091 6430
rect 50429 6490 50495 6493
rect 50797 6490 50863 6493
rect 50429 6488 50863 6490
rect 50429 6432 50434 6488
rect 50490 6432 50802 6488
rect 50858 6432 50863 6488
rect 50429 6430 50863 6432
rect 50429 6427 50495 6430
rect 50797 6427 50863 6430
rect 33869 6354 33935 6357
rect 31940 6352 33935 6354
rect 31940 6296 33874 6352
rect 33930 6296 33935 6352
rect 31940 6294 33935 6296
rect 28717 6291 28783 6294
rect 31477 6291 31543 6294
rect 33869 6291 33935 6294
rect 35617 6354 35683 6357
rect 55673 6354 55739 6357
rect 35617 6352 55739 6354
rect 35617 6296 35622 6352
rect 35678 6296 55678 6352
rect 55734 6296 55739 6352
rect 35617 6294 55739 6296
rect 35617 6291 35683 6294
rect 55673 6291 55739 6294
rect 13445 6218 13511 6221
rect 34237 6218 34303 6221
rect 13445 6216 34303 6218
rect 13445 6160 13450 6216
rect 13506 6160 34242 6216
rect 34298 6160 34303 6216
rect 13445 6158 34303 6160
rect 13445 6155 13511 6158
rect 34237 6155 34303 6158
rect 41873 6218 41939 6221
rect 44817 6218 44883 6221
rect 41873 6216 44883 6218
rect 41873 6160 41878 6216
rect 41934 6160 44822 6216
rect 44878 6160 44883 6216
rect 41873 6158 44883 6160
rect 41873 6155 41939 6158
rect 44817 6155 44883 6158
rect 48773 6218 48839 6221
rect 51901 6218 51967 6221
rect 48773 6216 51967 6218
rect 48773 6160 48778 6216
rect 48834 6160 51906 6216
rect 51962 6160 51967 6216
rect 48773 6158 51967 6160
rect 48773 6155 48839 6158
rect 51901 6155 51967 6158
rect 53005 6218 53071 6221
rect 55029 6218 55095 6221
rect 53005 6216 55095 6218
rect 53005 6160 53010 6216
rect 53066 6160 55034 6216
rect 55090 6160 55095 6216
rect 53005 6158 55095 6160
rect 53005 6155 53071 6158
rect 55029 6155 55095 6158
rect 10961 6082 11027 6085
rect 19241 6082 19307 6085
rect 10961 6080 19307 6082
rect 10961 6024 10966 6080
rect 11022 6024 19246 6080
rect 19302 6024 19307 6080
rect 10961 6022 19307 6024
rect 10961 6019 11027 6022
rect 19241 6019 19307 6022
rect 23105 6082 23171 6085
rect 24393 6082 24459 6085
rect 31477 6082 31543 6085
rect 31661 6082 31727 6085
rect 31937 6082 32003 6085
rect 23105 6080 31586 6082
rect 23105 6024 23110 6080
rect 23166 6024 24398 6080
rect 24454 6024 31482 6080
rect 31538 6024 31586 6080
rect 23105 6022 31586 6024
rect 23105 6019 23171 6022
rect 24393 6019 24459 6022
rect 31477 6019 31586 6022
rect 31661 6080 32003 6082
rect 31661 6024 31666 6080
rect 31722 6024 31942 6080
rect 31998 6024 32003 6080
rect 31661 6022 32003 6024
rect 31661 6019 31727 6022
rect 31937 6019 32003 6022
rect 40493 6082 40559 6085
rect 41689 6082 41755 6085
rect 42241 6082 42307 6085
rect 40493 6080 42307 6082
rect 40493 6024 40498 6080
rect 40554 6024 41694 6080
rect 41750 6024 42246 6080
rect 42302 6024 42307 6080
rect 40493 6022 42307 6024
rect 40493 6019 40559 6022
rect 41689 6019 41755 6022
rect 42241 6019 42307 6022
rect 21736 6016 22056 6017
rect 21736 5952 21744 6016
rect 21808 5952 21824 6016
rect 21888 5952 21904 6016
rect 21968 5952 21984 6016
rect 22048 5952 22056 6016
rect 21736 5951 22056 5952
rect 24209 5946 24275 5949
rect 27797 5946 27863 5949
rect 24209 5944 27863 5946
rect 24209 5888 24214 5944
rect 24270 5888 27802 5944
rect 27858 5888 27863 5944
rect 24209 5886 27863 5888
rect 24209 5883 24275 5886
rect 27797 5883 27863 5886
rect 29085 5946 29151 5949
rect 31385 5946 31451 5949
rect 29085 5944 31451 5946
rect 29085 5888 29090 5944
rect 29146 5888 31390 5944
rect 31446 5888 31451 5944
rect 29085 5886 31451 5888
rect 31526 5946 31586 6019
rect 42528 6016 42848 6017
rect 42528 5952 42536 6016
rect 42600 5952 42616 6016
rect 42680 5952 42696 6016
rect 42760 5952 42776 6016
rect 42840 5952 42848 6016
rect 42528 5951 42848 5952
rect 32029 5946 32095 5949
rect 31526 5944 32095 5946
rect 31526 5888 32034 5944
rect 32090 5888 32095 5944
rect 31526 5886 32095 5888
rect 29085 5883 29151 5886
rect 31385 5883 31451 5886
rect 32029 5883 32095 5886
rect 46790 5884 46796 5948
rect 46860 5946 46866 5948
rect 59997 5946 60063 5949
rect 46860 5944 60063 5946
rect 46860 5888 60002 5944
rect 60058 5888 60063 5944
rect 46860 5886 60063 5888
rect 46860 5884 46866 5886
rect 59997 5883 60063 5886
rect 21265 5810 21331 5813
rect 46422 5810 46428 5812
rect 21265 5808 46428 5810
rect 21265 5752 21270 5808
rect 21326 5752 46428 5808
rect 21265 5750 46428 5752
rect 21265 5747 21331 5750
rect 46422 5748 46428 5750
rect 46492 5748 46498 5812
rect 46790 5748 46796 5812
rect 46860 5810 46866 5812
rect 49141 5810 49207 5813
rect 46860 5808 49207 5810
rect 46860 5752 49146 5808
rect 49202 5752 49207 5808
rect 46860 5750 49207 5752
rect 46860 5748 46866 5750
rect 49141 5747 49207 5750
rect 20161 5674 20227 5677
rect 23197 5674 23263 5677
rect 20161 5672 23263 5674
rect 20161 5616 20166 5672
rect 20222 5616 23202 5672
rect 23258 5616 23263 5672
rect 20161 5614 23263 5616
rect 20161 5611 20227 5614
rect 23197 5611 23263 5614
rect 23933 5674 23999 5677
rect 26693 5674 26759 5677
rect 23933 5672 26759 5674
rect 23933 5616 23938 5672
rect 23994 5616 26698 5672
rect 26754 5616 26759 5672
rect 23933 5614 26759 5616
rect 23933 5611 23999 5614
rect 26693 5611 26759 5614
rect 31940 5643 56610 5674
rect 31940 5638 56659 5643
rect 31940 5614 56598 5638
rect 0 5538 800 5568
rect 4061 5538 4127 5541
rect 0 5536 4127 5538
rect 0 5480 4066 5536
rect 4122 5480 4127 5536
rect 0 5478 4127 5480
rect 0 5448 800 5478
rect 4061 5475 4127 5478
rect 16205 5538 16271 5541
rect 27521 5538 27587 5541
rect 31940 5538 32000 5614
rect 56550 5582 56598 5614
rect 56654 5582 56659 5638
rect 56550 5580 56659 5582
rect 56593 5577 56659 5580
rect 16205 5536 32000 5538
rect 16205 5480 16210 5536
rect 16266 5480 27526 5536
rect 27582 5480 32000 5536
rect 16205 5478 32000 5480
rect 39021 5538 39087 5541
rect 46289 5538 46355 5541
rect 39021 5536 46355 5538
rect 39021 5480 39026 5536
rect 39082 5480 46294 5536
rect 46350 5480 46355 5536
rect 39021 5478 46355 5480
rect 16205 5475 16271 5478
rect 27521 5475 27587 5478
rect 39021 5475 39087 5478
rect 46289 5475 46355 5478
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 32132 5472 32452 5473
rect 32132 5408 32140 5472
rect 32204 5408 32220 5472
rect 32284 5408 32300 5472
rect 32364 5408 32380 5472
rect 32444 5408 32452 5472
rect 32132 5407 32452 5408
rect 52924 5472 53244 5473
rect 52924 5408 52932 5472
rect 52996 5408 53012 5472
rect 53076 5408 53092 5472
rect 53156 5408 53172 5472
rect 53236 5408 53244 5472
rect 52924 5407 53244 5408
rect 15653 5402 15719 5405
rect 21173 5402 21239 5405
rect 15653 5400 21239 5402
rect 15653 5344 15658 5400
rect 15714 5344 21178 5400
rect 21234 5344 21239 5400
rect 15653 5342 21239 5344
rect 15653 5339 15719 5342
rect 21173 5339 21239 5342
rect 21909 5402 21975 5405
rect 22185 5402 22251 5405
rect 21909 5400 22251 5402
rect 21909 5344 21914 5400
rect 21970 5344 22190 5400
rect 22246 5344 22251 5400
rect 21909 5342 22251 5344
rect 21909 5339 21975 5342
rect 22185 5339 22251 5342
rect 22369 5402 22435 5405
rect 27981 5402 28047 5405
rect 28993 5404 29059 5405
rect 22369 5400 28047 5402
rect 22369 5344 22374 5400
rect 22430 5344 27986 5400
rect 28042 5344 28047 5400
rect 22369 5342 28047 5344
rect 22369 5339 22435 5342
rect 27981 5339 28047 5342
rect 28942 5340 28948 5404
rect 29012 5402 29059 5404
rect 29545 5402 29611 5405
rect 29012 5400 29611 5402
rect 29054 5344 29550 5400
rect 29606 5344 29611 5400
rect 29012 5342 29611 5344
rect 29012 5340 29059 5342
rect 28993 5339 29059 5340
rect 29545 5339 29611 5342
rect 33041 5402 33107 5405
rect 40953 5402 41019 5405
rect 33041 5400 41019 5402
rect 33041 5344 33046 5400
rect 33102 5344 40958 5400
rect 41014 5344 41019 5400
rect 33041 5342 41019 5344
rect 33041 5339 33107 5342
rect 40953 5339 41019 5342
rect 30373 5266 30439 5269
rect 27110 5264 30439 5266
rect 27110 5208 30378 5264
rect 30434 5208 30439 5264
rect 27110 5206 30439 5208
rect 8293 5130 8359 5133
rect 11881 5130 11947 5133
rect 8293 5128 11947 5130
rect 8293 5072 8298 5128
rect 8354 5072 11886 5128
rect 11942 5072 11947 5128
rect 8293 5070 11947 5072
rect 8293 5067 8359 5070
rect 11881 5067 11947 5070
rect 12157 5130 12223 5133
rect 19149 5130 19215 5133
rect 12157 5128 19215 5130
rect 12157 5072 12162 5128
rect 12218 5072 19154 5128
rect 19210 5072 19215 5128
rect 12157 5070 19215 5072
rect 12157 5067 12223 5070
rect 19149 5067 19215 5070
rect 20437 5130 20503 5133
rect 24485 5130 24551 5133
rect 20437 5128 24551 5130
rect 20437 5072 20442 5128
rect 20498 5072 24490 5128
rect 24546 5072 24551 5128
rect 20437 5070 24551 5072
rect 20437 5067 20503 5070
rect 24485 5067 24551 5070
rect 24669 5130 24735 5133
rect 27110 5130 27170 5206
rect 30373 5203 30439 5206
rect 32029 5266 32095 5269
rect 55305 5266 55371 5269
rect 56409 5266 56475 5269
rect 32029 5264 56475 5266
rect 32029 5208 32034 5264
rect 32090 5208 55310 5264
rect 55366 5208 56414 5264
rect 56470 5208 56475 5264
rect 32029 5206 56475 5208
rect 32029 5203 32095 5206
rect 55305 5203 55371 5206
rect 56409 5203 56475 5206
rect 24669 5128 27170 5130
rect 24669 5072 24674 5128
rect 24730 5072 27170 5128
rect 24669 5070 27170 5072
rect 27245 5130 27311 5133
rect 50889 5130 50955 5133
rect 27245 5128 50955 5130
rect 27245 5072 27250 5128
rect 27306 5072 50894 5128
rect 50950 5072 50955 5128
rect 27245 5070 50955 5072
rect 24669 5067 24735 5070
rect 27245 5067 27311 5070
rect 50889 5067 50955 5070
rect 2773 4994 2839 4997
rect 5809 4994 5875 4997
rect 8937 4994 9003 4997
rect 2773 4992 9003 4994
rect 2773 4936 2778 4992
rect 2834 4936 5814 4992
rect 5870 4936 8942 4992
rect 8998 4936 9003 4992
rect 2773 4934 9003 4936
rect 2773 4931 2839 4934
rect 5809 4931 5875 4934
rect 8937 4931 9003 4934
rect 29729 4994 29795 4997
rect 30649 4994 30715 4997
rect 29729 4992 30715 4994
rect 29729 4936 29734 4992
rect 29790 4936 30654 4992
rect 30710 4936 30715 4992
rect 29729 4934 30715 4936
rect 29729 4931 29795 4934
rect 30649 4931 30715 4934
rect 31201 4994 31267 4997
rect 31937 4994 32003 4997
rect 40677 4994 40743 4997
rect 31201 4992 32003 4994
rect 31201 4936 31206 4992
rect 31262 4936 31942 4992
rect 31998 4936 32003 4992
rect 31201 4934 32003 4936
rect 31201 4931 31267 4934
rect 31937 4931 32003 4934
rect 32078 4992 40743 4994
rect 32078 4936 40682 4992
rect 40738 4936 40743 4992
rect 32078 4934 40743 4936
rect 21736 4928 22056 4929
rect 21736 4864 21744 4928
rect 21808 4864 21824 4928
rect 21888 4864 21904 4928
rect 21968 4864 21984 4928
rect 22048 4864 22056 4928
rect 21736 4863 22056 4864
rect 10133 4858 10199 4861
rect 16573 4858 16639 4861
rect 19701 4858 19767 4861
rect 10133 4856 19767 4858
rect 10133 4800 10138 4856
rect 10194 4800 16578 4856
rect 16634 4800 19706 4856
rect 19762 4800 19767 4856
rect 10133 4798 19767 4800
rect 10133 4795 10199 4798
rect 16573 4795 16639 4798
rect 19701 4795 19767 4798
rect 25497 4858 25563 4861
rect 25865 4858 25931 4861
rect 32078 4858 32138 4934
rect 40677 4931 40743 4934
rect 42528 4928 42848 4929
rect 42528 4864 42536 4928
rect 42600 4864 42616 4928
rect 42680 4864 42696 4928
rect 42760 4864 42776 4928
rect 42840 4864 42848 4928
rect 42528 4863 42848 4864
rect 25497 4856 32138 4858
rect 25497 4800 25502 4856
rect 25558 4800 25870 4856
rect 25926 4800 32138 4856
rect 25497 4798 32138 4800
rect 32305 4858 32371 4861
rect 40309 4858 40375 4861
rect 32305 4856 40375 4858
rect 32305 4800 32310 4856
rect 32366 4800 40314 4856
rect 40370 4800 40375 4856
rect 32305 4798 40375 4800
rect 25497 4795 25563 4798
rect 25865 4795 25931 4798
rect 32305 4795 32371 4798
rect 40309 4795 40375 4798
rect 4521 4722 4587 4725
rect 24945 4722 25011 4725
rect 4521 4720 25011 4722
rect 4521 4664 4526 4720
rect 4582 4664 24950 4720
rect 25006 4664 25011 4720
rect 4521 4662 25011 4664
rect 4521 4659 4587 4662
rect 24945 4659 25011 4662
rect 28901 4722 28967 4725
rect 31569 4722 31635 4725
rect 28901 4720 31635 4722
rect 28901 4664 28906 4720
rect 28962 4664 31574 4720
rect 31630 4664 31635 4720
rect 28901 4662 31635 4664
rect 28901 4659 28967 4662
rect 31569 4659 31635 4662
rect 31702 4660 31708 4724
rect 31772 4722 31778 4724
rect 33133 4722 33199 4725
rect 36353 4722 36419 4725
rect 31772 4720 36419 4722
rect 31772 4664 33138 4720
rect 33194 4664 36358 4720
rect 36414 4664 36419 4720
rect 31772 4662 36419 4664
rect 31772 4660 31778 4662
rect 33133 4659 33199 4662
rect 36353 4659 36419 4662
rect 38745 4722 38811 4725
rect 42149 4722 42215 4725
rect 46657 4722 46723 4725
rect 38745 4720 46723 4722
rect 38745 4664 38750 4720
rect 38806 4664 42154 4720
rect 42210 4664 46662 4720
rect 46718 4664 46723 4720
rect 38745 4662 46723 4664
rect 38745 4659 38811 4662
rect 42149 4659 42215 4662
rect 46657 4659 46723 4662
rect 49601 4722 49667 4725
rect 51533 4722 51599 4725
rect 49601 4720 51599 4722
rect 49601 4664 49606 4720
rect 49662 4664 51538 4720
rect 51594 4664 51599 4720
rect 49601 4662 51599 4664
rect 49601 4659 49667 4662
rect 51533 4659 51599 4662
rect 15469 4586 15535 4589
rect 27429 4586 27495 4589
rect 30005 4586 30071 4589
rect 34605 4586 34671 4589
rect 54293 4586 54359 4589
rect 55029 4586 55095 4589
rect 15469 4584 27538 4586
rect 15469 4528 15474 4584
rect 15530 4528 27434 4584
rect 27490 4528 27538 4584
rect 15469 4526 27538 4528
rect 15469 4523 15535 4526
rect 27429 4523 27538 4526
rect 30005 4584 34671 4586
rect 30005 4528 30010 4584
rect 30066 4528 34610 4584
rect 34666 4528 34671 4584
rect 30005 4526 34671 4528
rect 30005 4523 30071 4526
rect 34605 4523 34671 4526
rect 51904 4584 55095 4586
rect 51904 4528 54298 4584
rect 54354 4528 55034 4584
rect 55090 4528 55095 4584
rect 51904 4526 55095 4528
rect 19425 4450 19491 4453
rect 23749 4450 23815 4453
rect 19425 4448 23815 4450
rect 19425 4392 19430 4448
rect 19486 4392 23754 4448
rect 23810 4392 23815 4448
rect 19425 4390 23815 4392
rect 27478 4450 27538 4523
rect 51904 4453 51964 4526
rect 54293 4523 54359 4526
rect 55029 4523 55095 4526
rect 32581 4450 32647 4453
rect 36629 4450 36695 4453
rect 27478 4390 31954 4450
rect 19425 4387 19491 4390
rect 23749 4387 23815 4390
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 12249 4314 12315 4317
rect 31702 4314 31708 4316
rect 12249 4312 31708 4314
rect 12249 4256 12254 4312
rect 12310 4256 31708 4312
rect 12249 4254 31708 4256
rect 12249 4251 12315 4254
rect 31702 4252 31708 4254
rect 31772 4252 31778 4316
rect 11145 4178 11211 4181
rect 12433 4178 12499 4181
rect 11145 4176 12499 4178
rect 11145 4120 11150 4176
rect 11206 4120 12438 4176
rect 12494 4120 12499 4176
rect 11145 4118 12499 4120
rect 11145 4115 11211 4118
rect 12433 4115 12499 4118
rect 13537 4178 13603 4181
rect 18781 4178 18847 4181
rect 13537 4176 18847 4178
rect 13537 4120 13542 4176
rect 13598 4120 18786 4176
rect 18842 4120 18847 4176
rect 13537 4118 18847 4120
rect 13537 4115 13603 4118
rect 18781 4115 18847 4118
rect 18965 4178 19031 4181
rect 21081 4178 21147 4181
rect 18965 4176 21147 4178
rect 18965 4120 18970 4176
rect 19026 4120 21086 4176
rect 21142 4120 21147 4176
rect 18965 4118 21147 4120
rect 18965 4115 19031 4118
rect 21081 4115 21147 4118
rect 22001 4178 22067 4181
rect 25865 4178 25931 4181
rect 22001 4176 25931 4178
rect 22001 4120 22006 4176
rect 22062 4120 25870 4176
rect 25926 4120 25931 4176
rect 22001 4118 25931 4120
rect 31894 4178 31954 4390
rect 32581 4448 36695 4450
rect 32581 4392 32586 4448
rect 32642 4392 36634 4448
rect 36690 4392 36695 4448
rect 32581 4390 36695 4392
rect 32581 4387 32647 4390
rect 36629 4387 36695 4390
rect 48497 4450 48563 4453
rect 51901 4450 51967 4453
rect 48497 4448 51967 4450
rect 48497 4392 48502 4448
rect 48558 4392 51906 4448
rect 51962 4392 51967 4448
rect 48497 4390 51967 4392
rect 48497 4387 48563 4390
rect 51901 4387 51967 4390
rect 32132 4384 32452 4385
rect 32132 4320 32140 4384
rect 32204 4320 32220 4384
rect 32284 4320 32300 4384
rect 32364 4320 32380 4384
rect 32444 4320 32452 4384
rect 32132 4319 32452 4320
rect 52924 4384 53244 4385
rect 52924 4320 52932 4384
rect 52996 4320 53012 4384
rect 53076 4320 53092 4384
rect 53156 4320 53172 4384
rect 53236 4320 53244 4384
rect 52924 4319 53244 4320
rect 33777 4314 33843 4317
rect 36813 4314 36879 4317
rect 33777 4312 36879 4314
rect 33777 4256 33782 4312
rect 33838 4256 36818 4312
rect 36874 4256 36879 4312
rect 33777 4254 36879 4256
rect 33777 4251 33843 4254
rect 36813 4251 36879 4254
rect 32029 4178 32095 4181
rect 35617 4178 35683 4181
rect 45645 4178 45711 4181
rect 47945 4178 48011 4181
rect 31894 4176 35683 4178
rect 31894 4120 32034 4176
rect 32090 4120 35622 4176
rect 35678 4120 35683 4176
rect 31894 4118 35683 4120
rect 22001 4115 22067 4118
rect 25865 4115 25931 4118
rect 32029 4115 32095 4118
rect 35617 4115 35683 4118
rect 41094 4118 43178 4178
rect 4061 4042 4127 4045
rect 41094 4042 41154 4118
rect 43118 4042 43178 4118
rect 45645 4176 48011 4178
rect 45645 4120 45650 4176
rect 45706 4120 47950 4176
rect 48006 4120 48011 4176
rect 45645 4118 48011 4120
rect 45645 4115 45711 4118
rect 47945 4115 48011 4118
rect 52177 4178 52243 4181
rect 54661 4178 54727 4181
rect 52177 4176 54727 4178
rect 52177 4120 52182 4176
rect 52238 4120 54666 4176
rect 54722 4120 54727 4176
rect 52177 4118 54727 4120
rect 52177 4115 52243 4118
rect 54661 4115 54727 4118
rect 49877 4042 49943 4045
rect 4061 4040 41154 4042
rect 4061 3984 4066 4040
rect 4122 3984 41154 4040
rect 4061 3982 41154 3984
rect 42382 3982 42994 4042
rect 43118 4040 49943 4042
rect 43118 3984 49882 4040
rect 49938 3984 49943 4040
rect 43118 3982 49943 3984
rect 4061 3979 4127 3982
rect 14825 3906 14891 3909
rect 2822 3904 14891 3906
rect 2822 3848 14830 3904
rect 14886 3848 14891 3904
rect 2822 3846 14891 3848
rect 2822 3498 2882 3846
rect 14825 3843 14891 3846
rect 16481 3906 16547 3909
rect 20529 3906 20595 3909
rect 20805 3906 20871 3909
rect 16481 3904 20871 3906
rect 16481 3848 16486 3904
rect 16542 3848 20534 3904
rect 20590 3848 20810 3904
rect 20866 3848 20871 3904
rect 16481 3846 20871 3848
rect 16481 3843 16547 3846
rect 20529 3843 20595 3846
rect 20805 3843 20871 3846
rect 22185 3906 22251 3909
rect 22921 3906 22987 3909
rect 23381 3906 23447 3909
rect 22185 3904 23447 3906
rect 22185 3848 22190 3904
rect 22246 3848 22926 3904
rect 22982 3848 23386 3904
rect 23442 3848 23447 3904
rect 22185 3846 23447 3848
rect 22185 3843 22251 3846
rect 22921 3843 22987 3846
rect 23381 3843 23447 3846
rect 23565 3906 23631 3909
rect 28441 3906 28507 3909
rect 23565 3904 28507 3906
rect 23565 3848 23570 3904
rect 23626 3848 28446 3904
rect 28502 3848 28507 3904
rect 23565 3846 28507 3848
rect 23565 3843 23631 3846
rect 28441 3843 28507 3846
rect 32213 3906 32279 3909
rect 32857 3906 32923 3909
rect 32213 3904 32923 3906
rect 32213 3848 32218 3904
rect 32274 3848 32862 3904
rect 32918 3848 32923 3904
rect 32213 3846 32923 3848
rect 32213 3843 32279 3846
rect 32857 3843 32923 3846
rect 33133 3906 33199 3909
rect 42382 3906 42442 3982
rect 33133 3904 42442 3906
rect 33133 3848 33138 3904
rect 33194 3848 42442 3904
rect 33133 3846 42442 3848
rect 42934 3906 42994 3982
rect 49877 3979 49943 3982
rect 50889 4042 50955 4045
rect 52545 4042 52611 4045
rect 50889 4040 52611 4042
rect 50889 3984 50894 4040
rect 50950 3984 52550 4040
rect 52606 3984 52611 4040
rect 50889 3982 52611 3984
rect 50889 3979 50955 3982
rect 52545 3979 52611 3982
rect 52729 4042 52795 4045
rect 55213 4042 55279 4045
rect 52729 4040 55279 4042
rect 52729 3984 52734 4040
rect 52790 3984 55218 4040
rect 55274 3984 55279 4040
rect 52729 3982 55279 3984
rect 52729 3979 52795 3982
rect 55213 3979 55279 3982
rect 54109 3906 54175 3909
rect 42934 3904 54175 3906
rect 42934 3848 54114 3904
rect 54170 3848 54175 3904
rect 42934 3846 54175 3848
rect 33133 3843 33199 3846
rect 54109 3843 54175 3846
rect 21736 3840 22056 3841
rect 21736 3776 21744 3840
rect 21808 3776 21824 3840
rect 21888 3776 21904 3840
rect 21968 3776 21984 3840
rect 22048 3776 22056 3840
rect 21736 3775 22056 3776
rect 42528 3840 42848 3841
rect 42528 3776 42536 3840
rect 42600 3776 42616 3840
rect 42680 3776 42696 3840
rect 42760 3776 42776 3840
rect 42840 3776 42848 3840
rect 42528 3775 42848 3776
rect 3417 3770 3483 3773
rect 13353 3770 13419 3773
rect 3417 3768 13419 3770
rect 3417 3712 3422 3768
rect 3478 3712 13358 3768
rect 13414 3712 13419 3768
rect 3417 3710 13419 3712
rect 3417 3707 3483 3710
rect 13353 3707 13419 3710
rect 26877 3770 26943 3773
rect 42241 3770 42307 3773
rect 26877 3768 42307 3770
rect 26877 3712 26882 3768
rect 26938 3712 42246 3768
rect 42302 3712 42307 3768
rect 26877 3710 42307 3712
rect 26877 3707 26943 3710
rect 42241 3707 42307 3710
rect 50429 3770 50495 3773
rect 51717 3770 51783 3773
rect 50429 3768 51783 3770
rect 50429 3712 50434 3768
rect 50490 3712 51722 3768
rect 51778 3712 51783 3768
rect 50429 3710 51783 3712
rect 50429 3707 50495 3710
rect 51717 3707 51783 3710
rect 4797 3634 4863 3637
rect 25313 3634 25379 3637
rect 30833 3634 30899 3637
rect 4797 3632 25379 3634
rect 4797 3576 4802 3632
rect 4858 3576 25318 3632
rect 25374 3576 25379 3632
rect 4797 3574 25379 3576
rect 4797 3571 4863 3574
rect 25313 3571 25379 3574
rect 27846 3632 30899 3634
rect 27846 3576 30838 3632
rect 30894 3576 30899 3632
rect 27846 3574 30899 3576
rect 2638 3438 2882 3498
rect 11605 3498 11671 3501
rect 23381 3498 23447 3501
rect 11605 3496 23447 3498
rect 11605 3440 11610 3496
rect 11666 3440 23386 3496
rect 23442 3440 23447 3496
rect 11605 3438 23447 3440
rect 0 3362 800 3392
rect 2638 3362 2698 3438
rect 11605 3435 11671 3438
rect 23381 3435 23447 3438
rect 24669 3498 24735 3501
rect 27846 3498 27906 3574
rect 30833 3571 30899 3574
rect 31385 3634 31451 3637
rect 47025 3634 47091 3637
rect 31385 3632 47091 3634
rect 31385 3576 31390 3632
rect 31446 3576 47030 3632
rect 47086 3576 47091 3632
rect 31385 3574 47091 3576
rect 31385 3571 31451 3574
rect 47025 3571 47091 3574
rect 24669 3496 27906 3498
rect 24669 3440 24674 3496
rect 24730 3440 27906 3496
rect 24669 3438 27906 3440
rect 27981 3498 28047 3501
rect 31845 3498 31911 3501
rect 27981 3496 31911 3498
rect 27981 3440 27986 3496
rect 28042 3440 31850 3496
rect 31906 3440 31911 3496
rect 27981 3438 31911 3440
rect 24669 3435 24735 3438
rect 27981 3435 28047 3438
rect 31845 3435 31911 3438
rect 32029 3498 32095 3501
rect 34881 3498 34947 3501
rect 43897 3498 43963 3501
rect 32029 3496 32644 3498
rect 32029 3440 32034 3496
rect 32090 3440 32644 3496
rect 32029 3438 32644 3440
rect 32029 3435 32095 3438
rect 0 3302 2698 3362
rect 13813 3362 13879 3365
rect 17769 3362 17835 3365
rect 25681 3362 25747 3365
rect 13813 3360 25747 3362
rect 13813 3304 13818 3360
rect 13874 3304 17774 3360
rect 17830 3304 25686 3360
rect 25742 3304 25747 3360
rect 13813 3302 25747 3304
rect 0 3272 800 3302
rect 13813 3299 13879 3302
rect 17769 3299 17835 3302
rect 25681 3299 25747 3302
rect 26141 3362 26207 3365
rect 26785 3362 26851 3365
rect 29269 3362 29335 3365
rect 31293 3362 31359 3365
rect 26141 3360 26851 3362
rect 26141 3304 26146 3360
rect 26202 3304 26790 3360
rect 26846 3304 26851 3360
rect 26141 3302 26851 3304
rect 26141 3299 26207 3302
rect 26785 3299 26851 3302
rect 28582 3360 31359 3362
rect 28582 3304 29274 3360
rect 29330 3304 31298 3360
rect 31354 3304 31359 3360
rect 28582 3302 31359 3304
rect 32584 3362 32644 3438
rect 34881 3496 43963 3498
rect 34881 3440 34886 3496
rect 34942 3440 43902 3496
rect 43958 3440 43963 3496
rect 34881 3438 43963 3440
rect 34881 3435 34947 3438
rect 43897 3435 43963 3438
rect 44173 3498 44239 3501
rect 46105 3498 46171 3501
rect 44173 3496 46171 3498
rect 44173 3440 44178 3496
rect 44234 3440 46110 3496
rect 46166 3440 46171 3496
rect 44173 3438 46171 3440
rect 44173 3435 44239 3438
rect 46105 3435 46171 3438
rect 48865 3498 48931 3501
rect 56317 3498 56383 3501
rect 48865 3496 56383 3498
rect 48865 3440 48870 3496
rect 48926 3440 56322 3496
rect 56378 3440 56383 3496
rect 48865 3438 56383 3440
rect 48865 3435 48931 3438
rect 56317 3435 56383 3438
rect 38009 3362 38075 3365
rect 32584 3360 38075 3362
rect 32584 3304 38014 3360
rect 38070 3304 38075 3360
rect 32584 3302 38075 3304
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 12893 3226 12959 3229
rect 18965 3226 19031 3229
rect 12893 3224 19031 3226
rect 12893 3168 12898 3224
rect 12954 3168 18970 3224
rect 19026 3168 19031 3224
rect 12893 3166 19031 3168
rect 12893 3163 12959 3166
rect 18965 3163 19031 3166
rect 19241 3226 19307 3229
rect 22829 3226 22895 3229
rect 28582 3226 28642 3302
rect 29269 3299 29335 3302
rect 31293 3299 31359 3302
rect 38009 3299 38075 3302
rect 38745 3362 38811 3365
rect 47669 3362 47735 3365
rect 38745 3360 47735 3362
rect 38745 3304 38750 3360
rect 38806 3304 47674 3360
rect 47730 3304 47735 3360
rect 38745 3302 47735 3304
rect 38745 3299 38811 3302
rect 47669 3299 47735 3302
rect 32132 3296 32452 3297
rect 32132 3232 32140 3296
rect 32204 3232 32220 3296
rect 32284 3232 32300 3296
rect 32364 3232 32380 3296
rect 32444 3232 32452 3296
rect 32132 3231 32452 3232
rect 52924 3296 53244 3297
rect 52924 3232 52932 3296
rect 52996 3232 53012 3296
rect 53076 3232 53092 3296
rect 53156 3232 53172 3296
rect 53236 3232 53244 3296
rect 52924 3231 53244 3232
rect 19241 3224 28642 3226
rect 19241 3168 19246 3224
rect 19302 3168 22834 3224
rect 22890 3168 28642 3224
rect 19241 3166 28642 3168
rect 28809 3226 28875 3229
rect 31477 3226 31543 3229
rect 28809 3224 31543 3226
rect 28809 3168 28814 3224
rect 28870 3168 31482 3224
rect 31538 3168 31543 3224
rect 28809 3166 31543 3168
rect 19241 3163 19307 3166
rect 22829 3163 22895 3166
rect 28809 3163 28875 3166
rect 31477 3163 31543 3166
rect 32765 3226 32831 3229
rect 39297 3226 39363 3229
rect 32765 3224 39363 3226
rect 32765 3168 32770 3224
rect 32826 3168 39302 3224
rect 39358 3168 39363 3224
rect 32765 3166 39363 3168
rect 32765 3163 32831 3166
rect 39297 3163 39363 3166
rect 40309 3226 40375 3229
rect 41965 3226 42031 3229
rect 40309 3224 42031 3226
rect 40309 3168 40314 3224
rect 40370 3168 41970 3224
rect 42026 3168 42031 3224
rect 40309 3166 42031 3168
rect 40309 3163 40375 3166
rect 41965 3163 42031 3166
rect 42241 3226 42307 3229
rect 43437 3226 43503 3229
rect 49509 3226 49575 3229
rect 42241 3224 43362 3226
rect 42241 3168 42246 3224
rect 42302 3168 43362 3224
rect 42241 3166 43362 3168
rect 42241 3163 42307 3166
rect 381 3090 447 3093
rect 24669 3090 24735 3093
rect 381 3088 24735 3090
rect 381 3032 386 3088
rect 442 3032 24674 3088
rect 24730 3032 24735 3088
rect 381 3030 24735 3032
rect 381 3027 447 3030
rect 24669 3027 24735 3030
rect 25129 3090 25195 3093
rect 32121 3090 32187 3093
rect 43161 3090 43227 3093
rect 25129 3088 31954 3090
rect 25129 3032 25134 3088
rect 25190 3032 31954 3088
rect 25129 3030 31954 3032
rect 25129 3027 25195 3030
rect 7833 2954 7899 2957
rect 11145 2954 11211 2957
rect 7833 2952 11211 2954
rect 7833 2896 7838 2952
rect 7894 2896 11150 2952
rect 11206 2896 11211 2952
rect 7833 2894 11211 2896
rect 7833 2891 7899 2894
rect 11145 2891 11211 2894
rect 15929 2954 15995 2957
rect 17769 2954 17835 2957
rect 15929 2952 17835 2954
rect 15929 2896 15934 2952
rect 15990 2896 17774 2952
rect 17830 2896 17835 2952
rect 15929 2894 17835 2896
rect 15929 2891 15995 2894
rect 17769 2891 17835 2894
rect 20345 2954 20411 2957
rect 22553 2954 22619 2957
rect 20345 2952 22619 2954
rect 20345 2896 20350 2952
rect 20406 2896 22558 2952
rect 22614 2896 22619 2952
rect 20345 2894 22619 2896
rect 20345 2891 20411 2894
rect 22553 2891 22619 2894
rect 24393 2954 24459 2957
rect 30925 2954 30991 2957
rect 24393 2952 30991 2954
rect 24393 2896 24398 2952
rect 24454 2896 30930 2952
rect 30986 2896 30991 2952
rect 24393 2894 30991 2896
rect 31894 2954 31954 3030
rect 32121 3088 43227 3090
rect 32121 3032 32126 3088
rect 32182 3032 43166 3088
rect 43222 3032 43227 3088
rect 32121 3030 43227 3032
rect 43302 3090 43362 3166
rect 43437 3224 49575 3226
rect 43437 3168 43442 3224
rect 43498 3168 49514 3224
rect 49570 3168 49575 3224
rect 43437 3166 49575 3168
rect 43437 3163 43503 3166
rect 49509 3163 49575 3166
rect 44909 3090 44975 3093
rect 43302 3088 44975 3090
rect 43302 3032 44914 3088
rect 44970 3032 44975 3088
rect 43302 3030 44975 3032
rect 32121 3027 32187 3030
rect 43161 3027 43227 3030
rect 44909 3027 44975 3030
rect 45093 3090 45159 3093
rect 47025 3090 47091 3093
rect 45093 3088 47091 3090
rect 45093 3032 45098 3088
rect 45154 3032 47030 3088
rect 47086 3032 47091 3088
rect 45093 3030 47091 3032
rect 45093 3027 45159 3030
rect 47025 3027 47091 3030
rect 33777 2954 33843 2957
rect 31894 2952 33843 2954
rect 31894 2896 33782 2952
rect 33838 2896 33843 2952
rect 31894 2894 33843 2896
rect 24393 2891 24459 2894
rect 30925 2891 30991 2894
rect 33777 2891 33843 2894
rect 33961 2954 34027 2957
rect 60273 2954 60339 2957
rect 33961 2952 60339 2954
rect 33961 2896 33966 2952
rect 34022 2896 60278 2952
rect 60334 2896 60339 2952
rect 33961 2894 60339 2896
rect 33961 2891 34027 2894
rect 60273 2891 60339 2894
rect 3693 2818 3759 2821
rect 12985 2818 13051 2821
rect 3693 2816 13051 2818
rect 3693 2760 3698 2816
rect 3754 2760 12990 2816
rect 13046 2760 13051 2816
rect 3693 2758 13051 2760
rect 3693 2755 3759 2758
rect 12985 2755 13051 2758
rect 29545 2818 29611 2821
rect 38745 2818 38811 2821
rect 29545 2816 38811 2818
rect 29545 2760 29550 2816
rect 29606 2760 38750 2816
rect 38806 2760 38811 2816
rect 29545 2758 38811 2760
rect 29545 2755 29611 2758
rect 38745 2755 38811 2758
rect 44817 2818 44883 2821
rect 46381 2818 46447 2821
rect 44817 2816 46447 2818
rect 44817 2760 44822 2816
rect 44878 2760 46386 2816
rect 46442 2760 46447 2816
rect 44817 2758 46447 2760
rect 44817 2755 44883 2758
rect 46381 2755 46447 2758
rect 21736 2752 22056 2753
rect 21736 2688 21744 2752
rect 21808 2688 21824 2752
rect 21888 2688 21904 2752
rect 21968 2688 21984 2752
rect 22048 2688 22056 2752
rect 21736 2687 22056 2688
rect 42528 2752 42848 2753
rect 42528 2688 42536 2752
rect 42600 2688 42616 2752
rect 42680 2688 42696 2752
rect 42760 2688 42776 2752
rect 42840 2688 42848 2752
rect 42528 2687 42848 2688
rect 10685 2682 10751 2685
rect 19057 2682 19123 2685
rect 10685 2680 19123 2682
rect 10685 2624 10690 2680
rect 10746 2624 19062 2680
rect 19118 2624 19123 2680
rect 10685 2622 19123 2624
rect 10685 2619 10751 2622
rect 19057 2619 19123 2622
rect 39021 2546 39087 2549
rect 45461 2546 45527 2549
rect 39021 2544 45527 2546
rect 39021 2488 39026 2544
rect 39082 2488 45466 2544
rect 45522 2488 45527 2544
rect 39021 2486 45527 2488
rect 39021 2483 39087 2486
rect 45461 2483 45527 2486
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 32132 2208 32452 2209
rect 32132 2144 32140 2208
rect 32204 2144 32220 2208
rect 32284 2144 32300 2208
rect 32364 2144 32380 2208
rect 32444 2144 32452 2208
rect 32132 2143 32452 2144
rect 52924 2208 53244 2209
rect 52924 2144 52932 2208
rect 52996 2144 53012 2208
rect 53076 2144 53092 2208
rect 53156 2144 53172 2208
rect 53236 2144 53244 2208
rect 52924 2143 53244 2144
rect 0 1186 800 1216
rect 4061 1186 4127 1189
rect 0 1184 4127 1186
rect 0 1128 4066 1184
rect 4122 1128 4127 1184
rect 0 1126 4127 1128
rect 0 1096 800 1126
rect 4061 1123 4127 1126
<< via3 >>
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 32140 17436 32204 17440
rect 32140 17380 32144 17436
rect 32144 17380 32200 17436
rect 32200 17380 32204 17436
rect 32140 17376 32204 17380
rect 32220 17436 32284 17440
rect 32220 17380 32224 17436
rect 32224 17380 32280 17436
rect 32280 17380 32284 17436
rect 32220 17376 32284 17380
rect 32300 17436 32364 17440
rect 32300 17380 32304 17436
rect 32304 17380 32360 17436
rect 32360 17380 32364 17436
rect 32300 17376 32364 17380
rect 32380 17436 32444 17440
rect 32380 17380 32384 17436
rect 32384 17380 32440 17436
rect 32440 17380 32444 17436
rect 32380 17376 32444 17380
rect 52932 17436 52996 17440
rect 52932 17380 52936 17436
rect 52936 17380 52992 17436
rect 52992 17380 52996 17436
rect 52932 17376 52996 17380
rect 53012 17436 53076 17440
rect 53012 17380 53016 17436
rect 53016 17380 53072 17436
rect 53072 17380 53076 17436
rect 53012 17376 53076 17380
rect 53092 17436 53156 17440
rect 53092 17380 53096 17436
rect 53096 17380 53152 17436
rect 53152 17380 53156 17436
rect 53092 17376 53156 17380
rect 53172 17436 53236 17440
rect 53172 17380 53176 17436
rect 53176 17380 53232 17436
rect 53232 17380 53236 17436
rect 53172 17376 53236 17380
rect 21744 16892 21808 16896
rect 21744 16836 21748 16892
rect 21748 16836 21804 16892
rect 21804 16836 21808 16892
rect 21744 16832 21808 16836
rect 21824 16892 21888 16896
rect 21824 16836 21828 16892
rect 21828 16836 21884 16892
rect 21884 16836 21888 16892
rect 21824 16832 21888 16836
rect 21904 16892 21968 16896
rect 21904 16836 21908 16892
rect 21908 16836 21964 16892
rect 21964 16836 21968 16892
rect 21904 16832 21968 16836
rect 21984 16892 22048 16896
rect 21984 16836 21988 16892
rect 21988 16836 22044 16892
rect 22044 16836 22048 16892
rect 21984 16832 22048 16836
rect 42536 16892 42600 16896
rect 42536 16836 42540 16892
rect 42540 16836 42596 16892
rect 42596 16836 42600 16892
rect 42536 16832 42600 16836
rect 42616 16892 42680 16896
rect 42616 16836 42620 16892
rect 42620 16836 42676 16892
rect 42676 16836 42680 16892
rect 42616 16832 42680 16836
rect 42696 16892 42760 16896
rect 42696 16836 42700 16892
rect 42700 16836 42756 16892
rect 42756 16836 42760 16892
rect 42696 16832 42760 16836
rect 42776 16892 42840 16896
rect 42776 16836 42780 16892
rect 42780 16836 42836 16892
rect 42836 16836 42840 16892
rect 42776 16832 42840 16836
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 32140 16348 32204 16352
rect 32140 16292 32144 16348
rect 32144 16292 32200 16348
rect 32200 16292 32204 16348
rect 32140 16288 32204 16292
rect 32220 16348 32284 16352
rect 32220 16292 32224 16348
rect 32224 16292 32280 16348
rect 32280 16292 32284 16348
rect 32220 16288 32284 16292
rect 32300 16348 32364 16352
rect 32300 16292 32304 16348
rect 32304 16292 32360 16348
rect 32360 16292 32364 16348
rect 32300 16288 32364 16292
rect 32380 16348 32444 16352
rect 32380 16292 32384 16348
rect 32384 16292 32440 16348
rect 32440 16292 32444 16348
rect 32380 16288 32444 16292
rect 52932 16348 52996 16352
rect 52932 16292 52936 16348
rect 52936 16292 52992 16348
rect 52992 16292 52996 16348
rect 52932 16288 52996 16292
rect 53012 16348 53076 16352
rect 53012 16292 53016 16348
rect 53016 16292 53072 16348
rect 53072 16292 53076 16348
rect 53012 16288 53076 16292
rect 53092 16348 53156 16352
rect 53092 16292 53096 16348
rect 53096 16292 53152 16348
rect 53152 16292 53156 16348
rect 53092 16288 53156 16292
rect 53172 16348 53236 16352
rect 53172 16292 53176 16348
rect 53176 16292 53232 16348
rect 53232 16292 53236 16348
rect 53172 16288 53236 16292
rect 21744 15804 21808 15808
rect 21744 15748 21748 15804
rect 21748 15748 21804 15804
rect 21804 15748 21808 15804
rect 21744 15744 21808 15748
rect 21824 15804 21888 15808
rect 21824 15748 21828 15804
rect 21828 15748 21884 15804
rect 21884 15748 21888 15804
rect 21824 15744 21888 15748
rect 21904 15804 21968 15808
rect 21904 15748 21908 15804
rect 21908 15748 21964 15804
rect 21964 15748 21968 15804
rect 21904 15744 21968 15748
rect 21984 15804 22048 15808
rect 21984 15748 21988 15804
rect 21988 15748 22044 15804
rect 22044 15748 22048 15804
rect 21984 15744 22048 15748
rect 42536 15804 42600 15808
rect 42536 15748 42540 15804
rect 42540 15748 42596 15804
rect 42596 15748 42600 15804
rect 42536 15744 42600 15748
rect 42616 15804 42680 15808
rect 42616 15748 42620 15804
rect 42620 15748 42676 15804
rect 42676 15748 42680 15804
rect 42616 15744 42680 15748
rect 42696 15804 42760 15808
rect 42696 15748 42700 15804
rect 42700 15748 42756 15804
rect 42756 15748 42760 15804
rect 42696 15744 42760 15748
rect 42776 15804 42840 15808
rect 42776 15748 42780 15804
rect 42780 15748 42836 15804
rect 42836 15748 42840 15804
rect 42776 15744 42840 15748
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 32140 15260 32204 15264
rect 32140 15204 32144 15260
rect 32144 15204 32200 15260
rect 32200 15204 32204 15260
rect 32140 15200 32204 15204
rect 32220 15260 32284 15264
rect 32220 15204 32224 15260
rect 32224 15204 32280 15260
rect 32280 15204 32284 15260
rect 32220 15200 32284 15204
rect 32300 15260 32364 15264
rect 32300 15204 32304 15260
rect 32304 15204 32360 15260
rect 32360 15204 32364 15260
rect 32300 15200 32364 15204
rect 32380 15260 32444 15264
rect 32380 15204 32384 15260
rect 32384 15204 32440 15260
rect 32440 15204 32444 15260
rect 32380 15200 32444 15204
rect 52932 15260 52996 15264
rect 52932 15204 52936 15260
rect 52936 15204 52992 15260
rect 52992 15204 52996 15260
rect 52932 15200 52996 15204
rect 53012 15260 53076 15264
rect 53012 15204 53016 15260
rect 53016 15204 53072 15260
rect 53072 15204 53076 15260
rect 53012 15200 53076 15204
rect 53092 15260 53156 15264
rect 53092 15204 53096 15260
rect 53096 15204 53152 15260
rect 53152 15204 53156 15260
rect 53092 15200 53156 15204
rect 53172 15260 53236 15264
rect 53172 15204 53176 15260
rect 53176 15204 53232 15260
rect 53232 15204 53236 15260
rect 53172 15200 53236 15204
rect 21744 14716 21808 14720
rect 21744 14660 21748 14716
rect 21748 14660 21804 14716
rect 21804 14660 21808 14716
rect 21744 14656 21808 14660
rect 21824 14716 21888 14720
rect 21824 14660 21828 14716
rect 21828 14660 21884 14716
rect 21884 14660 21888 14716
rect 21824 14656 21888 14660
rect 21904 14716 21968 14720
rect 21904 14660 21908 14716
rect 21908 14660 21964 14716
rect 21964 14660 21968 14716
rect 21904 14656 21968 14660
rect 21984 14716 22048 14720
rect 21984 14660 21988 14716
rect 21988 14660 22044 14716
rect 22044 14660 22048 14716
rect 21984 14656 22048 14660
rect 42536 14716 42600 14720
rect 42536 14660 42540 14716
rect 42540 14660 42596 14716
rect 42596 14660 42600 14716
rect 42536 14656 42600 14660
rect 42616 14716 42680 14720
rect 42616 14660 42620 14716
rect 42620 14660 42676 14716
rect 42676 14660 42680 14716
rect 42616 14656 42680 14660
rect 42696 14716 42760 14720
rect 42696 14660 42700 14716
rect 42700 14660 42756 14716
rect 42756 14660 42760 14716
rect 42696 14656 42760 14660
rect 42776 14716 42840 14720
rect 42776 14660 42780 14716
rect 42780 14660 42836 14716
rect 42836 14660 42840 14716
rect 42776 14656 42840 14660
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 32140 14172 32204 14176
rect 32140 14116 32144 14172
rect 32144 14116 32200 14172
rect 32200 14116 32204 14172
rect 32140 14112 32204 14116
rect 32220 14172 32284 14176
rect 32220 14116 32224 14172
rect 32224 14116 32280 14172
rect 32280 14116 32284 14172
rect 32220 14112 32284 14116
rect 32300 14172 32364 14176
rect 32300 14116 32304 14172
rect 32304 14116 32360 14172
rect 32360 14116 32364 14172
rect 32300 14112 32364 14116
rect 32380 14172 32444 14176
rect 32380 14116 32384 14172
rect 32384 14116 32440 14172
rect 32440 14116 32444 14172
rect 32380 14112 32444 14116
rect 52932 14172 52996 14176
rect 52932 14116 52936 14172
rect 52936 14116 52992 14172
rect 52992 14116 52996 14172
rect 52932 14112 52996 14116
rect 53012 14172 53076 14176
rect 53012 14116 53016 14172
rect 53016 14116 53072 14172
rect 53072 14116 53076 14172
rect 53012 14112 53076 14116
rect 53092 14172 53156 14176
rect 53092 14116 53096 14172
rect 53096 14116 53152 14172
rect 53152 14116 53156 14172
rect 53092 14112 53156 14116
rect 53172 14172 53236 14176
rect 53172 14116 53176 14172
rect 53176 14116 53232 14172
rect 53232 14116 53236 14172
rect 53172 14112 53236 14116
rect 21744 13628 21808 13632
rect 21744 13572 21748 13628
rect 21748 13572 21804 13628
rect 21804 13572 21808 13628
rect 21744 13568 21808 13572
rect 21824 13628 21888 13632
rect 21824 13572 21828 13628
rect 21828 13572 21884 13628
rect 21884 13572 21888 13628
rect 21824 13568 21888 13572
rect 21904 13628 21968 13632
rect 21904 13572 21908 13628
rect 21908 13572 21964 13628
rect 21964 13572 21968 13628
rect 21904 13568 21968 13572
rect 21984 13628 22048 13632
rect 21984 13572 21988 13628
rect 21988 13572 22044 13628
rect 22044 13572 22048 13628
rect 21984 13568 22048 13572
rect 42536 13628 42600 13632
rect 42536 13572 42540 13628
rect 42540 13572 42596 13628
rect 42596 13572 42600 13628
rect 42536 13568 42600 13572
rect 42616 13628 42680 13632
rect 42616 13572 42620 13628
rect 42620 13572 42676 13628
rect 42676 13572 42680 13628
rect 42616 13568 42680 13572
rect 42696 13628 42760 13632
rect 42696 13572 42700 13628
rect 42700 13572 42756 13628
rect 42756 13572 42760 13628
rect 42696 13568 42760 13572
rect 42776 13628 42840 13632
rect 42776 13572 42780 13628
rect 42780 13572 42836 13628
rect 42836 13572 42840 13628
rect 42776 13568 42840 13572
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 32140 13084 32204 13088
rect 32140 13028 32144 13084
rect 32144 13028 32200 13084
rect 32200 13028 32204 13084
rect 32140 13024 32204 13028
rect 32220 13084 32284 13088
rect 32220 13028 32224 13084
rect 32224 13028 32280 13084
rect 32280 13028 32284 13084
rect 32220 13024 32284 13028
rect 32300 13084 32364 13088
rect 32300 13028 32304 13084
rect 32304 13028 32360 13084
rect 32360 13028 32364 13084
rect 32300 13024 32364 13028
rect 32380 13084 32444 13088
rect 32380 13028 32384 13084
rect 32384 13028 32440 13084
rect 32440 13028 32444 13084
rect 32380 13024 32444 13028
rect 52932 13084 52996 13088
rect 52932 13028 52936 13084
rect 52936 13028 52992 13084
rect 52992 13028 52996 13084
rect 52932 13024 52996 13028
rect 53012 13084 53076 13088
rect 53012 13028 53016 13084
rect 53016 13028 53072 13084
rect 53072 13028 53076 13084
rect 53012 13024 53076 13028
rect 53092 13084 53156 13088
rect 53092 13028 53096 13084
rect 53096 13028 53152 13084
rect 53152 13028 53156 13084
rect 53092 13024 53156 13028
rect 53172 13084 53236 13088
rect 53172 13028 53176 13084
rect 53176 13028 53232 13084
rect 53232 13028 53236 13084
rect 53172 13024 53236 13028
rect 21744 12540 21808 12544
rect 21744 12484 21748 12540
rect 21748 12484 21804 12540
rect 21804 12484 21808 12540
rect 21744 12480 21808 12484
rect 21824 12540 21888 12544
rect 21824 12484 21828 12540
rect 21828 12484 21884 12540
rect 21884 12484 21888 12540
rect 21824 12480 21888 12484
rect 21904 12540 21968 12544
rect 21904 12484 21908 12540
rect 21908 12484 21964 12540
rect 21964 12484 21968 12540
rect 21904 12480 21968 12484
rect 21984 12540 22048 12544
rect 21984 12484 21988 12540
rect 21988 12484 22044 12540
rect 22044 12484 22048 12540
rect 21984 12480 22048 12484
rect 42536 12540 42600 12544
rect 42536 12484 42540 12540
rect 42540 12484 42596 12540
rect 42596 12484 42600 12540
rect 42536 12480 42600 12484
rect 42616 12540 42680 12544
rect 42616 12484 42620 12540
rect 42620 12484 42676 12540
rect 42676 12484 42680 12540
rect 42616 12480 42680 12484
rect 42696 12540 42760 12544
rect 42696 12484 42700 12540
rect 42700 12484 42756 12540
rect 42756 12484 42760 12540
rect 42696 12480 42760 12484
rect 42776 12540 42840 12544
rect 42776 12484 42780 12540
rect 42780 12484 42836 12540
rect 42836 12484 42840 12540
rect 42776 12480 42840 12484
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 32140 11996 32204 12000
rect 32140 11940 32144 11996
rect 32144 11940 32200 11996
rect 32200 11940 32204 11996
rect 32140 11936 32204 11940
rect 32220 11996 32284 12000
rect 32220 11940 32224 11996
rect 32224 11940 32280 11996
rect 32280 11940 32284 11996
rect 32220 11936 32284 11940
rect 32300 11996 32364 12000
rect 32300 11940 32304 11996
rect 32304 11940 32360 11996
rect 32360 11940 32364 11996
rect 32300 11936 32364 11940
rect 32380 11996 32444 12000
rect 32380 11940 32384 11996
rect 32384 11940 32440 11996
rect 32440 11940 32444 11996
rect 32380 11936 32444 11940
rect 52932 11996 52996 12000
rect 52932 11940 52936 11996
rect 52936 11940 52992 11996
rect 52992 11940 52996 11996
rect 52932 11936 52996 11940
rect 53012 11996 53076 12000
rect 53012 11940 53016 11996
rect 53016 11940 53072 11996
rect 53072 11940 53076 11996
rect 53012 11936 53076 11940
rect 53092 11996 53156 12000
rect 53092 11940 53096 11996
rect 53096 11940 53152 11996
rect 53152 11940 53156 11996
rect 53092 11936 53156 11940
rect 53172 11996 53236 12000
rect 53172 11940 53176 11996
rect 53176 11940 53232 11996
rect 53232 11940 53236 11996
rect 53172 11936 53236 11940
rect 21744 11452 21808 11456
rect 21744 11396 21748 11452
rect 21748 11396 21804 11452
rect 21804 11396 21808 11452
rect 21744 11392 21808 11396
rect 21824 11452 21888 11456
rect 21824 11396 21828 11452
rect 21828 11396 21884 11452
rect 21884 11396 21888 11452
rect 21824 11392 21888 11396
rect 21904 11452 21968 11456
rect 21904 11396 21908 11452
rect 21908 11396 21964 11452
rect 21964 11396 21968 11452
rect 21904 11392 21968 11396
rect 21984 11452 22048 11456
rect 21984 11396 21988 11452
rect 21988 11396 22044 11452
rect 22044 11396 22048 11452
rect 21984 11392 22048 11396
rect 42536 11452 42600 11456
rect 42536 11396 42540 11452
rect 42540 11396 42596 11452
rect 42596 11396 42600 11452
rect 42536 11392 42600 11396
rect 42616 11452 42680 11456
rect 42616 11396 42620 11452
rect 42620 11396 42676 11452
rect 42676 11396 42680 11452
rect 42616 11392 42680 11396
rect 42696 11452 42760 11456
rect 42696 11396 42700 11452
rect 42700 11396 42756 11452
rect 42756 11396 42760 11452
rect 42696 11392 42760 11396
rect 42776 11452 42840 11456
rect 42776 11396 42780 11452
rect 42780 11396 42836 11452
rect 42836 11396 42840 11452
rect 42776 11392 42840 11396
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 32140 10908 32204 10912
rect 32140 10852 32144 10908
rect 32144 10852 32200 10908
rect 32200 10852 32204 10908
rect 32140 10848 32204 10852
rect 32220 10908 32284 10912
rect 32220 10852 32224 10908
rect 32224 10852 32280 10908
rect 32280 10852 32284 10908
rect 32220 10848 32284 10852
rect 32300 10908 32364 10912
rect 32300 10852 32304 10908
rect 32304 10852 32360 10908
rect 32360 10852 32364 10908
rect 32300 10848 32364 10852
rect 32380 10908 32444 10912
rect 32380 10852 32384 10908
rect 32384 10852 32440 10908
rect 32440 10852 32444 10908
rect 32380 10848 32444 10852
rect 52932 10908 52996 10912
rect 52932 10852 52936 10908
rect 52936 10852 52992 10908
rect 52992 10852 52996 10908
rect 52932 10848 52996 10852
rect 53012 10908 53076 10912
rect 53012 10852 53016 10908
rect 53016 10852 53072 10908
rect 53072 10852 53076 10908
rect 53012 10848 53076 10852
rect 53092 10908 53156 10912
rect 53092 10852 53096 10908
rect 53096 10852 53152 10908
rect 53152 10852 53156 10908
rect 53092 10848 53156 10852
rect 53172 10908 53236 10912
rect 53172 10852 53176 10908
rect 53176 10852 53232 10908
rect 53232 10852 53236 10908
rect 53172 10848 53236 10852
rect 21744 10364 21808 10368
rect 21744 10308 21748 10364
rect 21748 10308 21804 10364
rect 21804 10308 21808 10364
rect 21744 10304 21808 10308
rect 21824 10364 21888 10368
rect 21824 10308 21828 10364
rect 21828 10308 21884 10364
rect 21884 10308 21888 10364
rect 21824 10304 21888 10308
rect 21904 10364 21968 10368
rect 21904 10308 21908 10364
rect 21908 10308 21964 10364
rect 21964 10308 21968 10364
rect 21904 10304 21968 10308
rect 21984 10364 22048 10368
rect 21984 10308 21988 10364
rect 21988 10308 22044 10364
rect 22044 10308 22048 10364
rect 21984 10304 22048 10308
rect 42536 10364 42600 10368
rect 42536 10308 42540 10364
rect 42540 10308 42596 10364
rect 42596 10308 42600 10364
rect 42536 10304 42600 10308
rect 42616 10364 42680 10368
rect 42616 10308 42620 10364
rect 42620 10308 42676 10364
rect 42676 10308 42680 10364
rect 42616 10304 42680 10308
rect 42696 10364 42760 10368
rect 42696 10308 42700 10364
rect 42700 10308 42756 10364
rect 42756 10308 42760 10364
rect 42696 10304 42760 10308
rect 42776 10364 42840 10368
rect 42776 10308 42780 10364
rect 42780 10308 42836 10364
rect 42836 10308 42840 10364
rect 42776 10304 42840 10308
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 32140 9820 32204 9824
rect 32140 9764 32144 9820
rect 32144 9764 32200 9820
rect 32200 9764 32204 9820
rect 32140 9760 32204 9764
rect 32220 9820 32284 9824
rect 32220 9764 32224 9820
rect 32224 9764 32280 9820
rect 32280 9764 32284 9820
rect 32220 9760 32284 9764
rect 32300 9820 32364 9824
rect 32300 9764 32304 9820
rect 32304 9764 32360 9820
rect 32360 9764 32364 9820
rect 32300 9760 32364 9764
rect 32380 9820 32444 9824
rect 32380 9764 32384 9820
rect 32384 9764 32440 9820
rect 32440 9764 32444 9820
rect 32380 9760 32444 9764
rect 52932 9820 52996 9824
rect 52932 9764 52936 9820
rect 52936 9764 52992 9820
rect 52992 9764 52996 9820
rect 52932 9760 52996 9764
rect 53012 9820 53076 9824
rect 53012 9764 53016 9820
rect 53016 9764 53072 9820
rect 53072 9764 53076 9820
rect 53012 9760 53076 9764
rect 53092 9820 53156 9824
rect 53092 9764 53096 9820
rect 53096 9764 53152 9820
rect 53152 9764 53156 9820
rect 53092 9760 53156 9764
rect 53172 9820 53236 9824
rect 53172 9764 53176 9820
rect 53176 9764 53232 9820
rect 53232 9764 53236 9820
rect 53172 9760 53236 9764
rect 21744 9276 21808 9280
rect 21744 9220 21748 9276
rect 21748 9220 21804 9276
rect 21804 9220 21808 9276
rect 21744 9216 21808 9220
rect 21824 9276 21888 9280
rect 21824 9220 21828 9276
rect 21828 9220 21884 9276
rect 21884 9220 21888 9276
rect 21824 9216 21888 9220
rect 21904 9276 21968 9280
rect 21904 9220 21908 9276
rect 21908 9220 21964 9276
rect 21964 9220 21968 9276
rect 21904 9216 21968 9220
rect 21984 9276 22048 9280
rect 21984 9220 21988 9276
rect 21988 9220 22044 9276
rect 22044 9220 22048 9276
rect 21984 9216 22048 9220
rect 42536 9276 42600 9280
rect 42536 9220 42540 9276
rect 42540 9220 42596 9276
rect 42596 9220 42600 9276
rect 42536 9216 42600 9220
rect 42616 9276 42680 9280
rect 42616 9220 42620 9276
rect 42620 9220 42676 9276
rect 42676 9220 42680 9276
rect 42616 9216 42680 9220
rect 42696 9276 42760 9280
rect 42696 9220 42700 9276
rect 42700 9220 42756 9276
rect 42756 9220 42760 9276
rect 42696 9216 42760 9220
rect 42776 9276 42840 9280
rect 42776 9220 42780 9276
rect 42780 9220 42836 9276
rect 42836 9220 42840 9276
rect 42776 9216 42840 9220
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 32140 8732 32204 8736
rect 32140 8676 32144 8732
rect 32144 8676 32200 8732
rect 32200 8676 32204 8732
rect 32140 8672 32204 8676
rect 32220 8732 32284 8736
rect 32220 8676 32224 8732
rect 32224 8676 32280 8732
rect 32280 8676 32284 8732
rect 32220 8672 32284 8676
rect 32300 8732 32364 8736
rect 32300 8676 32304 8732
rect 32304 8676 32360 8732
rect 32360 8676 32364 8732
rect 32300 8672 32364 8676
rect 32380 8732 32444 8736
rect 32380 8676 32384 8732
rect 32384 8676 32440 8732
rect 32440 8676 32444 8732
rect 32380 8672 32444 8676
rect 52932 8732 52996 8736
rect 52932 8676 52936 8732
rect 52936 8676 52992 8732
rect 52992 8676 52996 8732
rect 52932 8672 52996 8676
rect 53012 8732 53076 8736
rect 53012 8676 53016 8732
rect 53016 8676 53072 8732
rect 53072 8676 53076 8732
rect 53012 8672 53076 8676
rect 53092 8732 53156 8736
rect 53092 8676 53096 8732
rect 53096 8676 53152 8732
rect 53152 8676 53156 8732
rect 53092 8672 53156 8676
rect 53172 8732 53236 8736
rect 53172 8676 53176 8732
rect 53176 8676 53232 8732
rect 53232 8676 53236 8732
rect 53172 8672 53236 8676
rect 28948 8196 29012 8260
rect 21744 8188 21808 8192
rect 21744 8132 21748 8188
rect 21748 8132 21804 8188
rect 21804 8132 21808 8188
rect 21744 8128 21808 8132
rect 21824 8188 21888 8192
rect 21824 8132 21828 8188
rect 21828 8132 21884 8188
rect 21884 8132 21888 8188
rect 21824 8128 21888 8132
rect 21904 8188 21968 8192
rect 21904 8132 21908 8188
rect 21908 8132 21964 8188
rect 21964 8132 21968 8188
rect 21904 8128 21968 8132
rect 21984 8188 22048 8192
rect 21984 8132 21988 8188
rect 21988 8132 22044 8188
rect 22044 8132 22048 8188
rect 21984 8128 22048 8132
rect 42536 8188 42600 8192
rect 42536 8132 42540 8188
rect 42540 8132 42596 8188
rect 42596 8132 42600 8188
rect 42536 8128 42600 8132
rect 42616 8188 42680 8192
rect 42616 8132 42620 8188
rect 42620 8132 42676 8188
rect 42676 8132 42680 8188
rect 42616 8128 42680 8132
rect 42696 8188 42760 8192
rect 42696 8132 42700 8188
rect 42700 8132 42756 8188
rect 42756 8132 42760 8188
rect 42696 8128 42760 8132
rect 42776 8188 42840 8192
rect 42776 8132 42780 8188
rect 42780 8132 42836 8188
rect 42836 8132 42840 8188
rect 42776 8128 42840 8132
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 32140 7644 32204 7648
rect 32140 7588 32144 7644
rect 32144 7588 32200 7644
rect 32200 7588 32204 7644
rect 32140 7584 32204 7588
rect 32220 7644 32284 7648
rect 32220 7588 32224 7644
rect 32224 7588 32280 7644
rect 32280 7588 32284 7644
rect 32220 7584 32284 7588
rect 32300 7644 32364 7648
rect 32300 7588 32304 7644
rect 32304 7588 32360 7644
rect 32360 7588 32364 7644
rect 32300 7584 32364 7588
rect 32380 7644 32444 7648
rect 32380 7588 32384 7644
rect 32384 7588 32440 7644
rect 32440 7588 32444 7644
rect 32380 7584 32444 7588
rect 52932 7644 52996 7648
rect 52932 7588 52936 7644
rect 52936 7588 52992 7644
rect 52992 7588 52996 7644
rect 52932 7584 52996 7588
rect 53012 7644 53076 7648
rect 53012 7588 53016 7644
rect 53016 7588 53072 7644
rect 53072 7588 53076 7644
rect 53012 7584 53076 7588
rect 53092 7644 53156 7648
rect 53092 7588 53096 7644
rect 53096 7588 53152 7644
rect 53152 7588 53156 7644
rect 53092 7584 53156 7588
rect 53172 7644 53236 7648
rect 53172 7588 53176 7644
rect 53176 7588 53232 7644
rect 53232 7588 53236 7644
rect 53172 7584 53236 7588
rect 21744 7100 21808 7104
rect 21744 7044 21748 7100
rect 21748 7044 21804 7100
rect 21804 7044 21808 7100
rect 21744 7040 21808 7044
rect 21824 7100 21888 7104
rect 21824 7044 21828 7100
rect 21828 7044 21884 7100
rect 21884 7044 21888 7100
rect 21824 7040 21888 7044
rect 21904 7100 21968 7104
rect 21904 7044 21908 7100
rect 21908 7044 21964 7100
rect 21964 7044 21968 7100
rect 21904 7040 21968 7044
rect 21984 7100 22048 7104
rect 21984 7044 21988 7100
rect 21988 7044 22044 7100
rect 22044 7044 22048 7100
rect 21984 7040 22048 7044
rect 42536 7100 42600 7104
rect 42536 7044 42540 7100
rect 42540 7044 42596 7100
rect 42596 7044 42600 7100
rect 42536 7040 42600 7044
rect 42616 7100 42680 7104
rect 42616 7044 42620 7100
rect 42620 7044 42676 7100
rect 42676 7044 42680 7100
rect 42616 7040 42680 7044
rect 42696 7100 42760 7104
rect 42696 7044 42700 7100
rect 42700 7044 42756 7100
rect 42756 7044 42760 7100
rect 42696 7040 42760 7044
rect 42776 7100 42840 7104
rect 42776 7044 42780 7100
rect 42780 7044 42836 7100
rect 42836 7044 42840 7100
rect 42776 7040 42840 7044
rect 46796 6564 46860 6628
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 32140 6556 32204 6560
rect 32140 6500 32144 6556
rect 32144 6500 32200 6556
rect 32200 6500 32204 6556
rect 32140 6496 32204 6500
rect 32220 6556 32284 6560
rect 32220 6500 32224 6556
rect 32224 6500 32280 6556
rect 32280 6500 32284 6556
rect 32220 6496 32284 6500
rect 32300 6556 32364 6560
rect 32300 6500 32304 6556
rect 32304 6500 32360 6556
rect 32360 6500 32364 6556
rect 32300 6496 32364 6500
rect 32380 6556 32444 6560
rect 32380 6500 32384 6556
rect 32384 6500 32440 6556
rect 32440 6500 32444 6556
rect 32380 6496 32444 6500
rect 52932 6556 52996 6560
rect 52932 6500 52936 6556
rect 52936 6500 52992 6556
rect 52992 6500 52996 6556
rect 52932 6496 52996 6500
rect 53012 6556 53076 6560
rect 53012 6500 53016 6556
rect 53016 6500 53072 6556
rect 53072 6500 53076 6556
rect 53012 6496 53076 6500
rect 53092 6556 53156 6560
rect 53092 6500 53096 6556
rect 53096 6500 53152 6556
rect 53152 6500 53156 6556
rect 53092 6496 53156 6500
rect 53172 6556 53236 6560
rect 53172 6500 53176 6556
rect 53176 6500 53232 6556
rect 53232 6500 53236 6556
rect 53172 6496 53236 6500
rect 21744 6012 21808 6016
rect 21744 5956 21748 6012
rect 21748 5956 21804 6012
rect 21804 5956 21808 6012
rect 21744 5952 21808 5956
rect 21824 6012 21888 6016
rect 21824 5956 21828 6012
rect 21828 5956 21884 6012
rect 21884 5956 21888 6012
rect 21824 5952 21888 5956
rect 21904 6012 21968 6016
rect 21904 5956 21908 6012
rect 21908 5956 21964 6012
rect 21964 5956 21968 6012
rect 21904 5952 21968 5956
rect 21984 6012 22048 6016
rect 21984 5956 21988 6012
rect 21988 5956 22044 6012
rect 22044 5956 22048 6012
rect 21984 5952 22048 5956
rect 42536 6012 42600 6016
rect 42536 5956 42540 6012
rect 42540 5956 42596 6012
rect 42596 5956 42600 6012
rect 42536 5952 42600 5956
rect 42616 6012 42680 6016
rect 42616 5956 42620 6012
rect 42620 5956 42676 6012
rect 42676 5956 42680 6012
rect 42616 5952 42680 5956
rect 42696 6012 42760 6016
rect 42696 5956 42700 6012
rect 42700 5956 42756 6012
rect 42756 5956 42760 6012
rect 42696 5952 42760 5956
rect 42776 6012 42840 6016
rect 42776 5956 42780 6012
rect 42780 5956 42836 6012
rect 42836 5956 42840 6012
rect 42776 5952 42840 5956
rect 46796 5884 46860 5948
rect 46428 5748 46492 5812
rect 46796 5748 46860 5812
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 32140 5468 32204 5472
rect 32140 5412 32144 5468
rect 32144 5412 32200 5468
rect 32200 5412 32204 5468
rect 32140 5408 32204 5412
rect 32220 5468 32284 5472
rect 32220 5412 32224 5468
rect 32224 5412 32280 5468
rect 32280 5412 32284 5468
rect 32220 5408 32284 5412
rect 32300 5468 32364 5472
rect 32300 5412 32304 5468
rect 32304 5412 32360 5468
rect 32360 5412 32364 5468
rect 32300 5408 32364 5412
rect 32380 5468 32444 5472
rect 32380 5412 32384 5468
rect 32384 5412 32440 5468
rect 32440 5412 32444 5468
rect 32380 5408 32444 5412
rect 52932 5468 52996 5472
rect 52932 5412 52936 5468
rect 52936 5412 52992 5468
rect 52992 5412 52996 5468
rect 52932 5408 52996 5412
rect 53012 5468 53076 5472
rect 53012 5412 53016 5468
rect 53016 5412 53072 5468
rect 53072 5412 53076 5468
rect 53012 5408 53076 5412
rect 53092 5468 53156 5472
rect 53092 5412 53096 5468
rect 53096 5412 53152 5468
rect 53152 5412 53156 5468
rect 53092 5408 53156 5412
rect 53172 5468 53236 5472
rect 53172 5412 53176 5468
rect 53176 5412 53232 5468
rect 53232 5412 53236 5468
rect 53172 5408 53236 5412
rect 28948 5400 29012 5404
rect 28948 5344 28998 5400
rect 28998 5344 29012 5400
rect 28948 5340 29012 5344
rect 21744 4924 21808 4928
rect 21744 4868 21748 4924
rect 21748 4868 21804 4924
rect 21804 4868 21808 4924
rect 21744 4864 21808 4868
rect 21824 4924 21888 4928
rect 21824 4868 21828 4924
rect 21828 4868 21884 4924
rect 21884 4868 21888 4924
rect 21824 4864 21888 4868
rect 21904 4924 21968 4928
rect 21904 4868 21908 4924
rect 21908 4868 21964 4924
rect 21964 4868 21968 4924
rect 21904 4864 21968 4868
rect 21984 4924 22048 4928
rect 21984 4868 21988 4924
rect 21988 4868 22044 4924
rect 22044 4868 22048 4924
rect 21984 4864 22048 4868
rect 42536 4924 42600 4928
rect 42536 4868 42540 4924
rect 42540 4868 42596 4924
rect 42596 4868 42600 4924
rect 42536 4864 42600 4868
rect 42616 4924 42680 4928
rect 42616 4868 42620 4924
rect 42620 4868 42676 4924
rect 42676 4868 42680 4924
rect 42616 4864 42680 4868
rect 42696 4924 42760 4928
rect 42696 4868 42700 4924
rect 42700 4868 42756 4924
rect 42756 4868 42760 4924
rect 42696 4864 42760 4868
rect 42776 4924 42840 4928
rect 42776 4868 42780 4924
rect 42780 4868 42836 4924
rect 42836 4868 42840 4924
rect 42776 4864 42840 4868
rect 31708 4660 31772 4724
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 31708 4252 31772 4316
rect 32140 4380 32204 4384
rect 32140 4324 32144 4380
rect 32144 4324 32200 4380
rect 32200 4324 32204 4380
rect 32140 4320 32204 4324
rect 32220 4380 32284 4384
rect 32220 4324 32224 4380
rect 32224 4324 32280 4380
rect 32280 4324 32284 4380
rect 32220 4320 32284 4324
rect 32300 4380 32364 4384
rect 32300 4324 32304 4380
rect 32304 4324 32360 4380
rect 32360 4324 32364 4380
rect 32300 4320 32364 4324
rect 32380 4380 32444 4384
rect 32380 4324 32384 4380
rect 32384 4324 32440 4380
rect 32440 4324 32444 4380
rect 32380 4320 32444 4324
rect 52932 4380 52996 4384
rect 52932 4324 52936 4380
rect 52936 4324 52992 4380
rect 52992 4324 52996 4380
rect 52932 4320 52996 4324
rect 53012 4380 53076 4384
rect 53012 4324 53016 4380
rect 53016 4324 53072 4380
rect 53072 4324 53076 4380
rect 53012 4320 53076 4324
rect 53092 4380 53156 4384
rect 53092 4324 53096 4380
rect 53096 4324 53152 4380
rect 53152 4324 53156 4380
rect 53092 4320 53156 4324
rect 53172 4380 53236 4384
rect 53172 4324 53176 4380
rect 53176 4324 53232 4380
rect 53232 4324 53236 4380
rect 53172 4320 53236 4324
rect 21744 3836 21808 3840
rect 21744 3780 21748 3836
rect 21748 3780 21804 3836
rect 21804 3780 21808 3836
rect 21744 3776 21808 3780
rect 21824 3836 21888 3840
rect 21824 3780 21828 3836
rect 21828 3780 21884 3836
rect 21884 3780 21888 3836
rect 21824 3776 21888 3780
rect 21904 3836 21968 3840
rect 21904 3780 21908 3836
rect 21908 3780 21964 3836
rect 21964 3780 21968 3836
rect 21904 3776 21968 3780
rect 21984 3836 22048 3840
rect 21984 3780 21988 3836
rect 21988 3780 22044 3836
rect 22044 3780 22048 3836
rect 21984 3776 22048 3780
rect 42536 3836 42600 3840
rect 42536 3780 42540 3836
rect 42540 3780 42596 3836
rect 42596 3780 42600 3836
rect 42536 3776 42600 3780
rect 42616 3836 42680 3840
rect 42616 3780 42620 3836
rect 42620 3780 42676 3836
rect 42676 3780 42680 3836
rect 42616 3776 42680 3780
rect 42696 3836 42760 3840
rect 42696 3780 42700 3836
rect 42700 3780 42756 3836
rect 42756 3780 42760 3836
rect 42696 3776 42760 3780
rect 42776 3836 42840 3840
rect 42776 3780 42780 3836
rect 42780 3780 42836 3836
rect 42836 3780 42840 3836
rect 42776 3776 42840 3780
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 32140 3292 32204 3296
rect 32140 3236 32144 3292
rect 32144 3236 32200 3292
rect 32200 3236 32204 3292
rect 32140 3232 32204 3236
rect 32220 3292 32284 3296
rect 32220 3236 32224 3292
rect 32224 3236 32280 3292
rect 32280 3236 32284 3292
rect 32220 3232 32284 3236
rect 32300 3292 32364 3296
rect 32300 3236 32304 3292
rect 32304 3236 32360 3292
rect 32360 3236 32364 3292
rect 32300 3232 32364 3236
rect 32380 3292 32444 3296
rect 32380 3236 32384 3292
rect 32384 3236 32440 3292
rect 32440 3236 32444 3292
rect 32380 3232 32444 3236
rect 52932 3292 52996 3296
rect 52932 3236 52936 3292
rect 52936 3236 52992 3292
rect 52992 3236 52996 3292
rect 52932 3232 52996 3236
rect 53012 3292 53076 3296
rect 53012 3236 53016 3292
rect 53016 3236 53072 3292
rect 53072 3236 53076 3292
rect 53012 3232 53076 3236
rect 53092 3292 53156 3296
rect 53092 3236 53096 3292
rect 53096 3236 53152 3292
rect 53152 3236 53156 3292
rect 53092 3232 53156 3236
rect 53172 3292 53236 3296
rect 53172 3236 53176 3292
rect 53176 3236 53232 3292
rect 53232 3236 53236 3292
rect 53172 3232 53236 3236
rect 21744 2748 21808 2752
rect 21744 2692 21748 2748
rect 21748 2692 21804 2748
rect 21804 2692 21808 2748
rect 21744 2688 21808 2692
rect 21824 2748 21888 2752
rect 21824 2692 21828 2748
rect 21828 2692 21884 2748
rect 21884 2692 21888 2748
rect 21824 2688 21888 2692
rect 21904 2748 21968 2752
rect 21904 2692 21908 2748
rect 21908 2692 21964 2748
rect 21964 2692 21968 2748
rect 21904 2688 21968 2692
rect 21984 2748 22048 2752
rect 21984 2692 21988 2748
rect 21988 2692 22044 2748
rect 22044 2692 22048 2748
rect 21984 2688 22048 2692
rect 42536 2748 42600 2752
rect 42536 2692 42540 2748
rect 42540 2692 42596 2748
rect 42596 2692 42600 2748
rect 42536 2688 42600 2692
rect 42616 2748 42680 2752
rect 42616 2692 42620 2748
rect 42620 2692 42676 2748
rect 42676 2692 42680 2748
rect 42616 2688 42680 2692
rect 42696 2748 42760 2752
rect 42696 2692 42700 2748
rect 42700 2692 42756 2748
rect 42756 2692 42760 2748
rect 42696 2688 42760 2692
rect 42776 2748 42840 2752
rect 42776 2692 42780 2748
rect 42780 2692 42836 2748
rect 42836 2692 42840 2748
rect 42776 2688 42840 2692
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 32140 2204 32204 2208
rect 32140 2148 32144 2204
rect 32144 2148 32200 2204
rect 32200 2148 32204 2204
rect 32140 2144 32204 2148
rect 32220 2204 32284 2208
rect 32220 2148 32224 2204
rect 32224 2148 32280 2204
rect 32280 2148 32284 2204
rect 32220 2144 32284 2148
rect 32300 2204 32364 2208
rect 32300 2148 32304 2204
rect 32304 2148 32360 2204
rect 32360 2148 32364 2204
rect 32300 2144 32364 2148
rect 32380 2204 32444 2208
rect 32380 2148 32384 2204
rect 32384 2148 32440 2204
rect 32440 2148 32444 2204
rect 32380 2144 32444 2148
rect 52932 2204 52996 2208
rect 52932 2148 52936 2204
rect 52936 2148 52992 2204
rect 52992 2148 52996 2204
rect 52932 2144 52996 2148
rect 53012 2204 53076 2208
rect 53012 2148 53016 2204
rect 53016 2148 53072 2204
rect 53072 2148 53076 2204
rect 53012 2144 53076 2148
rect 53092 2204 53156 2208
rect 53092 2148 53096 2204
rect 53096 2148 53152 2204
rect 53152 2148 53156 2204
rect 53092 2144 53156 2148
rect 53172 2204 53236 2208
rect 53172 2148 53176 2204
rect 53176 2148 53232 2204
rect 53232 2148 53236 2204
rect 53172 2144 53236 2148
<< metal4 >>
rect 11340 17440 11660 17456
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 21736 16896 22056 17456
rect 21736 16832 21744 16896
rect 21808 16832 21824 16896
rect 21888 16832 21904 16896
rect 21968 16832 21984 16896
rect 22048 16832 22056 16896
rect 21736 15808 22056 16832
rect 21736 15744 21744 15808
rect 21808 15744 21824 15808
rect 21888 15744 21904 15808
rect 21968 15744 21984 15808
rect 22048 15744 22056 15808
rect 21736 14720 22056 15744
rect 21736 14656 21744 14720
rect 21808 14656 21824 14720
rect 21888 14656 21904 14720
rect 21968 14656 21984 14720
rect 22048 14656 22056 14720
rect 21736 13632 22056 14656
rect 21736 13568 21744 13632
rect 21808 13568 21824 13632
rect 21888 13568 21904 13632
rect 21968 13568 21984 13632
rect 22048 13568 22056 13632
rect 21736 12544 22056 13568
rect 21736 12480 21744 12544
rect 21808 12480 21824 12544
rect 21888 12480 21904 12544
rect 21968 12480 21984 12544
rect 22048 12480 22056 12544
rect 21736 11456 22056 12480
rect 21736 11392 21744 11456
rect 21808 11392 21824 11456
rect 21888 11392 21904 11456
rect 21968 11392 21984 11456
rect 22048 11392 22056 11456
rect 21736 10368 22056 11392
rect 21736 10304 21744 10368
rect 21808 10304 21824 10368
rect 21888 10304 21904 10368
rect 21968 10304 21984 10368
rect 22048 10304 22056 10368
rect 21736 9280 22056 10304
rect 21736 9216 21744 9280
rect 21808 9216 21824 9280
rect 21888 9216 21904 9280
rect 21968 9216 21984 9280
rect 22048 9216 22056 9280
rect 21736 8192 22056 9216
rect 32132 17440 32452 17456
rect 32132 17376 32140 17440
rect 32204 17376 32220 17440
rect 32284 17376 32300 17440
rect 32364 17376 32380 17440
rect 32444 17376 32452 17440
rect 32132 16352 32452 17376
rect 32132 16288 32140 16352
rect 32204 16288 32220 16352
rect 32284 16288 32300 16352
rect 32364 16288 32380 16352
rect 32444 16288 32452 16352
rect 32132 15264 32452 16288
rect 32132 15200 32140 15264
rect 32204 15200 32220 15264
rect 32284 15200 32300 15264
rect 32364 15200 32380 15264
rect 32444 15200 32452 15264
rect 32132 14176 32452 15200
rect 32132 14112 32140 14176
rect 32204 14112 32220 14176
rect 32284 14112 32300 14176
rect 32364 14112 32380 14176
rect 32444 14112 32452 14176
rect 32132 13088 32452 14112
rect 32132 13024 32140 13088
rect 32204 13024 32220 13088
rect 32284 13024 32300 13088
rect 32364 13024 32380 13088
rect 32444 13024 32452 13088
rect 32132 12000 32452 13024
rect 32132 11936 32140 12000
rect 32204 11936 32220 12000
rect 32284 11936 32300 12000
rect 32364 11936 32380 12000
rect 32444 11936 32452 12000
rect 32132 10912 32452 11936
rect 32132 10848 32140 10912
rect 32204 10848 32220 10912
rect 32284 10848 32300 10912
rect 32364 10848 32380 10912
rect 32444 10848 32452 10912
rect 32132 9824 32452 10848
rect 32132 9760 32140 9824
rect 32204 9760 32220 9824
rect 32284 9760 32300 9824
rect 32364 9760 32380 9824
rect 32444 9760 32452 9824
rect 32132 8736 32452 9760
rect 32132 8672 32140 8736
rect 32204 8672 32220 8736
rect 32284 8672 32300 8736
rect 32364 8672 32380 8736
rect 32444 8672 32452 8736
rect 28947 8260 29013 8261
rect 28947 8196 28948 8260
rect 29012 8196 29013 8260
rect 28947 8195 29013 8196
rect 21736 8128 21744 8192
rect 21808 8128 21824 8192
rect 21888 8128 21904 8192
rect 21968 8128 21984 8192
rect 22048 8128 22056 8192
rect 21736 7104 22056 8128
rect 21736 7040 21744 7104
rect 21808 7040 21824 7104
rect 21888 7040 21904 7104
rect 21968 7040 21984 7104
rect 22048 7040 22056 7104
rect 21736 6016 22056 7040
rect 21736 5952 21744 6016
rect 21808 5952 21824 6016
rect 21888 5952 21904 6016
rect 21968 5952 21984 6016
rect 22048 5952 22056 6016
rect 21736 4928 22056 5952
rect 28950 5405 29010 8195
rect 32132 7648 32452 8672
rect 32132 7584 32140 7648
rect 32204 7584 32220 7648
rect 32284 7584 32300 7648
rect 32364 7584 32380 7648
rect 32444 7584 32452 7648
rect 32132 6560 32452 7584
rect 32132 6496 32140 6560
rect 32204 6496 32220 6560
rect 32284 6496 32300 6560
rect 32364 6496 32380 6560
rect 32444 6496 32452 6560
rect 32132 5472 32452 6496
rect 32132 5408 32140 5472
rect 32204 5408 32220 5472
rect 32284 5408 32300 5472
rect 32364 5408 32380 5472
rect 32444 5408 32452 5472
rect 28947 5404 29013 5405
rect 28947 5340 28948 5404
rect 29012 5340 29013 5404
rect 28947 5339 29013 5340
rect 21736 4864 21744 4928
rect 21808 4864 21824 4928
rect 21888 4864 21904 4928
rect 21968 4864 21984 4928
rect 22048 4864 22056 4928
rect 21736 3840 22056 4864
rect 31707 4724 31773 4725
rect 31707 4660 31708 4724
rect 31772 4660 31773 4724
rect 31707 4659 31773 4660
rect 31710 4317 31770 4659
rect 32132 4384 32452 5408
rect 32132 4320 32140 4384
rect 32204 4320 32220 4384
rect 32284 4320 32300 4384
rect 32364 4320 32380 4384
rect 32444 4320 32452 4384
rect 31707 4316 31773 4317
rect 31707 4252 31708 4316
rect 31772 4252 31773 4316
rect 31707 4251 31773 4252
rect 21736 3776 21744 3840
rect 21808 3776 21824 3840
rect 21888 3776 21904 3840
rect 21968 3776 21984 3840
rect 22048 3776 22056 3840
rect 21736 2752 22056 3776
rect 21736 2688 21744 2752
rect 21808 2688 21824 2752
rect 21888 2688 21904 2752
rect 21968 2688 21984 2752
rect 22048 2688 22056 2752
rect 21736 2128 22056 2688
rect 32132 3296 32452 4320
rect 32132 3232 32140 3296
rect 32204 3232 32220 3296
rect 32284 3232 32300 3296
rect 32364 3232 32380 3296
rect 32444 3232 32452 3296
rect 32132 2208 32452 3232
rect 32132 2144 32140 2208
rect 32204 2144 32220 2208
rect 32284 2144 32300 2208
rect 32364 2144 32380 2208
rect 32444 2144 32452 2208
rect 32132 2128 32452 2144
rect 42528 16896 42848 17456
rect 42528 16832 42536 16896
rect 42600 16832 42616 16896
rect 42680 16832 42696 16896
rect 42760 16832 42776 16896
rect 42840 16832 42848 16896
rect 42528 15808 42848 16832
rect 42528 15744 42536 15808
rect 42600 15744 42616 15808
rect 42680 15744 42696 15808
rect 42760 15744 42776 15808
rect 42840 15744 42848 15808
rect 42528 14720 42848 15744
rect 42528 14656 42536 14720
rect 42600 14656 42616 14720
rect 42680 14656 42696 14720
rect 42760 14656 42776 14720
rect 42840 14656 42848 14720
rect 42528 13632 42848 14656
rect 42528 13568 42536 13632
rect 42600 13568 42616 13632
rect 42680 13568 42696 13632
rect 42760 13568 42776 13632
rect 42840 13568 42848 13632
rect 42528 12544 42848 13568
rect 42528 12480 42536 12544
rect 42600 12480 42616 12544
rect 42680 12480 42696 12544
rect 42760 12480 42776 12544
rect 42840 12480 42848 12544
rect 42528 11456 42848 12480
rect 42528 11392 42536 11456
rect 42600 11392 42616 11456
rect 42680 11392 42696 11456
rect 42760 11392 42776 11456
rect 42840 11392 42848 11456
rect 42528 10368 42848 11392
rect 42528 10304 42536 10368
rect 42600 10304 42616 10368
rect 42680 10304 42696 10368
rect 42760 10304 42776 10368
rect 42840 10304 42848 10368
rect 42528 9280 42848 10304
rect 42528 9216 42536 9280
rect 42600 9216 42616 9280
rect 42680 9216 42696 9280
rect 42760 9216 42776 9280
rect 42840 9216 42848 9280
rect 42528 8192 42848 9216
rect 42528 8128 42536 8192
rect 42600 8128 42616 8192
rect 42680 8128 42696 8192
rect 42760 8128 42776 8192
rect 42840 8128 42848 8192
rect 42528 7104 42848 8128
rect 42528 7040 42536 7104
rect 42600 7040 42616 7104
rect 42680 7040 42696 7104
rect 42760 7040 42776 7104
rect 42840 7040 42848 7104
rect 42528 6016 42848 7040
rect 52924 17440 53244 17456
rect 52924 17376 52932 17440
rect 52996 17376 53012 17440
rect 53076 17376 53092 17440
rect 53156 17376 53172 17440
rect 53236 17376 53244 17440
rect 52924 16352 53244 17376
rect 52924 16288 52932 16352
rect 52996 16288 53012 16352
rect 53076 16288 53092 16352
rect 53156 16288 53172 16352
rect 53236 16288 53244 16352
rect 52924 15264 53244 16288
rect 52924 15200 52932 15264
rect 52996 15200 53012 15264
rect 53076 15200 53092 15264
rect 53156 15200 53172 15264
rect 53236 15200 53244 15264
rect 52924 14176 53244 15200
rect 52924 14112 52932 14176
rect 52996 14112 53012 14176
rect 53076 14112 53092 14176
rect 53156 14112 53172 14176
rect 53236 14112 53244 14176
rect 52924 13088 53244 14112
rect 52924 13024 52932 13088
rect 52996 13024 53012 13088
rect 53076 13024 53092 13088
rect 53156 13024 53172 13088
rect 53236 13024 53244 13088
rect 52924 12000 53244 13024
rect 52924 11936 52932 12000
rect 52996 11936 53012 12000
rect 53076 11936 53092 12000
rect 53156 11936 53172 12000
rect 53236 11936 53244 12000
rect 52924 10912 53244 11936
rect 52924 10848 52932 10912
rect 52996 10848 53012 10912
rect 53076 10848 53092 10912
rect 53156 10848 53172 10912
rect 53236 10848 53244 10912
rect 52924 9824 53244 10848
rect 52924 9760 52932 9824
rect 52996 9760 53012 9824
rect 53076 9760 53092 9824
rect 53156 9760 53172 9824
rect 53236 9760 53244 9824
rect 52924 8736 53244 9760
rect 52924 8672 52932 8736
rect 52996 8672 53012 8736
rect 53076 8672 53092 8736
rect 53156 8672 53172 8736
rect 53236 8672 53244 8736
rect 52924 7648 53244 8672
rect 52924 7584 52932 7648
rect 52996 7584 53012 7648
rect 53076 7584 53092 7648
rect 53156 7584 53172 7648
rect 53236 7584 53244 7648
rect 46795 6628 46861 6629
rect 46795 6564 46796 6628
rect 46860 6564 46861 6628
rect 46795 6563 46861 6564
rect 42528 5952 42536 6016
rect 42600 5952 42616 6016
rect 42680 5952 42696 6016
rect 42760 5952 42776 6016
rect 42840 5952 42848 6016
rect 42528 4928 42848 5952
rect 46798 5949 46858 6563
rect 52924 6560 53244 7584
rect 52924 6496 52932 6560
rect 52996 6496 53012 6560
rect 53076 6496 53092 6560
rect 53156 6496 53172 6560
rect 53236 6496 53244 6560
rect 46795 5948 46861 5949
rect 46795 5884 46796 5948
rect 46860 5884 46861 5948
rect 46795 5883 46861 5884
rect 46427 5812 46493 5813
rect 46427 5748 46428 5812
rect 46492 5810 46493 5812
rect 46795 5812 46861 5813
rect 46795 5810 46796 5812
rect 46492 5750 46796 5810
rect 46492 5748 46493 5750
rect 46427 5747 46493 5748
rect 46795 5748 46796 5750
rect 46860 5748 46861 5812
rect 46795 5747 46861 5748
rect 42528 4864 42536 4928
rect 42600 4864 42616 4928
rect 42680 4864 42696 4928
rect 42760 4864 42776 4928
rect 42840 4864 42848 4928
rect 42528 3840 42848 4864
rect 42528 3776 42536 3840
rect 42600 3776 42616 3840
rect 42680 3776 42696 3840
rect 42760 3776 42776 3840
rect 42840 3776 42848 3840
rect 42528 2752 42848 3776
rect 42528 2688 42536 2752
rect 42600 2688 42616 2752
rect 42680 2688 42696 2752
rect 42760 2688 42776 2752
rect 42840 2688 42848 2752
rect 42528 2128 42848 2688
rect 52924 5472 53244 6496
rect 52924 5408 52932 5472
rect 52996 5408 53012 5472
rect 53076 5408 53092 5472
rect 53156 5408 53172 5472
rect 53236 5408 53244 5472
rect 52924 4384 53244 5408
rect 52924 4320 52932 4384
rect 52996 4320 53012 4384
rect 53076 4320 53092 4384
rect 53156 4320 53172 4384
rect 53236 4320 53244 4384
rect 52924 3296 53244 4320
rect 52924 3232 52932 3296
rect 52996 3232 53012 3296
rect 53076 3232 53092 3296
rect 53156 3232 53172 3296
rect 53236 3232 53244 3296
rect 52924 2208 53244 3232
rect 52924 2144 52932 2208
rect 52996 2144 53012 2208
rect 53076 2144 53092 2208
rect 53156 2144 53172 2208
rect 53236 2144 53244 2208
rect 52924 2128 53244 2144
use sky130_fd_sc_hd__decap_4  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 1380 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1607721120
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 2024 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 1748 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12
timestamp 1607721120
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9
timestamp 1607721120
transform 1 0 1932 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1417__CLK $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1416__CLK
timestamp 1607721120
transform 1 0 1840 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1415__CLK
timestamp 1607721120
transform 1 0 2208 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_18
timestamp 1607721120
transform 1 0 2760 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_14
timestamp 1607721120
transform 1 0 2392 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16
timestamp 1607721120
transform 1 0 2576 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1414__CLK
timestamp 1607721120
transform 1 0 2392 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1412__CLK
timestamp 1607721120
transform 1 0 2760 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__B
timestamp 1607721120
transform 1 0 2944 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__A
timestamp 1607721120
transform 1 0 2576 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0676_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 2944 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_22
timestamp 1607721120
transform 1 0 3128 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32
timestamp 1607721120
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27
timestamp 1607721120
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23
timestamp 1607721120
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1415__D
timestamp 1607721120
transform 1 0 3496 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1414__D
timestamp 1607721120
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__A
timestamp 1607721120
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1415_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 3680 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1414_
timestamp 1607721120
transform 1 0 4324 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1607721120
transform 1 0 6072 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_51
timestamp 1607721120
transform 1 0 5796 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_47
timestamp 1607721120
transform 1 0 5428 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1607721120
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__B1
timestamp 1607721120
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__A1
timestamp 1607721120
transform 1 0 6256 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__C1
timestamp 1607721120
transform 1 0 5888 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_58
timestamp 1607721120
transform 1 0 6440 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63
timestamp 1607721120
transform 1 0 6900 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58
timestamp 1607721120
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1412__D
timestamp 1607721120
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1607721120
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1607721120
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1412_
timestamp 1607721120
transform 1 0 7176 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__a211o_4  _1023_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 6808 0 1 2720
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_1_80
timestamp 1607721120
transform 1 0 8464 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_76
timestamp 1607721120
transform 1 0 8096 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89
timestamp 1607721120
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1607721120
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__B1
timestamp 1607721120
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__A
timestamp 1607721120
transform 1 0 8648 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__C1
timestamp 1607721120
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__B
timestamp 1607721120
transform 1 0 8280 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1034_
timestamp 1607721120
transform 1 0 8832 0 1 2720
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_1_98
timestamp 1607721120
transform 1 0 10120 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_99
timestamp 1607721120
transform 1 0 10212 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_94
timestamp 1607721120
transform 1 0 9752 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__C
timestamp 1607721120
transform 1 0 10028 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__B
timestamp 1607721120
transform 1 0 10396 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__A1
timestamp 1607721120
transform 1 0 10304 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1607721120
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_102
timestamp 1607721120
transform 1 0 10488 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103
timestamp 1607721120
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__A
timestamp 1607721120
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__A1
timestamp 1607721120
transform 1 0 10764 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1022_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 10948 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1008_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 10948 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_1_114
timestamp 1607721120
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_118
timestamp 1607721120
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_116
timestamp 1607721120
transform 1 0 11776 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__B
timestamp 1607721120
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_123
timestamp 1607721120
transform 1 0 12420 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_123
timestamp 1607721120
transform 1 0 12420 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_120
timestamp 1607721120
transform 1 0 12144 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__B1
timestamp 1607721120
transform 1 0 12236 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__B2
timestamp 1607721120
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1607721120
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_125
timestamp 1607721120
transform 1 0 12604 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1607721120
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_129
timestamp 1607721120
transform 1 0 12972 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__B1
timestamp 1607721120
transform 1 0 13340 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__A1_N
timestamp 1607721120
transform 1 0 12788 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1009_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 12696 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_4  _0992_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 13524 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_146
timestamp 1607721120
transform 1 0 14536 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_142
timestamp 1607721120
transform 1 0 14168 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_138
timestamp 1607721120
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_147
timestamp 1607721120
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__B1
timestamp 1607721120
transform 1 0 14720 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__A2
timestamp 1607721120
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__A1
timestamp 1607721120
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_151
timestamp 1607721120
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__A1
timestamp 1607721120
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1417__D
timestamp 1607721120
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1607721120
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1417_
timestamp 1607721120
transform 1 0 15456 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__a211o_4  _1001_
timestamp 1607721120
transform 1 0 14904 0 1 2720
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_1_164
timestamp 1607721120
transform 1 0 16192 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_168
timestamp 1607721120
transform 1 0 16560 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__B1
timestamp 1607721120
transform 1 0 16376 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_172
timestamp 1607721120
transform 1 0 16928 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__A2
timestamp 1607721120
transform 1 0 16744 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_179
timestamp 1607721120
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_176
timestamp 1607721120
transform 1 0 17296 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_179
timestamp 1607721120
transform 1 0 17572 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_175
timestamp 1607721120
transform 1 0 17204 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__A
timestamp 1607721120
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_182
timestamp 1607721120
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__C
timestamp 1607721120
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__B
timestamp 1607721120
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__B
timestamp 1607721120
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1607721120
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1607721120
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1090_
timestamp 1607721120
transform 1 0 18308 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and3_4  _0999_
timestamp 1607721120
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_197
timestamp 1607721120
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_193
timestamp 1607721120
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1607721120
transform 1 0 18952 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__B
timestamp 1607721120
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__A
timestamp 1607721120
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_201
timestamp 1607721120
transform 1 0 19596 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_198
timestamp 1607721120
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__B
timestamp 1607721120
transform 1 0 19504 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__B
timestamp 1607721120
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1036_
timestamp 1607721120
transform 1 0 19688 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and3_4  _1007_
timestamp 1607721120
transform 1 0 19872 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_213
timestamp 1607721120
transform 1 0 20700 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_213
timestamp 1607721120
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_209
timestamp 1607721120
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1411__D
timestamp 1607721120
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__A
timestamp 1607721120
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_220
timestamp 1607721120
transform 1 0 21344 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_217
timestamp 1607721120
transform 1 0 21068 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_218
timestamp 1607721120
transform 1 0 21160 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1416__D
timestamp 1607721120
transform 1 0 21160 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1607721120
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1411_
timestamp 1607721120
transform 1 0 21436 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__a211o_4  _1039_
timestamp 1607721120
transform 1 0 21528 0 1 2720
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_1_236
timestamp 1607721120
transform 1 0 22816 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__A1
timestamp 1607721120
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_240
timestamp 1607721120
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_244
timestamp 1607721120
transform 1 0 23552 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_240
timestamp 1607721120
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__B1_N
timestamp 1607721120
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__A
timestamp 1607721120
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1032__A2
timestamp 1607721120
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1607721120
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1607721120
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1038_
timestamp 1607721120
transform 1 0 24012 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_4  _1037_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 23644 0 1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_1_258
timestamp 1607721120
transform 1 0 24840 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_258
timestamp 1607721120
transform 1 0 24840 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__A2
timestamp 1607721120
transform 1 0 25024 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_265
timestamp 1607721120
transform 1 0 25484 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_262
timestamp 1607721120
transform 1 0 25208 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_262
timestamp 1607721120
transform 1 0 25208 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__B
timestamp 1607721120
transform 1 0 25392 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__A
timestamp 1607721120
transform 1 0 25300 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_269
timestamp 1607721120
transform 1 0 25852 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_270
timestamp 1607721120
transform 1 0 25944 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1032__B1
timestamp 1607721120
transform 1 0 25668 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0917_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 25576 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_273
timestamp 1607721120
transform 1 0 26220 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_274
timestamp 1607721120
transform 1 0 26312 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__C
timestamp 1607721120
transform 1 0 26036 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__A
timestamp 1607721120
transform 1 0 26128 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_295
timestamp 1607721120
transform 1 0 28244 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_291
timestamp 1607721120
transform 1 0 27876 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__B1
timestamp 1607721120
transform 1 0 26404 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1410__D
timestamp 1607721120
transform 1 0 26588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__A1
timestamp 1607721120
transform 1 0 28336 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1607721120
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1410_
timestamp 1607721120
transform 1 0 26864 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__a211o_4  _1045_
timestamp 1607721120
transform 1 0 26588 0 1 2720
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_1_302
timestamp 1607721120
transform 1 0 28888 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_298
timestamp 1607721120
transform 1 0 28520 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_303
timestamp 1607721120
transform 1 0 28980 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_299
timestamp 1607721120
transform 1 0 28612 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__B1
timestamp 1607721120
transform 1 0 28796 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__A1
timestamp 1607721120
transform 1 0 28704 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_311
timestamp 1607721120
transform 1 0 29716 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_307
timestamp 1607721120
transform 1 0 29348 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__A3
timestamp 1607721120
transform 1 0 29164 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1607721120
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1607721120
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1040_
timestamp 1607721120
transform 1 0 29256 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_1_317
timestamp 1607721120
transform 1 0 30268 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_313
timestamp 1607721120
transform 1 0 29900 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_316
timestamp 1607721120
transform 1 0 30176 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__B1
timestamp 1607721120
transform 1 0 29992 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__A2
timestamp 1607721120
transform 1 0 30360 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__A
timestamp 1607721120
transform 1 0 30452 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1040__A
timestamp 1607721120
transform 1 0 30084 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_339
timestamp 1607721120
transform 1 0 32292 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_334
timestamp 1607721120
transform 1 0 31832 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1607721120
transform 1 0 32108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_333
timestamp 1607721120
transform 1 0 31740 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__B
timestamp 1607721120
transform 1 0 32292 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__A1
timestamp 1607721120
transform 1 0 31924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__A
timestamp 1607721120
transform 1 0 32108 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__D
timestamp 1607721120
transform 1 0 32476 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1607721120
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1425_
timestamp 1607721120
transform 1 0 32568 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__a21oi_4  _0930_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 30544 0 -1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _0929_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 30636 0 1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_1_347
timestamp 1607721120
transform 1 0 33028 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_343
timestamp 1607721120
transform 1 0 32660 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1425__D
timestamp 1607721120
transform 1 0 32844 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0913_
timestamp 1607721120
transform 1 0 33212 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_362
timestamp 1607721120
transform 1 0 34408 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_358
timestamp 1607721120
transform 1 0 34040 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_361
timestamp 1607721120
transform 1 0 34316 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__B
timestamp 1607721120
transform 1 0 34224 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1607721120
transform 1 0 34684 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__A1
timestamp 1607721120
transform 1 0 34500 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__A2
timestamp 1607721120
transform 1 0 34592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_375
timestamp 1607721120
transform 1 0 35604 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_371
timestamp 1607721120
transform 1 0 35236 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_373
timestamp 1607721120
transform 1 0 35420 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_369
timestamp 1607721120
transform 1 0 35052 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__A
timestamp 1607721120
transform 1 0 34868 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__B
timestamp 1607721120
transform 1 0 35696 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1607721120
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1607721120
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1041_
timestamp 1607721120
transform 1 0 34868 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_378
timestamp 1607721120
transform 1 0 35880 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0695__A
timestamp 1607721120
transform 1 0 35788 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0702_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 36064 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_4  _0695_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 35972 0 -1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_1_393
timestamp 1607721120
transform 1 0 37260 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_389
timestamp 1607721120
transform 1 0 36892 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_392
timestamp 1607721120
transform 1 0 37168 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__D
timestamp 1607721120
transform 1 0 37076 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_397
timestamp 1607721120
transform 1 0 37628 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_396
timestamp 1607721120
transform 1 0 37536 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0695__B
timestamp 1607721120
transform 1 0 37352 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_400
timestamp 1607721120
transform 1 0 37904 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1199__C
timestamp 1607721120
transform 1 0 37720 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0695__C
timestamp 1607721120
transform 1 0 37720 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1158_
timestamp 1607721120
transform 1 0 37904 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_404
timestamp 1607721120
transform 1 0 38272 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_404
timestamp 1607721120
transform 1 0 38272 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__B
timestamp 1607721120
transform 1 0 38456 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1607721120
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1161_
timestamp 1607721120
transform 1 0 38364 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_408
timestamp 1607721120
transform 1 0 38640 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_409
timestamp 1607721120
transform 1 0 38732 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1161__A
timestamp 1607721120
transform 1 0 38916 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__A
timestamp 1607721120
transform 1 0 38824 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_419
timestamp 1607721120
transform 1 0 39652 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_413
timestamp 1607721120
transform 1 0 39100 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1199__A
timestamp 1607721120
transform 1 0 39284 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1193__A
timestamp 1607721120
transform 1 0 39836 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1199_
timestamp 1607721120
transform 1 0 39468 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1193_
timestamp 1607721120
transform 1 0 39008 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_1_423
timestamp 1607721120
transform 1 0 40020 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_433
timestamp 1607721120
transform 1 0 40940 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_430
timestamp 1607721120
transform 1 0 40664 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_426
timestamp 1607721120
transform 1 0 40296 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__C1
timestamp 1607721120
transform 1 0 40204 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1386__D
timestamp 1607721120
transform 1 0 40756 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1607721120
transform 1 0 40388 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1386_
timestamp 1607721120
transform 1 0 40480 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_0_439
timestamp 1607721120
transform 1 0 41492 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_435
timestamp 1607721120
transform 1 0 41124 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__D
timestamp 1607721120
transform 1 0 41584 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1607721120
transform 1 0 41032 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0675_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 41768 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_451
timestamp 1607721120
transform 1 0 42596 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_447
timestamp 1607721120
transform 1 0 42228 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_451
timestamp 1607721120
transform 1 0 42596 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1196__C1
timestamp 1607721120
transform 1 0 42780 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__C
timestamp 1607721120
transform 1 0 42412 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__A
timestamp 1607721120
transform 1 0 42780 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_455
timestamp 1607721120
transform 1 0 42964 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0674_
timestamp 1607721120
transform 1 0 42964 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_465
timestamp 1607721120
transform 1 0 43884 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_462
timestamp 1607721120
transform 1 0 43608 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_458
timestamp 1607721120
transform 1 0 43240 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_466
timestamp 1607721120
transform 1 0 43976 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_459
timestamp 1607721120
transform 1 0 43332 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__B
timestamp 1607721120
transform 1 0 43148 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1387__D
timestamp 1607721120
transform 1 0 43700 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__D
timestamp 1607721120
transform 1 0 43700 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1607721120
transform 1 0 43884 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1387_
timestamp 1607721120
transform 1 0 44252 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__a211o_4  _1196_
timestamp 1607721120
transform 1 0 43976 0 1 2720
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_1_484
timestamp 1607721120
transform 1 0 45632 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_480
timestamp 1607721120
transform 1 0 45264 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_488
timestamp 1607721120
transform 1 0 46000 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1388__D
timestamp 1607721120
transform 1 0 46184 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__A
timestamp 1607721120
transform 1 0 45816 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__B
timestamp 1607721120
transform 1 0 45448 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1607721120
transform 1 0 46000 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_502
timestamp 1607721120
transform 1 0 47288 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 1607721120
transform 1 0 47196 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_492
timestamp 1607721120
transform 1 0 46368 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__A
timestamp 1607721120
transform 1 0 46552 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1607721120
transform 1 0 46736 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1174_
timestamp 1607721120
transform 1 0 46828 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_4  _1194_
timestamp 1607721120
transform 1 0 46092 0 1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_1_510
timestamp 1607721120
transform 1 0 48024 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_506
timestamp 1607721120
transform 1 0 47656 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_506
timestamp 1607721120
transform 1 0 47656 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__A2
timestamp 1607721120
transform 1 0 47840 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__A1
timestamp 1607721120
transform 1 0 47472 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__C
timestamp 1607721120
transform 1 0 47472 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__D
timestamp 1607721120
transform 1 0 47840 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0685_
timestamp 1607721120
transform 1 0 48024 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_520
timestamp 1607721120
transform 1 0 48944 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_516
timestamp 1607721120
transform 1 0 48576 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_523
timestamp 1607721120
transform 1 0 49220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_519
timestamp 1607721120
transform 1 0 48852 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__B1_N
timestamp 1607721120
transform 1 0 48760 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__A
timestamp 1607721120
transform 1 0 49128 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__C
timestamp 1607721120
transform 1 0 49404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__A
timestamp 1607721120
transform 1 0 48392 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__B
timestamp 1607721120
transform 1 0 49036 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__nor4_4  _0682_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 49312 0 1 2720
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_0_528
timestamp 1607721120
transform 1 0 49680 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__B
timestamp 1607721120
transform 1 0 49864 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1607721120
transform 1 0 49588 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0705_
timestamp 1607721120
transform 1 0 50048 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_541
timestamp 1607721120
transform 1 0 50876 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_541
timestamp 1607721120
transform 1 0 50876 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__C
timestamp 1607721120
transform 1 0 51060 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__A
timestamp 1607721120
transform 1 0 51060 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_545
timestamp 1607721120
transform 1 0 51244 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_545
timestamp 1607721120
transform 1 0 51244 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__D
timestamp 1607721120
transform 1 0 51428 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__D
timestamp 1607721120
transform 1 0 51428 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_550
timestamp 1607721120
transform 1 0 51704 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_554
timestamp 1607721120
transform 1 0 52072 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_549
timestamp 1607721120
transform 1 0 51612 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__B
timestamp 1607721120
transform 1 0 51888 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__D
timestamp 1607721120
transform 1 0 52256 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__C
timestamp 1607721120
transform 1 0 52072 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1607721120
transform 1 0 51612 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0688_
timestamp 1607721120
transform 1 0 52256 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_565
timestamp 1607721120
transform 1 0 53084 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_563
timestamp 1607721120
transform 1 0 52900 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_559
timestamp 1607721120
transform 1 0 52532 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__B
timestamp 1607721120
transform 1 0 52992 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__A
timestamp 1607721120
transform 1 0 53268 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1607721120
transform 1 0 52440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0679_
timestamp 1607721120
transform 1 0 53176 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_569
timestamp 1607721120
transform 1 0 53452 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_579
timestamp 1607721120
transform 1 0 54372 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_575
timestamp 1607721120
transform 1 0 54004 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__C
timestamp 1607721120
transform 1 0 53636 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__A
timestamp 1607721120
transform 1 0 54188 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1179_
timestamp 1607721120
transform 1 0 53820 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_582
timestamp 1607721120
transform 1 0 54648 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_583
timestamp 1607721120
transform 1 0 54740 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__A
timestamp 1607721120
transform 1 0 54556 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_586
timestamp 1607721120
transform 1 0 55016 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__C
timestamp 1607721120
transform 1 0 54924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__B
timestamp 1607721120
transform 1 0 54832 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_587
timestamp 1607721120
transform 1 0 55108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__A
timestamp 1607721120
transform 1 0 55200 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1607721120
transform 1 0 55292 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_590
timestamp 1607721120
transform 1 0 55384 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_590
timestamp 1607721120
transform 1 0 55384 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1154__B
timestamp 1607721120
transform 1 0 55568 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__B
timestamp 1607721120
transform 1 0 55568 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_594
timestamp 1607721120
transform 1 0 55752 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_598
timestamp 1607721120
transform 1 0 56120 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_594
timestamp 1607721120
transform 1 0 55752 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1387__CLK
timestamp 1607721120
transform 1 0 55936 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1154__C
timestamp 1607721120
transform 1 0 55936 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1152_
timestamp 1607721120
transform 1 0 56120 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_602
timestamp 1607721120
transform 1 0 56488 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_602
timestamp 1607721120
transform 1 0 56488 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1388__CLK
timestamp 1607721120
transform 1 0 56304 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1390__CLK
timestamp 1607721120
transform 1 0 56672 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1165__B
timestamp 1607721120
transform 1 0 56672 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_615
timestamp 1607721120
transform 1 0 57684 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_611
timestamp 1607721120
transform 1 0 57316 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_606
timestamp 1607721120
transform 1 0 56856 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1165__A
timestamp 1607721120
transform 1 0 57040 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__B1
timestamp 1607721120
transform 1 0 57500 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1607721120
transform 1 0 57224 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_606 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 56856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_619
timestamp 1607721120
transform 1 0 58052 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1391__CLK
timestamp 1607721120
transform 1 0 57960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__B
timestamp 1607721120
transform 1 0 57868 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1607721120
transform 1 0 58144 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_623
timestamp 1607721120
transform 1 0 58420 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_621
timestamp 1607721120
transform 1 0 58236 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__C
timestamp 1607721120
transform 1 0 58512 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__C1
timestamp 1607721120
transform 1 0 58236 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_626
timestamp 1607721120
transform 1 0 58696 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__A
timestamp 1607721120
transform 1 0 58604 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__D
timestamp 1607721120
transform 1 0 58880 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_630
timestamp 1607721120
transform 1 0 59064 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__B
timestamp 1607721120
transform 1 0 59248 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0681_
timestamp 1607721120
transform 1 0 59432 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _1176_
timestamp 1607721120
transform 1 0 58788 0 1 2720
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_1_645
timestamp 1607721120
transform 1 0 60444 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_641
timestamp 1607721120
transform 1 0 60076 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_647
timestamp 1607721120
transform 1 0 60628 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_643
timestamp 1607721120
transform 1 0 60260 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__C
timestamp 1607721120
transform 1 0 60812 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1172__A
timestamp 1607721120
transform 1 0 60260 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__D
timestamp 1607721120
transform 1 0 60628 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__A
timestamp 1607721120
transform 1 0 60444 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0690_
timestamp 1607721120
transform 1 0 60812 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_658
timestamp 1607721120
transform 1 0 61640 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_659
timestamp 1607721120
transform 1 0 61732 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_655
timestamp 1607721120
transform 1 0 61364 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0680__A
timestamp 1607721120
transform 1 0 61548 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1607721120
transform 1 0 60996 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0680_
timestamp 1607721120
transform 1 0 61088 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_662
timestamp 1607721120
transform 1 0 62008 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__A
timestamp 1607721120
transform 1 0 61824 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_666
timestamp 1607721120
transform 1 0 62376 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_666
timestamp 1607721120
transform 1 0 62376 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__A1
timestamp 1607721120
transform 1 0 62192 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0689_
timestamp 1607721120
transform 1 0 62100 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_670
timestamp 1607721120
transform 1 0 62744 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_670
timestamp 1607721120
transform 1 0 62744 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__A
timestamp 1607721120
transform 1 0 62560 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1607721120
transform 1 0 62836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_672
timestamp 1607721120
transform 1 0 62928 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_674
timestamp 1607721120
transform 1 0 63112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1607721120
transform -1 0 63480 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1607721120
transform -1 0 63480 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_15
timestamp 1607721120
transform 1 0 2484 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1607721120
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1607721120
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _1015_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 2576 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1607721120
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_23
timestamp 1607721120
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__A
timestamp 1607721120
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__A1
timestamp 1607721120
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1607721120
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0677_
timestamp 1607721120
transform 1 0 4048 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_43
timestamp 1607721120
transform 1 0 5060 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_39
timestamp 1607721120
transform 1 0 4692 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_35
timestamp 1607721120
transform 1 0 4324 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__A2
timestamp 1607721120
transform 1 0 4876 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__A
timestamp 1607721120
transform 1 0 4508 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1016_
timestamp 1607721120
transform 1 0 5244 0 -1 3808
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_2_63
timestamp 1607721120
transform 1 0 6900 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_59
timestamp 1607721120
transform 1 0 6532 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__B1
timestamp 1607721120
transform 1 0 7084 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__A2
timestamp 1607721120
transform 1 0 6716 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  _1017_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 7268 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_88
timestamp 1607721120
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_84
timestamp 1607721120
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_80
timestamp 1607721120
transform 1 0 8464 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_76
timestamp 1607721120
transform 1 0 8096 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__B1
timestamp 1607721120
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__A2
timestamp 1607721120
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__A2
timestamp 1607721120
transform 1 0 8648 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__C1
timestamp 1607721120
transform 1 0 8280 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_111
timestamp 1607721120
transform 1 0 11316 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_93
timestamp 1607721120
transform 1 0 9660 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__A2
timestamp 1607721120
transform 1 0 11500 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__D
timestamp 1607721120
transform 1 0 10028 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1607721120
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1033_
timestamp 1607721120
transform 1 0 10212 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_135
timestamp 1607721120
transform 1 0 13524 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_115
timestamp 1607721120
transform 1 0 11684 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__A2_N
timestamp 1607721120
transform 1 0 11868 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__B1
timestamp 1607721120
transform 1 0 13708 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1014_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 12052 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_149
timestamp 1607721120
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_143
timestamp 1607721120
transform 1 0 14260 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_139
timestamp 1607721120
transform 1 0 13892 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__C
timestamp 1607721120
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__A2
timestamp 1607721120
transform 1 0 14076 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__C1
timestamp 1607721120
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1607721120
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _0998_
timestamp 1607721120
transform 1 0 15272 0 -1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_2_182
timestamp 1607721120
transform 1 0 17848 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_171
timestamp 1607721120
transform 1 0 16836 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_167
timestamp 1607721120
transform 1 0 16468 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__B
timestamp 1607721120
transform 1 0 17020 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__A2
timestamp 1607721120
transform 1 0 16652 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _0982_
timestamp 1607721120
transform 1 0 17204 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_2_194
timestamp 1607721120
transform 1 0 18952 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_190
timestamp 1607721120
transform 1 0 18584 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_186
timestamp 1607721120
transform 1 0 18216 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__B
timestamp 1607721120
transform 1 0 19044 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__C
timestamp 1607721120
transform 1 0 18400 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__A
timestamp 1607721120
transform 1 0 18032 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  _1004_
timestamp 1607721120
transform 1 0 19228 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_210
timestamp 1607721120
transform 1 0 20424 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_206
timestamp 1607721120
transform 1 0 20056 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__A
timestamp 1607721120
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__A
timestamp 1607721120
transform 1 0 20240 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1607721120
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1416_
timestamp 1607721120
transform 1 0 20884 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_2_238
timestamp 1607721120
transform 1 0 23000 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_234
timestamp 1607721120
transform 1 0 22632 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__C1
timestamp 1607721120
transform 1 0 23184 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__A2
timestamp 1607721120
transform 1 0 22816 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1032_
timestamp 1607721120
transform 1 0 23368 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_254
timestamp 1607721120
transform 1 0 24472 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__A1
timestamp 1607721120
transform 1 0 24656 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_258
timestamp 1607721120
transform 1 0 24840 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1032__A1
timestamp 1607721120
transform 1 0 25024 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_262
timestamp 1607721120
transform 1 0 25208 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0925_
timestamp 1607721120
transform 1 0 25300 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_267
timestamp 1607721120
transform 1 0 25668 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__B
timestamp 1607721120
transform 1 0 25852 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_271
timestamp 1607721120
transform 1 0 26036 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__C1
timestamp 1607721120
transform 1 0 26220 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_284
timestamp 1607721120
transform 1 0 27232 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_280
timestamp 1607721120
transform 1 0 26864 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__A
timestamp 1607721120
transform 1 0 27048 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__A2
timestamp 1607721120
transform 1 0 27416 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1607721120
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__a41o_4  _0996_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 27600 0 -1 3808
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_2  _0912_
timestamp 1607721120
transform 1 0 26496 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_309
timestamp 1607721120
transform 1 0 29532 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_305
timestamp 1607721120
transform 1 0 29164 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__A4
timestamp 1607721120
transform 1 0 29716 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__A2
timestamp 1607721120
transform 1 0 29348 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  _1042_
timestamp 1607721120
transform 1 0 29900 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_332
timestamp 1607721120
transform 1 0 31648 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_328
timestamp 1607721120
transform 1 0 31280 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_322
timestamp 1607721120
transform 1 0 30728 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__B1
timestamp 1607721120
transform 1 0 31464 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__A2
timestamp 1607721120
transform 1 0 31096 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__C
timestamp 1607721120
transform 1 0 31832 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1607721120
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _0926_
timestamp 1607721120
transform 1 0 32108 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_2_354
timestamp 1607721120
transform 1 0 33672 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_350
timestamp 1607721120
transform 1 0 33304 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_346
timestamp 1607721120
transform 1 0 32936 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__A
timestamp 1607721120
transform 1 0 33120 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__C
timestamp 1607721120
transform 1 0 33488 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _0914_
timestamp 1607721120
transform 1 0 33764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_386
timestamp 1607721120
transform 1 0 36616 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_382
timestamp 1607721120
transform 1 0 36248 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_371
timestamp 1607721120
transform 1 0 35236 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_367
timestamp 1607721120
transform 1 0 34868 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__B1
timestamp 1607721120
transform 1 0 35052 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__A
timestamp 1607721120
transform 1 0 35420 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__B
timestamp 1607721120
transform 1 0 36800 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__A
timestamp 1607721120
transform 1 0 36432 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0911_
timestamp 1607721120
transform 1 0 35604 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_2_402
timestamp 1607721120
transform 1 0 38088 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_398
timestamp 1607721120
transform 1 0 37720 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_394
timestamp 1607721120
transform 1 0 37352 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_390
timestamp 1607721120
transform 1 0 36984 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1199__B
timestamp 1607721120
transform 1 0 38456 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1158__A
timestamp 1607721120
transform 1 0 37904 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__C
timestamp 1607721120
transform 1 0 37168 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1607721120
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1197_
timestamp 1607721120
transform 1 0 38640 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_2_419
timestamp 1607721120
transform 1 0 39652 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_415
timestamp 1607721120
transform 1 0 39284 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__C
timestamp 1607721120
transform 1 0 39836 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1193__B
timestamp 1607721120
transform 1 0 39468 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1200_
timestamp 1607721120
transform 1 0 40020 0 -1 3808
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_2_453
timestamp 1607721120
transform 1 0 42780 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_449
timestamp 1607721120
transform 1 0 42412 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_441
timestamp 1607721120
transform 1 0 41676 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_437
timestamp 1607721120
transform 1 0 41308 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__A2
timestamp 1607721120
transform 1 0 42596 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__B1
timestamp 1607721120
transform 1 0 41860 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__A1
timestamp 1607721120
transform 1 0 41492 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__A
timestamp 1607721120
transform 1 0 42964 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0750_
timestamp 1607721120
transform 1 0 42044 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_476
timestamp 1607721120
transform 1 0 44896 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_472
timestamp 1607721120
transform 1 0 44528 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_459
timestamp 1607721120
transform 1 0 43332 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_457
timestamp 1607721120
transform 1 0 43148 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1196__A2
timestamp 1607721120
transform 1 0 43516 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1196__A1
timestamp 1607721120
transform 1 0 45080 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__C
timestamp 1607721120
transform 1 0 44712 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1607721120
transform 1 0 43240 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0686_
timestamp 1607721120
transform 1 0 43700 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_499
timestamp 1607721120
transform 1 0 47012 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1189__B1_N
timestamp 1607721120
transform 1 0 47196 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1388_
timestamp 1607721120
transform 1 0 45264 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_2_503
timestamp 1607721120
transform 1 0 47380 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__A2
timestamp 1607721120
transform 1 0 47564 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1003_
timestamp 1607721120
transform 1 0 47748 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_511
timestamp 1607721120
transform 1 0 48116 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_515
timestamp 1607721120
transform 1 0 48484 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1003__A
timestamp 1607721120
transform 1 0 48300 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__D
timestamp 1607721120
transform 1 0 48668 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1607721120
transform 1 0 48852 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0744_
timestamp 1607721120
transform 1 0 48944 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_524
timestamp 1607721120
transform 1 0 49312 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_545
timestamp 1607721120
transform 1 0 51244 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_528
timestamp 1607721120
transform 1 0 49680 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__D
timestamp 1607721120
transform 1 0 51428 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__B
timestamp 1607721120
transform 1 0 49864 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__A
timestamp 1607721120
transform 1 0 49496 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__nor3_4  _0691_
timestamp 1607721120
transform 1 0 50048 0 -1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  FILLER_2_570
timestamp 1607721120
transform 1 0 53544 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_566
timestamp 1607721120
transform 1 0 53176 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_562
timestamp 1607721120
transform 1 0 52808 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_549
timestamp 1607721120
transform 1 0 51612 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__B
timestamp 1607721120
transform 1 0 53360 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__A
timestamp 1607721120
transform 1 0 51796 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__B
timestamp 1607721120
transform 1 0 52992 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _0707_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 51980 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_581
timestamp 1607721120
transform 1 0 54556 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_579
timestamp 1607721120
transform 1 0 54372 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_575
timestamp 1607721120
transform 1 0 54004 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0744__A
timestamp 1607721120
transform 1 0 54740 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__C
timestamp 1607721120
transform 1 0 54188 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__A
timestamp 1607721120
transform 1 0 53820 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1607721120
transform 1 0 54464 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _1182_
timestamp 1607721120
transform 1 0 54924 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_613
timestamp 1607721120
transform 1 0 57500 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_609
timestamp 1607721120
transform 1 0 57132 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_600
timestamp 1607721120
transform 1 0 56304 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_594
timestamp 1607721120
transform 1 0 55752 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1154__A
timestamp 1607721120
transform 1 0 57316 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1152__A
timestamp 1607721120
transform 1 0 56120 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1165_
timestamp 1607721120
transform 1 0 56488 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_2_637
timestamp 1607721120
transform 1 0 59708 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_633
timestamp 1607721120
transform 1 0 59340 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_620
timestamp 1607721120
transform 1 0 58144 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_617
timestamp 1607721120
transform 1 0 57868 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__A2
timestamp 1607721120
transform 1 0 57960 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1166__A2
timestamp 1607721120
transform 1 0 58328 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1172__B
timestamp 1607721120
transform 1 0 59892 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1166__B1
timestamp 1607721120
transform 1 0 59524 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _1171_
timestamp 1607721120
transform 1 0 58512 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_2_658
timestamp 1607721120
transform 1 0 61640 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_654
timestamp 1607721120
transform 1 0 61272 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_649
timestamp 1607721120
transform 1 0 60812 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__C
timestamp 1607721120
transform 1 0 61456 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__B
timestamp 1607721120
transform 1 0 61088 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1607721120
transform 1 0 60076 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1172_
timestamp 1607721120
transform 1 0 60168 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_2_674
timestamp 1607721120
transform 1 0 63112 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_670
timestamp 1607721120
transform 1 0 62744 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1607721120
transform -1 0 63480 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1607721120
transform 1 0 1380 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1607721120
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_12
timestamp 1607721120
transform 1 0 2208 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_9
timestamp 1607721120
transform 1 0 1932 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__A
timestamp 1607721120
transform 1 0 2024 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_20
timestamp 1607721120
transform 1 0 2944 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_16
timestamp 1607721120
transform 1 0 2576 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__B
timestamp 1607721120
transform 1 0 2392 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__A
timestamp 1607721120
transform 1 0 2760 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__D
timestamp 1607721120
transform 1 0 3128 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_37
timestamp 1607721120
transform 1 0 4508 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_33
timestamp 1607721120
transform 1 0 4140 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__B1
timestamp 1607721120
transform 1 0 4692 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__B
timestamp 1607721120
transform 1 0 4324 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1024_
timestamp 1607721120
transform 1 0 4876 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _0678_
timestamp 1607721120
transform 1 0 3312 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_62
timestamp 1607721120
transform 1 0 6808 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1607721120
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_53
timestamp 1607721120
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__A2
timestamp 1607721120
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__A1
timestamp 1607721120
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__A1
timestamp 1607721120
transform 1 0 7176 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1607721120
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _0986_
timestamp 1607721120
transform 1 0 7360 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_89
timestamp 1607721120
transform 1 0 9292 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_85
timestamp 1607721120
transform 1 0 8924 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_81
timestamp 1607721120
transform 1 0 8556 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_77
timestamp 1607721120
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__C
timestamp 1607721120
transform 1 0 9108 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__D
timestamp 1607721120
transform 1 0 9476 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__B2
timestamp 1607721120
transform 1 0 8740 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__B1
timestamp 1607721120
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_114
timestamp 1607721120
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_106
timestamp 1607721120
transform 1 0 10856 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_102
timestamp 1607721120
transform 1 0 10488 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__C
timestamp 1607721120
transform 1 0 11040 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__B
timestamp 1607721120
transform 1 0 10672 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0985_
timestamp 1607721120
transform 1 0 11224 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _0983_
timestamp 1607721120
transform 1 0 9660 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_136
timestamp 1607721120
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_132
timestamp 1607721120
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_118
timestamp 1607721120
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__B
timestamp 1607721120
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__B
timestamp 1607721120
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__A
timestamp 1607721120
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1607721120
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0984_
timestamp 1607721120
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_158
timestamp 1607721120
transform 1 0 15640 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_154
timestamp 1607721120
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_140
timestamp 1607721120
transform 1 0 13984 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1287__C
timestamp 1607721120
transform 1 0 15456 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__A
timestamp 1607721120
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__nor3_4  _1287_
timestamp 1607721120
transform 1 0 14076 0 1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_3_182
timestamp 1607721120
transform 1 0 17848 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_178
timestamp 1607721120
transform 1 0 17480 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_174
timestamp 1607721120
transform 1 0 17112 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_162
timestamp 1607721120
transform 1 0 16008 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__B1
timestamp 1607721120
transform 1 0 16100 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__A2
timestamp 1607721120
transform 1 0 17664 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__A1
timestamp 1607721120
transform 1 0 17296 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0987_
timestamp 1607721120
transform 1 0 16284 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_201
timestamp 1607721120
transform 1 0 19596 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_197
timestamp 1607721120
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_184
timestamp 1607721120
transform 1 0 18032 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__C
timestamp 1607721120
transform 1 0 19780 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1006__B
timestamp 1607721120
transform 1 0 18400 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1006__A
timestamp 1607721120
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1607721120
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1010_
timestamp 1607721120
transform 1 0 19964 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _1006_
timestamp 1607721120
transform 1 0 18584 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1607721120
transform 1 0 21804 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_221
timestamp 1607721120
transform 1 0 21436 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_217
timestamp 1607721120
transform 1 0 21068 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1063__B
timestamp 1607721120
transform 1 0 21988 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__A1
timestamp 1607721120
transform 1 0 21620 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__A
timestamp 1607721120
transform 1 0 21252 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_236
timestamp 1607721120
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1075_
timestamp 1607721120
transform 1 0 22172 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_3_240
timestamp 1607721120
transform 1 0 23184 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1063__A
timestamp 1607721120
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__A
timestamp 1607721120
transform 1 0 23000 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1607721120
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_249
timestamp 1607721120
transform 1 0 24012 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_245
timestamp 1607721120
transform 1 0 23644 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__A
timestamp 1607721120
transform 1 0 24196 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__A
timestamp 1607721120
transform 1 0 23828 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_267
timestamp 1607721120
transform 1 0 25668 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_263
timestamp 1607721120
transform 1 0 25300 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_253
timestamp 1607721120
transform 1 0 24380 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__B1
timestamp 1607721120
transform 1 0 25852 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1345__B
timestamp 1607721120
transform 1 0 25484 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1345_
timestamp 1607721120
transform 1 0 24656 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _1074_
timestamp 1607721120
transform 1 0 26036 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_284
timestamp 1607721120
transform 1 0 27232 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_280
timestamp 1607721120
transform 1 0 26864 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__A1
timestamp 1607721120
transform 1 0 27048 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__A2
timestamp 1607721120
transform 1 0 27416 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1043_
timestamp 1607721120
transform 1 0 27600 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_301
timestamp 1607721120
transform 1 0 28796 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_297
timestamp 1607721120
transform 1 0 28428 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__A
timestamp 1607721120
transform 1 0 28980 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__A4
timestamp 1607721120
transform 1 0 28612 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_312
timestamp 1607721120
transform 1 0 29808 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_306
timestamp 1607721120
transform 1 0 29256 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__A
timestamp 1607721120
transform 1 0 29624 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1607721120
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__C
timestamp 1607721120
transform 1 0 29992 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0696_
timestamp 1607721120
transform 1 0 30176 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_3_339
timestamp 1607721120
transform 1 0 32292 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_335
timestamp 1607721120
transform 1 0 31924 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_327
timestamp 1607721120
transform 1 0 31188 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_323
timestamp 1607721120
transform 1 0 30820 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__B1
timestamp 1607721120
transform 1 0 32476 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1040__B
timestamp 1607721120
transform 1 0 31372 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__A
timestamp 1607721120
transform 1 0 32108 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__A
timestamp 1607721120
transform 1 0 31004 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0995_
timestamp 1607721120
transform 1 0 31556 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_346
timestamp 1607721120
transform 1 0 32936 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0700_
timestamp 1607721120
transform 1 0 32660 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_350
timestamp 1607721120
transform 1 0 33304 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__A
timestamp 1607721120
transform 1 0 33488 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__A
timestamp 1607721120
transform 1 0 33120 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0994_
timestamp 1607721120
transform 1 0 33672 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_358
timestamp 1607721120
transform 1 0 34040 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__A
timestamp 1607721120
transform 1 0 34224 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_362
timestamp 1607721120
transform 1 0 34408 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1160__A1
timestamp 1607721120
transform 1 0 34592 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1607721120
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__a41oi_4  _1157_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 34868 0 1 3808
box -38 -48 2062 592
use sky130_fd_sc_hd__fill_2  FILLER_3_393
timestamp 1607721120
transform 1 0 37260 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_389
timestamp 1607721120
transform 1 0 36892 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1160__A2
timestamp 1607721120
transform 1 0 37444 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__A3
timestamp 1607721120
transform 1 0 37076 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1005_
timestamp 1607721120
transform 1 0 37628 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1607721120
transform 1 0 38364 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_401
timestamp 1607721120
transform 1 0 37996 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__A
timestamp 1607721120
transform 1 0 38548 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__A
timestamp 1607721120
transform 1 0 38180 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_409
timestamp 1607721120
transform 1 0 38732 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1163_
timestamp 1607721120
transform 1 0 38824 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_423
timestamp 1607721120
transform 1 0 40020 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_419
timestamp 1607721120
transform 1 0 39652 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__A2
timestamp 1607721120
transform 1 0 40204 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__C1
timestamp 1607721120
transform 1 0 39836 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1607721120
transform 1 0 40388 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1198_
timestamp 1607721120
transform 1 0 40480 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_453
timestamp 1607721120
transform 1 0 42780 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_449
timestamp 1607721120
transform 1 0 42412 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_441
timestamp 1607721120
transform 1 0 41676 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_437
timestamp 1607721120
transform 1 0 41308 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__A1
timestamp 1607721120
transform 1 0 41860 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__A
timestamp 1607721120
transform 1 0 42596 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1198__A
timestamp 1607721120
transform 1 0 41492 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1144_
timestamp 1607721120
transform 1 0 42044 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_464
timestamp 1607721120
transform 1 0 43792 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_460
timestamp 1607721120
transform 1 0 43424 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_457
timestamp 1607721120
transform 1 0 43148 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1196__B1
timestamp 1607721120
transform 1 0 43240 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__B1
timestamp 1607721120
transform 1 0 43608 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1002__A
timestamp 1607721120
transform 1 0 43976 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1190_
timestamp 1607721120
transform 1 0 44160 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_502
timestamp 1607721120
transform 1 0 47288 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_484
timestamp 1607721120
transform 1 0 45632 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_480
timestamp 1607721120
transform 1 0 45264 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__A2
timestamp 1607721120
transform 1 0 45816 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__A1
timestamp 1607721120
transform 1 0 45448 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1607721120
transform 1 0 46000 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_4  _1189_
timestamp 1607721120
transform 1 0 46092 0 1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_3_522
timestamp 1607721120
transform 1 0 49128 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_506
timestamp 1607721120
transform 1 0 47656 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1116__A
timestamp 1607721120
transform 1 0 49312 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1189__A2
timestamp 1607721120
transform 1 0 47840 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1189__A1
timestamp 1607721120
transform 1 0 47472 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1191_
timestamp 1607721120
transform 1 0 48024 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_545
timestamp 1607721120
transform 1 0 51244 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_541
timestamp 1607721120
transform 1 0 50876 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_537
timestamp 1607721120
transform 1 0 50508 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_526
timestamp 1607721120
transform 1 0 49496 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__C
timestamp 1607721120
transform 1 0 51428 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__B
timestamp 1607721120
transform 1 0 51060 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0687__B
timestamp 1607721120
transform 1 0 49680 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0687__A
timestamp 1607721120
transform 1 0 50692 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _0687_
timestamp 1607721120
transform 1 0 49864 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_3_561
timestamp 1607721120
transform 1 0 52716 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_557
timestamp 1607721120
transform 1 0 52348 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__B
timestamp 1607721120
transform 1 0 52900 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__C
timestamp 1607721120
transform 1 0 52532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1607721120
transform 1 0 51612 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1180_
timestamp 1607721120
transform 1 0 51704 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _1177_
timestamp 1607721120
transform 1 0 53084 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_591
timestamp 1607721120
transform 1 0 55476 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_578
timestamp 1607721120
transform 1 0 54280 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_574
timestamp 1607721120
transform 1 0 53912 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1154__D
timestamp 1607721120
transform 1 0 55660 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__A
timestamp 1607721120
transform 1 0 54464 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__A
timestamp 1607721120
transform 1 0 54096 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _1154_
timestamp 1607721120
transform 1 0 54648 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_599
timestamp 1607721120
transform 1 0 56212 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_595
timestamp 1607721120
transform 1 0 55844 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__B
timestamp 1607721120
transform 1 0 56396 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1390__D
timestamp 1607721120
transform 1 0 56028 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_607
timestamp 1607721120
transform 1 0 56948 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_603
timestamp 1607721120
transform 1 0 56580 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__B
timestamp 1607721120
transform 1 0 57040 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_611
timestamp 1607721120
transform 1 0 57316 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1607721120
transform 1 0 57224 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1175_
timestamp 1607721120
transform 1 0 57408 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_3_623
timestamp 1607721120
transform 1 0 58420 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_619
timestamp 1607721120
transform 1 0 58052 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1166__A1
timestamp 1607721120
transform 1 0 58604 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__A
timestamp 1607721120
transform 1 0 58236 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1391_
timestamp 1607721120
transform 1 0 58788 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_3_662
timestamp 1607721120
transform 1 0 62008 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_658
timestamp 1607721120
transform 1 0 61640 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_653
timestamp 1607721120
transform 1 0 61180 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_650
timestamp 1607721120
transform 1 0 60904 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_646
timestamp 1607721120
transform 1 0 60536 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__A2
timestamp 1607721120
transform 1 0 61824 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__A1
timestamp 1607721120
transform 1 0 60996 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0713_
timestamp 1607721120
transform 1 0 61272 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_672
timestamp 1607721120
transform 1 0 62928 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_670
timestamp 1607721120
transform 1 0 62744 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_666
timestamp 1607721120
transform 1 0 62376 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__B1
timestamp 1607721120
transform 1 0 62192 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1607721120
transform 1 0 62836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1607721120
transform -1 0 63480 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_15
timestamp 1607721120
transform 1 0 2484 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1607721120
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1607721120
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1029_
timestamp 1607721120
transform 1 0 2576 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_4_44
timestamp 1607721120
transform 1 0 5152 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_28
timestamp 1607721120
transform 1 0 3680 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_23
timestamp 1607721120
transform 1 0 3220 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__C
timestamp 1607721120
transform 1 0 3496 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1607721120
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1030_
timestamp 1607721120
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_52
timestamp 1607721120
transform 1 0 5888 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_48
timestamp 1607721120
transform 1 0 5520 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__B1
timestamp 1607721120
transform 1 0 5704 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__A
timestamp 1607721120
transform 1 0 6164 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__A1
timestamp 1607721120
transform 1 0 5336 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _1028_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 6348 0 -1 4896
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_4_86
timestamp 1607721120
transform 1 0 9016 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1607721120
transform 1 0 8648 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_75
timestamp 1607721120
transform 1 0 8004 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_71
timestamp 1607721120
transform 1 0 7636 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__D
timestamp 1607721120
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__A
timestamp 1607721120
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__A2
timestamp 1607721120
transform 1 0 8188 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1018__A
timestamp 1607721120
transform 1 0 7820 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1027_
timestamp 1607721120
transform 1 0 8372 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_112
timestamp 1607721120
transform 1 0 11408 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_106
timestamp 1607721120
transform 1 0 10856 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_93
timestamp 1607721120
transform 1 0 9660 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__A
timestamp 1607721120
transform 1 0 11224 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1276__B
timestamp 1607721120
transform 1 0 9844 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1607721120
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _1026_
timestamp 1607721120
transform 1 0 10028 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1021_
timestamp 1607721120
transform 1 0 11592 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_4_125
timestamp 1607721120
transform 1 0 12604 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_121
timestamp 1607721120
transform 1 0 12236 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__B
timestamp 1607721120
transform 1 0 12788 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__D
timestamp 1607721120
transform 1 0 12420 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  _1019_
timestamp 1607721120
transform 1 0 12972 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1607721120
transform 1 0 13800 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__B
timestamp 1607721120
transform 1 0 13984 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_142
timestamp 1607721120
transform 1 0 14168 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__D
timestamp 1607721120
transform 1 0 14536 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_148
timestamp 1607721120
transform 1 0 14720 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1287__B
timestamp 1607721120
transform 1 0 14904 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_152
timestamp 1607721120
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1607721120
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0920_
timestamp 1607721120
transform 1 0 15272 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_158
timestamp 1607721120
transform 1 0 15640 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_180
timestamp 1607721120
transform 1 0 17664 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_166
timestamp 1607721120
transform 1 0 16376 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_162
timestamp 1607721120
transform 1 0 16008 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1059__C
timestamp 1607721120
transform 1 0 17848 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__A2
timestamp 1607721120
transform 1 0 16192 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__C1
timestamp 1607721120
transform 1 0 15824 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_4  _0989_
timestamp 1607721120
transform 1 0 16468 0 -1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  FILLER_4_205
timestamp 1607721120
transform 1 0 19964 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_201
timestamp 1607721120
transform 1 0 19596 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1607721120
transform 1 0 19228 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_184
timestamp 1607721120
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__B
timestamp 1607721120
transform 1 0 19780 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1091__B1_N
timestamp 1607721120
transform 1 0 19412 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__A
timestamp 1607721120
transform 1 0 18216 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1096_
timestamp 1607721120
transform 1 0 18400 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_228
timestamp 1607721120
transform 1 0 22080 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_224
timestamp 1607721120
transform 1 0 21712 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_210
timestamp 1607721120
transform 1 0 20424 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__A2
timestamp 1607721120
transform 1 0 20240 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__B
timestamp 1607721120
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1607721120
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _1011_
timestamp 1607721120
transform 1 0 20884 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_251
timestamp 1607721120
transform 1 0 24196 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_243
timestamp 1607721120
transform 1 0 23460 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_239
timestamp 1607721120
transform 1 0 23092 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_231
timestamp 1607721120
transform 1 0 22356 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__B1
timestamp 1607721120
transform 1 0 23644 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__A
timestamp 1607721120
transform 1 0 23276 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__B
timestamp 1607721120
transform 1 0 22172 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1063_
timestamp 1607721120
transform 1 0 22448 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0927_
timestamp 1607721120
transform 1 0 23828 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_255
timestamp 1607721120
transform 1 0 24564 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__B
timestamp 1607721120
transform 1 0 24380 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_259
timestamp 1607721120
transform 1 0 24932 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__C
timestamp 1607721120
transform 1 0 24748 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__A
timestamp 1607721120
transform 1 0 25116 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0991_
timestamp 1607721120
transform 1 0 25300 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_267
timestamp 1607721120
transform 1 0 25668 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__A
timestamp 1607721120
transform 1 0 25852 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_271
timestamp 1607721120
transform 1 0 26036 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__C
timestamp 1607721120
transform 1 0 26220 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1607721120
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__a41oi_4  _0990_
timestamp 1607721120
transform 1 0 26496 0 -1 4896
box -38 -48 2062 592
use sky130_fd_sc_hd__fill_2  FILLER_4_319
timestamp 1607721120
transform 1 0 30452 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_308
timestamp 1607721120
transform 1 0 29440 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_302
timestamp 1607721120
transform 1 0 28888 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_298
timestamp 1607721120
transform 1 0 28520 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__A2
timestamp 1607721120
transform 1 0 29256 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__A3
timestamp 1607721120
transform 1 0 28704 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0931_
timestamp 1607721120
transform 1 0 29624 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_323
timestamp 1607721120
transform 1 0 30820 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__B
timestamp 1607721120
transform 1 0 30636 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_327
timestamp 1607721120
transform 1 0 31188 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__B
timestamp 1607721120
transform 1 0 31004 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_331
timestamp 1607721120
transform 1 0 31556 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__B1
timestamp 1607721120
transform 1 0 31372 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_335
timestamp 1607721120
transform 1 0 31924 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__B1
timestamp 1607721120
transform 1 0 31740 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_337
timestamp 1607721120
transform 1 0 32108 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1607721120
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_341
timestamp 1607721120
transform 1 0 32476 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__A1
timestamp 1607721120
transform 1 0 32292 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_355
timestamp 1607721120
transform 1 0 33764 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_350
timestamp 1607721120
transform 1 0 33304 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__A
timestamp 1607721120
transform 1 0 32752 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1160__B1
timestamp 1607721120
transform 1 0 33580 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1160__A4
timestamp 1607721120
transform 1 0 33948 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__a41o_4  _1160_
timestamp 1607721120
transform 1 0 34132 0 -1 4896
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_2  _1020_
timestamp 1607721120
transform 1 0 32936 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_388
timestamp 1607721120
transform 1 0 36800 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_380
timestamp 1607721120
transform 1 0 36064 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_376
timestamp 1607721120
transform 1 0 35696 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__A1
timestamp 1607721120
transform 1 0 36248 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1160__A3
timestamp 1607721120
transform 1 0 35880 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0958_
timestamp 1607721120
transform 1 0 36432 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_392
timestamp 1607721120
transform 1 0 37168 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__A2
timestamp 1607721120
transform 1 0 36984 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_396
timestamp 1607721120
transform 1 0 37536 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__A4
timestamp 1607721120
transform 1 0 37352 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1607721120
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_398
timestamp 1607721120
transform 1 0 37720 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0981_
timestamp 1607721120
transform 1 0 37904 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_404
timestamp 1607721120
transform 1 0 38272 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_410
timestamp 1607721120
transform 1 0 38824 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__A
timestamp 1607721120
transform 1 0 38640 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_432
timestamp 1607721120
transform 1 0 40848 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_428
timestamp 1607721120
transform 1 0 40480 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__B
timestamp 1607721120
transform 1 0 39008 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1198__B
timestamp 1607721120
transform 1 0 40664 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1164_
timestamp 1607721120
transform 1 0 39192 0 -1 4896
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_4_452
timestamp 1607721120
transform 1 0 42688 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_448
timestamp 1607721120
transform 1 0 42320 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__B
timestamp 1607721120
transform 1 0 43056 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__B1
timestamp 1607721120
transform 1 0 41032 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__A2
timestamp 1607721120
transform 1 0 42504 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1159_
timestamp 1607721120
transform 1 0 41216 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_476
timestamp 1607721120
transform 1 0 44896 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_470
timestamp 1607721120
transform 1 0 44344 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_463
timestamp 1607721120
transform 1 0 43700 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_459
timestamp 1607721120
transform 1 0 43332 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__A
timestamp 1607721120
transform 1 0 43516 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__B1
timestamp 1607721120
transform 1 0 44712 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1607721120
transform 1 0 43240 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1192_
timestamp 1607721120
transform 1 0 45080 0 -1 4896
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _1002_
timestamp 1607721120
transform 1 0 43976 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_496
timestamp 1607721120
transform 1 0 46736 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_492
timestamp 1607721120
transform 1 0 46368 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__A1
timestamp 1607721120
transform 1 0 46920 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__C1
timestamp 1607721120
transform 1 0 46552 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _1155_
timestamp 1607721120
transform 1 0 47104 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_524
timestamp 1607721120
transform 1 0 49312 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_520
timestamp 1607721120
transform 1 0 48944 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_515
timestamp 1607721120
transform 1 0 48484 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_509
timestamp 1607721120
transform 1 0 47932 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__A2
timestamp 1607721120
transform 1 0 48300 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__B1
timestamp 1607721120
transform 1 0 48668 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__A1
timestamp 1607721120
transform 1 0 49128 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1607721120
transform 1 0 48852 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_544
timestamp 1607721120
transform 1 0 51152 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_540
timestamp 1607721120
transform 1 0 50784 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_528
timestamp 1607721120
transform 1 0 49680 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__B
timestamp 1607721120
transform 1 0 51336 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1116__C
timestamp 1607721120
transform 1 0 49772 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1116__B
timestamp 1607721120
transform 1 0 50968 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1150_
timestamp 1607721120
transform 1 0 51520 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _1116_
timestamp 1607721120
transform 1 0 49956 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_561
timestamp 1607721120
transform 1 0 52716 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_557
timestamp 1607721120
transform 1 0 52348 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__A1
timestamp 1607721120
transform 1 0 52900 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__A
timestamp 1607721120
transform 1 0 52532 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1178_
timestamp 1607721120
transform 1 0 53084 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_4_572
timestamp 1607721120
transform 1 0 53728 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__A
timestamp 1607721120
transform 1 0 53912 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_576
timestamp 1607721120
transform 1 0 54096 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__B1
timestamp 1607721120
transform 1 0 54280 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1607721120
transform 1 0 54464 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_585
timestamp 1607721120
transform 1 0 54924 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1035_
timestamp 1607721120
transform 1 0 54556 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_589
timestamp 1607721120
transform 1 0 55292 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1181__A2
timestamp 1607721120
transform 1 0 55384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_592
timestamp 1607721120
transform 1 0 55568 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_613
timestamp 1607721120
transform 1 0 57500 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1390_
timestamp 1607721120
transform 1 0 55752 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_4_637
timestamp 1607721120
transform 1 0 59708 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_633
timestamp 1607721120
transform 1 0 59340 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_620
timestamp 1607721120
transform 1 0 58144 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_617
timestamp 1607721120
transform 1 0 57868 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1173__B1
timestamp 1607721120
transform 1 0 59892 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__A2
timestamp 1607721120
transform 1 0 57960 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1391__D
timestamp 1607721120
transform 1 0 59524 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1166_
timestamp 1607721120
transform 1 0 58236 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_658
timestamp 1607721120
transform 1 0 61640 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_654
timestamp 1607721120
transform 1 0 61272 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0713__A
timestamp 1607721120
transform 1 0 61456 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1607721120
transform 1 0 60076 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1167_
timestamp 1607721120
transform 1 0 60168 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_674
timestamp 1607721120
transform 1 0 63112 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_670
timestamp 1607721120
transform 1 0 62744 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1607721120
transform -1 0 63480 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_18
timestamp 1607721120
transform 1 0 2760 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_14
timestamp 1607721120
transform 1 0 2392 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_11
timestamp 1607721120
transform 1 0 2116 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 1380 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__B
timestamp 1607721120
transform 1 0 2208 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__A
timestamp 1607721120
transform 1 0 2576 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1607721120
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1413_
timestamp 1607721120
transform 1 0 2944 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_5_43
timestamp 1607721120
transform 1 0 5060 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_39
timestamp 1607721120
transform 1 0 4692 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__A2
timestamp 1607721120
transform 1 0 5244 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__B1
timestamp 1607721120
transform 1 0 4876 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1607721120
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_53
timestamp 1607721120
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_47
timestamp 1607721120
transform 1 0 5428 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__C
timestamp 1607721120
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0950__A
timestamp 1607721120
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1607721120
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1018_
timestamp 1607721120
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0881_
timestamp 1607721120
transform 1 0 5612 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_75
timestamp 1607721120
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_71
timestamp 1607721120
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0949__B
timestamp 1607721120
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0949__A
timestamp 1607721120
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__a21bo_4  _1031_
timestamp 1607721120
transform 1 0 8372 0 1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_5_111
timestamp 1607721120
transform 1 0 11316 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_107
timestamp 1607721120
transform 1 0 10948 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_96
timestamp 1607721120
transform 1 0 9936 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_92
timestamp 1607721120
transform 1 0 9568 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1268__A
timestamp 1607721120
transform 1 0 11500 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1276__A
timestamp 1607721120
transform 1 0 10120 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__A1
timestamp 1607721120
transform 1 0 9752 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1282__A
timestamp 1607721120
transform 1 0 11132 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1282_
timestamp 1607721120
transform 1 0 10304 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_5_119
timestamp 1607721120
transform 1 0 12052 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_115
timestamp 1607721120
transform 1 0 11684 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1268__B
timestamp 1607721120
transform 1 0 11868 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1607721120
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1409_
timestamp 1607721120
transform 1 0 12420 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_5_146
timestamp 1607721120
transform 1 0 14536 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_142
timestamp 1607721120
transform 1 0 14168 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__B1
timestamp 1607721120
transform 1 0 14720 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1286__C
timestamp 1607721120
transform 1 0 14352 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1060_
timestamp 1607721120
transform 1 0 14904 0 1 4896
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_5_179
timestamp 1607721120
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_176
timestamp 1607721120
transform 1 0 17296 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_172
timestamp 1607721120
transform 1 0 16928 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_168
timestamp 1607721120
transform 1 0 16560 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_164
timestamp 1607721120
transform 1 0 16192 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1059__A
timestamp 1607721120
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__A2
timestamp 1607721120
transform 1 0 16744 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1059__B
timestamp 1607721120
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__B1
timestamp 1607721120
transform 1 0 16376 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_205
timestamp 1607721120
transform 1 0 19964 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_197
timestamp 1607721120
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_193
timestamp 1607721120
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__A
timestamp 1607721120
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1091__A1
timestamp 1607721120
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1607721120
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1059_
timestamp 1607721120
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0997_
timestamp 1607721120
transform 1 0 19596 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_228
timestamp 1607721120
transform 1 0 22080 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_224
timestamp 1607721120
transform 1 0 21712 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_209
timestamp 1607721120
transform 1 0 20332 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__C
timestamp 1607721120
transform 1 0 20700 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__A
timestamp 1607721120
transform 1 0 21896 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__A
timestamp 1607721120
transform 1 0 20148 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  _1062_
timestamp 1607721120
transform 1 0 20884 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__B1
timestamp 1607721120
transform 1 0 22264 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0904_
timestamp 1607721120
transform 1 0 22448 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_236
timestamp 1607721120
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__A
timestamp 1607721120
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_240
timestamp 1607721120
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1064__C
timestamp 1607721120
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1607721120
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1044_
timestamp 1607721120
transform 1 0 23644 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_249
timestamp 1607721120
transform 1 0 24012 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1044__A
timestamp 1607721120
transform 1 0 24196 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_253
timestamp 1607721120
transform 1 0 24380 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__A
timestamp 1607721120
transform 1 0 24564 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1408_
timestamp 1607721120
transform 1 0 24748 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_5_296
timestamp 1607721120
transform 1 0 28336 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_282
timestamp 1607721120
transform 1 0 27048 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_276
timestamp 1607721120
transform 1 0 26496 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__B
timestamp 1607721120
transform 1 0 26864 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1078_
timestamp 1607721120
transform 1 0 27232 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_301
timestamp 1607721120
transform 1 0 28796 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__A1
timestamp 1607721120
transform 1 0 28612 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__A3
timestamp 1607721120
transform 1 0 28980 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1607721120
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__a41o_4  _1056_
timestamp 1607721120
transform 1 0 29256 0 1 4896
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_5_339
timestamp 1607721120
transform 1 0 32292 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_335
timestamp 1607721120
transform 1 0 31924 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_327
timestamp 1607721120
transform 1 0 31188 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_323
timestamp 1607721120
transform 1 0 30820 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__A2
timestamp 1607721120
transform 1 0 32476 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__A
timestamp 1607721120
transform 1 0 32108 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__A4
timestamp 1607721120
transform 1 0 31372 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__A
timestamp 1607721120
transform 1 0 31004 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0993_
timestamp 1607721120
transform 1 0 31556 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_346
timestamp 1607721120
transform 1 0 32936 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0701_
timestamp 1607721120
transform 1 0 32660 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_350
timestamp 1607721120
transform 1 0 33304 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__A
timestamp 1607721120
transform 1 0 33488 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__A
timestamp 1607721120
transform 1 0 33120 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0965_
timestamp 1607721120
transform 1 0 33672 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_358
timestamp 1607721120
transform 1 0 34040 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__A
timestamp 1607721120
transform 1 0 34224 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_362
timestamp 1607721120
transform 1 0 34408 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__A
timestamp 1607721120
transform 1 0 34592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_388
timestamp 1607721120
transform 1 0 36800 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_377
timestamp 1607721120
transform 1 0 35788 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_373
timestamp 1607721120
transform 1 0 35420 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_367
timestamp 1607721120
transform 1 0 34868 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__A2
timestamp 1607721120
transform 1 0 35972 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__A3
timestamp 1607721120
transform 1 0 35604 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1607721120
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1153_
timestamp 1607721120
transform 1 0 36156 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0820_
timestamp 1607721120
transform 1 0 35052 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_396
timestamp 1607721120
transform 1 0 37536 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_392
timestamp 1607721120
transform 1 0 37168 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__A4
timestamp 1607721120
transform 1 0 37352 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__A
timestamp 1607721120
transform 1 0 36984 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_4  _1162_
timestamp 1607721120
transform 1 0 37812 0 1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_5_412
timestamp 1607721120
transform 1 0 39008 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__B1
timestamp 1607721120
transform 1 0 39192 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_420
timestamp 1607721120
transform 1 0 39744 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_416
timestamp 1607721120
transform 1 0 39376 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1393__D
timestamp 1607721120
transform 1 0 39560 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_424
timestamp 1607721120
transform 1 0 40112 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__A
timestamp 1607721120
transform 1 0 39928 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_428
timestamp 1607721120
transform 1 0 40480 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1607721120
transform 1 0 40388 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0936_
timestamp 1607721120
transform 1 0 40572 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_433
timestamp 1607721120
transform 1 0 40940 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_454
timestamp 1607721120
transform 1 0 42872 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_450
timestamp 1607721120
transform 1 0 42504 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_437
timestamp 1607721120
transform 1 0 41308 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__B
timestamp 1607721120
transform 1 0 41492 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__A
timestamp 1607721120
transform 1 0 41124 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__A
timestamp 1607721120
transform 1 0 43056 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__A
timestamp 1607721120
transform 1 0 42688 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  _1147_
timestamp 1607721120
transform 1 0 41676 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_467
timestamp 1607721120
transform 1 0 44068 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_463
timestamp 1607721120
transform 1 0 43700 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_458
timestamp 1607721120
transform 1 0 43240 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__B
timestamp 1607721120
transform 1 0 44252 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__A
timestamp 1607721120
transform 1 0 43884 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1195_
timestamp 1607721120
transform 1 0 44436 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0959_
timestamp 1607721120
transform 1 0 43332 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_489
timestamp 1607721120
transform 1 0 46092 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_484
timestamp 1607721120
transform 1 0 45632 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_480
timestamp 1607721120
transform 1 0 45264 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__B
timestamp 1607721120
transform 1 0 45816 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__A
timestamp 1607721120
transform 1 0 45448 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1156__B1
timestamp 1607721120
transform 1 0 46276 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1607721120
transform 1 0 46000 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1156_
timestamp 1607721120
transform 1 0 46460 0 1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  FILLER_5_514
timestamp 1607721120
transform 1 0 48392 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_510
timestamp 1607721120
transform 1 0 48024 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_506
timestamp 1607721120
transform 1 0 47656 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1156__A2
timestamp 1607721120
transform 1 0 48208 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1168__A
timestamp 1607721120
transform 1 0 47840 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _1186_
timestamp 1607721120
transform 1 0 48668 0 1 4896
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_5_547
timestamp 1607721120
transform 1 0 51428 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_543
timestamp 1607721120
transform 1 0 51060 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_539
timestamp 1607721120
transform 1 0 50692 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_535
timestamp 1607721120
transform 1 0 50324 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_531
timestamp 1607721120
transform 1 0 49956 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__B
timestamp 1607721120
transform 1 0 51244 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__A
timestamp 1607721120
transform 1 0 50876 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__A2
timestamp 1607721120
transform 1 0 50508 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__A1
timestamp 1607721120
transform 1 0 50140 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_554
timestamp 1607721120
transform 1 0 52072 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_550
timestamp 1607721120
transform 1 0 51704 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__D
timestamp 1607721120
transform 1 0 51888 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__B1
timestamp 1607721120
transform 1 0 52348 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1607721120
transform 1 0 51612 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1184_
timestamp 1607721120
transform 1 0 52532 0 1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_5_593
timestamp 1607721120
transform 1 0 55660 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_580
timestamp 1607721120
transform 1 0 54464 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_576
timestamp 1607721120
transform 1 0 54096 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_572
timestamp 1607721120
transform 1 0 53728 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__A2
timestamp 1607721120
transform 1 0 54280 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__B1
timestamp 1607721120
transform 1 0 53912 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1181_
timestamp 1607721120
transform 1 0 54556 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_606
timestamp 1607721120
transform 1 0 56856 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_601
timestamp 1607721120
transform 1 0 56396 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_597
timestamp 1607721120
transform 1 0 56028 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1151__D
timestamp 1607721120
transform 1 0 56212 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__C
timestamp 1607721120
transform 1 0 56672 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__B
timestamp 1607721120
transform 1 0 57040 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1151__B
timestamp 1607721120
transform 1 0 55844 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1607721120
transform 1 0 57224 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _1120_
timestamp 1607721120
transform 1 0 57316 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_624
timestamp 1607721120
transform 1 0 58512 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_620
timestamp 1607721120
transform 1 0 58144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__A
timestamp 1607721120
transform 1 0 58328 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__A
timestamp 1607721120
transform 1 0 58880 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1173_
timestamp 1607721120
transform 1 0 59064 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_5_658
timestamp 1607721120
transform 1 0 61640 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_654
timestamp 1607721120
transform 1 0 61272 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_650
timestamp 1607721120
transform 1 0 60904 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_646
timestamp 1607721120
transform 1 0 60536 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1392__CLK
timestamp 1607721120
transform 1 0 61456 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1173__A2_N
timestamp 1607721120
transform 1 0 61088 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1392__D
timestamp 1607721120
transform 1 0 60720 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_672
timestamp 1607721120
transform 1 0 62928 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_670
timestamp 1607721120
transform 1 0 62744 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1607721120
transform 1 0 62836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1607721120
transform -1 0 63480 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_11
timestamp 1607721120
transform 1 0 2116 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp 1607721120
transform 1 0 1380 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1607721120
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1607721120
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_22
timestamp 1607721120
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_18
timestamp 1607721120
transform 1 0 2760 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_15
timestamp 1607721120
transform 1 0 2484 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1421__CLK
timestamp 1607721120
transform 1 0 2576 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1413__CLK
timestamp 1607721120
transform 1 0 2944 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1409__CLK
timestamp 1607721120
transform 1 0 2392 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1274_
timestamp 1607721120
transform 1 0 2576 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1607721120
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_32
timestamp 1607721120
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_27
timestamp 1607721120
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_23
timestamp 1607721120
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0881__A
timestamp 1607721120
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1413__D
timestamp 1607721120
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1607721120
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_42
timestamp 1607721120
transform 1 0 4968 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1424__D
timestamp 1607721120
transform 1 0 5152 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1421_
timestamp 1607721120
transform 1 0 3220 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _0951_
timestamp 1607721120
transform 1 0 4232 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_53
timestamp 1607721120
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_50
timestamp 1607721120
transform 1 0 5704 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_46
timestamp 1607721120
transform 1 0 5336 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_50
timestamp 1607721120
transform 1 0 5704 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_46
timestamp 1607721120
transform 1 0 5336 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__B
timestamp 1607721120
transform 1 0 5888 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__B
timestamp 1607721120
transform 1 0 5796 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__A1
timestamp 1607721120
transform 1 0 5520 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1607721120
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_58
timestamp 1607721120
transform 1 0 6440 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__A
timestamp 1607721120
transform 1 0 6624 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__D
timestamp 1607721120
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__B
timestamp 1607721120
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1607721120
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0950_
timestamp 1607721120
transform 1 0 6072 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_66
timestamp 1607721120
transform 1 0 7176 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_62
timestamp 1607721120
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1018__B
timestamp 1607721120
transform 1 0 6992 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1013_
timestamp 1607721120
transform 1 0 6808 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _0949_
timestamp 1607721120
transform 1 0 7268 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_7_73
timestamp 1607721120
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_69
timestamp 1607721120
transform 1 0 7452 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_74
timestamp 1607721120
transform 1 0 7912 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__A
timestamp 1607721120
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1278__A
timestamp 1607721120
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_84
timestamp 1607721120
transform 1 0 8832 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_84
timestamp 1607721120
transform 1 0 8832 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_80
timestamp 1607721120
transform 1 0 8464 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__B1_N
timestamp 1607721120
transform 1 0 8648 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__B
timestamp 1607721120
transform 1 0 8280 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1272_
timestamp 1607721120
transform 1 0 8188 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_7_88
timestamp 1607721120
transform 1 0 9200 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1607721120
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_88
timestamp 1607721120
transform 1 0 9200 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__A2
timestamp 1607721120
transform 1 0 9292 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__B
timestamp 1607721120
transform 1 0 9384 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__A
timestamp 1607721120
transform 1 0 9016 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_99
timestamp 1607721120
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1607721120
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1280_
timestamp 1607721120
transform 1 0 9568 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1276_
timestamp 1607721120
transform 1 0 9660 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_7_103
timestamp 1607721120
transform 1 0 10580 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_104
timestamp 1607721120
transform 1 0 10672 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_100
timestamp 1607721120
transform 1 0 10304 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1282__B
timestamp 1607721120
transform 1 0 10488 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1385__D
timestamp 1607721120
transform 1 0 10764 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__A
timestamp 1607721120
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1270_
timestamp 1607721120
transform 1 0 10948 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_7_114
timestamp 1607721120
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_110
timestamp 1607721120
transform 1 0 11224 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1270__B
timestamp 1607721120
transform 1 0 11040 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1268_
timestamp 1607721120
transform 1 0 11500 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_7_123
timestamp 1607721120
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_118
timestamp 1607721120
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_124
timestamp 1607721120
transform 1 0 12512 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_120
timestamp 1607721120
transform 1 0 12144 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__A
timestamp 1607721120
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__A
timestamp 1607721120
transform 1 0 12328 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1270__A
timestamp 1607721120
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1607721120
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_136
timestamp 1607721120
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_132
timestamp 1607721120
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_128
timestamp 1607721120
transform 1 0 12880 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_128
timestamp 1607721120
transform 1 0 12880 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__A
timestamp 1607721120
transform 1 0 12696 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__C
timestamp 1607721120
transform 1 0 13064 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__B1
timestamp 1607721120
transform 1 0 13064 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__A2
timestamp 1607721120
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1409__D
timestamp 1607721120
transform 1 0 12696 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__nor3_4  _1286_
timestamp 1607721120
transform 1 0 13248 0 -1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_7_140
timestamp 1607721120
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_145
timestamp 1607721120
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1286__B
timestamp 1607721120
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__C1
timestamp 1607721120
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_158
timestamp 1607721120
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_154
timestamp 1607721120
transform 1 0 15272 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_154
timestamp 1607721120
transform 1 0 15272 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_149
timestamp 1607721120
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__B
timestamp 1607721120
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__A1
timestamp 1607721120
transform 1 0 15456 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1607721120
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1058_
timestamp 1607721120
transform 1 0 15364 0 -1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_4  _1055_
timestamp 1607721120
transform 1 0 14168 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_168
timestamp 1607721120
transform 1 0 16560 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__A2
timestamp 1607721120
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_179
timestamp 1607721120
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_175
timestamp 1607721120
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_174
timestamp 1607721120
transform 1 0 17112 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__A2
timestamp 1607721120
transform 1 0 16928 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__A1
timestamp 1607721120
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__A1
timestamp 1607721120
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__a21bo_4  _1091_
timestamp 1607721120
transform 1 0 17296 0 -1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__a21bo_4  _1086_
timestamp 1607721120
transform 1 0 16008 0 1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_6_193
timestamp 1607721120
transform 1 0 18860 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_189
timestamp 1607721120
transform 1 0 18492 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1091__A2
timestamp 1607721120
transform 1 0 18676 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1607721120
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_200
timestamp 1607721120
transform 1 0 19504 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_196
timestamp 1607721120
transform 1 0 19136 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1087__A2
timestamp 1607721120
transform 1 0 19044 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__A1
timestamp 1607721120
transform 1 0 19688 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1087__A1
timestamp 1607721120
transform 1 0 19320 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  _1095_
timestamp 1607721120
transform 1 0 19872 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _1092_
timestamp 1607721120
transform 1 0 19228 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_4  _1087_
timestamp 1607721120
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_213
timestamp 1607721120
transform 1 0 20700 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_215
timestamp 1607721120
transform 1 0 20884 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_210
timestamp 1607721120
transform 1 0 20424 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_206
timestamp 1607721120
transform 1 0 20056 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__A2
timestamp 1607721120
transform 1 0 20240 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__B
timestamp 1607721120
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1607721120
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_219
timestamp 1607721120
transform 1 0 21252 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1607721120
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1069__B
timestamp 1607721120
transform 1 0 21068 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1069__A
timestamp 1607721120
transform 1 0 21068 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1064_
timestamp 1607721120
transform 1 0 21344 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1049_
timestamp 1607721120
transform 1 0 21436 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_7_228
timestamp 1607721120
transform 1 0 22080 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_232
timestamp 1607721120
transform 1 0 22448 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_233
timestamp 1607721120
transform 1 0 22540 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_229
timestamp 1607721120
transform 1 0 22172 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1064__A
timestamp 1607721120
transform 1 0 22356 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__A
timestamp 1607721120
transform 1 0 22264 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_236
timestamp 1607721120
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1345__A
timestamp 1607721120
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1064__B
timestamp 1607721120
transform 1 0 22724 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__A
timestamp 1607721120
transform 1 0 22632 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1000_
timestamp 1607721120
transform 1 0 22908 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_245
timestamp 1607721120
transform 1 0 23644 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_240
timestamp 1607721120
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_246
timestamp 1607721120
transform 1 0 23736 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_241
timestamp 1607721120
transform 1 0 23276 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__A
timestamp 1607721120
transform 1 0 23552 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__B1
timestamp 1607721120
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__C
timestamp 1607721120
transform 1 0 23920 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1048__A
timestamp 1607721120
transform 1 0 23828 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1607721120
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_249
timestamp 1607721120
transform 1 0 24012 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _1068_
timestamp 1607721120
transform 1 0 24104 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_259
timestamp 1607721120
transform 1 0 24932 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1076__A
timestamp 1607721120
transform 1 0 24288 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1408__D
timestamp 1607721120
transform 1 0 25116 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_263
timestamp 1607721120
transform 1 0 25300 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__A2
timestamp 1607721120
transform 1 0 25484 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_266
timestamp 1607721120
transform 1 0 25576 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_267
timestamp 1607721120
transform 1 0 25668 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__A1
timestamp 1607721120
transform 1 0 25760 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_270
timestamp 1607721120
transform 1 0 25944 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_271
timestamp 1607721120
transform 1 0 26036 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__A1
timestamp 1607721120
transform 1 0 25852 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__D
timestamp 1607721120
transform 1 0 26220 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1070__B2
timestamp 1607721120
transform 1 0 26128 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1067_
timestamp 1607721120
transform 1 0 24472 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_4  _1066_
timestamp 1607721120
transform 1 0 26312 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_276
timestamp 1607721120
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1607721120
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _1047_
timestamp 1607721120
transform 1 0 26588 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_290
timestamp 1607721120
transform 1 0 27784 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_286
timestamp 1607721120
transform 1 0 27416 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_292
timestamp 1607721120
transform 1 0 27968 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_286
timestamp 1607721120
transform 1 0 27416 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__B
timestamp 1607721120
transform 1 0 27784 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__B1
timestamp 1607721120
transform 1 0 27968 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__A1
timestamp 1607721120
transform 1 0 27600 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0928_
timestamp 1607721120
transform 1 0 28152 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__a41oi_4  _1053_
timestamp 1607721120
transform 1 0 28244 0 -1 5984
box -38 -48 2062 592
use sky130_fd_sc_hd__fill_2  FILLER_7_301
timestamp 1607721120
transform 1 0 28796 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_297
timestamp 1607721120
transform 1 0 28428 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_317
timestamp 1607721120
transform 1 0 30268 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__B1
timestamp 1607721120
transform 1 0 28980 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__A
timestamp 1607721120
transform 1 0 28612 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__A3
timestamp 1607721120
transform 1 0 30452 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1607721120
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1406_
timestamp 1607721120
transform 1 0 29256 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_7_329
timestamp 1607721120
transform 1 0 31372 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_325
timestamp 1607721120
transform 1 0 31004 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_328
timestamp 1607721120
transform 1 0 31280 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_321
timestamp 1607721120
transform 1 0 30636 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__A2
timestamp 1607721120
transform 1 0 30820 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__A
timestamp 1607721120
transform 1 0 31188 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0924_
timestamp 1607721120
transform 1 0 31004 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_332
timestamp 1607721120
transform 1 0 31648 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__C
timestamp 1607721120
transform 1 0 31832 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__A
timestamp 1607721120
transform 1 0 31556 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__A4
timestamp 1607721120
transform 1 0 31464 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1607721120
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _1079_
timestamp 1607721120
transform 1 0 31740 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1054_
timestamp 1607721120
transform 1 0 32108 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_342
timestamp 1607721120
transform 1 0 32568 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_341
timestamp 1607721120
transform 1 0 32476 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_346
timestamp 1607721120
transform 1 0 32936 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_345
timestamp 1607721120
transform 1 0 32844 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__A1
timestamp 1607721120
transform 1 0 32660 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__A
timestamp 1607721120
transform 1 0 33028 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__A
timestamp 1607721120
transform 1 0 32752 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_350
timestamp 1607721120
transform 1 0 33304 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__B1
timestamp 1607721120
transform 1 0 33120 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__A
timestamp 1607721120
transform 1 0 33488 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0966_
timestamp 1607721120
transform 1 0 33212 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_353
timestamp 1607721120
transform 1 0 33580 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_362
timestamp 1607721120
transform 1 0 34408 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_358
timestamp 1607721120
transform 1 0 34040 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_357
timestamp 1607721120
transform 1 0 33948 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__A1
timestamp 1607721120
transform 1 0 33764 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__B1
timestamp 1607721120
transform 1 0 34592 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__A1
timestamp 1607721120
transform 1 0 34132 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1384__D
timestamp 1607721120
transform 1 0 34224 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0967_
timestamp 1607721120
transform 1 0 33672 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_4  _1109_
timestamp 1607721120
transform 1 0 34316 0 -1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_6_382
timestamp 1607721120
transform 1 0 36248 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_378
timestamp 1607721120
transform 1 0 35880 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__A
timestamp 1607721120
transform 1 0 36432 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1250__A
timestamp 1607721120
transform 1 0 36064 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1607721120
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__a41oi_4  _1106_
timestamp 1607721120
transform 1 0 34868 0 1 5984
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 1607721120
transform 1 0 36616 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_393
timestamp 1607721120
transform 1 0 37260 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_389
timestamp 1607721120
transform 1 0 36892 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_393
timestamp 1607721120
transform 1 0 37260 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_389
timestamp 1607721120
transform 1 0 36892 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__A1
timestamp 1607721120
transform 1 0 37444 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__B
timestamp 1607721120
transform 1 0 37076 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__A4
timestamp 1607721120
transform 1 0 37444 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__A3
timestamp 1607721120
transform 1 0 37076 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_402
timestamp 1607721120
transform 1 0 38088 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_397
timestamp 1607721120
transform 1 0 37628 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_402
timestamp 1607721120
transform 1 0 38088 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1607721120
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1097_
timestamp 1607721120
transform 1 0 37720 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0935_
timestamp 1607721120
transform 1 0 37720 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_406
timestamp 1607721120
transform 1 0 38456 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_410
timestamp 1607721120
transform 1 0 38824 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_406
timestamp 1607721120
transform 1 0 38456 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__A2
timestamp 1607721120
transform 1 0 38640 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__A2
timestamp 1607721120
transform 1 0 38272 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__B
timestamp 1607721120
transform 1 0 38640 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__A
timestamp 1607721120
transform 1 0 38272 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1099_
timestamp 1607721120
transform 1 0 38824 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_7_421
timestamp 1607721120
transform 1 0 39836 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_417
timestamp 1607721120
transform 1 0 39468 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__B1
timestamp 1607721120
transform 1 0 39100 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1141__B
timestamp 1607721120
transform 1 0 40204 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__A
timestamp 1607721120
transform 1 0 39652 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1607721120
transform 1 0 40388 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1393_
timestamp 1607721120
transform 1 0 39284 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_4  _1141_
timestamp 1607721120
transform 1 0 40480 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_7_439
timestamp 1607721120
transform 1 0 41492 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_435
timestamp 1607721120
transform 1 0 41124 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_438
timestamp 1607721120
transform 1 0 41400 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_434
timestamp 1607721120
transform 1 0 41032 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1148__C
timestamp 1607721120
transform 1 0 41216 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1148__B
timestamp 1607721120
transform 1 0 41584 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1148__A
timestamp 1607721120
transform 1 0 41676 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1141__A
timestamp 1607721120
transform 1 0 41308 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1146_
timestamp 1607721120
transform 1 0 41768 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_6_453
timestamp 1607721120
transform 1 0 42780 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_449
timestamp 1607721120
transform 1 0 42412 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__B1
timestamp 1607721120
transform 1 0 42964 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__B
timestamp 1607721120
transform 1 0 42596 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1149_
timestamp 1607721120
transform 1 0 41860 0 1 5984
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_7_461
timestamp 1607721120
transform 1 0 43516 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_457
timestamp 1607721120
transform 1 0 43148 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_467
timestamp 1607721120
transform 1 0 44068 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_459
timestamp 1607721120
transform 1 0 43332 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_457
timestamp 1607721120
transform 1 0 43148 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1138__B1
timestamp 1607721120
transform 1 0 43700 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__A1
timestamp 1607721120
transform 1 0 43332 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1607721120
transform 1 0 43240 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1169_
timestamp 1607721120
transform 1 0 43424 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_7_477
timestamp 1607721120
transform 1 0 44988 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_471
timestamp 1607721120
transform 1 0 44436 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__B1_N
timestamp 1607721120
transform 1 0 44252 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1138__A2
timestamp 1607721120
transform 1 0 44620 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__A1
timestamp 1607721120
transform 1 0 45172 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1143_
timestamp 1607721120
transform 1 0 44804 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_4  _1138_
timestamp 1607721120
transform 1 0 43884 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_489
timestamp 1607721120
transform 1 0 46092 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_485
timestamp 1607721120
transform 1 0 45724 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_481
timestamp 1607721120
transform 1 0 45356 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_488
timestamp 1607721120
transform 1 0 46000 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_484
timestamp 1607721120
transform 1 0 45632 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__C
timestamp 1607721120
transform 1 0 45816 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1138__A1
timestamp 1607721120
transform 1 0 45540 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1607721120
transform 1 0 46000 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_499
timestamp 1607721120
transform 1 0 47012 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__A
timestamp 1607721120
transform 1 0 46184 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1170_
timestamp 1607721120
transform 1 0 46184 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1168_
timestamp 1607721120
transform 1 0 46368 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_501
timestamp 1607721120
transform 1 0 47196 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1185__B
timestamp 1607721120
transform 1 0 47196 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_503
timestamp 1607721120
transform 1 0 47380 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_505
timestamp 1607721120
transform 1 0 47564 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1156__A1
timestamp 1607721120
transform 1 0 47748 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1168__B
timestamp 1607721120
transform 1 0 47380 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1185__D
timestamp 1607721120
transform 1 0 47564 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0988_
timestamp 1607721120
transform 1 0 47748 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_511
timestamp 1607721120
transform 1 0 48116 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_509
timestamp 1607721120
transform 1 0 47932 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__B
timestamp 1607721120
transform 1 0 48116 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_513
timestamp 1607721120
transform 1 0 48300 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__A
timestamp 1607721120
transform 1 0 48300 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_515
timestamp 1607721120
transform 1 0 48484 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_524
timestamp 1607721120
transform 1 0 49312 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__B2
timestamp 1607721120
transform 1 0 48668 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__A2
timestamp 1607721120
transform 1 0 48852 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1607721120
transform 1 0 48852 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1012_
timestamp 1607721120
transform 1 0 48944 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1105_
timestamp 1607721120
transform 1 0 49036 0 1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_7_534
timestamp 1607721120
transform 1 0 50232 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_532
timestamp 1607721120
transform 1 0 50048 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_528
timestamp 1607721120
transform 1 0 49680 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__A1
timestamp 1607721120
transform 1 0 49864 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__A
timestamp 1607721120
transform 1 0 49496 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  _1114_
timestamp 1607721120
transform 1 0 50232 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_542
timestamp 1607721120
transform 1 0 50968 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_538
timestamp 1607721120
transform 1 0 50600 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_543
timestamp 1607721120
transform 1 0 51060 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1100__B
timestamp 1607721120
transform 1 0 51152 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1100__C
timestamp 1607721120
transform 1 0 50784 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1395__D
timestamp 1607721120
transform 1 0 50416 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_546
timestamp 1607721120
transform 1 0 51336 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_547
timestamp 1607721120
transform 1 0 51428 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__C
timestamp 1607721120
transform 1 0 51244 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_556
timestamp 1607721120
transform 1 0 52256 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_550
timestamp 1607721120
transform 1 0 51704 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_558
timestamp 1607721120
transform 1 0 52440 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_552
timestamp 1607721120
transform 1 0 51888 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__C
timestamp 1607721120
transform 1 0 51704 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__B
timestamp 1607721120
transform 1 0 52256 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1025__A
timestamp 1607721120
transform 1 0 52440 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1607721120
transform 1 0 51612 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1025_
timestamp 1607721120
transform 1 0 51888 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_560
timestamp 1607721120
transform 1 0 52624 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__A
timestamp 1607721120
transform 1 0 52808 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1389_
timestamp 1607721120
transform 1 0 52992 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__a21o_4  _1188_
timestamp 1607721120
transform 1 0 52532 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_579
timestamp 1607721120
transform 1 0 54372 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_575
timestamp 1607721120
transform 1 0 54004 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_571
timestamp 1607721120
transform 1 0 53636 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__A1
timestamp 1607721120
transform 1 0 54188 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__A2
timestamp 1607721120
transform 1 0 53820 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1607721120
transform 1 0 54464 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_587
timestamp 1607721120
transform 1 0 55108 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_583
timestamp 1607721120
transform 1 0 54740 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_588
timestamp 1607721120
transform 1 0 55200 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_584
timestamp 1607721120
transform 1 0 54832 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1181__B1
timestamp 1607721120
transform 1 0 55292 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1183__A
timestamp 1607721120
transform 1 0 55016 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1181__A1
timestamp 1607721120
transform 1 0 55384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1107__A
timestamp 1607721120
transform 1 0 54924 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1183_
timestamp 1607721120
transform 1 0 54556 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_591
timestamp 1607721120
transform 1 0 55476 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__A
timestamp 1607721120
transform 1 0 55660 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1151_
timestamp 1607721120
transform 1 0 55568 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_602
timestamp 1607721120
transform 1 0 56488 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_605
timestamp 1607721120
transform 1 0 56764 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_601
timestamp 1607721120
transform 1 0 56396 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1151__C
timestamp 1607721120
transform 1 0 56580 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__A
timestamp 1607721120
transform 1 0 56672 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1121_
timestamp 1607721120
transform 1 0 55844 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_7_615
timestamp 1607721120
transform 1 0 57684 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_611
timestamp 1607721120
transform 1 0 57316 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_606
timestamp 1607721120
transform 1 0 56856 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__B1
timestamp 1607721120
transform 1 0 56948 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__B
timestamp 1607721120
transform 1 0 57040 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__B1
timestamp 1607721120
transform 1 0 57500 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1607721120
transform 1 0 57224 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1119_
timestamp 1607721120
transform 1 0 57132 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_625
timestamp 1607721120
transform 1 0 58604 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_621
timestamp 1607721120
transform 1 0 58236 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__A2
timestamp 1607721120
transform 1 0 58788 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__A1
timestamp 1607721120
transform 1 0 58420 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1400__D
timestamp 1607721120
transform 1 0 57868 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_638
timestamp 1607721120
transform 1 0 59800 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_637
timestamp 1607721120
transform 1 0 59708 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_633
timestamp 1607721120
transform 1 0 59340 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1173__A1_N
timestamp 1607721120
transform 1 0 59892 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1173__B2
timestamp 1607721120
transform 1 0 59524 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0960_
timestamp 1607721120
transform 1 0 58972 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1400_
timestamp 1607721120
transform 1 0 58052 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_7_642
timestamp 1607721120
transform 1 0 60168 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1252__A
timestamp 1607721120
transform 1 0 59984 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1254__A
timestamp 1607721120
transform 1 0 60352 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1607721120
transform 1 0 60076 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1254_
timestamp 1607721120
transform 1 0 60536 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_7_659
timestamp 1607721120
transform 1 0 61732 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_653
timestamp 1607721120
transform 1 0 61180 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1256__B
timestamp 1607721120
transform 1 0 61916 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1256__A
timestamp 1607721120
transform 1 0 61548 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_661
timestamp 1607721120
transform 1 0 61916 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1392_
timestamp 1607721120
transform 1 0 60168 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_7_672
timestamp 1607721120
transform 1 0 62928 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_663
timestamp 1607721120
transform 1 0 62100 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_673
timestamp 1607721120
transform 1 0 63020 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1607721120
transform 1 0 62836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1607721120
transform -1 0 63480 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1607721120
transform -1 0 63480 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_21
timestamp 1607721120
transform 1 0 3036 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_15
timestamp 1607721120
transform 1 0 2484 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1607721120
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1424__CLK
timestamp 1607721120
transform 1 0 3128 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1607721120
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_28
timestamp 1607721120
transform 1 0 3680 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_24
timestamp 1607721120
transform 1 0 3312 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1421__D
timestamp 1607721120
transform 1 0 3496 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1607721120
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1424_
timestamp 1607721120
transform 1 0 4048 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_8_68
timestamp 1607721120
transform 1 0 7360 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_55
timestamp 1607721120
transform 1 0 6164 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_51
timestamp 1607721120
transform 1 0 5796 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0942__A1
timestamp 1607721120
transform 1 0 5980 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__C
timestamp 1607721120
transform 1 0 6348 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0939_
timestamp 1607721120
transform 1 0 6532 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_8_87
timestamp 1607721120
transform 1 0 9108 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_83
timestamp 1607721120
transform 1 0 8740 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_75
timestamp 1607721120
transform 1 0 8004 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_72
timestamp 1607721120
transform 1 0 7728 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_wb_clk_i_A
timestamp 1607721120
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1201__A1
timestamp 1607721120
transform 1 0 7820 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1278__B
timestamp 1607721120
transform 1 0 8924 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1278_
timestamp 1607721120
transform 1 0 8096 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_8_93
timestamp 1607721120
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1266__B
timestamp 1607721120
transform 1 0 9844 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1607721120
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1385_
timestamp 1607721120
transform 1 0 10028 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_8_127
timestamp 1607721120
transform 1 0 12788 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_123
timestamp 1607721120
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_120
timestamp 1607721120
transform 1 0 12144 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_116
timestamp 1607721120
transform 1 0 11776 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__A1
timestamp 1607721120
transform 1 0 12236 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1286__A
timestamp 1607721120
transform 1 0 12604 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__A1
timestamp 1607721120
transform 1 0 12972 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1089_
timestamp 1607721120
transform 1 0 13156 0 -1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_8_158
timestamp 1607721120
transform 1 0 15640 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_154
timestamp 1607721120
transform 1 0 15272 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_149
timestamp 1607721120
transform 1 0 14812 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_145
timestamp 1607721120
transform 1 0 14444 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__B1
timestamp 1607721120
transform 1 0 15732 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__A1
timestamp 1607721120
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__B1
timestamp 1607721120
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1607721120
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_179
timestamp 1607721120
transform 1 0 17572 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_161
timestamp 1607721120
transform 1 0 15916 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__B1_N
timestamp 1607721120
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__C1
timestamp 1607721120
transform 1 0 17756 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1093_
timestamp 1607721120
transform 1 0 16284 0 -1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_8_205
timestamp 1607721120
transform 1 0 19964 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_201
timestamp 1607721120
transform 1 0 19596 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_183
timestamp 1607721120
transform 1 0 17940 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1087__B1
timestamp 1607721120
transform 1 0 18124 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1098_
timestamp 1607721120
transform 1 0 18308 0 -1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1607721120
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_208
timestamp 1607721120
transform 1 0 20240 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__B
timestamp 1607721120
transform 1 0 20056 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__A
timestamp 1607721120
transform 1 0 20516 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1607721120
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1069_
timestamp 1607721120
transform 1 0 20884 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_8_226
timestamp 1607721120
transform 1 0 21896 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_222
timestamp 1607721120
transform 1 0 21528 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__B1
timestamp 1607721120
transform 1 0 22080 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__B
timestamp 1607721120
transform 1 0 21712 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1607721120
transform 1 0 24104 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_242
timestamp 1607721120
transform 1 0 23368 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_238
timestamp 1607721120
transform 1 0 23000 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_230
timestamp 1607721120
transform 1 0 22264 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1408__CLK
timestamp 1607721120
transform 1 0 23552 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1403__CLK
timestamp 1607721120
transform 1 0 23184 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__C1
timestamp 1607721120
transform 1 0 22448 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1057_
timestamp 1607721120
transform 1 0 22632 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1048_
timestamp 1607721120
transform 1 0 23736 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_271
timestamp 1607721120
transform 1 0 26036 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_267
timestamp 1607721120
transform 1 0 25668 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_254
timestamp 1607721120
transform 1 0 24472 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1076__C
timestamp 1607721120
transform 1 0 24288 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1076__B
timestamp 1607721120
transform 1 0 24656 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__A2
timestamp 1607721120
transform 1 0 25852 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1070__B1
timestamp 1607721120
transform 1 0 26220 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1076_
timestamp 1607721120
transform 1 0 24840 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_296
timestamp 1607721120
transform 1 0 28336 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_292
timestamp 1607721120
transform 1 0 27968 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__B1
timestamp 1607721120
transform 1 0 28152 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1607721120
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1070_
timestamp 1607721120
transform 1 0 26496 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_317
timestamp 1607721120
transform 1 0 30268 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_313
timestamp 1607721120
transform 1 0 29900 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__A2
timestamp 1607721120
transform 1 0 30452 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__A1
timestamp 1607721120
transform 1 0 28520 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1406__D
timestamp 1607721120
transform 1 0 30084 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_4  _1052_
timestamp 1607721120
transform 1 0 28704 0 -1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_8_341
timestamp 1607721120
transform 1 0 32476 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_333
timestamp 1607721120
transform 1 0 31740 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_329
timestamp 1607721120
transform 1 0 31372 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_325
timestamp 1607721120
transform 1 0 31004 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__A
timestamp 1607721120
transform 1 0 31188 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__B
timestamp 1607721120
transform 1 0 31832 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1607721120
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1071_
timestamp 1607721120
transform 1 0 32108 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0937_
timestamp 1607721120
transform 1 0 30636 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_349
timestamp 1607721120
transform 1 0 33212 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_345
timestamp 1607721120
transform 1 0 32844 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__B
timestamp 1607721120
transform 1 0 33028 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__A
timestamp 1607721120
transform 1 0 32660 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1384_
timestamp 1607721120
transform 1 0 33488 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_8_386
timestamp 1607721120
transform 1 0 36616 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_376
timestamp 1607721120
transform 1 0 35696 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_371
timestamp 1607721120
transform 1 0 35236 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1250__B
timestamp 1607721120
transform 1 0 36800 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__A1
timestamp 1607721120
transform 1 0 35512 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1250_
timestamp 1607721120
transform 1 0 35972 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_8_398
timestamp 1607721120
transform 1 0 37720 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_394
timestamp 1607721120
transform 1 0 37352 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_390
timestamp 1607721120
transform 1 0 36984 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1285__A
timestamp 1607721120
transform 1 0 37168 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1607721120
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1111_
timestamp 1607721120
transform 1 0 37812 0 -1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_8_433
timestamp 1607721120
transform 1 0 40940 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_429
timestamp 1607721120
transform 1 0 40572 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_416
timestamp 1607721120
transform 1 0 39376 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_412
timestamp 1607721120
transform 1 0 39008 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__A2
timestamp 1607721120
transform 1 0 39560 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__B
timestamp 1607721120
transform 1 0 40756 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__B1
timestamp 1607721120
transform 1 0 39192 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1112_
timestamp 1607721120
transform 1 0 39744 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_456
timestamp 1607721120
transform 1 0 43056 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_452
timestamp 1607721120
transform 1 0 42688 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_447
timestamp 1607721120
transform 1 0 42228 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_437
timestamp 1607721120
transform 1 0 41308 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__C1
timestamp 1607721120
transform 1 0 42504 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__C
timestamp 1607721120
transform 1 0 41124 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__A2
timestamp 1607721120
transform 1 0 42872 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1148_
timestamp 1607721120
transform 1 0 41400 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_464
timestamp 1607721120
transform 1 0 43792 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_459
timestamp 1607721120
transform 1 0 43332 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1185__C
timestamp 1607721120
transform 1 0 43608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__C
timestamp 1607721120
transform 1 0 43976 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1607721120
transform 1 0 43240 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_4  _1142_
timestamp 1607721120
transform 1 0 44160 0 -1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_8_502
timestamp 1607721120
transform 1 0 47288 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_492
timestamp 1607721120
transform 1 0 46368 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_489
timestamp 1607721120
transform 1 0 46092 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_485
timestamp 1607721120
transform 1 0 45724 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_481
timestamp 1607721120
transform 1 0 45356 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__A
timestamp 1607721120
transform 1 0 46184 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__A2
timestamp 1607721120
transform 1 0 45540 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1185_
timestamp 1607721120
transform 1 0 46460 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_506
timestamp 1607721120
transform 1 0 47656 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__B1
timestamp 1607721120
transform 1 0 47472 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_510
timestamp 1607721120
transform 1 0 48024 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__B2
timestamp 1607721120
transform 1 0 47840 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__C
timestamp 1607721120
transform 1 0 48208 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_514
timestamp 1607721120
transform 1 0 48392 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__C
timestamp 1607721120
transform 1 0 48576 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_520
timestamp 1607721120
transform 1 0 48944 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_518
timestamp 1607721120
transform 1 0 48760 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1607721120
transform 1 0 48852 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_524
timestamp 1607721120
transform 1 0 49312 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__B1
timestamp 1607721120
transform 1 0 49128 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_548
timestamp 1607721120
transform 1 0 51520 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__C1
timestamp 1607721120
transform 1 0 49588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1395_
timestamp 1607721120
transform 1 0 49772 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_8_569
timestamp 1607721120
transform 1 0 53452 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_563
timestamp 1607721120
transform 1 0 52900 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_552
timestamp 1607721120
transform 1 0 51888 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1100__A
timestamp 1607721120
transform 1 0 52072 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__A
timestamp 1607721120
transform 1 0 51704 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1389__D
timestamp 1607721120
transform 1 0 53268 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1187_
timestamp 1607721120
transform 1 0 52256 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_8_573
timestamp 1607721120
transform 1 0 53820 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__A
timestamp 1607721120
transform 1 0 54004 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__B
timestamp 1607721120
transform 1 0 53636 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_577
timestamp 1607721120
transform 1 0 54188 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1607721120
transform 1 0 54464 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_581
timestamp 1607721120
transform 1 0 54556 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1389__CLK
timestamp 1607721120
transform 1 0 54740 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1107_
timestamp 1607721120
transform 1 0 54924 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_589
timestamp 1607721120
transform 1 0 55292 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_593
timestamp 1607721120
transform 1 0 55660 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1151__A
timestamp 1607721120
transform 1 0 55476 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_610
timestamp 1607721120
transform 1 0 57224 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_606
timestamp 1607721120
transform 1 0 56856 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__C
timestamp 1607721120
transform 1 0 57040 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__A1
timestamp 1607721120
transform 1 0 57408 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__B
timestamp 1607721120
transform 1 0 55844 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1129_
timestamp 1607721120
transform 1 0 56028 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_4  _1118_
timestamp 1607721120
transform 1 0 57592 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_638
timestamp 1607721120
transform 1 0 59800 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_634
timestamp 1607721120
transform 1 0 59432 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_630
timestamp 1607721120
transform 1 0 59064 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_626
timestamp 1607721120
transform 1 0 58696 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__A2
timestamp 1607721120
transform 1 0 59248 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1252__B
timestamp 1607721120
transform 1 0 59892 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__A1
timestamp 1607721120
transform 1 0 58880 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_653
timestamp 1607721120
transform 1 0 61180 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_649
timestamp 1607721120
transform 1 0 60812 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1400__CLK
timestamp 1607721120
transform 1 0 61364 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1254__B
timestamp 1607721120
transform 1 0 60996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1607721120
transform 1 0 60076 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1256_
timestamp 1607721120
transform 1 0 61548 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1252_
timestamp 1607721120
transform 1 0 60168 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_8_672
timestamp 1607721120
transform 1 0 62928 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_664
timestamp 1607721120
transform 1 0 62192 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1607721120
transform -1 0 63480 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1607721120
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1607721120
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1607721120
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_37
timestamp 1607721120
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_33
timestamp 1607721120
transform 1 0 4140 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_29
timestamp 1607721120
transform 1 0 3772 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1423__CLK
timestamp 1607721120
transform 1 0 3588 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1404__CLK
timestamp 1607721120
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1385__CLK
timestamp 1607721120
transform 1 0 4692 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1423__D
timestamp 1607721120
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _0942_
timestamp 1607721120
transform 1 0 4876 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1607721120
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_53
timestamp 1607721120
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0942__A2
timestamp 1607721120
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__B1
timestamp 1607721120
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1607721120
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1201_
timestamp 1607721120
transform 1 0 6808 0 1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_9_88
timestamp 1607721120
transform 1 0 9200 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_84
timestamp 1607721120
transform 1 0 8832 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_80
timestamp 1607721120
transform 1 0 8464 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_76
timestamp 1607721120
transform 1 0 8096 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1201__B2
timestamp 1607721120
transform 1 0 9016 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1201__A2
timestamp 1607721120
transform 1 0 8648 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1201__B1
timestamp 1607721120
transform 1 0 8280 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_114
timestamp 1607721120
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_92
timestamp 1607721120
transform 1 0 9568 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1404__D
timestamp 1607721120
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1404_
timestamp 1607721120
transform 1 0 9844 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_9_118
timestamp 1607721120
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__A
timestamp 1607721120
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__A1
timestamp 1607721120
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1607721120
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0932_
timestamp 1607721120
transform 1 0 12420 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_127
timestamp 1607721120
transform 1 0 12788 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_131
timestamp 1607721120
transform 1 0 13156 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__A
timestamp 1607721120
transform 1 0 13340 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__B
timestamp 1607721120
transform 1 0 12972 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_135
timestamp 1607721120
transform 1 0 13524 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1287__A
timestamp 1607721120
transform 1 0 13892 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1403_
timestamp 1607721120
transform 1 0 14076 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_9_179
timestamp 1607721120
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_175
timestamp 1607721120
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp 1607721120
transform 1 0 16284 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_160
timestamp 1607721120
transform 1 0 15824 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__A2
timestamp 1607721120
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__A1
timestamp 1607721120
transform 1 0 16100 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__A
timestamp 1607721120
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0946_
timestamp 1607721120
transform 1 0 16560 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_9_188
timestamp 1607721120
transform 1 0 18400 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_184
timestamp 1607721120
transform 1 0 18032 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__C
timestamp 1607721120
transform 1 0 18768 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1402__D
timestamp 1607721120
transform 1 0 18216 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1607721120
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1083_
timestamp 1607721120
transform 1 0 18952 0 1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_9_227
timestamp 1607721120
transform 1 0 21988 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_223
timestamp 1607721120
transform 1 0 21620 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_212
timestamp 1607721120
transform 1 0 20608 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_208
timestamp 1607721120
transform 1 0 20240 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1083__A2
timestamp 1607721120
transform 1 0 20792 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__A
timestamp 1607721120
transform 1 0 21804 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1083__A1
timestamp 1607721120
transform 1 0 20424 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1094_
timestamp 1607721120
transform 1 0 20976 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_9_231
timestamp 1607721120
transform 1 0 22356 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__B
timestamp 1607721120
transform 1 0 22172 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1061_
timestamp 1607721120
transform 1 0 22448 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_236
timestamp 1607721120
transform 1 0 22816 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__A
timestamp 1607721120
transform 1 0 23000 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_240
timestamp 1607721120
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__A
timestamp 1607721120
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_245
timestamp 1607721120
transform 1 0 23644 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__B
timestamp 1607721120
transform 1 0 23828 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1607721120
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_249
timestamp 1607721120
transform 1 0 24012 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__D
timestamp 1607721120
transform 1 0 24196 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_264
timestamp 1607721120
transform 1 0 25392 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_260
timestamp 1607721120
transform 1 0 25024 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1073__C1
timestamp 1607721120
transform 1 0 25576 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1072__A
timestamp 1607721120
transform 1 0 25208 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1073_
timestamp 1607721120
transform 1 0 25760 0 1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_4  _1072_
timestamp 1607721120
transform 1 0 24380 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_9_286
timestamp 1607721120
transform 1 0 27416 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_282
timestamp 1607721120
transform 1 0 27048 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1070__A1_N
timestamp 1607721120
transform 1 0 27600 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1407__D
timestamp 1607721120
transform 1 0 27232 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1065_
timestamp 1607721120
transform 1 0 27784 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_9_319
timestamp 1607721120
transform 1 0 30452 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_315
timestamp 1607721120
transform 1 0 30084 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_301
timestamp 1607721120
transform 1 0 28796 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_297
timestamp 1607721120
transform 1 0 28428 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__D
timestamp 1607721120
transform 1 0 30268 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1070__A2_N
timestamp 1607721120
transform 1 0 28980 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__B
timestamp 1607721120
transform 1 0 28612 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1607721120
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _1051_
timestamp 1607721120
transform 1 0 29256 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__D
timestamp 1607721120
transform 1 0 30636 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0887_
timestamp 1607721120
transform 1 0 30820 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_327
timestamp 1607721120
transform 1 0 31188 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__A
timestamp 1607721120
transform 1 0 31372 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_331
timestamp 1607721120
transform 1 0 31556 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__B
timestamp 1607721120
transform 1 0 31740 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_339
timestamp 1607721120
transform 1 0 32292 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_335
timestamp 1607721120
transform 1 0 31924 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__A
timestamp 1607721120
transform 1 0 32384 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1206_
timestamp 1607721120
transform 1 0 32568 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_362
timestamp 1607721120
transform 1 0 34408 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_358
timestamp 1607721120
transform 1 0 34040 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_350
timestamp 1607721120
transform 1 0 33304 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_346
timestamp 1607721120
transform 1 0 32936 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__A
timestamp 1607721120
transform 1 0 33120 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0944__A
timestamp 1607721120
transform 1 0 33488 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__B
timestamp 1607721120
transform 1 0 34592 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__A
timestamp 1607721120
transform 1 0 34224 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0944_
timestamp 1607721120
transform 1 0 33672 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_382
timestamp 1607721120
transform 1 0 36248 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_378
timestamp 1607721120
transform 1 0 35880 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_374
timestamp 1607721120
transform 1 0 35512 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__A2
timestamp 1607721120
transform 1 0 36064 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1244__A
timestamp 1607721120
transform 1 0 35696 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1607721120
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _1285_
timestamp 1607721120
transform 1 0 36524 0 1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_4  _1244_
timestamp 1607721120
transform 1 0 34868 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_9_402
timestamp 1607721120
transform 1 0 38088 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_398
timestamp 1607721120
transform 1 0 37720 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__B1
timestamp 1607721120
transform 1 0 38364 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1285__C
timestamp 1607721120
transform 1 0 37904 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1108_
timestamp 1607721120
transform 1 0 38548 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_423
timestamp 1607721120
transform 1 0 40020 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_419
timestamp 1607721120
transform 1 0 39652 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__A1
timestamp 1607721120
transform 1 0 40204 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__C1
timestamp 1607721120
transform 1 0 39836 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1607721120
transform 1 0 40388 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1128_
timestamp 1607721120
transform 1 0 40480 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1607721120
transform 1 0 42228 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_443
timestamp 1607721120
transform 1 0 41860 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_439
timestamp 1607721120
transform 1 0 41492 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_435
timestamp 1607721120
transform 1 0 41124 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0806__A
timestamp 1607721120
transform 1 0 42044 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0806__B
timestamp 1607721120
transform 1 0 41676 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__A
timestamp 1607721120
transform 1 0 41308 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1394_
timestamp 1607721120
transform 1 0 42320 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_9_479
timestamp 1607721120
transform 1 0 45172 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_471
timestamp 1607721120
transform 1 0 44436 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_467
timestamp 1607721120
transform 1 0 44068 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__A
timestamp 1607721120
transform 1 0 44252 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__B1
timestamp 1607721120
transform 1 0 44620 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0805_
timestamp 1607721120
transform 1 0 44804 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_499
timestamp 1607721120
transform 1 0 47012 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_489
timestamp 1607721120
transform 1 0 46092 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_487
timestamp 1607721120
transform 1 0 45908 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_483
timestamp 1607721120
transform 1 0 45540 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__A1
timestamp 1607721120
transform 1 0 45724 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__C1
timestamp 1607721120
transform 1 0 45356 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1132__B
timestamp 1607721120
transform 1 0 47196 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1607721120
transform 1 0 46000 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _1132_
timestamp 1607721120
transform 1 0 46184 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_520
timestamp 1607721120
transform 1 0 48944 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_516
timestamp 1607721120
transform 1 0 48576 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_503
timestamp 1607721120
transform 1 0 47380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1115__B
timestamp 1607721120
transform 1 0 48760 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1115__A
timestamp 1607721120
transform 1 0 49128 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__A1
timestamp 1607721120
transform 1 0 47564 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1145_
timestamp 1607721120
transform 1 0 49312 0 1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__and4_4  _1104_
timestamp 1607721120
transform 1 0 47748 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_9_546
timestamp 1607721120
transform 1 0 51336 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_542
timestamp 1607721120
transform 1 0 50968 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_538
timestamp 1607721120
transform 1 0 50600 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__A2
timestamp 1607721120
transform 1 0 51152 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__A1
timestamp 1607721120
transform 1 0 50784 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1607721120
transform 1 0 51612 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0796_
timestamp 1607721120
transform 1 0 51704 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_554
timestamp 1607721120
transform 1 0 52072 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__A
timestamp 1607721120
transform 1 0 52256 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_558
timestamp 1607721120
transform 1 0 52440 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__B
timestamp 1607721120
transform 1 0 52624 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0934_
timestamp 1607721120
transform 1 0 52808 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_566
timestamp 1607721120
transform 1 0 53176 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_570
timestamp 1607721120
transform 1 0 53544 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__A
timestamp 1607721120
transform 1 0 53360 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_578
timestamp 1607721120
transform 1 0 54280 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__A
timestamp 1607721120
transform 1 0 54464 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1102__A
timestamp 1607721120
transform 1 0 53728 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1110_
timestamp 1607721120
transform 1 0 53912 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_589
timestamp 1607721120
transform 1 0 55292 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_586
timestamp 1607721120
transform 1 0 55016 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_582
timestamp 1607721120
transform 1 0 54648 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__A1
timestamp 1607721120
transform 1 0 55108 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1125__B
timestamp 1607721120
transform 1 0 55476 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  _1125_
timestamp 1607721120
transform 1 0 55660 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_611
timestamp 1607721120
transform 1 0 57316 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_606
timestamp 1607721120
transform 1 0 56856 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_602
timestamp 1607721120
transform 1 0 56488 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__B1
timestamp 1607721120
transform 1 0 56672 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__B2
timestamp 1607721120
transform 1 0 57040 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1607721120
transform 1 0 57224 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1122_
timestamp 1607721120
transform 1 0 57408 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_632
timestamp 1607721120
transform 1 0 59248 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_628
timestamp 1607721120
transform 1 0 58880 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__A2_N
timestamp 1607721120
transform 1 0 59432 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__A1_N
timestamp 1607721120
transform 1 0 59064 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  _1127_
timestamp 1607721120
transform 1 0 59616 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_9_653
timestamp 1607721120
transform 1 0 61180 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_649
timestamp 1607721120
transform 1 0 60812 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_645
timestamp 1607721120
transform 1 0 60444 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1126__A
timestamp 1607721120
transform 1 0 60996 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__A
timestamp 1607721120
transform 1 0 60628 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_672
timestamp 1607721120
transform 1 0 62928 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_665
timestamp 1607721120
transform 1 0 62284 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1607721120
transform 1 0 62836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1607721120
transform -1 0 63480 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1607721120
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1607721120
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1607721120
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1607721120
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1607721120
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1423_
timestamp 1607721120
transform 1 0 4048 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_10_55
timestamp 1607721120
transform 1 0 6164 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_51
timestamp 1607721120
transform 1 0 5796 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__B2
timestamp 1607721120
transform 1 0 6348 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0942__B1
timestamp 1607721120
transform 1 0 5980 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _1202_
timestamp 1607721120
transform 1 0 6532 0 -1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_10_89
timestamp 1607721120
transform 1 0 9292 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1607721120
transform 1 0 8924 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_81
timestamp 1607721120
transform 1 0 8556 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_77
timestamp 1607721120
transform 1 0 8188 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_73
timestamp 1607721120
transform 1 0 7820 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__A1
timestamp 1607721120
transform 1 0 9108 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0948__A1
timestamp 1607721120
transform 1 0 8740 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1279__A1
timestamp 1607721120
transform 1 0 8372 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__A2
timestamp 1607721120
transform 1 0 8004 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_106
timestamp 1607721120
transform 1 0 10856 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_102
timestamp 1607721120
transform 1 0 10488 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1281__A2
timestamp 1607721120
transform 1 0 11040 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1266__A
timestamp 1607721120
transform 1 0 10672 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1607721120
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1266_
timestamp 1607721120
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _0940_
timestamp 1607721120
transform 1 0 11224 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_10_134
timestamp 1607721120
transform 1 0 13432 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_125
timestamp 1607721120
transform 1 0 12604 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_121
timestamp 1607721120
transform 1 0 12236 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_117
timestamp 1607721120
transform 1 0 11868 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__A
timestamp 1607721120
transform 1 0 13616 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__B
timestamp 1607721120
transform 1 0 12052 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0932__A
timestamp 1607721120
transform 1 0 12420 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0882_
timestamp 1607721120
transform 1 0 12788 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_10_150
timestamp 1607721120
transform 1 0 14904 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_146
timestamp 1607721120
transform 1 0 14536 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_142
timestamp 1607721120
transform 1 0 14168 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1607721120
transform 1 0 13800 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__B1
timestamp 1607721120
transform 1 0 13984 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__A1
timestamp 1607721120
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1403__D
timestamp 1607721120
transform 1 0 14352 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1607721120
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1088_
timestamp 1607721120
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_177
timestamp 1607721120
transform 1 0 17388 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_171
timestamp 1607721120
transform 1 0 16836 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_166
timestamp 1607721120
transform 1 0 16376 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__B
timestamp 1607721120
transform 1 0 16652 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0861__A
timestamp 1607721120
transform 1 0 17204 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1402_
timestamp 1607721120
transform 1 0 17572 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_10_203
timestamp 1607721120
transform 1 0 19780 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_198
timestamp 1607721120
transform 1 0 19320 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1083__B1
timestamp 1607721120
transform 1 0 19964 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1083__B2
timestamp 1607721120
transform 1 0 19596 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_226
timestamp 1607721120
transform 1 0 21896 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_222
timestamp 1607721120
transform 1 0 21528 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_211
timestamp 1607721120
transform 1 0 20516 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_207
timestamp 1607721120
transform 1 0 20148 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__B
timestamp 1607721120
transform 1 0 22080 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__A
timestamp 1607721120
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__B
timestamp 1607721120
transform 1 0 21712 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1607721120
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1084_
timestamp 1607721120
transform 1 0 20884 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_10_248
timestamp 1607721120
transform 1 0 23920 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_242
timestamp 1607721120
transform 1 0 23368 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_238
timestamp 1607721120
transform 1 0 23000 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_234
timestamp 1607721120
transform 1 0 22632 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1407__CLK
timestamp 1607721120
transform 1 0 23736 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1402__CLK
timestamp 1607721120
transform 1 0 23184 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__C
timestamp 1607721120
transform 1 0 24104 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__A
timestamp 1607721120
transform 1 0 22816 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0860_
timestamp 1607721120
transform 1 0 22264 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_271
timestamp 1607721120
transform 1 0 26036 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_267
timestamp 1607721120
transform 1 0 25668 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_256
timestamp 1607721120
transform 1 0 24656 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_252
timestamp 1607721120
transform 1 0 24288 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1072__B
timestamp 1607721120
transform 1 0 24472 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1073__A2
timestamp 1607721120
transform 1 0 25852 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1073__A1
timestamp 1607721120
transform 1 0 26220 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1046_
timestamp 1607721120
transform 1 0 24840 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_295
timestamp 1607721120
transform 1 0 28244 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1607721120
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1407_
timestamp 1607721120
transform 1 0 26496 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_10_316
timestamp 1607721120
transform 1 0 30176 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_312
timestamp 1607721120
transform 1 0 29808 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_299
timestamp 1607721120
transform 1 0 28612 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__C
timestamp 1607721120
transform 1 0 30360 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__C
timestamp 1607721120
transform 1 0 29992 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__A1
timestamp 1607721120
transform 1 0 28796 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1073__B1
timestamp 1607721120
transform 1 0 28428 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _1050_
timestamp 1607721120
transform 1 0 28980 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_324
timestamp 1607721120
transform 1 0 30912 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0826_
timestamp 1607721120
transform 1 0 30544 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_328
timestamp 1607721120
transform 1 0 31280 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__A
timestamp 1607721120
transform 1 0 31096 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_332
timestamp 1607721120
transform 1 0 31648 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__A
timestamp 1607721120
transform 1 0 31832 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__B
timestamp 1607721120
transform 1 0 31464 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_337
timestamp 1607721120
transform 1 0 32108 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1607721120
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0938_
timestamp 1607721120
transform 1 0 32384 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_362
timestamp 1607721120
transform 1 0 34408 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_353
timestamp 1607721120
transform 1 0 33580 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_348
timestamp 1607721120
transform 1 0 33120 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_344
timestamp 1607721120
transform 1 0 32752 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1347__A
timestamp 1607721120
transform 1 0 32936 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1245__B1
timestamp 1607721120
transform 1 0 34592 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1230__B
timestamp 1607721120
transform 1 0 33396 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0933_
timestamp 1607721120
transform 1 0 33764 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_10_387
timestamp 1607721120
transform 1 0 36708 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_383
timestamp 1607721120
transform 1 0 36340 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_366
timestamp 1607721120
transform 1 0 34776 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1284__C
timestamp 1607721120
transform 1 0 36524 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1244__B
timestamp 1607721120
transform 1 0 34960 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__nor3_4  _1284_
timestamp 1607721120
transform 1 0 35144 0 -1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_10_398
timestamp 1607721120
transform 1 0 37720 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_396
timestamp 1607721120
transform 1 0 37536 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_391
timestamp 1607721120
transform 1 0 37076 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1284__B
timestamp 1607721120
transform 1 0 36892 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1285__B
timestamp 1607721120
transform 1 0 37352 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1607721120
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_402
timestamp 1607721120
transform 1 0 38088 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1284__A
timestamp 1607721120
transform 1 0 37904 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__B1
timestamp 1607721120
transform 1 0 38364 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1113_
timestamp 1607721120
transform 1 0 38548 0 -1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_10_430
timestamp 1607721120
transform 1 0 40664 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_425
timestamp 1607721120
transform 1 0 40204 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_421
timestamp 1607721120
transform 1 0 39836 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__A1
timestamp 1607721120
transform 1 0 40848 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__A2
timestamp 1607721120
transform 1 0 40020 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__B
timestamp 1607721120
transform 1 0 40480 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_453
timestamp 1607721120
transform 1 0 42780 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_448
timestamp 1607721120
transform 1 0 42320 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_444
timestamp 1607721120
transform 1 0 41952 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_434
timestamp 1607721120
transform 1 0 41032 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__A
timestamp 1607721120
transform 1 0 42964 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__A
timestamp 1607721120
transform 1 0 42136 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1394__D
timestamp 1607721120
transform 1 0 42596 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0806_
timestamp 1607721120
transform 1 0 41308 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_10_463
timestamp 1607721120
transform 1 0 43700 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_459
timestamp 1607721120
transform 1 0 43332 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_457
timestamp 1607721120
transform 1 0 43148 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1132__A
timestamp 1607721120
transform 1 0 43976 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1234__B
timestamp 1607721120
transform 1 0 43516 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1607721120
transform 1 0 43240 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1140_
timestamp 1607721120
transform 1 0 44160 0 -1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_10_492
timestamp 1607721120
transform 1 0 46368 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_486
timestamp 1607721120
transform 1 0 45816 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_482
timestamp 1607721120
transform 1 0 45448 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__A2
timestamp 1607721120
transform 1 0 45632 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1132__D
timestamp 1607721120
transform 1 0 46184 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _1134_
timestamp 1607721120
transform 1 0 46644 0 -1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_10_517
timestamp 1607721120
transform 1 0 48668 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_513
timestamp 1607721120
transform 1 0 48300 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_509
timestamp 1607721120
transform 1 0 47932 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__D
timestamp 1607721120
transform 1 0 48484 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__A2
timestamp 1607721120
transform 1 0 48116 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1607721120
transform 1 0 48852 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1115_
timestamp 1607721120
transform 1 0 48944 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_10_548
timestamp 1607721120
transform 1 0 51520 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_544
timestamp 1607721120
transform 1 0 51152 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_532
timestamp 1607721120
transform 1 0 50048 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_527
timestamp 1607721120
transform 1 0 49588 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1261__A1
timestamp 1607721120
transform 1 0 51336 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__B1
timestamp 1607721120
transform 1 0 49864 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1100_
timestamp 1607721120
transform 1 0 50324 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_563
timestamp 1607721120
transform 1 0 52900 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_559
timestamp 1607721120
transform 1 0 52532 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__A
timestamp 1607721120
transform 1 0 53084 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__A
timestamp 1607721120
transform 1 0 52716 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1100__D
timestamp 1607721120
transform 1 0 51704 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1260_
timestamp 1607721120
transform 1 0 51888 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1102_
timestamp 1607721120
transform 1 0 53268 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_581
timestamp 1607721120
transform 1 0 54556 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_579
timestamp 1607721120
transform 1 0 54372 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_575
timestamp 1607721120
transform 1 0 54004 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_571
timestamp 1607721120
transform 1 0 53636 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1395__CLK
timestamp 1607721120
transform 1 0 54188 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1361__CLK
timestamp 1607721120
transform 1 0 53820 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1607721120
transform 1 0 54464 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_589
timestamp 1607721120
transform 1 0 55292 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_585
timestamp 1607721120
transform 1 0 54924 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1397__CLK
timestamp 1607721120
transform 1 0 55108 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__A
timestamp 1607721120
transform 1 0 54740 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__A2
timestamp 1607721120
transform 1 0 55476 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1136_
timestamp 1607721120
transform 1 0 55660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_609
timestamp 1607721120
transform 1 0 57132 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_605
timestamp 1607721120
transform 1 0 56764 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__B1
timestamp 1607721120
transform 1 0 57316 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1125__A
timestamp 1607721120
transform 1 0 56948 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1124_
timestamp 1607721120
transform 1 0 57500 0 -1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_10_635
timestamp 1607721120
transform 1 0 59524 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_631
timestamp 1607721120
transform 1 0 59156 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_627
timestamp 1607721120
transform 1 0 58788 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__B
timestamp 1607721120
transform 1 0 59800 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__B
timestamp 1607721120
transform 1 0 59340 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__C1
timestamp 1607721120
transform 1 0 58972 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_655
timestamp 1607721120
transform 1 0 61364 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_651
timestamp 1607721120
transform 1 0 60996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_640
timestamp 1607721120
transform 1 0 59984 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1126__B
timestamp 1607721120
transform 1 0 61180 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1607721120
transform 1 0 60076 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1126_
timestamp 1607721120
transform 1 0 60168 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_667
timestamp 1607721120
transform 1 0 62468 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1607721120
transform -1 0 63480 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_22
timestamp 1607721120
transform 1 0 3128 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_18
timestamp 1607721120
transform 1 0 2760 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_15
timestamp 1607721120
transform 1 0 2484 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1607721120
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1283__B1
timestamp 1607721120
transform 1 0 2576 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1283__A2
timestamp 1607721120
transform 1 0 2944 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1607721120
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_26
timestamp 1607721120
transform 1 0 3496 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1283__A1
timestamp 1607721120
transform 1 0 3312 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1422__D
timestamp 1607721120
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1422_
timestamp 1607721120
transform 1 0 4232 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1607721120
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_53
timestamp 1607721120
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__A2
timestamp 1607721120
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__B1
timestamp 1607721120
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1607721120
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _0948_
timestamp 1607721120
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_91
timestamp 1607721120
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_78
timestamp 1607721120
transform 1 0 8280 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_74
timestamp 1607721120
transform 1 0 7912 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0948__A2
timestamp 1607721120
transform 1 0 8464 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0948__B1
timestamp 1607721120
transform 1 0 8096 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1203_
timestamp 1607721120
transform 1 0 8648 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_114
timestamp 1607721120
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_95
timestamp 1607721120
transform 1 0 9844 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1203__B
timestamp 1607721120
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0941__B1
timestamp 1607721120
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_4  _0941_
timestamp 1607721120
transform 1 0 10396 0 1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_11_123
timestamp 1607721120
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_118
timestamp 1607721120
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__A2
timestamp 1607721120
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__A1
timestamp 1607721120
transform 1 0 12604 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0941__A1
timestamp 1607721120
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1607721120
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_131
timestamp 1607721120
transform 1 0 13156 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_127
timestamp 1607721120
transform 1 0 12788 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__B
timestamp 1607721120
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1210_
timestamp 1607721120
transform 1 0 13432 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_154
timestamp 1607721120
transform 1 0 15272 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_150
timestamp 1607721120
transform 1 0 14904 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_146
timestamp 1607721120
transform 1 0 14536 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__A1
timestamp 1607721120
transform 1 0 15088 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__A2
timestamp 1607721120
transform 1 0 14720 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0852_
timestamp 1607721120
transform 1 0 15456 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_179
timestamp 1607721120
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_175
timestamp 1607721120
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_164
timestamp 1607721120
transform 1 0 16192 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_160
timestamp 1607721120
transform 1 0 15824 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__A2
timestamp 1607721120
transform 1 0 16376 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0861__B
timestamp 1607721120
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__B
timestamp 1607721120
transform 1 0 16008 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1224__A
timestamp 1607721120
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1224_
timestamp 1607721120
transform 1 0 16560 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_11_203
timestamp 1607721120
transform 1 0 19780 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_199
timestamp 1607721120
transform 1 0 19412 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_195
timestamp 1607721120
transform 1 0 19044 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_184
timestamp 1607721120
transform 1 0 18032 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__D
timestamp 1607721120
transform 1 0 19596 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__B
timestamp 1607721120
transform 1 0 19228 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1607721120
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _1082_
timestamp 1607721120
transform 1 0 18216 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_219
timestamp 1607721120
transform 1 0 21252 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_215
timestamp 1607721120
transform 1 0 20884 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__A
timestamp 1607721120
transform 1 0 21436 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__A
timestamp 1607721120
transform 1 0 21068 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1228_
timestamp 1607721120
transform 1 0 21620 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _1212_
timestamp 1607721120
transform 1 0 20056 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_230
timestamp 1607721120
transform 1 0 22264 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1220__A
timestamp 1607721120
transform 1 0 22448 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_238
timestamp 1607721120
transform 1 0 23000 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_234
timestamp 1607721120
transform 1 0 22632 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1220__B
timestamp 1607721120
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1405__CLK
timestamp 1607721120
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_245
timestamp 1607721120
transform 1 0 23644 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1607721120
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_250
timestamp 1607721120
transform 1 0 24104 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__A1
timestamp 1607721120
transform 1 0 23920 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_262
timestamp 1607721120
transform 1 0 25208 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_257
timestamp 1607721120
transform 1 0 24748 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__B1
timestamp 1607721120
transform 1 0 24288 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__B1
timestamp 1607721120
transform 1 0 25024 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_4  _1081_
timestamp 1607721120
transform 1 0 25484 0 1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1080_
timestamp 1607721120
transform 1 0 24472 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_295
timestamp 1607721120
transform 1 0 28244 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_284
timestamp 1607721120
transform 1 0 27232 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_278
timestamp 1607721120
transform 1 0 26680 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__B1
timestamp 1607721120
transform 1 0 27048 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _0961_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 27416 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_303
timestamp 1607721120
transform 1 0 28980 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_299
timestamp 1607721120
transform 1 0 28612 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__B
timestamp 1607721120
transform 1 0 28796 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__B
timestamp 1607721120
transform 1 0 28428 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1607721120
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1077_
timestamp 1607721120
transform 1 0 29256 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_11_317
timestamp 1607721120
transform 1 0 30268 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_313
timestamp 1607721120
transform 1 0 29900 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__A
timestamp 1607721120
transform 1 0 30452 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__B
timestamp 1607721120
transform 1 0 30084 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_341
timestamp 1607721120
transform 1 0 32476 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_329
timestamp 1607721120
transform 1 0 31372 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_325
timestamp 1607721120
transform 1 0 31004 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1246__B
timestamp 1607721120
transform 1 0 31648 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__A
timestamp 1607721120
transform 1 0 31188 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1246_
timestamp 1607721120
transform 1 0 31832 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0853_
timestamp 1607721120
transform 1 0 30636 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_362
timestamp 1607721120
transform 1 0 34408 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_358
timestamp 1607721120
transform 1 0 34040 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_345
timestamp 1607721120
transform 1 0 32844 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1245__A2
timestamp 1607721120
transform 1 0 34592 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1347__B
timestamp 1607721120
transform 1 0 33028 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1230__A
timestamp 1607721120
transform 1 0 34224 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1246__A
timestamp 1607721120
transform 1 0 32660 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  _1230_
timestamp 1607721120
transform 1 0 33212 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_11_388
timestamp 1607721120
transform 1 0 36800 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_384
timestamp 1607721120
transform 1 0 36432 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_380
timestamp 1607721120
transform 1 0 36064 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_376
timestamp 1607721120
transform 1 0 35696 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1245__A1
timestamp 1607721120
transform 1 0 36616 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1248__A
timestamp 1607721120
transform 1 0 36248 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__A
timestamp 1607721120
transform 1 0 35880 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1607721120
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1248_
timestamp 1607721120
transform 1 0 34868 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_411
timestamp 1607721120
transform 1 0 38916 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_407
timestamp 1607721120
transform 1 0 38548 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_402
timestamp 1607721120
transform 1 0 38088 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_398
timestamp 1607721120
transform 1 0 37720 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1262__B
timestamp 1607721120
transform 1 0 38364 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1401__D
timestamp 1607721120
transform 1 0 38732 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1240__A
timestamp 1607721120
transform 1 0 37904 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1240_
timestamp 1607721120
transform 1 0 37076 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_11_423
timestamp 1607721120
transform 1 0 40020 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_419
timestamp 1607721120
transform 1 0 39652 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__A1
timestamp 1607721120
transform 1 0 40204 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1262__A
timestamp 1607721120
transform 1 0 39836 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1607721120
transform 1 0 40388 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1262_
timestamp 1607721120
transform 1 0 39008 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1232_
timestamp 1607721120
transform 1 0 40480 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_11_455
timestamp 1607721120
transform 1 0 42964 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_451
timestamp 1607721120
transform 1 0 42596 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_439
timestamp 1607721120
transform 1 0 41492 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_435
timestamp 1607721120
transform 1 0 41124 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__B
timestamp 1607721120
transform 1 0 41768 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__B
timestamp 1607721120
transform 1 0 42780 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1232__A
timestamp 1607721120
transform 1 0 41308 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0797_
timestamp 1607721120
transform 1 0 41952 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_11_476
timestamp 1607721120
transform 1 0 44896 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_461
timestamp 1607721120
transform 1 0 43516 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1396__D
timestamp 1607721120
transform 1 0 45080 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1234__A
timestamp 1607721120
transform 1 0 43332 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1139_
timestamp 1607721120
transform 1 0 43792 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_502
timestamp 1607721120
transform 1 0 47288 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_484
timestamp 1607721120
transform 1 0 45632 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_480
timestamp 1607721120
transform 1 0 45264 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__B1_N
timestamp 1607721120
transform 1 0 45816 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__A1
timestamp 1607721120
transform 1 0 45448 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1607721120
transform 1 0 46000 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_4  _1137_
timestamp 1607721120
transform 1 0 46092 0 1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_11_524
timestamp 1607721120
transform 1 0 49312 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_514
timestamp 1607721120
transform 1 0 48392 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_510
timestamp 1607721120
transform 1 0 48024 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_506
timestamp 1607721120
transform 1 0 47656 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1258__B
timestamp 1607721120
transform 1 0 48484 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__A
timestamp 1607721120
transform 1 0 47840 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__A1
timestamp 1607721120
transform 1 0 47472 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1258_
timestamp 1607721120
transform 1 0 48668 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_11_545
timestamp 1607721120
transform 1 0 51244 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_541
timestamp 1607721120
transform 1 0 50876 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_528
timestamp 1607721120
transform 1 0 49680 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1261__B1
timestamp 1607721120
transform 1 0 49864 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1261__A2
timestamp 1607721120
transform 1 0 51060 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__B
timestamp 1607721120
transform 1 0 51428 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1258__A
timestamp 1607721120
transform 1 0 49496 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _1103_
timestamp 1607721120
transform 1 0 50048 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_567
timestamp 1607721120
transform 1 0 53268 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_563
timestamp 1607721120
transform 1 0 52900 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_559
timestamp 1607721120
transform 1 0 52532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__C
timestamp 1607721120
transform 1 0 53084 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1133__A
timestamp 1607721120
transform 1 0 53452 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__B
timestamp 1607721120
transform 1 0 52716 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1607721120
transform 1 0 51612 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _1101_
timestamp 1607721120
transform 1 0 51704 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_586
timestamp 1607721120
transform 1 0 55016 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_582
timestamp 1607721120
transform 1 0 54648 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_571
timestamp 1607721120
transform 1 0 53636 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__B1
timestamp 1607721120
transform 1 0 55200 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__B
timestamp 1607721120
transform 1 0 53820 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__B
timestamp 1607721120
transform 1 0 54832 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1135_
timestamp 1607721120
transform 1 0 54004 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_4  _1131_
timestamp 1607721120
transform 1 0 55384 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_606
timestamp 1607721120
transform 1 0 56856 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_602
timestamp 1607721120
transform 1 0 56488 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__A1
timestamp 1607721120
transform 1 0 57040 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1397__D
timestamp 1607721120
transform 1 0 56672 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1607721120
transform 1 0 57224 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1117_
timestamp 1607721120
transform 1 0 57316 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_11_622
timestamp 1607721120
transform 1 0 58328 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_618
timestamp 1607721120
transform 1 0 57960 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__B
timestamp 1607721120
transform 1 0 58144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__A
timestamp 1607721120
transform 1 0 58604 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1399_
timestamp 1607721120
transform 1 0 58788 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_11_662
timestamp 1607721120
transform 1 0 62008 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_658
timestamp 1607721120
transform 1 0 61640 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_653
timestamp 1607721120
transform 1 0 61180 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_650
timestamp 1607721120
transform 1 0 60904 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_646
timestamp 1607721120
transform 1 0 60536 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1255__A1
timestamp 1607721120
transform 1 0 61824 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1255__A2
timestamp 1607721120
transform 1 0 60996 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0771_
timestamp 1607721120
transform 1 0 61272 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_672
timestamp 1607721120
transform 1 0 62928 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_670
timestamp 1607721120
transform 1 0 62744 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_666
timestamp 1607721120
transform 1 0 62376 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1399__CLK
timestamp 1607721120
transform 1 0 62192 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1607721120
transform 1 0 62836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1607721120
transform -1 0 63480 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3
timestamp 1607721120
transform 1 0 1380 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1607721120
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_4  _1283_
timestamp 1607721120
transform 1 0 2116 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_36
timestamp 1607721120
transform 1 0 4416 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_32
timestamp 1607721120
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_23
timestamp 1607721120
transform 1 0 3220 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1422__CLK
timestamp 1607721120
transform 1 0 4232 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1353__D
timestamp 1607721120
transform 1 0 4692 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1607721120
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _0945_
timestamp 1607721120
transform 1 0 4876 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_57
timestamp 1607721120
transform 1 0 6348 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_53
timestamp 1607721120
transform 1 0 5980 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__A1
timestamp 1607721120
transform 1 0 6164 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1279__B1
timestamp 1607721120
transform 1 0 6532 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1279_
timestamp 1607721120
transform 1 0 6716 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_88
timestamp 1607721120
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_84
timestamp 1607721120
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_81
timestamp 1607721120
transform 1 0 8556 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_77
timestamp 1607721120
transform 1 0 8188 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_73
timestamp 1607721120
transform 1 0 7820 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1281__B1
timestamp 1607721120
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1279__A2
timestamp 1607721120
transform 1 0 8004 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1203__C
timestamp 1607721120
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1203__A
timestamp 1607721120
transform 1 0 8648 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_110
timestamp 1607721120
transform 1 0 11224 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_105
timestamp 1607721120
transform 1 0 10764 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0941__A2
timestamp 1607721120
transform 1 0 11040 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1607721120
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1281_
timestamp 1607721120
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_4  _1208_
timestamp 1607721120
transform 1 0 11500 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_129
timestamp 1607721120
transform 1 0 12972 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_125
timestamp 1607721120
transform 1 0 12604 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_wb_clk_i_A
timestamp 1607721120
transform 1 0 13156 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__B1
timestamp 1607721120
transform 1 0 12788 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 13340 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _0874_
timestamp 1607721120
transform 1 0 13616 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_12_147
timestamp 1607721120
transform 1 0 14628 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_143
timestamp 1607721120
transform 1 0 14260 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__A
timestamp 1607721120
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__B1
timestamp 1607721120
transform 1 0 14444 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1607721120
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0866_
timestamp 1607721120
transform 1 0 15272 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_12_182
timestamp 1607721120
transform 1 0 17848 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_174
timestamp 1607721120
transform 1 0 17112 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_165
timestamp 1607721120
transform 1 0 16284 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_161
timestamp 1607721120
transform 1 0 15916 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__A
timestamp 1607721120
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1224__B
timestamp 1607721120
transform 1 0 16652 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_wb_clk_i
timestamp 1607721120
transform 1 0 16836 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _0861_
timestamp 1607721120
transform 1 0 17204 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_12_202
timestamp 1607721120
transform 1 0 19688 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_188
timestamp 1607721120
transform 1 0 18400 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1227__A2
timestamp 1607721120
transform 1 0 19872 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__B
timestamp 1607721120
transform 1 0 18216 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1227_
timestamp 1607721120
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_210
timestamp 1607721120
transform 1 0 20424 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_206
timestamp 1607721120
transform 1 0 20056 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1227__A1
timestamp 1607721120
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__B
timestamp 1607721120
transform 1 0 20240 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1607721120
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1214_
timestamp 1607721120
transform 1 0 20884 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_12_226
timestamp 1607721120
transform 1 0 21896 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_222
timestamp 1607721120
transform 1 0 21528 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1228__B
timestamp 1607721120
transform 1 0 22080 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1228__A
timestamp 1607721120
transform 1 0 21712 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_251
timestamp 1607721120
transform 1 0 24196 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_245
timestamp 1607721120
transform 1 0 23644 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_241
timestamp 1607721120
transform 1 0 23276 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_237
timestamp 1607721120
transform 1 0 22908 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_wb_clk_i_A
timestamp 1607721120
transform 1 0 23460 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1080__A
timestamp 1607721120
transform 1 0 24012 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__A
timestamp 1607721120
transform 1 0 23092 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1220_
timestamp 1607721120
transform 1 0 22264 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_12_271
timestamp 1607721120
transform 1 0 26036 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_267
timestamp 1607721120
transform 1 0 25668 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__A2
timestamp 1607721120
transform 1 0 24380 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__A2
timestamp 1607721120
transform 1 0 26220 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__A1
timestamp 1607721120
transform 1 0 25852 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1085_
timestamp 1607721120
transform 1 0 24564 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_292
timestamp 1607721120
transform 1 0 27968 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_288
timestamp 1607721120
transform 1 0 27600 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__A
timestamp 1607721120
transform 1 0 28152 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__A2
timestamp 1607721120
transform 1 0 27784 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1607721120
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1207_
timestamp 1607721120
transform 1 0 26496 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _0832_
timestamp 1607721120
transform 1 0 28336 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_12_312
timestamp 1607721120
transform 1 0 29808 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_308
timestamp 1607721120
transform 1 0 29440 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_303
timestamp 1607721120
transform 1 0 28980 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1077__B
timestamp 1607721120
transform 1 0 29624 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1077__A
timestamp 1607721120
transform 1 0 29256 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0813_
timestamp 1607721120
transform 1 0 29900 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_12_324
timestamp 1607721120
transform 1 0 30912 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_320
timestamp 1607721120
transform 1 0 30544 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1410__CLK
timestamp 1607721120
transform 1 0 31096 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__A
timestamp 1607721120
transform 1 0 30728 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_332
timestamp 1607721120
transform 1 0 31648 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_328
timestamp 1607721120
transform 1 0 31280 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1401__CLK
timestamp 1607721120
transform 1 0 31464 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1384__CLK
timestamp 1607721120
transform 1 0 31832 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_337
timestamp 1607721120
transform 1 0 32108 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1607721120
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1347_
timestamp 1607721120
transform 1 0 32292 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_12_353
timestamp 1607721120
transform 1 0 33580 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_350
timestamp 1607721120
transform 1 0 33304 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_346
timestamp 1607721120
transform 1 0 32936 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1366__D
timestamp 1607721120
transform 1 0 33396 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1245_
timestamp 1607721120
transform 1 0 33672 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_385
timestamp 1607721120
transform 1 0 36524 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_381
timestamp 1607721120
transform 1 0 36156 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_371
timestamp 1607721120
transform 1 0 35236 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_366
timestamp 1607721120
transform 1 0 34776 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1247__B1
timestamp 1607721120
transform 1 0 36708 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1248__B
timestamp 1607721120
transform 1 0 35052 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__B
timestamp 1607721120
transform 1 0 36340 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0943_
timestamp 1607721120
transform 1 0 35512 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_12_402
timestamp 1607721120
transform 1 0 38088 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_398
timestamp 1607721120
transform 1 0 37720 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_394
timestamp 1607721120
transform 1 0 37352 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_389
timestamp 1607721120
transform 1 0 36892 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1301__B
timestamp 1607721120
transform 1 0 38272 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1303__B
timestamp 1607721120
transform 1 0 37904 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1240__B
timestamp 1607721120
transform 1 0 37168 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1607721120
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1401_
timestamp 1607721120
transform 1 0 38456 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_12_431
timestamp 1607721120
transform 1 0 40756 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_425
timestamp 1607721120
transform 1 0 40204 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1232__B
timestamp 1607721120
transform 1 0 40572 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_453
timestamp 1607721120
transform 1 0 42780 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_449
timestamp 1607721120
transform 1 0 42412 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_438
timestamp 1607721120
transform 1 0 41400 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_435
timestamp 1607721120
transform 1 0 41124 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1360__CLK
timestamp 1607721120
transform 1 0 42964 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1263__A1
timestamp 1607721120
transform 1 0 41584 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1263__B1
timestamp 1607721120
transform 1 0 41216 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__A
timestamp 1607721120
transform 1 0 42596 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0791_
timestamp 1607721120
transform 1 0 41768 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_12_470
timestamp 1607721120
transform 1 0 44344 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_466
timestamp 1607721120
transform 1 0 43976 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_457
timestamp 1607721120
transform 1 0 43148 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__B1
timestamp 1607721120
transform 1 0 44160 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__A2
timestamp 1607721120
transform 1 0 44528 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1607721120
transform 1 0 43240 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1396_
timestamp 1607721120
transform 1 0 44712 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1234_
timestamp 1607721120
transform 1 0 43332 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_12_497
timestamp 1607721120
transform 1 0 46828 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_493
timestamp 1607721120
transform 1 0 46460 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1132__C
timestamp 1607721120
transform 1 0 46644 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__A2
timestamp 1607721120
transform 1 0 47012 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1264_
timestamp 1607721120
transform 1 0 47196 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_12_524
timestamp 1607721120
transform 1 0 49312 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_516
timestamp 1607721120
transform 1 0 48576 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_512
timestamp 1607721120
transform 1 0 48208 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_508
timestamp 1607721120
transform 1 0 47840 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__A
timestamp 1607721120
transform 1 0 48668 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__B
timestamp 1607721120
transform 1 0 48024 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1607721120
transform 1 0 48852 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0751_
timestamp 1607721120
transform 1 0 48944 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_546
timestamp 1607721120
transform 1 0 51336 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_528
timestamp 1607721120
transform 1 0 49680 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__D
timestamp 1607721120
transform 1 0 50048 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0745__A
timestamp 1607721120
transform 1 0 51520 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__A
timestamp 1607721120
transform 1 0 49496 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1261_
timestamp 1607721120
transform 1 0 50232 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_566
timestamp 1607721120
transform 1 0 53176 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_561
timestamp 1607721120
transform 1 0 52716 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_550
timestamp 1607721120
transform 1 0 51704 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__B1
timestamp 1607721120
transform 1 0 52992 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__D
timestamp 1607721120
transform 1 0 51888 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1133_
timestamp 1607721120
transform 1 0 53452 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _0698_
timestamp 1607721120
transform 1 0 52072 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_12_592
timestamp 1607721120
transform 1 0 55568 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_588
timestamp 1607721120
transform 1 0 55200 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_579
timestamp 1607721120
transform 1 0 54372 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_576
timestamp 1607721120
transform 1 0 54096 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_572
timestamp 1607721120
transform 1 0 53728 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__A
timestamp 1607721120
transform 1 0 55384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__A
timestamp 1607721120
transform 1 0 54188 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1607721120
transform 1 0 54464 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0736_
timestamp 1607721120
transform 1 0 54556 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__A2
timestamp 1607721120
transform 1 0 55936 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1397_
timestamp 1607721120
transform 1 0 56120 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_12_636
timestamp 1607721120
transform 1 0 59616 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_632
timestamp 1607721120
transform 1 0 59248 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_621
timestamp 1607721120
transform 1 0 58236 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_617
timestamp 1607721120
transform 1 0 57868 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__A
timestamp 1607721120
transform 1 0 59800 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__B1
timestamp 1607721120
transform 1 0 58052 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1130__C1
timestamp 1607721120
transform 1 0 58420 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1399__D
timestamp 1607721120
transform 1 0 59432 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1123_
timestamp 1607721120
transform 1 0 58604 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_12_662
timestamp 1607721120
transform 1 0 62008 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_658
timestamp 1607721120
transform 1 0 61640 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_654
timestamp 1607721120
transform 1 0 61272 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_640
timestamp 1607721120
transform 1 0 59984 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__A
timestamp 1607721120
transform 1 0 61824 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1255__B1
timestamp 1607721120
transform 1 0 61456 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1607721120
transform 1 0 60076 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1255_
timestamp 1607721120
transform 1 0 60168 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_674
timestamp 1607721120
transform 1 0 63112 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1607721120
transform -1 0 63480 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1607721120
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1607721120
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_22
timestamp 1607721120
transform 1 0 3128 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_15
timestamp 1607721120
transform 1 0 2484 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1607721120
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1607721120
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1607721120
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1267_
timestamp 1607721120
transform 1 0 2760 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_32
timestamp 1607721120
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1607721120
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_26
timestamp 1607721120
transform 1 0 3496 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1351__CLK
timestamp 1607721120
transform 1 0 3680 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1267__A
timestamp 1607721120
transform 1 0 3312 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1351__D
timestamp 1607721120
transform 1 0 4232 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1607721120
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1353_
timestamp 1607721120
transform 1 0 4416 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1351_
timestamp 1607721120
transform 1 0 3864 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_14_55
timestamp 1607721120
transform 1 0 6164 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1607721120
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_53
timestamp 1607721120
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_49
timestamp 1607721120
transform 1 0 5612 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1357__CLK
timestamp 1607721120
transform 1 0 6348 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1353__CLK
timestamp 1607721120
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1352__CLK
timestamp 1607721120
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_59
timestamp 1607721120
transform 1 0 6532 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1273__A1
timestamp 1607721120
transform 1 0 6716 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1352__D
timestamp 1607721120
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1607721120
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1352_
timestamp 1607721120
transform 1 0 6808 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__a21o_4  _1277_
timestamp 1607721120
transform 1 0 6900 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_75
timestamp 1607721120
transform 1 0 8004 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_83
timestamp 1607721120
transform 1 0 8740 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_79
timestamp 1607721120
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_81
timestamp 1607721120
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1277__A1
timestamp 1607721120
transform 1 0 8556 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1277__B1
timestamp 1607721120
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1277__A2
timestamp 1607721120
transform 1 0 8188 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_88
timestamp 1607721120
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_85
timestamp 1607721120
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__A
timestamp 1607721120
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__A
timestamp 1607721120
transform 1 0 9108 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__B
timestamp 1607721120
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0888_
timestamp 1607721120
transform 1 0 9292 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_14_100
timestamp 1607721120
transform 1 0 10304 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_100
timestamp 1607721120
transform 1 0 10304 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_96
timestamp 1607721120
transform 1 0 9936 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1281__A1
timestamp 1607721120
transform 1 0 10488 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__B
timestamp 1607721120
transform 1 0 10120 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1607721120
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0899_
timestamp 1607721120
transform 1 0 9660 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_14_110
timestamp 1607721120
transform 1 0 11224 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_104
timestamp 1607721120
transform 1 0 10672 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_114
timestamp 1607721120
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_104
timestamp 1607721120
transform 1 0 10672 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0905__A
timestamp 1607721120
transform 1 0 10764 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0905__B
timestamp 1607721120
transform 1 0 11040 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0905_
timestamp 1607721120
transform 1 0 10948 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_4  _1357_
timestamp 1607721120
transform 1 0 11408 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_13_118
timestamp 1607721120
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1271__A1
timestamp 1607721120
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1357__D
timestamp 1607721120
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1607721120
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_135
timestamp 1607721120
transform 1 0 13524 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_131
timestamp 1607721120
transform 1 0 13156 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_135
timestamp 1607721120
transform 1 0 13524 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1269__B1
timestamp 1607721120
transform 1 0 13340 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1269__A2
timestamp 1607721120
transform 1 0 13708 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1269_
timestamp 1607721120
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_140
timestamp 1607721120
transform 1 0 13984 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_139
timestamp 1607721120
transform 1 0 13892 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1269__A1
timestamp 1607721120
transform 1 0 14076 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__C
timestamp 1607721120
transform 1 0 13800 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_144
timestamp 1607721120
transform 1 0 14352 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_143
timestamp 1607721120
transform 1 0 14260 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__A
timestamp 1607721120
transform 1 0 14536 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__A
timestamp 1607721120
transform 1 0 14536 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__D
timestamp 1607721120
transform 1 0 14168 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_148
timestamp 1607721120
transform 1 0 14720 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_148
timestamp 1607721120
transform 1 0 14720 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0875__A
timestamp 1607721120
transform 1 0 14904 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__A
timestamp 1607721120
transform 1 0 14904 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_152
timestamp 1607721120
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_155
timestamp 1607721120
transform 1 0 15364 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_wb_clk_i
timestamp 1607721120
transform 1 0 15088 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1607721120
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0947_
timestamp 1607721120
transform 1 0 15456 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0846_
timestamp 1607721120
transform 1 0 15272 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_158
timestamp 1607721120
transform 1 0 15640 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_166
timestamp 1607721120
transform 1 0 16376 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_162
timestamp 1607721120
transform 1 0 16008 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_164
timestamp 1607721120
transform 1 0 16192 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_160
timestamp 1607721120
transform 1 0 15824 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_wb_clk_i_A
timestamp 1607721120
transform 1 0 16192 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__C
timestamp 1607721120
transform 1 0 16376 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__C
timestamp 1607721120
transform 1 0 15824 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0846__A
timestamp 1607721120
transform 1 0 16008 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_171
timestamp 1607721120
transform 1 0 16836 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_175
timestamp 1607721120
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__B
timestamp 1607721120
transform 1 0 16652 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1226_
timestamp 1607721120
transform 1 0 16928 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1218_
timestamp 1607721120
transform 1 0 16560 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_14_179
timestamp 1607721120
transform 1 0 17572 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_179
timestamp 1607721120
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__B
timestamp 1607721120
transform 1 0 17756 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__A
timestamp 1607721120
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__A
timestamp 1607721120
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_183
timestamp 1607721120
transform 1 0 17940 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_192
timestamp 1607721120
transform 1 0 18768 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_184
timestamp 1607721120
transform 1 0 18032 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__A
timestamp 1607721120
transform 1 0 18124 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1376__D
timestamp 1607721120
transform 1 0 18952 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1607721120
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0854_
timestamp 1607721120
transform 1 0 18124 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_13_196
timestamp 1607721120
transform 1 0 19136 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1227__B1
timestamp 1607721120
transform 1 0 19320 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1376_
timestamp 1607721120
transform 1 0 18308 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__a21o_4  _1225_
timestamp 1607721120
transform 1 0 19504 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_210
timestamp 1607721120
transform 1 0 20424 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_206
timestamp 1607721120
transform 1 0 20056 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_216
timestamp 1607721120
transform 1 0 20976 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_212
timestamp 1607721120
transform 1 0 20608 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__B1
timestamp 1607721120
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__A2
timestamp 1607721120
transform 1 0 20792 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__B
timestamp 1607721120
transform 1 0 20240 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1607721120
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_227
timestamp 1607721120
transform 1 0 21988 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_227
timestamp 1607721120
transform 1 0 21988 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__B
timestamp 1607721120
transform 1 0 21160 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1216_
timestamp 1607721120
transform 1 0 21344 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_4  _1229_
timestamp 1607721120
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_231
timestamp 1607721120
transform 1 0 22356 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_231
timestamp 1607721120
transform 1 0 22356 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1229__A1
timestamp 1607721120
transform 1 0 22540 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1229__B1
timestamp 1607721120
transform 1 0 22172 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1229__A2
timestamp 1607721120
transform 1 0 22540 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__A
timestamp 1607721120
transform 1 0 22172 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_238
timestamp 1607721120
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_wb_clk_i
timestamp 1607721120
transform 1 0 22724 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0821_
timestamp 1607721120
transform 1 0 22724 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_239
timestamp 1607721120
transform 1 0 23092 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_242
timestamp 1607721120
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0971__A
timestamp 1607721120
transform 1 0 23276 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__A
timestamp 1607721120
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_243
timestamp 1607721120
transform 1 0 23460 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_245
timestamp 1607721120
transform 1 0 23644 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__A
timestamp 1607721120
transform 1 0 23736 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__A1
timestamp 1607721120
transform 1 0 23828 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1607721120
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1302_
timestamp 1607721120
transform 1 0 23920 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0957_
timestamp 1607721120
transform 1 0 24012 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_256
timestamp 1607721120
transform 1 0 24656 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_252
timestamp 1607721120
transform 1 0 24288 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_256
timestamp 1607721120
transform 1 0 24656 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_252
timestamp 1607721120
transform 1 0 24288 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1302__A
timestamp 1607721120
transform 1 0 24472 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__B
timestamp 1607721120
transform 1 0 24840 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__A
timestamp 1607721120
transform 1 0 24472 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1405__D
timestamp 1607721120
transform 1 0 24840 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0847_
timestamp 1607721120
transform 1 0 25024 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_14_271
timestamp 1607721120
transform 1 0 26036 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_267
timestamp 1607721120
transform 1 0 25668 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__A
timestamp 1607721120
transform 1 0 26220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__B
timestamp 1607721120
transform 1 0 25852 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1405_
timestamp 1607721120
transform 1 0 25024 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_14_280
timestamp 1607721120
transform 1 0 26864 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_276
timestamp 1607721120
transform 1 0 26496 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_279
timestamp 1607721120
transform 1 0 26772 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__A2
timestamp 1607721120
transform 1 0 26956 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0827__A
timestamp 1607721120
transform 1 0 26956 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1607721120
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_283
timestamp 1607721120
transform 1 0 27140 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_283
timestamp 1607721120
transform 1 0 27140 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0827__B
timestamp 1607721120
transform 1 0 27324 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0827_
timestamp 1607721120
transform 1 0 27232 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _0819_
timestamp 1607721120
transform 1 0 27508 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_14_295
timestamp 1607721120
transform 1 0 28244 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_291
timestamp 1607721120
transform 1 0 27876 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_294
timestamp 1607721120
transform 1 0 28152 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__B1
timestamp 1607721120
transform 1 0 28060 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__B
timestamp 1607721120
transform 1 0 28336 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_302
timestamp 1607721120
transform 1 0 28888 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_298
timestamp 1607721120
transform 1 0 28520 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__A
timestamp 1607721120
transform 1 0 28428 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__B
timestamp 1607721120
transform 1 0 28704 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0840_
timestamp 1607721120
transform 1 0 28612 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_14_310
timestamp 1607721120
transform 1 0 29624 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_306
timestamp 1607721120
transform 1 0 29256 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_310
timestamp 1607721120
transform 1 0 29624 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_306
timestamp 1607721120
transform 1 0 29256 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1406__CLK
timestamp 1607721120
transform 1 0 29808 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__A
timestamp 1607721120
transform 1 0 29440 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__A
timestamp 1607721120
transform 1 0 29716 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1607721120
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_318
timestamp 1607721120
transform 1 0 30360 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_317
timestamp 1607721120
transform 1 0 30268 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0818_
timestamp 1607721120
transform 1 0 29992 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0697_
timestamp 1607721120
transform 1 0 29900 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_322
timestamp 1607721120
transform 1 0 30728 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_324
timestamp 1607721120
transform 1 0 30912 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1425__CLK
timestamp 1607721120
transform 1 0 30912 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__A
timestamp 1607721120
transform 1 0 30544 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0784_
timestamp 1607721120
transform 1 0 30544 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_326
timestamp 1607721120
transform 1 0 31096 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_328
timestamp 1607721120
transform 1 0 31280 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__A
timestamp 1607721120
transform 1 0 31280 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__A
timestamp 1607721120
transform 1 0 31096 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_330
timestamp 1607721120
transform 1 0 31464 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1251__A1
timestamp 1607721120
transform 1 0 31464 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_340
timestamp 1607721120
transform 1 0 32384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_334
timestamp 1607721120
transform 1 0 31832 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1348__B
timestamp 1607721120
transform 1 0 32568 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_wb_clk_i_A
timestamp 1607721120
transform 1 0 31648 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1607721120
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0964_
timestamp 1607721120
transform 1 0 32108 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 31648 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_14_344
timestamp 1607721120
transform 1 0 32752 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_364
timestamp 1607721120
transform 1 0 34592 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1251__B1
timestamp 1607721120
transform 1 0 32936 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1366_
timestamp 1607721120
transform 1 0 33120 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__a21o_4  _1251_
timestamp 1607721120
transform 1 0 33488 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_372
timestamp 1607721120
transform 1 0 35328 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_367
timestamp 1607721120
transform 1 0 34868 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_376
timestamp 1607721120
transform 1 0 35696 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_367
timestamp 1607721120
transform 1 0 34868 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1242__B
timestamp 1607721120
transform 1 0 35144 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1607721120
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1242_
timestamp 1607721120
transform 1 0 35052 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_14_387
timestamp 1607721120
transform 1 0 36708 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_380
timestamp 1607721120
transform 1 0 36064 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1247__A2
timestamp 1607721120
transform 1 0 36248 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1242__A
timestamp 1607721120
transform 1 0 35880 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1247_
timestamp 1607721120
transform 1 0 35604 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_4  _1243_
timestamp 1607721120
transform 1 0 36432 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_398
timestamp 1607721120
transform 1 0 37720 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_395
timestamp 1607721120
transform 1 0 37444 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_391
timestamp 1607721120
transform 1 0 37076 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_396
timestamp 1607721120
transform 1 0 37536 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1247__A1
timestamp 1607721120
transform 1 0 37260 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1243__B1
timestamp 1607721120
transform 1 0 36892 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1243__A2
timestamp 1607721120
transform 1 0 37720 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1607721120
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_402
timestamp 1607721120
transform 1 0 38088 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_408
timestamp 1607721120
transform 1 0 38640 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_400
timestamp 1607721120
transform 1 0 37904 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1243__A1
timestamp 1607721120
transform 1 0 37904 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1241__B1
timestamp 1607721120
transform 1 0 38088 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__A
timestamp 1607721120
transform 1 0 38824 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0703_
timestamp 1607721120
transform 1 0 38272 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _1241_
timestamp 1607721120
transform 1 0 38180 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_419
timestamp 1607721120
transform 1 0 39652 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_415
timestamp 1607721120
transform 1 0 39284 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_420
timestamp 1607721120
transform 1 0 39744 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_416
timestamp 1607721120
transform 1 0 39376 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_412
timestamp 1607721120
transform 1 0 39008 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1315__A2
timestamp 1607721120
transform 1 0 39836 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1241__A1
timestamp 1607721120
transform 1 0 39560 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__A
timestamp 1607721120
transform 1 0 39468 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1241__A2
timestamp 1607721120
transform 1 0 39192 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_433
timestamp 1607721120
transform 1 0 40940 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_423
timestamp 1607721120
transform 1 0 40020 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_428
timestamp 1607721120
transform 1 0 40480 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_424
timestamp 1607721120
transform 1 0 40112 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__A
timestamp 1607721120
transform 1 0 40204 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1607721120
transform 1 0 40388 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1238_
timestamp 1607721120
transform 1 0 40296 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_4  _1263_
timestamp 1607721120
transform 1 0 40756 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_437
timestamp 1607721120
transform 1 0 41308 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_443
timestamp 1607721120
transform 1 0 41860 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1233__B1
timestamp 1607721120
transform 1 0 41492 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__B
timestamp 1607721120
transform 1 0 41124 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0785__B
timestamp 1607721120
transform 1 0 42044 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0785_
timestamp 1607721120
transform 1 0 41676 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_14_456
timestamp 1607721120
transform 1 0 43056 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_452
timestamp 1607721120
transform 1 0 42688 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_448
timestamp 1607721120
transform 1 0 42320 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_447
timestamp 1607721120
transform 1 0 42228 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0785__A
timestamp 1607721120
transform 1 0 42504 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1263__A2
timestamp 1607721120
transform 1 0 42412 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1360__D
timestamp 1607721120
transform 1 0 42872 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1360_
timestamp 1607721120
transform 1 0 42596 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_14_463
timestamp 1607721120
transform 1 0 43700 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_459
timestamp 1607721120
transform 1 0 43332 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1386__CLK
timestamp 1607721120
transform 1 0 43516 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_wb_clk_i_A
timestamp 1607721120
transform 1 0 43884 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_wb_clk_i
timestamp 1607721120
transform 1 0 44068 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1607721120
transform 1 0 43240 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_477
timestamp 1607721120
transform 1 0 44988 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_474
timestamp 1607721120
transform 1 0 44712 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_470
timestamp 1607721120
transform 1 0 44344 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1235__B1
timestamp 1607721120
transform 1 0 44804 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1235__A2
timestamp 1607721120
transform 1 0 45172 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1235_
timestamp 1607721120
transform 1 0 44344 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_482
timestamp 1607721120
transform 1 0 45448 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_481
timestamp 1607721120
transform 1 0 45356 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1235__A1
timestamp 1607721120
transform 1 0 45540 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_489
timestamp 1607721120
transform 1 0 46092 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_486
timestamp 1607721120
transform 1 0 45816 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_489
timestamp 1607721120
transform 1 0 46092 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_wb_clk_i_A
timestamp 1607721120
transform 1 0 45908 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_wb_clk_i
timestamp 1607721120
transform 1 0 45724 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1607721120
transform 1 0 46000 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_493
timestamp 1607721120
transform 1 0 46460 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1185__A
timestamp 1607721120
transform 1 0 46460 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__A
timestamp 1607721120
transform 1 0 46276 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__A
timestamp 1607721120
transform 1 0 46644 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0753_
timestamp 1607721120
transform 1 0 46828 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0742_
timestamp 1607721120
transform 1 0 46644 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_499
timestamp 1607721120
transform 1 0 47012 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_501
timestamp 1607721120
transform 1 0 47196 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__A
timestamp 1607721120
transform 1 0 47196 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_511
timestamp 1607721120
transform 1 0 48116 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_503
timestamp 1607721120
transform 1 0 47380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_509
timestamp 1607721120
transform 1 0 47932 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_505
timestamp 1607721120
transform 1 0 47564 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__B
timestamp 1607721120
transform 1 0 47564 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__A
timestamp 1607721120
transform 1 0 47380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__A
timestamp 1607721120
transform 1 0 47748 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1359__D
timestamp 1607721120
transform 1 0 48300 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0733_
timestamp 1607721120
transform 1 0 47748 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_515
timestamp 1607721120
transform 1 0 48484 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__B1
timestamp 1607721120
transform 1 0 48668 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1607721120
transform 1 0 48852 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0758_
timestamp 1607721120
transform 1 0 48944 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_4  _1359_
timestamp 1607721120
transform 1 0 48024 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_14_531
timestamp 1607721120
transform 1 0 49956 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_527
timestamp 1607721120
transform 1 0 49588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_533
timestamp 1607721120
transform 1 0 50140 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_529
timestamp 1607721120
transform 1 0 49772 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__B
timestamp 1607721120
transform 1 0 49956 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__A
timestamp 1607721120
transform 1 0 50140 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__B
timestamp 1607721120
transform 1 0 49772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_538
timestamp 1607721120
transform 1 0 50600 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__A
timestamp 1607721120
transform 1 0 50784 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__C
timestamp 1607721120
transform 1 0 50324 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_wb_clk_i
timestamp 1607721120
transform 1 0 50324 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0714_
timestamp 1607721120
transform 1 0 50508 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_542
timestamp 1607721120
transform 1 0 50968 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_545
timestamp 1607721120
transform 1 0 51244 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_541
timestamp 1607721120
transform 1 0 50876 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0745__B
timestamp 1607721120
transform 1 0 51428 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__A
timestamp 1607721120
transform 1 0 51060 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0745_
timestamp 1607721120
transform 1 0 51152 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_14_555
timestamp 1607721120
transform 1 0 52164 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_551
timestamp 1607721120
transform 1 0 51796 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_569
timestamp 1607721120
transform 1 0 53452 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_wb_clk_i_A
timestamp 1607721120
transform 1 0 52348 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1361__D
timestamp 1607721120
transform 1 0 51980 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1607721120
transform 1 0 51612 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1361_
timestamp 1607721120
transform 1 0 51704 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__a21o_4  _1259_
timestamp 1607721120
transform 1 0 52532 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_575
timestamp 1607721120
transform 1 0 54004 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_571
timestamp 1607721120
transform 1 0 53636 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_577
timestamp 1607721120
transform 1 0 54188 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_573
timestamp 1607721120
transform 1 0 53820 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1359__CLK
timestamp 1607721120
transform 1 0 53820 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__A
timestamp 1607721120
transform 1 0 54280 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__A1
timestamp 1607721120
transform 1 0 54004 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__A2
timestamp 1607721120
transform 1 0 53636 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_581
timestamp 1607721120
transform 1 0 54556 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__A
timestamp 1607721120
transform 1 0 54372 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__B
timestamp 1607721120
transform 1 0 54740 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1607721120
transform 1 0 54464 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0727_
timestamp 1607721120
transform 1 0 54556 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _0726_
timestamp 1607721120
transform 1 0 54924 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_14_592
timestamp 1607721120
transform 1 0 55568 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_592
timestamp 1607721120
transform 1 0 55568 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_588
timestamp 1607721120
transform 1 0 55200 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__B
timestamp 1607721120
transform 1 0 55384 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_596
timestamp 1607721120
transform 1 0 55936 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_599
timestamp 1607721120
transform 1 0 56212 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__A
timestamp 1607721120
transform 1 0 55752 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__A
timestamp 1607721120
transform 1 0 55752 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__D
timestamp 1607721120
transform 1 0 56212 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0921_
timestamp 1607721120
transform 1 0 55936 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_603
timestamp 1607721120
transform 1 0 56580 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__B
timestamp 1607721120
transform 1 0 56764 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__A
timestamp 1607721120
transform 1 0 56396 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0715_
timestamp 1607721120
transform 1 0 56396 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_14_612
timestamp 1607721120
transform 1 0 57408 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_608
timestamp 1607721120
transform 1 0 57040 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1607721120
transform 1 0 57684 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_611
timestamp 1607721120
transform 1 0 57316 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_607
timestamp 1607721120
transform 1 0 56948 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__A
timestamp 1607721120
transform 1 0 57592 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1130__B1
timestamp 1607721120
transform 1 0 57776 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__B
timestamp 1607721120
transform 1 0 57224 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1607721120
transform 1 0 57224 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1130_
timestamp 1607721120
transform 1 0 57776 0 -1 10336
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_14_638
timestamp 1607721120
transform 1 0 59800 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_634
timestamp 1607721120
transform 1 0 59432 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_630
timestamp 1607721120
transform 1 0 59064 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_618
timestamp 1607721120
transform 1 0 57960 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1130__A1
timestamp 1607721120
transform 1 0 59616 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1130__A2
timestamp 1607721120
transform 1 0 59248 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1398__D
timestamp 1607721120
transform 1 0 58144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1398_
timestamp 1607721120
transform 1 0 58328 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_13_647
timestamp 1607721120
transform 1 0 60628 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_641
timestamp 1607721120
transform 1 0 60076 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1364__CLK
timestamp 1607721120
transform 1 0 60812 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1364__D
timestamp 1607721120
transform 1 0 60444 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1607721120
transform 1 0 60076 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_651
timestamp 1607721120
transform 1 0 60996 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1398__CLK
timestamp 1607721120
transform 1 0 61180 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_661
timestamp 1607721120
transform 1 0 61916 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_655
timestamp 1607721120
transform 1 0 61364 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1364_
timestamp 1607721120
transform 1 0 60168 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_14_673
timestamp 1607721120
transform 1 0 63020 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_672
timestamp 1607721120
transform 1 0 62928 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_667
timestamp 1607721120
transform 1 0 62468 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1607721120
transform 1 0 62836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1607721120
transform -1 0 63480 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1607721120
transform -1 0 63480 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1607721120
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1607721120
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1607721120
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_30
timestamp 1607721120
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_27
timestamp 1607721120
transform 1 0 3588 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1356__D
timestamp 1607721120
transform 1 0 3680 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1354__D
timestamp 1607721120
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1356_
timestamp 1607721120
transform 1 0 4232 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1607721120
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_53
timestamp 1607721120
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1354__CLK
timestamp 1607721120
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__C
timestamp 1607721120
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1607721120
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1273_
timestamp 1607721120
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_89
timestamp 1607721120
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_78
timestamp 1607721120
transform 1 0 8280 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_74
timestamp 1607721120
transform 1 0 7912 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__D
timestamp 1607721120
transform 1 0 8464 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__B
timestamp 1607721120
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__A
timestamp 1607721120
transform 1 0 8096 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0894_
timestamp 1607721120
transform 1 0 8648 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_15_114
timestamp 1607721120
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_101
timestamp 1607721120
transform 1 0 10396 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_97
timestamp 1607721120
transform 1 0 10028 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_93
timestamp 1607721120
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0883__A
timestamp 1607721120
transform 1 0 10764 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__A
timestamp 1607721120
transform 1 0 10212 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__B
timestamp 1607721120
transform 1 0 9844 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0883_
timestamp 1607721120
transform 1 0 10948 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_15_118
timestamp 1607721120
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1271__A2
timestamp 1607721120
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0883__B
timestamp 1607721120
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1607721120
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1358_
timestamp 1607721120
transform 1 0 12420 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_15_157
timestamp 1607721120
transform 1 0 15548 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_146
timestamp 1607721120
transform 1 0 14536 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_142
timestamp 1607721120
transform 1 0 14168 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__B
timestamp 1607721120
transform 1 0 14720 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__A
timestamp 1607721120
transform 1 0 15732 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__A
timestamp 1607721120
transform 1 0 14352 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0875_
timestamp 1607721120
transform 1 0 14904 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_15_161
timestamp 1607721120
transform 1 0 15916 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__B
timestamp 1607721120
transform 1 0 16100 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_169
timestamp 1607721120
transform 1 0 16652 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_165
timestamp 1607721120
transform 1 0 16284 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__D
timestamp 1607721120
transform 1 0 16468 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__A
timestamp 1607721120
transform 1 0 17020 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_179
timestamp 1607721120
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_175
timestamp 1607721120
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__B
timestamp 1607721120
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__B
timestamp 1607721120
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_195
timestamp 1607721120
transform 1 0 19044 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_191
timestamp 1607721120
transform 1 0 18676 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__A
timestamp 1607721120
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__A
timestamp 1607721120
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1607721120
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1375_
timestamp 1607721120
transform 1 0 19596 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1222_
timestamp 1607721120
transform 1 0 18032 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_15_224
timestamp 1607721120
transform 1 0 21712 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_220
timestamp 1607721120
transform 1 0 21344 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__B
timestamp 1607721120
transform 1 0 21896 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__A
timestamp 1607721120
transform 1 0 21528 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1325_
timestamp 1607721120
transform 1 0 22080 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_15_249
timestamp 1607721120
transform 1 0 24012 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_239
timestamp 1607721120
transform 1 0 23092 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_235
timestamp 1607721120
transform 1 0 22724 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__B
timestamp 1607721120
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1325__A
timestamp 1607721120
transform 1 0 22908 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__A
timestamp 1607721120
transform 1 0 24196 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1607721120
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0855_
timestamp 1607721120
transform 1 0 23644 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_269
timestamp 1607721120
transform 1 0 25852 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_265
timestamp 1607721120
transform 1 0 25484 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_253
timestamp 1607721120
transform 1 0 24380 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__A3
timestamp 1607721120
transform 1 0 26036 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__A
timestamp 1607721120
transform 1 0 24656 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__A
timestamp 1607721120
transform 1 0 25668 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0963_
timestamp 1607721120
transform 1 0 24840 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_4  _0962_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 26220 0 1 10336
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_15_294
timestamp 1607721120
transform 1 0 28152 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_290
timestamp 1607721120
transform 1 0 27784 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__B2
timestamp 1607721120
transform 1 0 28336 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1420__D
timestamp 1607721120
transform 1 0 27968 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_317
timestamp 1607721120
transform 1 0 30268 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_313
timestamp 1607721120
transform 1 0 29900 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_302
timestamp 1607721120
transform 1 0 28888 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_298
timestamp 1607721120
transform 1 0 28520 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1366__CLK
timestamp 1607721120
transform 1 0 30452 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__A
timestamp 1607721120
transform 1 0 28704 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0956__A
timestamp 1607721120
transform 1 0 30084 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1607721120
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0956_
timestamp 1607721120
transform 1 0 29256 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_15_335
timestamp 1607721120
transform 1 0 31924 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_329
timestamp 1607721120
transform 1 0 31372 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_325
timestamp 1607721120
transform 1 0 31004 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1313__B
timestamp 1607721120
transform 1 0 31740 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0889__A
timestamp 1607721120
transform 1 0 31188 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1368__D
timestamp 1607721120
transform 1 0 32108 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1368_
timestamp 1607721120
transform 1 0 32292 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1209_
timestamp 1607721120
transform 1 0 30636 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_362
timestamp 1607721120
transform 1 0 34408 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_358
timestamp 1607721120
transform 1 0 34040 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1251__A2
timestamp 1607721120
transform 1 0 34592 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1367__D
timestamp 1607721120
transform 1 0 34224 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_380
timestamp 1607721120
transform 1 0 36064 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_376
timestamp 1607721120
transform 1 0 35696 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_367
timestamp 1607721120
transform 1 0 34868 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1301__A
timestamp 1607721120
transform 1 0 36248 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1313__A
timestamp 1607721120
transform 1 0 35880 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1607721120
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1369_
timestamp 1607721120
transform 1 0 36432 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_4  _1313_
timestamp 1607721120
transform 1 0 35052 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_15_407
timestamp 1607721120
transform 1 0 38548 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_403
timestamp 1607721120
transform 1 0 38180 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__A
timestamp 1607721120
transform 1 0 38364 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1370__D
timestamp 1607721120
transform 1 0 38732 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1314_
timestamp 1607721120
transform 1 0 38916 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_15_428
timestamp 1607721120
transform 1 0 40480 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_426
timestamp 1607721120
transform 1 0 40296 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_422
timestamp 1607721120
transform 1 0 39928 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_418
timestamp 1607721120
transform 1 0 39560 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1314__B
timestamp 1607721120
transform 1 0 40112 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1314__A
timestamp 1607721120
transform 1 0 39744 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1607721120
transform 1 0 40388 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0918_
timestamp 1607721120
transform 1 0 40664 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_438
timestamp 1607721120
transform 1 0 41400 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_434
timestamp 1607721120
transform 1 0 41032 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1233__A2
timestamp 1607721120
transform 1 0 41584 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0918__A
timestamp 1607721120
transform 1 0 41216 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1374_
timestamp 1607721120
transform 1 0 41768 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_15_476
timestamp 1607721120
transform 1 0 44896 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_465
timestamp 1607721120
transform 1 0 43884 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_461
timestamp 1607721120
transform 1 0 43516 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1393__CLK
timestamp 1607721120
transform 1 0 44068 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__A
timestamp 1607721120
transform 1 0 43700 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1236__A
timestamp 1607721120
transform 1 0 45080 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1236_
timestamp 1607721120
transform 1 0 44252 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_15_484
timestamp 1607721120
transform 1 0 45632 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_480
timestamp 1607721120
transform 1 0 45264 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1373__D
timestamp 1607721120
transform 1 0 45448 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_489
timestamp 1607721120
transform 1 0 46092 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_wb_clk_i_A
timestamp 1607721120
transform 1 0 45816 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1607721120
transform 1 0 46000 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_494
timestamp 1607721120
transform 1 0 46552 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0741_
timestamp 1607721120
transform 1 0 46184 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_498
timestamp 1607721120
transform 1 0 46920 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__A
timestamp 1607721120
transform 1 0 46736 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__B
timestamp 1607721120
transform 1 0 47196 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_522
timestamp 1607721120
transform 1 0 49128 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_506
timestamp 1607721120
transform 1 0 47656 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__B
timestamp 1607721120
transform 1 0 49312 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__A
timestamp 1607721120
transform 1 0 47840 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_wb_clk_i
timestamp 1607721120
transform 1 0 47380 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_4  _1265_
timestamp 1607721120
transform 1 0 48024 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_545
timestamp 1607721120
transform 1 0 51244 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_541
timestamp 1607721120
transform 1 0 50876 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_537
timestamp 1607721120
transform 1 0 50508 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_526
timestamp 1607721120
transform 1 0 49496 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__A
timestamp 1607721120
transform 1 0 51060 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0704__A
timestamp 1607721120
transform 1 0 51428 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__A
timestamp 1607721120
transform 1 0 49680 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__B
timestamp 1607721120
transform 1 0 50692 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0772_
timestamp 1607721120
transform 1 0 49864 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_15_558
timestamp 1607721120
transform 1 0 52440 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_554
timestamp 1607721120
transform 1 0 52072 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0704__B
timestamp 1607721120
transform 1 0 52256 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1362__D
timestamp 1607721120
transform 1 0 52808 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1607721120
transform 1 0 51612 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1362_
timestamp 1607721120
transform 1 0 52992 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _0706_
timestamp 1607721120
transform 1 0 51704 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_589
timestamp 1607721120
transform 1 0 55292 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_583
timestamp 1607721120
transform 1 0 54740 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__B
timestamp 1607721120
transform 1 0 55108 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__C
timestamp 1607721120
transform 1 0 55660 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_607
timestamp 1607721120
transform 1 0 56948 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_602
timestamp 1607721120
transform 1 0 56488 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__A
timestamp 1607721120
transform 1 0 56764 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1607721120
transform 1 0 57224 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0722_
timestamp 1607721120
transform 1 0 57316 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _0721_
timestamp 1607721120
transform 1 0 55844 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_15_628
timestamp 1607721120
transform 1 0 58880 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_622
timestamp 1607721120
transform 1 0 58328 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_618
timestamp 1607721120
transform 1 0 57960 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__B1
timestamp 1607721120
transform 1 0 58696 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__A2
timestamp 1607721120
transform 1 0 59064 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__B
timestamp 1607721120
transform 1 0 58144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1365_
timestamp 1607721120
transform 1 0 59248 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_15_659
timestamp 1607721120
transform 1 0 61732 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_655
timestamp 1607721120
transform 1 0 61364 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_651
timestamp 1607721120
transform 1 0 60996 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1365__CLK
timestamp 1607721120
transform 1 0 61916 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1363__CLK
timestamp 1607721120
transform 1 0 61548 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1363__D
timestamp 1607721120
transform 1 0 61180 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_672
timestamp 1607721120
transform 1 0 62928 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_663
timestamp 1607721120
transform 1 0 62100 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1607721120
transform 1 0 62836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1607721120
transform -1 0 63480 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_15
timestamp 1607721120
transform 1 0 2484 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1607721120
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1355__CLK
timestamp 1607721120
transform 1 0 3036 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1607721120
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_36
timestamp 1607721120
transform 1 0 4416 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_32
timestamp 1607721120
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_23
timestamp 1607721120
transform 1 0 3220 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1356__CLK
timestamp 1607721120
transform 1 0 4232 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1607721120
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1354_
timestamp 1607721120
transform 1 0 4600 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_16_63
timestamp 1607721120
transform 1 0 6900 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_57
timestamp 1607721120
transform 1 0 6348 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1273__B1
timestamp 1607721120
transform 1 0 6716 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1273__A2
timestamp 1607721120
transform 1 0 7084 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0901_
timestamp 1607721120
transform 1 0 7268 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1607721120
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_86
timestamp 1607721120
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 1607721120
transform 1 0 8464 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_76
timestamp 1607721120
transform 1 0 8096 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__A
timestamp 1607721120
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__A
timestamp 1607721120
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__B
timestamp 1607721120
transform 1 0 8280 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_110
timestamp 1607721120
transform 1 0 11224 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_106
timestamp 1607721120
transform 1 0 10856 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_100
timestamp 1607721120
transform 1 0 10304 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0907__D
timestamp 1607721120
transform 1 0 10672 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__C
timestamp 1607721120
transform 1 0 11040 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1607721120
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1271_
timestamp 1607721120
transform 1 0 11500 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _0900_
timestamp 1607721120
transform 1 0 9660 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_16_133
timestamp 1607721120
transform 1 0 13340 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_129
timestamp 1607721120
transform 1 0 12972 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_125
timestamp 1607721120
transform 1 0 12604 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1271__B1
timestamp 1607721120
transform 1 0 13156 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1358__D
timestamp 1607721120
transform 1 0 12788 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0876_
timestamp 1607721120
transform 1 0 13616 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_149
timestamp 1607721120
transform 1 0 14812 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_145
timestamp 1607721120
transform 1 0 14444 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__A
timestamp 1607721120
transform 1 0 14628 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0875__B
timestamp 1607721120
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1607721120
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0868_
timestamp 1607721120
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_167
timestamp 1607721120
transform 1 0 16468 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_163
timestamp 1607721120
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_wb_clk_i_A
timestamp 1607721120
transform 1 0 16284 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_175
timestamp 1607721120
transform 1 0 17204 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_171
timestamp 1607721120
transform 1 0 16836 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__A1
timestamp 1607721120
transform 1 0 17020 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1328__B
timestamp 1607721120
transform 1 0 16652 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_179
timestamp 1607721120
transform 1 0 17572 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__A
timestamp 1607721120
transform 1 0 17664 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0862_
timestamp 1607721120
transform 1 0 17848 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_16_193
timestamp 1607721120
transform 1 0 18860 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_189
timestamp 1607721120
transform 1 0 18492 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__D
timestamp 1607721120
transform 1 0 18676 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__C
timestamp 1607721120
transform 1 0 19044 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0857_
timestamp 1607721120
transform 1 0 19228 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_228
timestamp 1607721120
transform 1 0 22080 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_224
timestamp 1607721120
transform 1 0 21712 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_210
timestamp 1607721120
transform 1 0 20424 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_206
timestamp 1607721120
transform 1 0 20056 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__D
timestamp 1607721120
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__C
timestamp 1607721120
transform 1 0 21896 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1375__D
timestamp 1607721120
transform 1 0 20240 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1607721120
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0849_
timestamp 1607721120
transform 1 0 20884 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1607721120
transform 1 0 24104 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_239
timestamp 1607721120
transform 1 0 23092 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_235
timestamp 1607721120
transform 1 0 22724 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__A1
timestamp 1607721120
transform 1 0 23276 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1325__B
timestamp 1607721120
transform 1 0 22264 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1323__B
timestamp 1607721120
transform 1 0 22908 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _0976_
timestamp 1607721120
transform 1 0 23460 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1607721120
transform 1 0 22448 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_271
timestamp 1607721120
transform 1 0 26036 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_267
timestamp 1607721120
transform 1 0 25668 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_254
timestamp 1607721120
transform 1 0 24472 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__C
timestamp 1607721120
transform 1 0 26220 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__A
timestamp 1607721120
transform 1 0 24288 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__B
timestamp 1607721120
transform 1 0 25852 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__B
timestamp 1607721120
transform 1 0 24656 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0980_
timestamp 1607721120
transform 1 0 24840 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_16_285
timestamp 1607721120
transform 1 0 27324 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_280
timestamp 1607721120
transform 1 0 26864 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__A1
timestamp 1607721120
transform 1 0 27140 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1607721120
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1420_
timestamp 1607721120
transform 1 0 27600 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _0977_
timestamp 1607721120
transform 1 0 26496 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_319
timestamp 1607721120
transform 1 0 30452 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_315
timestamp 1607721120
transform 1 0 30084 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_311
timestamp 1607721120
transform 1 0 29716 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_307
timestamp 1607721120
transform 1 0 29348 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1367__CLK
timestamp 1607721120
transform 1 0 30268 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1420__CLK
timestamp 1607721120
transform 1 0 29900 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0956__B
timestamp 1607721120
transform 1 0 29532 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_323
timestamp 1607721120
transform 1 0 30820 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__A
timestamp 1607721120
transform 1 0 30636 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0889_
timestamp 1607721120
transform 1 0 30912 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_332
timestamp 1607721120
transform 1 0 31648 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_328
timestamp 1607721120
transform 1 0 31280 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1295__B
timestamp 1607721120
transform 1 0 31464 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1348__A
timestamp 1607721120
transform 1 0 31832 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_337
timestamp 1607721120
transform 1 0 32108 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1607721120
transform 1 0 32016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1348_
timestamp 1607721120
transform 1 0 32384 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_16_351
timestamp 1607721120
transform 1 0 33396 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_347
timestamp 1607721120
transform 1 0 33028 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1317__A3
timestamp 1607721120
transform 1 0 33212 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1305__B1
timestamp 1607721120
transform 1 0 33580 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1367_
timestamp 1607721120
transform 1 0 33764 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_16_378
timestamp 1607721120
transform 1 0 35880 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_374
timestamp 1607721120
transform 1 0 35512 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__D
timestamp 1607721120
transform 1 0 35696 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__A
timestamp 1607721120
transform 1 0 36064 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1301_
timestamp 1607721120
transform 1 0 36248 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_16_398
timestamp 1607721120
transform 1 0 37720 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_393
timestamp 1607721120
transform 1 0 37260 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_389
timestamp 1607721120
transform 1 0 36892 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1303__A
timestamp 1607721120
transform 1 0 37444 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1369__D
timestamp 1607721120
transform 1 0 37076 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1607721120
transform 1 0 37628 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_402
timestamp 1607721120
transform 1 0 38088 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1316__B1
timestamp 1607721120
transform 1 0 37904 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1312__A
timestamp 1607721120
transform 1 0 38272 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1370_
timestamp 1607721120
transform 1 0 38456 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_16_429
timestamp 1607721120
transform 1 0 40572 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_425
timestamp 1607721120
transform 1 0 40204 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1312__B
timestamp 1607721120
transform 1 0 40388 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__C
timestamp 1607721120
transform 1 0 40940 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_455
timestamp 1607721120
transform 1 0 42964 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_451
timestamp 1607721120
transform 1 0 42596 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_447
timestamp 1607721120
transform 1 0 42228 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1233__A1
timestamp 1607721120
transform 1 0 42780 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1374__D
timestamp 1607721120
transform 1 0 42412 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1233_
timestamp 1607721120
transform 1 0 41124 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_472
timestamp 1607721120
transform 1 0 44528 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_467
timestamp 1607721120
transform 1 0 44068 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_463
timestamp 1607721120
transform 1 0 43700 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1394__CLK
timestamp 1607721120
transform 1 0 43884 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1236__B
timestamp 1607721120
transform 1 0 44344 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1607721120
transform 1 0 43240 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1373_
timestamp 1607721120
transform 1 0 44620 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _0786_
timestamp 1607721120
transform 1 0 43332 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_499
timestamp 1607721120
transform 1 0 47012 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_496
timestamp 1607721120
transform 1 0 46736 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_492
timestamp 1607721120
transform 1 0 46368 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__A
timestamp 1607721120
transform 1 0 47196 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__A
timestamp 1607721120
transform 1 0 46828 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_515
timestamp 1607721120
transform 1 0 48484 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_511
timestamp 1607721120
transform 1 0 48116 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_503
timestamp 1607721120
transform 1 0 47380 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__A1
timestamp 1607721120
transform 1 0 48300 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__A2
timestamp 1607721120
transform 1 0 48668 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1607721120
transform 1 0 48852 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0763_
timestamp 1607721120
transform 1 0 48944 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _0752_
timestamp 1607721120
transform 1 0 47472 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_16_547
timestamp 1607721120
transform 1 0 51428 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_542
timestamp 1607721120
transform 1 0 50968 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_533
timestamp 1607721120
transform 1 0 50140 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_527
timestamp 1607721120
transform 1 0 49588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1293__B1
timestamp 1607721120
transform 1 0 51244 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__B
timestamp 1607721120
transform 1 0 49956 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0779_
timestamp 1607721120
transform 1 0 50324 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_16_563
timestamp 1607721120
transform 1 0 52900 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_559
timestamp 1607721120
transform 1 0 52532 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1293__A2
timestamp 1607721120
transform 1 0 52716 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__A
timestamp 1607721120
transform 1 0 53084 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__A
timestamp 1607721120
transform 1 0 51704 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0709_
timestamp 1607721120
transform 1 0 53268 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _0704_
timestamp 1607721120
transform 1 0 51888 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_16_575
timestamp 1607721120
transform 1 0 54004 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_571
timestamp 1607721120
transform 1 0 53636 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__D
timestamp 1607721120
transform 1 0 54188 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__A
timestamp 1607721120
transform 1 0 53820 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_581
timestamp 1607721120
transform 1 0 54556 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_579
timestamp 1607721120
transform 1 0 54372 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__C
timestamp 1607721120
transform 1 0 54832 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1607721120
transform 1 0 54464 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0717_
timestamp 1607721120
transform 1 0 55016 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_16_593
timestamp 1607721120
transform 1 0 55660 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_614
timestamp 1607721120
transform 1 0 57592 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_610
timestamp 1607721120
transform 1 0 57224 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_598
timestamp 1607721120
transform 1 0 56120 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__B
timestamp 1607721120
transform 1 0 55936 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__A1
timestamp 1607721120
transform 1 0 57684 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0718_
timestamp 1607721120
transform 1 0 56396 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_637
timestamp 1607721120
transform 1 0 59708 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_633
timestamp 1607721120
transform 1 0 59340 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_617
timestamp 1607721120
transform 1 0 57868 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__A1
timestamp 1607721120
transform 1 0 59892 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__A
timestamp 1607721120
transform 1 0 58052 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1365__D
timestamp 1607721120
transform 1 0 59524 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1257_
timestamp 1607721120
transform 1 0 58236 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_661
timestamp 1607721120
transform 1 0 61916 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1607721120
transform 1 0 60076 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1363_
timestamp 1607721120
transform 1 0 60168 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_16_673
timestamp 1607721120
transform 1 0 63020 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1607721120
transform -1 0 63480 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_20
timestamp 1607721120
transform 1 0 2944 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_16
timestamp 1607721120
transform 1 0 2576 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_11
timestamp 1607721120
transform 1 0 2116 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_3
timestamp 1607721120
transform 1 0 1380 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1337__B
timestamp 1607721120
transform 1 0 2392 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1337__A
timestamp 1607721120
transform 1 0 2760 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1607721120
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1355_
timestamp 1607721120
transform 1 0 3036 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_17_45
timestamp 1607721120
transform 1 0 5244 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_40
timestamp 1607721120
transform 1 0 4784 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1275__B1
timestamp 1607721120
transform 1 0 5060 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_62
timestamp 1607721120
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_53
timestamp 1607721120
transform 1 0 5980 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_49
timestamp 1607721120
transform 1 0 5612 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1275__A1
timestamp 1607721120
transform 1 0 5796 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1275__A2
timestamp 1607721120
transform 1 0 5428 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0891__D
timestamp 1607721120
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__B
timestamp 1607721120
transform 1 0 7084 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1607721120
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0896_
timestamp 1607721120
transform 1 0 7268 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_91
timestamp 1607721120
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_80
timestamp 1607721120
transform 1 0 8464 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_76
timestamp 1607721120
transform 1 0 8096 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0891__B
timestamp 1607721120
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__A
timestamp 1607721120
transform 1 0 8280 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0895_
timestamp 1607721120
transform 1 0 8832 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_17_114
timestamp 1607721120
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_101
timestamp 1607721120
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_95
timestamp 1607721120
transform 1 0 9844 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__B
timestamp 1607721120
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0907__B
timestamp 1607721120
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__A
timestamp 1607721120
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _1205_
timestamp 1607721120
transform 1 0 10764 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_136
timestamp 1607721120
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_123
timestamp 1607721120
transform 1 0 12420 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_118
timestamp 1607721120
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0907__C
timestamp 1607721120
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__B
timestamp 1607721120
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0879__A
timestamp 1607721120
transform 1 0 12604 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1607721120
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1204_
timestamp 1607721120
transform 1 0 12788 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_155
timestamp 1607721120
transform 1 0 15364 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_151
timestamp 1607721120
transform 1 0 14996 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_140
timestamp 1607721120
transform 1 0 13984 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1333__A
timestamp 1607721120
transform 1 0 15548 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1335__B1
timestamp 1607721120
transform 1 0 14168 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__B
timestamp 1607721120
transform 1 0 13800 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__B
timestamp 1607721120
transform 1 0 15180 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0867_
timestamp 1607721120
transform 1 0 14352 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0845_
timestamp 1607721120
transform 1 0 15732 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_179
timestamp 1607721120
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_175
timestamp 1607721120
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_167
timestamp 1607721120
transform 1 0 16468 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_163
timestamp 1607721120
transform 1 0 16100 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1328__A
timestamp 1607721120
transform 1 0 16652 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1213__A
timestamp 1607721120
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__B
timestamp 1607721120
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__A
timestamp 1607721120
transform 1 0 16284 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1213_
timestamp 1607721120
transform 1 0 16836 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_199
timestamp 1607721120
transform 1 0 19412 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_194
timestamp 1607721120
transform 1 0 18952 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_184
timestamp 1607721120
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__A
timestamp 1607721120
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1607721120
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1377_
timestamp 1607721120
transform 1 0 19688 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _0856_
timestamp 1607721120
transform 1 0 18308 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_17_226
timestamp 1607721120
transform 1 0 21896 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_221
timestamp 1607721120
transform 1 0 21436 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__A2
timestamp 1607721120
transform 1 0 21712 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_236
timestamp 1607721120
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0848_
timestamp 1607721120
transform 1 0 22172 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_17_240
timestamp 1607721120
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1323__A
timestamp 1607721120
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0848__B
timestamp 1607721120
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1607721120
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_249
timestamp 1607721120
transform 1 0 24012 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_245
timestamp 1607721120
transform 1 0 23644 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1323__C
timestamp 1607721120
transform 1 0 23828 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _0979_
timestamp 1607721120
transform 1 0 24104 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_17_262
timestamp 1607721120
transform 1 0 25208 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_257
timestamp 1607721120
transform 1 0 24748 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__A
timestamp 1607721120
transform 1 0 25024 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1418_
timestamp 1607721120
transform 1 0 25484 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_17_296
timestamp 1607721120
transform 1 0 28336 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_288
timestamp 1607721120
transform 1 0 27600 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_284
timestamp 1607721120
transform 1 0 27232 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0969__B1
timestamp 1607721120
transform 1 0 27784 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0969__A2_N
timestamp 1607721120
transform 1 0 27416 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0953_
timestamp 1607721120
transform 1 0 27968 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_317
timestamp 1607721120
transform 1 0 30268 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_313
timestamp 1607721120
transform 1 0 29900 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_300
timestamp 1607721120
transform 1 0 28704 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__A
timestamp 1607721120
transform 1 0 30452 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__B
timestamp 1607721120
transform 1 0 28980 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__A
timestamp 1607721120
transform 1 0 30084 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0953__A
timestamp 1607721120
transform 1 0 28520 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1607721120
transform 1 0 29164 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0955_
timestamp 1607721120
transform 1 0 29256 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_17_340
timestamp 1607721120
transform 1 0 32384 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_329
timestamp 1607721120
transform 1 0 31372 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_325
timestamp 1607721120
transform 1 0 31004 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1295__A
timestamp 1607721120
transform 1 0 31556 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1249__A
timestamp 1607721120
transform 1 0 31188 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__B
timestamp 1607721120
transform 1 0 32568 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1295_
timestamp 1607721120
transform 1 0 31740 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1249_
timestamp 1607721120
transform 1 0 30636 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_363
timestamp 1607721120
transform 1 0 34500 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_357
timestamp 1607721120
transform 1 0 33948 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_344
timestamp 1607721120
transform 1 0 32752 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1297__C
timestamp 1607721120
transform 1 0 32936 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1305__C1
timestamp 1607721120
transform 1 0 34316 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1297_
timestamp 1607721120
transform 1 0 33120 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_385
timestamp 1607721120
transform 1 0 36524 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_371
timestamp 1607721120
transform 1 0 35236 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_367
timestamp 1607721120
transform 1 0 34868 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1305__A1
timestamp 1607721120
transform 1 0 35052 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__C
timestamp 1607721120
transform 1 0 35512 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__B
timestamp 1607721120
transform 1 0 36708 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1607721120
transform 1 0 34776 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1304_
timestamp 1607721120
transform 1 0 35696 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_406
timestamp 1607721120
transform 1 0 38456 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_400
timestamp 1607721120
transform 1 0 37904 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_389
timestamp 1607721120
transform 1 0 36892 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1304__A
timestamp 1607721120
transform 1 0 37076 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1315__B1
timestamp 1607721120
transform 1 0 38272 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1312_
timestamp 1607721120
transform 1 0 38640 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _1303_
timestamp 1607721120
transform 1 0 37260 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_17_433
timestamp 1607721120
transform 1 0 40940 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_428
timestamp 1607721120
transform 1 0 40480 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_421
timestamp 1607721120
transform 1 0 39836 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_415
timestamp 1607721120
transform 1 0 39284 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__D
timestamp 1607721120
transform 1 0 40204 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__B
timestamp 1607721120
transform 1 0 40756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__A
timestamp 1607721120
transform 1 0 39652 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1607721120
transform 1 0 40388 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_453
timestamp 1607721120
transform 1 0 42780 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_449
timestamp 1607721120
transform 1 0 42412 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__A1
timestamp 1607721120
transform 1 0 42964 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__A2
timestamp 1607721120
transform 1 0 42596 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__A
timestamp 1607721120
transform 1 0 41124 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1239_
timestamp 1607721120
transform 1 0 41308 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_464
timestamp 1607721120
transform 1 0 43792 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_461
timestamp 1607721120
transform 1 0 43516 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_457
timestamp 1607721120
transform 1 0 43148 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1396__CLK
timestamp 1607721120
transform 1 0 43608 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1372__D
timestamp 1607721120
transform 1 0 43976 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1237_
timestamp 1607721120
transform 1 0 44160 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_484
timestamp 1607721120
transform 1 0 45632 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_480
timestamp 1607721120
transform 1 0 45264 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1237__B1
timestamp 1607721120
transform 1 0 45816 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1237__A2
timestamp 1607721120
transform 1 0 45448 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_493
timestamp 1607721120
transform 1 0 46460 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_489
timestamp 1607721120
transform 1 0 46092 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1237__A1
timestamp 1607721120
transform 1 0 46276 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__B
timestamp 1607721120
transform 1 0 46644 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1607721120
transform 1 0 46000 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0764_
timestamp 1607721120
transform 1 0 46828 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_17_515
timestamp 1607721120
transform 1 0 48484 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_512
timestamp 1607721120
transform 1 0 48208 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_508
timestamp 1607721120
transform 1 0 47840 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_504
timestamp 1607721120
transform 1 0 47472 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1299__A
timestamp 1607721120
transform 1 0 48300 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__C
timestamp 1607721120
transform 1 0 48668 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__B
timestamp 1607721120
transform 1 0 47656 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1299_
timestamp 1607721120
transform 1 0 48852 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_17_545
timestamp 1607721120
transform 1 0 51244 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_541
timestamp 1607721120
transform 1 0 50876 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_530
timestamp 1607721120
transform 1 0 49864 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_526
timestamp 1607721120
transform 1 0 49496 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1299__B
timestamp 1607721120
transform 1 0 50048 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1293__A1
timestamp 1607721120
transform 1 0 51428 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__B
timestamp 1607721120
transform 1 0 49680 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__B
timestamp 1607721120
transform 1 0 51060 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0746_
timestamp 1607721120
transform 1 0 50232 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_17_567
timestamp 1607721120
transform 1 0 53268 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_563
timestamp 1607721120
transform 1 0 52900 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_550
timestamp 1607721120
transform 1 0 51704 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__B
timestamp 1607721120
transform 1 0 53452 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__D
timestamp 1607721120
transform 1 0 51888 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__A
timestamp 1607721120
transform 1 0 53084 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1607721120
transform 1 0 51612 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0710_
timestamp 1607721120
transform 1 0 52072 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_589
timestamp 1607721120
transform 1 0 55292 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_585
timestamp 1607721120
transform 1 0 54924 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_571
timestamp 1607721120
transform 1 0 53636 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__C
timestamp 1607721120
transform 1 0 53912 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__A
timestamp 1607721120
transform 1 0 55476 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__A
timestamp 1607721120
transform 1 0 55108 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0738_
timestamp 1607721120
transform 1 0 54096 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _0723_
timestamp 1607721120
transform 1 0 55660 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_606
timestamp 1607721120
transform 1 0 56856 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_602
timestamp 1607721120
transform 1 0 56488 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__C
timestamp 1607721120
transform 1 0 57040 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__A
timestamp 1607721120
transform 1 0 56672 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1607721120
transform 1 0 57224 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _0923_
timestamp 1607721120
transform 1 0 57316 0 1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_17_628
timestamp 1607721120
transform 1 0 58880 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_624
timestamp 1607721120
transform 1 0 58512 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__C
timestamp 1607721120
transform 1 0 59064 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__B
timestamp 1607721120
transform 1 0 58696 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1253_
timestamp 1607721120
transform 1 0 59248 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_656
timestamp 1607721120
transform 1 0 61456 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_652
timestamp 1607721120
transform 1 0 61088 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_648
timestamp 1607721120
transform 1 0 60720 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_644
timestamp 1607721120
transform 1 0 60352 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1253__A1
timestamp 1607721120
transform 1 0 61272 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1253__A2
timestamp 1607721120
transform 1 0 60904 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__B
timestamp 1607721120
transform 1 0 60536 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_672
timestamp 1607721120
transform 1 0 62928 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_668
timestamp 1607721120
transform 1 0 62560 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1607721120
transform 1 0 62836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1607721120
transform -1 0 63480 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_15
timestamp 1607721120
transform 1 0 2484 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1607721120
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1607721120
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1337_
timestamp 1607721120
transform 1 0 2576 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_18_32
timestamp 1607721120
transform 1 0 4048 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1607721120
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_23
timestamp 1607721120
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1355__D
timestamp 1607721120
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1607721120
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1275_
timestamp 1607721120
transform 1 0 4600 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_64
timestamp 1607721120
transform 1 0 6992 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_60
timestamp 1607721120
transform 1 0 6624 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_50
timestamp 1607721120
transform 1 0 5704 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1343__C1
timestamp 1607721120
transform 1 0 6440 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__D
timestamp 1607721120
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0891__C
timestamp 1607721120
transform 1 0 7176 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0891_
timestamp 1607721120
transform 1 0 7360 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1607721120
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_86
timestamp 1607721120
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_81
timestamp 1607721120
transform 1 0 8556 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_77
timestamp 1607721120
transform 1 0 8188 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1336__B2
timestamp 1607721120
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1336__B1
timestamp 1607721120
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0891__A
timestamp 1607721120
transform 1 0 8372 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_113
timestamp 1607721120
transform 1 0 11500 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_100
timestamp 1607721120
transform 1 0 10304 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_97
timestamp 1607721120
transform 1 0 10028 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_93
timestamp 1607721120
transform 1 0 9660 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1342__D
timestamp 1607721120
transform 1 0 10120 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__D
timestamp 1607721120
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1607721120
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0907_
timestamp 1607721120
transform 1 0 10672 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_129
timestamp 1607721120
transform 1 0 12972 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_125
timestamp 1607721120
transform 1 0 12604 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_117
timestamp 1607721120
transform 1 0 11868 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__A
timestamp 1607721120
transform 1 0 12052 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0884__D
timestamp 1607721120
transform 1 0 13156 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0884__C
timestamp 1607721120
transform 1 0 12788 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0907__A
timestamp 1607721120
transform 1 0 11684 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1335_
timestamp 1607721120
transform 1 0 13340 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0879_
timestamp 1607721120
transform 1 0 12236 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_149
timestamp 1607721120
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_145
timestamp 1607721120
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1335__A2
timestamp 1607721120
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1335__A1
timestamp 1607721120
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1607721120
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1333_
timestamp 1607721120
transform 1 0 15272 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_18_180
timestamp 1607721120
transform 1 0 17664 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_176
timestamp 1607721120
transform 1 0 17296 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_165
timestamp 1607721120
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_161
timestamp 1607721120
transform 1 0 15916 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1333__B
timestamp 1607721120
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1324__B1
timestamp 1607721120
transform 1 0 16468 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1321__A
timestamp 1607721120
transform 1 0 17848 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__A2
timestamp 1607721120
transform 1 0 17480 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1328_
timestamp 1607721120
transform 1 0 16652 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_18_202
timestamp 1607721120
transform 1 0 19688 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_187
timestamp 1607721120
transform 1 0 18308 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__B
timestamp 1607721120
transform 1 0 18676 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1377__D
timestamp 1607721120
transform 1 0 19964 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_wb_clk_i
timestamp 1607721120
transform 1 0 18032 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _0863_
timestamp 1607721120
transform 1 0 18860 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_227
timestamp 1607721120
transform 1 0 21988 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_213
timestamp 1607721120
transform 1 0 20700 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_207
timestamp 1607721120
transform 1 0 20148 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_wb_clk_i
timestamp 1607721120
transform 1 0 20424 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1607721120
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1215_
timestamp 1607721120
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_248
timestamp 1607721120
transform 1 0 23920 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_244
timestamp 1607721120
transform 1 0 23552 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_231
timestamp 1607721120
transform 1 0 22356 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0848__A
timestamp 1607721120
transform 1 0 23736 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1319__B
timestamp 1607721120
transform 1 0 22540 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__B1
timestamp 1607721120
transform 1 0 22172 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__B
timestamp 1607721120
transform 1 0 24104 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1323_
timestamp 1607721120
transform 1 0 22724 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_271
timestamp 1607721120
transform 1 0 26036 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_267
timestamp 1607721120
transform 1 0 25668 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_256
timestamp 1607721120
transform 1 0 24656 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_252
timestamp 1607721120
transform 1 0 24288 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__A
timestamp 1607721120
transform 1 0 24472 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0969__B2
timestamp 1607721120
transform 1 0 26220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1418__D
timestamp 1607721120
transform 1 0 25852 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _0973_
timestamp 1607721120
transform 1 0 24840 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_296
timestamp 1607721120
transform 1 0 28336 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_292
timestamp 1607721120
transform 1 0 27968 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0842__C
timestamp 1607721120
transform 1 0 28152 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1607721120
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0969_
timestamp 1607721120
transform 1 0 26496 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_319
timestamp 1607721120
transform 1 0 30452 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_311
timestamp 1607721120
transform 1 0 29716 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_307
timestamp 1607721120
transform 1 0 29348 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1418__CLK
timestamp 1607721120
transform 1 0 29900 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__B
timestamp 1607721120
transform 1 0 29532 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0969__A1_N
timestamp 1607721120
transform 1 0 28520 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0954_
timestamp 1607721120
transform 1 0 28704 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0952_
timestamp 1607721120
transform 1 0 30084 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_323
timestamp 1607721120
transform 1 0 30820 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__A
timestamp 1607721120
transform 1 0 30636 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1296__B
timestamp 1607721120
transform 1 0 31096 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_332
timestamp 1607721120
transform 1 0 31648 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_328
timestamp 1607721120
transform 1 0 31280 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__A
timestamp 1607721120
transform 1 0 31464 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1317__B1
timestamp 1607721120
transform 1 0 31832 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_337
timestamp 1607721120
transform 1 0 32108 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1607721120
transform 1 0 32016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0910_
timestamp 1607721120
transform 1 0 32292 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_18_350
timestamp 1607721120
transform 1 0 33304 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_346
timestamp 1607721120
transform 1 0 32936 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1297__B
timestamp 1607721120
transform 1 0 33488 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1297__A
timestamp 1607721120
transform 1 0 33120 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1305_
timestamp 1607721120
transform 1 0 33672 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_18_385
timestamp 1607721120
transform 1 0 36524 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_372
timestamp 1607721120
transform 1 0 35328 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_368
timestamp 1607721120
transform 1 0 34960 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1304__C
timestamp 1607721120
transform 1 0 35512 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1304__B
timestamp 1607721120
transform 1 0 36708 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1305__A2
timestamp 1607721120
transform 1 0 35144 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0915_
timestamp 1607721120
transform 1 0 35696 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_410
timestamp 1607721120
transform 1 0 38824 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_394
timestamp 1607721120
transform 1 0 37352 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_389
timestamp 1607721120
transform 1 0 36892 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1316__A1
timestamp 1607721120
transform 1 0 37168 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1607721120
transform 1 0 37628 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1315_
timestamp 1607721120
transform 1 0 37720 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_427
timestamp 1607721120
transform 1 0 40388 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_423
timestamp 1607721120
transform 1 0 40020 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_414
timestamp 1607721120
transform 1 0 39192 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1315__A1
timestamp 1607721120
transform 1 0 39008 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__C
timestamp 1607721120
transform 1 0 39468 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__B
timestamp 1607721120
transform 1 0 40204 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__D
timestamp 1607721120
transform 1 0 40572 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0799_
timestamp 1607721120
transform 1 0 40756 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0778_
timestamp 1607721120
transform 1 0 39652 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_452
timestamp 1607721120
transform 1 0 42688 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_448
timestamp 1607721120
transform 1 0 42320 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_444
timestamp 1607721120
transform 1 0 41952 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_440
timestamp 1607721120
transform 1 0 41584 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_wb_clk_i_A
timestamp 1607721120
transform 1 0 42964 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__B1
timestamp 1607721120
transform 1 0 42504 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__C
timestamp 1607721120
transform 1 0 42136 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__B
timestamp 1607721120
transform 1 0 41768 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_463
timestamp 1607721120
transform 1 0 43700 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_459
timestamp 1607721120
transform 1 0 43332 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_457
timestamp 1607721120
transform 1 0 43148 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1370__CLK
timestamp 1607721120
transform 1 0 43516 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1307__B
timestamp 1607721120
transform 1 0 43976 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1607721120
transform 1 0 43240 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1372_
timestamp 1607721120
transform 1 0 44160 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_18_502
timestamp 1607721120
transform 1 0 47288 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_491
timestamp 1607721120
transform 1 0 46276 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_487
timestamp 1607721120
transform 1 0 45908 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__A
timestamp 1607721120
transform 1 0 46460 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1350__B
timestamp 1607721120
transform 1 0 46092 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0759_
timestamp 1607721120
transform 1 0 46644 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_18_515
timestamp 1607721120
transform 1 0 48484 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_511
timestamp 1607721120
transform 1 0 48116 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_506
timestamp 1607721120
transform 1 0 47656 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__D
timestamp 1607721120
transform 1 0 47932 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__D
timestamp 1607721120
transform 1 0 47472 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__D
timestamp 1607721120
transform 1 0 48300 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__B
timestamp 1607721120
transform 1 0 48668 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1607721120
transform 1 0 48852 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0754_
timestamp 1607721120
transform 1 0 48944 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_18_537
timestamp 1607721120
transform 1 0 50508 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_533
timestamp 1607721120
transform 1 0 50140 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_527
timestamp 1607721120
transform 1 0 49588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__D
timestamp 1607721120
transform 1 0 49956 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__B
timestamp 1607721120
transform 1 0 50324 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1293_
timestamp 1607721120
transform 1 0 50692 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_563
timestamp 1607721120
transform 1 0 52900 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_559
timestamp 1607721120
transform 1 0 52532 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_555
timestamp 1607721120
transform 1 0 52164 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_551
timestamp 1607721120
transform 1 0 51796 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__A
timestamp 1607721120
transform 1 0 51980 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__C
timestamp 1607721120
transform 1 0 52716 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__B
timestamp 1607721120
transform 1 0 52348 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0737_
timestamp 1607721120
transform 1 0 53084 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_18_585
timestamp 1607721120
transform 1 0 54924 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_581
timestamp 1607721120
transform 1 0 54556 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_576
timestamp 1607721120
transform 1 0 54096 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_572
timestamp 1607721120
transform 1 0 53728 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1362__CLK
timestamp 1607721120
transform 1 0 53912 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__D
timestamp 1607721120
transform 1 0 54280 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__B
timestamp 1607721120
transform 1 0 54740 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1607721120
transform 1 0 54464 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0728_
timestamp 1607721120
transform 1 0 55108 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_604
timestamp 1607721120
transform 1 0 56672 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_600
timestamp 1607721120
transform 1 0 56304 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_596
timestamp 1607721120
transform 1 0 55936 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__B1
timestamp 1607721120
transform 1 0 56856 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__B
timestamp 1607721120
transform 1 0 56488 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__B
timestamp 1607721120
transform 1 0 56120 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_4  _0919_
timestamp 1607721120
transform 1 0 57040 0 -1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_18_639
timestamp 1607721120
transform 1 0 59892 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_633
timestamp 1607721120
transform 1 0 59340 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_629
timestamp 1607721120
transform 1 0 58972 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_625
timestamp 1607721120
transform 1 0 58604 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_621
timestamp 1607721120
transform 1 0 58236 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1253__B1
timestamp 1607721120
transform 1 0 59708 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0719__C
timestamp 1607721120
transform 1 0 59156 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0719__B
timestamp 1607721120
transform 1 0 58788 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__A2
timestamp 1607721120
transform 1 0 58420 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_653
timestamp 1607721120
transform 1 0 61180 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_649
timestamp 1607721120
transform 1 0 60812 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__A
timestamp 1607721120
transform 1 0 60996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1607721120
transform 1 0 60076 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0922_
timestamp 1607721120
transform 1 0 60168 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_18_673
timestamp 1607721120
transform 1 0 63020 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_665
timestamp 1607721120
transform 1 0 62284 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1607721120
transform -1 0 63480 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_11
timestamp 1607721120
transform 1 0 2116 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 1607721120
transform 1 0 1380 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_11
timestamp 1607721120
transform 1 0 2116 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1607721120
transform 1 0 1380 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1607721120
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1607721120
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_21
timestamp 1607721120
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1340__B
timestamp 1607721120
transform 1 0 2392 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1340_
timestamp 1607721120
transform 1 0 2392 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_20_16
timestamp 1607721120
transform 1 0 2576 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_32
timestamp 1607721120
transform 1 0 4048 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_28
timestamp 1607721120
transform 1 0 3680 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_25
timestamp 1607721120
transform 1 0 3404 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1332__B
timestamp 1607721120
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1340__A
timestamp 1607721120
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1607721120
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1332_
timestamp 1607721120
transform 1 0 3772 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_20_38
timestamp 1607721120
transform 1 0 4600 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_40
timestamp 1607721120
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_36
timestamp 1607721120
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0890__A
timestamp 1607721120
transform 1 0 4692 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1332__A
timestamp 1607721120
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0890__B
timestamp 1607721120
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0890_
timestamp 1607721120
transform 1 0 4876 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and3_4  _1339_
timestamp 1607721120
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_52
timestamp 1607721120
transform 1 0 5888 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_48
timestamp 1607721120
transform 1 0 5520 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1607721120
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_53
timestamp 1607721120
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1339__C
timestamp 1607721120
transform 1 0 6072 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1339__B
timestamp 1607721120
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1339__A
timestamp 1607721120
transform 1 0 5704 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_67
timestamp 1607721120
transform 1 0 7268 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_62
timestamp 1607721120
transform 1 0 6808 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1343__A2
timestamp 1607721120
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1343__A1
timestamp 1607721120
transform 1 0 7084 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1607721120
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1343_
timestamp 1607721120
transform 1 0 6256 0 -1 13600
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_20_78
timestamp 1607721120
transform 1 0 8280 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_74
timestamp 1607721120
transform 1 0 7912 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_70
timestamp 1607721120
transform 1 0 7544 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__C
timestamp 1607721120
transform 1 0 8096 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__C
timestamp 1607721120
transform 1 0 7452 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__B
timestamp 1607721120
transform 1 0 7728 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_86
timestamp 1607721120
transform 1 0 9016 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1607721120
transform 1 0 8648 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_88
timestamp 1607721120
transform 1 0 9200 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1336__A3
timestamp 1607721120
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1336__A2
timestamp 1607721120
transform 1 0 8464 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1341__A
timestamp 1607721120
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1336__A1
timestamp 1607721120
transform 1 0 9384 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _1336_
timestamp 1607721120
transform 1 0 7636 0 1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_20_100
timestamp 1607721120
transform 1 0 10304 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_92
timestamp 1607721120
transform 1 0 9568 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__B
timestamp 1607721120
transform 1 0 9752 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1607721120
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _1342_
timestamp 1607721120
transform 1 0 9936 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _0906_
timestamp 1607721120
transform 1 0 9660 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_20_110
timestamp 1607721120
transform 1 0 11224 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_104
timestamp 1607721120
transform 1 0 10672 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_109
timestamp 1607721120
transform 1 0 11132 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_105
timestamp 1607721120
transform 1 0 10764 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1342__C
timestamp 1607721120
transform 1 0 11316 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1342__B
timestamp 1607721120
transform 1 0 10948 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1342__A
timestamp 1607721120
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__C
timestamp 1607721120
transform 1 0 11040 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_114
timestamp 1607721120
transform 1 0 11592 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_113
timestamp 1607721120
transform 1 0 11500 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1341__B
timestamp 1607721120
transform 1 0 11408 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_118
timestamp 1607721120
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__A2
timestamp 1607721120
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__B1
timestamp 1607721120
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1607721120
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0884_
timestamp 1607721120
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_135
timestamp 1607721120
transform 1 0 13524 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_131
timestamp 1607721120
transform 1 0 13156 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_127
timestamp 1607721120
transform 1 0 12788 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_136
timestamp 1607721120
transform 1 0 13616 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_132
timestamp 1607721120
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0884__B
timestamp 1607721120
transform 1 0 13340 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0884__A
timestamp 1607721120
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__A1
timestamp 1607721120
transform 1 0 12972 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _0903_
timestamp 1607721120
transform 1 0 11684 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_145
timestamp 1607721120
transform 1 0 14444 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_142
timestamp 1607721120
transform 1 0 14168 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1329__C
timestamp 1607721120
transform 1 0 14352 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1327__A
timestamp 1607721120
transform 1 0 13984 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1329_
timestamp 1607721120
transform 1 0 14536 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1327_
timestamp 1607721120
transform 1 0 13800 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_20_149
timestamp 1607721120
transform 1 0 14812 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_155
timestamp 1607721120
transform 1 0 15364 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1329__B
timestamp 1607721120
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1329__A
timestamp 1607721120
transform 1 0 14628 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1607721120
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0880_
timestamp 1607721120
transform 1 0 15272 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_158
timestamp 1607721120
transform 1 0 15640 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_159
timestamp 1607721120
transform 1 0 15732 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0880__A
timestamp 1607721120
transform 1 0 15548 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_169
timestamp 1607721120
transform 1 0 16652 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_162
timestamp 1607721120
transform 1 0 16008 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1327__B
timestamp 1607721120
transform 1 0 16192 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1330__A2
timestamp 1607721120
transform 1 0 15824 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__B1
timestamp 1607721120
transform 1 0 15916 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_wb_clk_i
timestamp 1607721120
transform 1 0 16376 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_179
timestamp 1607721120
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_175
timestamp 1607721120
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1324__A1
timestamp 1607721120
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1324__C1
timestamp 1607721120
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1324_
timestamp 1607721120
transform 1 0 16744 0 -1 13600
box -38 -48 1326 592
use sky130_fd_sc_hd__a21o_4  _1219_
timestamp 1607721120
transform 1 0 16100 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_191
timestamp 1607721120
transform 1 0 18676 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_188
timestamp 1607721120
transform 1 0 18400 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_184
timestamp 1607721120
transform 1 0 18032 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_193
timestamp 1607721120
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_184
timestamp 1607721120
transform 1 0 18032 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1223__B1
timestamp 1607721120
transform 1 0 18492 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1607721120
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1321_
timestamp 1607721120
transform 1 0 18216 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_19_197
timestamp 1607721120
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__D
timestamp 1607721120
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__C
timestamp 1607721120
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1382_
timestamp 1607721120
transform 1 0 19596 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1320_
timestamp 1607721120
transform 1 0 18952 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_215
timestamp 1607721120
transform 1 0 20884 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_210
timestamp 1607721120
transform 1 0 20424 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_206
timestamp 1607721120
transform 1 0 20056 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1320__A1
timestamp 1607721120
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1382__D
timestamp 1607721120
transform 1 0 20240 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1607721120
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1607721120
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_227
timestamp 1607721120
transform 1 0 21988 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_224
timestamp 1607721120
transform 1 0 21712 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_220
timestamp 1607721120
transform 1 0 21344 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1320__A2
timestamp 1607721120
transform 1 0 21068 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1221__B1
timestamp 1607721120
transform 1 0 21804 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1319_
timestamp 1607721120
transform 1 0 22080 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_4  _1221_
timestamp 1607721120
transform 1 0 21344 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_236
timestamp 1607721120
transform 1 0 22816 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_232
timestamp 1607721120
transform 1 0 22448 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_239
timestamp 1607721120
transform 1 0 23092 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_235
timestamp 1607721120
transform 1 0 22724 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1221__A1
timestamp 1607721120
transform 1 0 23000 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1319__A
timestamp 1607721120
transform 1 0 22632 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1221__A2
timestamp 1607721120
transform 1 0 22908 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_248
timestamp 1607721120
transform 1 0 23920 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1326__A2
timestamp 1607721120
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1326__A1
timestamp 1607721120
transform 1 0 24104 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1607721120
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0970_
timestamp 1607721120
transform 1 0 23644 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _1326_
timestamp 1607721120
transform 1 0 23184 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_259
timestamp 1607721120
transform 1 0 24932 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_256
timestamp 1607721120
transform 1 0 24656 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_252
timestamp 1607721120
transform 1 0 24288 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_252
timestamp 1607721120
transform 1 0 24288 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0833__A
timestamp 1607721120
transform 1 0 25116 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1326__B1
timestamp 1607721120
transform 1 0 24472 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__B
timestamp 1607721120
transform 1 0 24748 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0974_
timestamp 1607721120
transform 1 0 24656 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_20_271
timestamp 1607721120
transform 1 0 26036 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_267
timestamp 1607721120
transform 1 0 25668 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_267
timestamp 1607721120
transform 1 0 25668 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_263
timestamp 1607721120
transform 1 0 25300 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__A
timestamp 1607721120
transform 1 0 25852 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1290__A
timestamp 1607721120
transform 1 0 25852 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__A
timestamp 1607721120
transform 1 0 25484 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0842__D
timestamp 1607721120
transform 1 0 26220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1290_
timestamp 1607721120
transform 1 0 25300 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1419_
timestamp 1607721120
transform 1 0 26036 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_20_280
timestamp 1607721120
transform 1 0 26864 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_276
timestamp 1607721120
transform 1 0 26496 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1419__D
timestamp 1607721120
transform 1 0 26680 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1607721120
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0842_
timestamp 1607721120
transform 1 0 27140 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_292
timestamp 1607721120
transform 1 0 27968 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_290
timestamp 1607721120
transform 1 0 27784 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0842__A
timestamp 1607721120
transform 1 0 27968 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_296
timestamp 1607721120
transform 1 0 28336 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_294
timestamp 1607721120
transform 1 0 28152 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0842__B
timestamp 1607721120
transform 1 0 28336 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__A
timestamp 1607721120
transform 1 0 28152 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_298
timestamp 1607721120
transform 1 0 28520 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__C
timestamp 1607721120
transform 1 0 28520 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__A
timestamp 1607721120
transform 1 0 28704 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0812_
timestamp 1607721120
transform 1 0 28704 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_304
timestamp 1607721120
transform 1 0 29072 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_302
timestamp 1607721120
transform 1 0 28888 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__D
timestamp 1607721120
transform 1 0 29256 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1607721120
transform 1 0 29164 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0968_
timestamp 1607721120
transform 1 0 29256 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_308
timestamp 1607721120
transform 1 0 29440 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_310
timestamp 1607721120
transform 1 0 29624 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__A
timestamp 1607721120
transform 1 0 29624 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_316
timestamp 1607721120
transform 1 0 30176 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_314
timestamp 1607721120
transform 1 0 29992 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__A
timestamp 1607721120
transform 1 0 30176 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__A
timestamp 1607721120
transform 1 0 29808 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0975_
timestamp 1607721120
transform 1 0 29808 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_318
timestamp 1607721120
transform 1 0 30360 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__B
timestamp 1607721120
transform 1 0 30452 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_328
timestamp 1607721120
transform 1 0 31280 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_321
timestamp 1607721120
transform 1 0 30636 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_326
timestamp 1607721120
transform 1 0 31096 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_322
timestamp 1607721120
transform 1 0 30728 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1308__B
timestamp 1607721120
transform 1 0 30544 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1306__C
timestamp 1607721120
transform 1 0 31464 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__A
timestamp 1607721120
transform 1 0 30912 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1308_
timestamp 1607721120
transform 1 0 31188 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0811_
timestamp 1607721120
transform 1 0 30912 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_332
timestamp 1607721120
transform 1 0 31648 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_338
timestamp 1607721120
transform 1 0 32200 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_334
timestamp 1607721120
transform 1 0 31832 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1306__B
timestamp 1607721120
transform 1 0 31832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1306__A
timestamp 1607721120
transform 1 0 32384 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1308__A
timestamp 1607721120
transform 1 0 32016 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1607721120
transform 1 0 32016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1306_
timestamp 1607721120
transform 1 0 32108 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _1298_
timestamp 1607721120
transform 1 0 32568 0 1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_20_350
timestamp 1607721120
transform 1 0 33304 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_346
timestamp 1607721120
transform 1 0 32936 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_360
timestamp 1607721120
transform 1 0 34224 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_356
timestamp 1607721120
transform 1 0 33856 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1298__A2
timestamp 1607721120
transform 1 0 33120 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1298__A1
timestamp 1607721120
transform 1 0 33488 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1317__A1
timestamp 1607721120
transform 1 0 34592 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1298__C1
timestamp 1607721120
transform 1 0 34040 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _1317_
timestamp 1607721120
transform 1 0 33672 0 -1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_20_375
timestamp 1607721120
transform 1 0 35604 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_371
timestamp 1607721120
transform 1 0 35236 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_374
timestamp 1607721120
transform 1 0 35512 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1317__B2
timestamp 1607721120
transform 1 0 35420 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1296__A
timestamp 1607721120
transform 1 0 35696 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1607721120
transform 1 0 34776 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1296_
timestamp 1607721120
transform 1 0 34868 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_20_388
timestamp 1607721120
transform 1 0 36800 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_378
timestamp 1607721120
transform 1 0 35880 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1309__D
timestamp 1607721120
transform 1 0 35788 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1349__B
timestamp 1607721120
transform 1 0 36064 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1349_
timestamp 1607721120
transform 1 0 35972 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_4  _1316_
timestamp 1607721120
transform 1 0 36248 0 1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_20_392
timestamp 1607721120
transform 1 0 37168 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__C
timestamp 1607721120
transform 1 0 37444 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1349__A
timestamp 1607721120
transform 1 0 36984 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_398
timestamp 1607721120
transform 1 0 37720 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_399
timestamp 1607721120
transform 1 0 37812 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__B
timestamp 1607721120
transform 1 0 38088 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1607721120
transform 1 0 37628 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0798_
timestamp 1607721120
transform 1 0 37996 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_20_408
timestamp 1607721120
transform 1 0 38640 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_408
timestamp 1607721120
transform 1 0 38640 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_404
timestamp 1607721120
transform 1 0 38272 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__D
timestamp 1607721120
transform 1 0 38456 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__C
timestamp 1607721120
transform 1 0 38824 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_415
timestamp 1607721120
transform 1 0 39284 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_412
timestamp 1607721120
transform 1 0 39008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_419
timestamp 1607721120
transform 1 0 39652 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__B
timestamp 1607721120
transform 1 0 39100 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0800_
timestamp 1607721120
transform 1 0 39376 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _0792_
timestamp 1607721120
transform 1 0 39008 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_20_429
timestamp 1607721120
transform 1 0 40572 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_425
timestamp 1607721120
transform 1 0 40204 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_423
timestamp 1607721120
transform 1 0 40020 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__C
timestamp 1607721120
transform 1 0 40204 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__A2
timestamp 1607721120
transform 1 0 40388 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__A
timestamp 1607721120
transform 1 0 39836 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1607721120
transform 1 0 40388 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0769_
timestamp 1607721120
transform 1 0 40480 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_432
timestamp 1607721120
transform 1 0 40848 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__D
timestamp 1607721120
transform 1 0 40756 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0788_
timestamp 1607721120
transform 1 0 40940 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_442
timestamp 1607721120
transform 1 0 41768 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_436
timestamp 1607721120
transform 1 0 41216 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__A
timestamp 1607721120
transform 1 0 41400 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__A
timestamp 1607721120
transform 1 0 41032 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1371__D
timestamp 1607721120
transform 1 0 41952 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_456
timestamp 1607721120
transform 1 0 43056 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_450
timestamp 1607721120
transform 1 0 42504 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_446
timestamp 1607721120
transform 1 0 42136 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__B
timestamp 1607721120
transform 1 0 42320 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_wb_clk_i
timestamp 1607721120
transform 1 0 42780 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1371_
timestamp 1607721120
transform 1 0 41584 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_20_466
timestamp 1607721120
transform 1 0 43976 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_463
timestamp 1607721120
transform 1 0 43700 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_459
timestamp 1607721120
transform 1 0 43332 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__A
timestamp 1607721120
transform 1 0 43884 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__B
timestamp 1607721120
transform 1 0 43516 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1607721120
transform 1 0 43240 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0780_
timestamp 1607721120
transform 1 0 43332 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_20_474
timestamp 1607721120
transform 1 0 44712 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_470
timestamp 1607721120
transform 1 0 44344 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_476
timestamp 1607721120
transform 1 0 44896 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_467
timestamp 1607721120
transform 1 0 44068 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1307__A
timestamp 1607721120
transform 1 0 44528 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__D
timestamp 1607721120
transform 1 0 44160 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1307_
timestamp 1607721120
transform 1 0 44252 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1350__C
timestamp 1607721120
transform 1 0 44988 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1350__A
timestamp 1607721120
transform 1 0 45172 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1350_
timestamp 1607721120
transform 1 0 45172 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_488
timestamp 1607721120
transform 1 0 46000 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_489
timestamp 1607721120
transform 1 0 46092 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_487
timestamp 1607721120
transform 1 0 45908 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_481
timestamp 1607721120
transform 1 0 45356 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_wb_clk_i
timestamp 1607721120
transform 1 0 45632 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1607721120
transform 1 0 46000 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_492
timestamp 1607721120
transform 1 0 46368 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_494
timestamp 1607721120
transform 1 0 46552 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__D
timestamp 1607721120
transform 1 0 46184 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__C
timestamp 1607721120
transform 1 0 46552 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__C
timestamp 1607721120
transform 1 0 46368 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__B
timestamp 1607721120
transform 1 0 46736 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0773_
timestamp 1607721120
transform 1 0 46736 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _0760_
timestamp 1607721120
transform 1 0 46920 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_507
timestamp 1607721120
transform 1 0 47748 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_503
timestamp 1607721120
transform 1 0 47380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_511
timestamp 1607721120
transform 1 0 48116 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_507
timestamp 1607721120
transform 1 0 47748 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__C
timestamp 1607721120
transform 1 0 47932 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__B
timestamp 1607721120
transform 1 0 47564 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__A
timestamp 1607721120
transform 1 0 47932 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_wb_clk_i
timestamp 1607721120
transform 1 0 48116 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_518
timestamp 1607721120
transform 1 0 48760 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_514
timestamp 1607721120
transform 1 0 48392 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__A
timestamp 1607721120
transform 1 0 48300 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__A
timestamp 1607721120
transform 1 0 48576 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1607721120
transform 1 0 48852 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0765_
timestamp 1607721120
transform 1 0 48944 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _0755_
timestamp 1607721120
transform 1 0 48484 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_524
timestamp 1607721120
transform 1 0 49312 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_536
timestamp 1607721120
transform 1 0 50416 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_533
timestamp 1607721120
transform 1 0 50140 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_529
timestamp 1607721120
transform 1 0 49772 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_528
timestamp 1607721120
transform 1 0 49680 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__B
timestamp 1607721120
transform 1 0 49864 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__A
timestamp 1607721120
transform 1 0 49496 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__B
timestamp 1607721120
transform 1 0 50232 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0747_
timestamp 1607721120
transform 1 0 50048 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_545
timestamp 1607721120
transform 1 0 51244 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_541
timestamp 1607721120
transform 1 0 50876 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__C
timestamp 1607721120
transform 1 0 51428 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__A
timestamp 1607721120
transform 1 0 51060 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1300_
timestamp 1607721120
transform 1 0 50508 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_553
timestamp 1607721120
transform 1 0 51980 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_549
timestamp 1607721120
transform 1 0 51612 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1292__A
timestamp 1607721120
transform 1 0 52164 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1300__A1
timestamp 1607721120
transform 1 0 51796 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1607721120
transform 1 0 51612 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1292_
timestamp 1607721120
transform 1 0 51704 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_20_561
timestamp 1607721120
transform 1 0 52716 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_561
timestamp 1607721120
transform 1 0 52716 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_557
timestamp 1607721120
transform 1 0 52348 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1300__A2
timestamp 1607721120
transform 1 0 52900 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1292__B
timestamp 1607721120
transform 1 0 52900 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__A
timestamp 1607721120
transform 1 0 52532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0708_
timestamp 1607721120
transform 1 0 52348 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_570
timestamp 1607721120
transform 1 0 53544 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_565
timestamp 1607721120
transform 1 0 53084 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_565
timestamp 1607721120
transform 1 0 53084 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__B
timestamp 1607721120
transform 1 0 53360 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1211_
timestamp 1607721120
transform 1 0 53268 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_20_574
timestamp 1607721120
transform 1 0 53912 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_578
timestamp 1607721120
transform 1 0 54280 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_574
timestamp 1607721120
transform 1 0 53912 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_wb_clk_i_A
timestamp 1607721120
transform 1 0 53728 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__A
timestamp 1607721120
transform 1 0 54464 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__A
timestamp 1607721120
transform 1 0 54096 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1607721120
transform 1 0 54464 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_589
timestamp 1607721120
transform 1 0 55292 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_585
timestamp 1607721120
transform 1 0 54924 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__A
timestamp 1607721120
transform 1 0 55108 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0731_
timestamp 1607721120
transform 1 0 54556 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__and3_4  _0729_
timestamp 1607721120
transform 1 0 54648 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_593
timestamp 1607721120
transform 1 0 55660 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_591
timestamp 1607721120
transform 1 0 55476 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__B
timestamp 1607721120
transform 1 0 55476 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__D
timestamp 1607721120
transform 1 0 55660 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_603
timestamp 1607721120
transform 1 0 56580 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_599
timestamp 1607721120
transform 1 0 56212 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_595
timestamp 1607721120
transform 1 0 55844 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1383__CLK
timestamp 1607721120
transform 1 0 56764 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__C
timestamp 1607721120
transform 1 0 56396 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1383__D
timestamp 1607721120
transform 1 0 56028 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_613
timestamp 1607721120
transform 1 0 57500 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_615
timestamp 1607721120
transform 1 0 57684 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_607
timestamp 1607721120
transform 1 0 56948 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1455__CLK
timestamp 1607721120
transform 1 0 57684 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1607721120
transform 1 0 57224 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0743_
timestamp 1607721120
transform 1 0 57316 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1383_
timestamp 1607721120
transform 1 0 55752 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_20_617
timestamp 1607721120
transform 1 0 57868 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_623
timestamp 1607721120
transform 1 0 58420 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_619
timestamp 1607721120
transform 1 0 58052 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1426__CLK
timestamp 1607721120
transform 1 0 58052 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__A
timestamp 1607721120
transform 1 0 57868 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0719__A
timestamp 1607721120
transform 1 0 58236 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0719_
timestamp 1607721120
transform 1 0 58236 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_20_634
timestamp 1607721120
transform 1 0 59432 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_630
timestamp 1607721120
transform 1 0 59064 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1426__D
timestamp 1607721120
transform 1 0 59248 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1426_
timestamp 1607721120
transform 1 0 58604 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_20_654
timestamp 1607721120
transform 1 0 61272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_642
timestamp 1607721120
transform 1 0 60168 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_640
timestamp 1607721120
transform 1 0 59984 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_656
timestamp 1607721120
transform 1 0 61456 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_644
timestamp 1607721120
transform 1 0 60352 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1607721120
transform 1 0 60076 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_674
timestamp 1607721120
transform 1 0 63112 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_666
timestamp 1607721120
transform 1 0 62376 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_672
timestamp 1607721120
transform 1 0 62928 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_668
timestamp 1607721120
transform 1 0 62560 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1607721120
transform 1 0 62836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1607721120
transform -1 0 63480 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1607721120
transform -1 0 63480 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1607721120
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1607721120
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1607721120
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_42
timestamp 1607721120
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_38
timestamp 1607721120
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_27
timestamp 1607721120
transform 1 0 3588 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1338__B
timestamp 1607721120
transform 1 0 3772 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1334__B
timestamp 1607721120
transform 1 0 5152 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1338__A
timestamp 1607721120
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1338_
timestamp 1607721120
transform 1 0 3956 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_21_53
timestamp 1607721120
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1334_
timestamp 1607721120
transform 1 0 5336 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1607721120
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__B
timestamp 1607721120
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__A
timestamp 1607721120
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1607721120
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_66
timestamp 1607721120
transform 1 0 7176 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_62
timestamp 1607721120
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1343__B1
timestamp 1607721120
transform 1 0 6992 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__A
timestamp 1607721120
transform 1 0 7360 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_83
timestamp 1607721120
transform 1 0 8740 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_79
timestamp 1607721120
transform 1 0 8372 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__A1
timestamp 1607721120
transform 1 0 8924 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__B1
timestamp 1607721120
transform 1 0 8556 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0972_
timestamp 1607721120
transform 1 0 9108 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and3_4  _0897_
timestamp 1607721120
transform 1 0 7544 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_114
timestamp 1607721120
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_102
timestamp 1607721120
transform 1 0 10488 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_98
timestamp 1607721120
transform 1 0 10120 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_94
timestamp 1607721120
transform 1 0 9752 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__A
timestamp 1607721120
transform 1 0 9936 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__B
timestamp 1607721120
transform 1 0 10580 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0908_
timestamp 1607721120
transform 1 0 10764 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_134
timestamp 1607721120
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_123
timestamp 1607721120
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1607721120
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1331__B
timestamp 1607721120
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1331__A
timestamp 1607721120
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1380__D
timestamp 1607721120
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1607721120
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1331_
timestamp 1607721120
transform 1 0 12604 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_156
timestamp 1607721120
transform 1 0 15456 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_138
timestamp 1607721120
transform 1 0 13800 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1330__C1
timestamp 1607721120
transform 1 0 15640 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__A
timestamp 1607721120
transform 1 0 13984 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1330_
timestamp 1607721120
transform 1 0 14168 0 1 13600
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_21_160
timestamp 1607721120
transform 1 0 15824 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1330__A1
timestamp 1607721120
transform 1 0 16008 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1289_
timestamp 1607721120
transform 1 0 16192 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_168
timestamp 1607721120
transform 1 0 16560 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_172
timestamp 1607721120
transform 1 0 16928 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1289__A
timestamp 1607721120
transform 1 0 16744 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1378__D
timestamp 1607721120
transform 1 0 17112 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_176
timestamp 1607721120
transform 1 0 17296 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_180
timestamp 1607721120
transform 1 0 17664 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1324__A2
timestamp 1607721120
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_200
timestamp 1607721120
transform 1 0 19504 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_196
timestamp 1607721120
transform 1 0 19136 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1320__B1
timestamp 1607721120
transform 1 0 19688 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1223__A2
timestamp 1607721120
transform 1 0 19320 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1607721120
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1322_
timestamp 1607721120
transform 1 0 19872 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_4  _1223_
timestamp 1607721120
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_215
timestamp 1607721120
transform 1 0 20884 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_211
timestamp 1607721120
transform 1 0 20516 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__B1
timestamp 1607721120
transform 1 0 21068 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1322__A
timestamp 1607721120
transform 1 0 20700 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1217_
timestamp 1607721120
transform 1 0 21252 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_231
timestamp 1607721120
transform 1 0 22356 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1379__D
timestamp 1607721120
transform 1 0 22540 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_235
timestamp 1607721120
transform 1 0 22724 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__A2
timestamp 1607721120
transform 1 0 22908 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_239
timestamp 1607721120
transform 1 0 23092 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__A1
timestamp 1607721120
transform 1 0 23276 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_243
timestamp 1607721120
transform 1 0 23460 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1607721120
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0978_
timestamp 1607721120
transform 1 0 23644 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_249
timestamp 1607721120
transform 1 0 24012 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__A
timestamp 1607721120
transform 1 0 24196 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_269
timestamp 1607721120
transform 1 0 25852 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_265
timestamp 1607721120
transform 1 0 25484 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_253
timestamp 1607721120
transform 1 0 24380 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__B
timestamp 1607721120
transform 1 0 26036 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0833__B
timestamp 1607721120
transform 1 0 24656 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0841__B
timestamp 1607721120
transform 1 0 25668 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0841_
timestamp 1607721120
transform 1 0 24840 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _0828_
timestamp 1607721120
transform 1 0 26220 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_21_284
timestamp 1607721120
transform 1 0 27232 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_280
timestamp 1607721120
transform 1 0 26864 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__C
timestamp 1607721120
transform 1 0 27048 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__B
timestamp 1607721120
transform 1 0 27416 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0834_
timestamp 1607721120
transform 1 0 27600 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_310
timestamp 1607721120
transform 1 0 29624 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_306
timestamp 1607721120
transform 1 0 29256 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_301
timestamp 1607721120
transform 1 0 28796 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_297
timestamp 1607721120
transform 1 0 28428 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__D
timestamp 1607721120
transform 1 0 28980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__C
timestamp 1607721120
transform 1 0 29716 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__A
timestamp 1607721120
transform 1 0 28612 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1607721120
transform 1 0 29164 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0814_
timestamp 1607721120
transform 1 0 29900 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_21_332
timestamp 1607721120
transform 1 0 31648 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_328
timestamp 1607721120
transform 1 0 31280 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_324
timestamp 1607721120
transform 1 0 30912 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_320
timestamp 1607721120
transform 1 0 30544 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1318__B1
timestamp 1607721120
transform 1 0 32016 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__D
timestamp 1607721120
transform 1 0 31464 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__A
timestamp 1607721120
transform 1 0 31096 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__B
timestamp 1607721120
transform 1 0 30728 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1318_
timestamp 1607721120
transform 1 0 32200 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_362
timestamp 1607721120
transform 1 0 34408 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_358
timestamp 1607721120
transform 1 0 34040 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_354
timestamp 1607721120
transform 1 0 33672 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_350
timestamp 1607721120
transform 1 0 33304 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1309__C
timestamp 1607721120
transform 1 0 34224 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1298__B1
timestamp 1607721120
transform 1 0 33856 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1309__B
timestamp 1607721120
transform 1 0 34592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1427__D
timestamp 1607721120
transform 1 0 33488 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_388
timestamp 1607721120
transform 1 0 36800 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_384
timestamp 1607721120
transform 1 0 36432 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_380
timestamp 1607721120
transform 1 0 36064 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_376
timestamp 1607721120
transform 1 0 35696 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1317__A2
timestamp 1607721120
transform 1 0 36616 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__B
timestamp 1607721120
transform 1 0 36248 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__A
timestamp 1607721120
transform 1 0 35880 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1607721120
transform 1 0 34776 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _1309_
timestamp 1607721120
transform 1 0 34868 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_406
timestamp 1607721120
transform 1 0 38456 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_402
timestamp 1607721120
transform 1 0 38088 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_392
timestamp 1607721120
transform 1 0 37168 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__B
timestamp 1607721120
transform 1 0 37260 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__B
timestamp 1607721120
transform 1 0 38640 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__A
timestamp 1607721120
transform 1 0 38272 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0807_
timestamp 1607721120
transform 1 0 37444 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _0793_
timestamp 1607721120
transform 1 0 38824 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_21_424
timestamp 1607721120
transform 1 0 40112 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_419
timestamp 1607721120
transform 1 0 39652 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__B1
timestamp 1607721120
transform 1 0 39928 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1607721120
transform 1 0 40388 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0787_
timestamp 1607721120
transform 1 0 40480 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_21_453
timestamp 1607721120
transform 1 0 42780 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_442
timestamp 1607721120
transform 1 0 41768 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_439
timestamp 1607721120
transform 1 0 41492 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_435
timestamp 1607721120
transform 1 0 41124 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__C
timestamp 1607721120
transform 1 0 42964 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__A
timestamp 1607721120
transform 1 0 41584 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0781_
timestamp 1607721120
transform 1 0 41952 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_478
timestamp 1607721120
transform 1 0 45080 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_474
timestamp 1607721120
transform 1 0 44712 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_470
timestamp 1607721120
transform 1 0 44344 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_457
timestamp 1607721120
transform 1 0 43148 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__B
timestamp 1607721120
transform 1 0 44896 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__A
timestamp 1607721120
transform 1 0 44528 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__A
timestamp 1607721120
transform 1 0 43332 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0808_
timestamp 1607721120
transform 1 0 43516 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_501
timestamp 1607721120
transform 1 0 47196 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_484
timestamp 1607721120
transform 1 0 45632 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_wb_clk_i_A
timestamp 1607721120
transform 1 0 45448 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1458__D
timestamp 1607721120
transform 1 0 45816 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1607721120
transform 1 0 46000 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1346_
timestamp 1607721120
transform 1 0 46092 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_523
timestamp 1607721120
transform 1 0 49220 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_519
timestamp 1607721120
transform 1 0 48852 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_509
timestamp 1607721120
transform 1 0 47932 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_505
timestamp 1607721120
transform 1 0 47564 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1346__A1
timestamp 1607721120
transform 1 0 47748 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__A
timestamp 1607721120
transform 1 0 49036 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1346__B1
timestamp 1607721120
transform 1 0 47380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0774_
timestamp 1607721120
transform 1 0 48024 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_545
timestamp 1607721120
transform 1 0 51244 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_541
timestamp 1607721120
transform 1 0 50876 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_528
timestamp 1607721120
transform 1 0 49680 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1300__B1
timestamp 1607721120
transform 1 0 51428 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__C
timestamp 1607721120
transform 1 0 49496 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__A
timestamp 1607721120
transform 1 0 49864 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1457__D
timestamp 1607721120
transform 1 0 51060 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0711_
timestamp 1607721120
transform 1 0 50048 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_554
timestamp 1607721120
transform 1 0 52072 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__A
timestamp 1607721120
transform 1 0 52256 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1607721120
transform 1 0 51612 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0683_
timestamp 1607721120
transform 1 0 51704 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_558
timestamp 1607721120
transform 1 0 52440 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__A
timestamp 1607721120
transform 1 0 52624 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0692_
timestamp 1607721120
transform 1 0 52808 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_570
timestamp 1607721120
transform 1 0 53544 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_566
timestamp 1607721120
transform 1 0 53176 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0692__A
timestamp 1607721120
transform 1 0 53360 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_580
timestamp 1607721120
transform 1 0 54464 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1454__CLK
timestamp 1607721120
transform 1 0 54280 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1454__D
timestamp 1607721120
transform 1 0 54648 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _0725_
timestamp 1607721120
transform 1 0 54832 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_604
timestamp 1607721120
transform 1 0 56672 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_600
timestamp 1607721120
transform 1 0 56304 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_596
timestamp 1607721120
transform 1 0 55936 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__A1
timestamp 1607721120
transform 1 0 56488 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1455__D
timestamp 1607721120
transform 1 0 57040 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__B1
timestamp 1607721120
transform 1 0 56120 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1607721120
transform 1 0 57224 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _0712_
timestamp 1607721120
transform 1 0 57316 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_631
timestamp 1607721120
transform 1 0 59156 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_627
timestamp 1607721120
transform 1 0 58788 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_623
timestamp 1607721120
transform 1 0 58420 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__A1
timestamp 1607721120
transform 1 0 58972 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__B1
timestamp 1607721120
transform 1 0 58604 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_655
timestamp 1607721120
transform 1 0 61364 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_643
timestamp 1607721120
transform 1 0 60260 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_672
timestamp 1607721120
transform 1 0 62928 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_667
timestamp 1607721120
transform 1 0 62468 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1607721120
transform 1 0 62836 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1607721120
transform -1 0 63480 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1607721120
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1607721120
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1607721120
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_44
timestamp 1607721120
transform 1 0 5152 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1607721120
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1607721120
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1607721120
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_64
timestamp 1607721120
transform 1 0 6992 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_60
timestamp 1607721120
transform 1 0 6624 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_50
timestamp 1607721120
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1334__A
timestamp 1607721120
transform 1 0 5520 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__C
timestamp 1607721120
transform 1 0 6808 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0902_
timestamp 1607721120
transform 1 0 5796 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_4  _0898_
timestamp 1607721120
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_90
timestamp 1607721120
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_84
timestamp 1607721120
transform 1 0 8832 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_80
timestamp 1607721120
transform 1 0 8464 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__B
timestamp 1607721120
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__A2
timestamp 1607721120
transform 1 0 8648 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_111
timestamp 1607721120
transform 1 0 11316 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_107
timestamp 1607721120
transform 1 0 10948 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_104
timestamp 1607721120
transform 1 0 10672 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_100
timestamp 1607721120
transform 1 0 10304 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__A2
timestamp 1607721120
transform 1 0 11132 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__A
timestamp 1607721120
transform 1 0 10764 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1607721120
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1380_
timestamp 1607721120
transform 1 0 11500 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_4  _1341_
timestamp 1607721120
transform 1 0 9660 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_22_136
timestamp 1607721120
transform 1 0 13616 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_132
timestamp 1607721120
transform 1 0 13248 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__A2
timestamp 1607721120
transform 1 0 13432 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_158
timestamp 1607721120
transform 1 0 15640 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_150
timestamp 1607721120
transform 1 0 14904 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_144
timestamp 1607721120
transform 1 0 14352 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1330__B1
timestamp 1607721120
transform 1 0 14720 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__C
timestamp 1607721120
transform 1 0 13800 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1607721120
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1294_
timestamp 1607721120
transform 1 0 15272 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0672_
timestamp 1607721120
transform 1 0 13984 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_167
timestamp 1607721120
transform 1 0 16468 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_162
timestamp 1607721120
transform 1 0 16008 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_wb_clk_i_A
timestamp 1607721120
transform 1 0 16284 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1321__B
timestamp 1607721120
transform 1 0 16652 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1294__A
timestamp 1607721120
transform 1 0 15824 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1378_
timestamp 1607721120
transform 1 0 16836 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_22_202
timestamp 1607721120
transform 1 0 19688 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_198
timestamp 1607721120
transform 1 0 19320 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1607721120
transform 1 0 18952 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_190
timestamp 1607721120
transform 1 0 18584 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1223__A1
timestamp 1607721120
transform 1 0 19504 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1322__B
timestamp 1607721120
transform 1 0 19872 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__C
timestamp 1607721120
transform 1 0 19136 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__B
timestamp 1607721120
transform 1 0 18768 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_215
timestamp 1607721120
transform 1 0 20884 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_212
timestamp 1607721120
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_206
timestamp 1607721120
transform 1 0 20056 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__A2
timestamp 1607721120
transform 1 0 20424 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1607721120
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_223
timestamp 1607721120
transform 1 0 21620 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_219
timestamp 1607721120
transform 1 0 21252 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1411__CLK
timestamp 1607721120
transform 1 0 21436 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_wb_clk_i_A
timestamp 1607721120
transform 1 0 21068 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1379_
timestamp 1607721120
transform 1 0 21804 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_22_249
timestamp 1607721120
transform 1 0 24012 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_244
timestamp 1607721120
transform 1 0 23552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__C
timestamp 1607721120
transform 1 0 24196 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__B
timestamp 1607721120
transform 1 0 23828 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_271
timestamp 1607721120
transform 1 0 26036 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_267
timestamp 1607721120
transform 1 0 25668 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_257
timestamp 1607721120
transform 1 0 24748 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_253
timestamp 1607721120
transform 1 0 24380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1291__A
timestamp 1607721120
transform 1 0 25852 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__A
timestamp 1607721120
transform 1 0 26220 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0841__A
timestamp 1607721120
transform 1 0 24840 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0833_
timestamp 1607721120
transform 1 0 25024 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_22_285
timestamp 1607721120
transform 1 0 27324 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_281
timestamp 1607721120
transform 1 0 26956 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_276
timestamp 1607721120
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__B
timestamp 1607721120
transform 1 0 27140 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__D
timestamp 1607721120
transform 1 0 27508 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1607721120
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1291_
timestamp 1607721120
transform 1 0 26588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _0823_
timestamp 1607721120
transform 1 0 27692 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_22_313
timestamp 1607721120
transform 1 0 29900 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1607721120
transform 1 0 29532 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_306
timestamp 1607721120
transform 1 0 29256 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_302
timestamp 1607721120
transform 1 0 28888 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_298
timestamp 1607721120
transform 1 0 28520 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__C
timestamp 1607721120
transform 1 0 29716 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__B
timestamp 1607721120
transform 1 0 28704 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__A1
timestamp 1607721120
transform 1 0 29348 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0815_
timestamp 1607721120
transform 1 0 30176 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_22_341
timestamp 1607721120
transform 1 0 32476 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_337
timestamp 1607721120
transform 1 0 32108 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_332
timestamp 1607721120
transform 1 0 31648 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_329
timestamp 1607721120
transform 1 0 31372 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_325
timestamp 1607721120
transform 1 0 31004 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1318__A2
timestamp 1607721120
transform 1 0 31464 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1318__A1
timestamp 1607721120
transform 1 0 31832 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__B
timestamp 1607721120
transform 1 0 32292 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1607721120
transform 1 0 32016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_363
timestamp 1607721120
transform 1 0 34500 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__C
timestamp 1607721120
transform 1 0 34684 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1427_
timestamp 1607721120
transform 1 0 32752 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_22_388
timestamp 1607721120
transform 1 0 36800 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_384
timestamp 1607721120
transform 1 0 36432 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_380
timestamp 1607721120
transform 1 0 36064 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_367
timestamp 1607721120
transform 1 0 34868 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1316__A3
timestamp 1607721120
transform 1 0 36616 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1309__A
timestamp 1607721120
transform 1 0 35052 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__C
timestamp 1607721120
transform 1 0 36248 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0916_
timestamp 1607721120
transform 1 0 35236 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_409
timestamp 1607721120
transform 1 0 38732 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_398
timestamp 1607721120
transform 1 0 37720 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_392
timestamp 1607721120
transform 1 0 37168 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1316__A2
timestamp 1607721120
transform 1 0 36984 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__B
timestamp 1607721120
transform 1 0 37444 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__A
timestamp 1607721120
transform 1 0 38916 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1607721120
transform 1 0 37628 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0794_
timestamp 1607721120
transform 1 0 37904 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_22_433
timestamp 1607721120
transform 1 0 40940 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_429
timestamp 1607721120
transform 1 0 40572 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_413
timestamp 1607721120
transform 1 0 39100 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__A
timestamp 1607721120
transform 1 0 39284 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__A1
timestamp 1607721120
transform 1 0 40756 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _0795_
timestamp 1607721120
transform 1 0 39468 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_453
timestamp 1607721120
transform 1 0 42780 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_449
timestamp 1607721120
transform 1 0 42412 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_437
timestamp 1607721120
transform 1 0 41308 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__A
timestamp 1607721120
transform 1 0 41400 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__A1
timestamp 1607721120
transform 1 0 42964 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__A1
timestamp 1607721120
transform 1 0 42596 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0775_
timestamp 1607721120
transform 1 0 41584 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_22_457
timestamp 1607721120
transform 1 0 43148 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1607721120
transform 1 0 43240 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0777_
timestamp 1607721120
transform 1 0 43332 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_463
timestamp 1607721120
transform 1 0 43700 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__B
timestamp 1607721120
transform 1 0 43884 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_471
timestamp 1607721120
transform 1 0 44436 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_467
timestamp 1607721120
transform 1 0 44068 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__C
timestamp 1607721120
transform 1 0 44252 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_475
timestamp 1607721120
transform 1 0 44804 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1372__CLK
timestamp 1607721120
transform 1 0 44620 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_479
timestamp 1607721120
transform 1 0 45172 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1373__CLK
timestamp 1607721120
transform 1 0 44988 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_502
timestamp 1607721120
transform 1 0 47288 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1458__CLK
timestamp 1607721120
transform 1 0 45356 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1458_
timestamp 1607721120
transform 1 0 45540 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_22_506
timestamp 1607721120
transform 1 0 47656 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1346__A2
timestamp 1607721120
transform 1 0 47472 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_510
timestamp 1607721120
transform 1 0 48024 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__B
timestamp 1607721120
transform 1 0 48116 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_513
timestamp 1607721120
transform 1 0 48300 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__A2
timestamp 1607721120
transform 1 0 48484 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_517
timestamp 1607721120
transform 1 0 48668 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1607721120
transform 1 0 48852 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0673_
timestamp 1607721120
transform 1 0 48944 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_524
timestamp 1607721120
transform 1 0 49312 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_532
timestamp 1607721120
transform 1 0 50048 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_528
timestamp 1607721120
transform 1 0 49680 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__C
timestamp 1607721120
transform 1 0 49864 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__A
timestamp 1607721120
transform 1 0 49496 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1457_
timestamp 1607721120
transform 1 0 50140 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_22_568
timestamp 1607721120
transform 1 0 53360 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_564
timestamp 1607721120
transform 1 0 52992 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_556
timestamp 1607721120
transform 1 0 52256 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_552
timestamp 1607721120
transform 1 0 51888 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1457__CLK
timestamp 1607721120
transform 1 0 52072 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__C
timestamp 1607721120
transform 1 0 53544 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__B
timestamp 1607721120
transform 1 0 53176 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0716_
timestamp 1607721120
transform 1 0 52624 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_572
timestamp 1607721120
transform 1 0 53728 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1607721120
transform 1 0 54464 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1454_
timestamp 1607721120
transform 1 0 54556 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_22_604
timestamp 1607721120
transform 1 0 56672 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_600
timestamp 1607721120
transform 1 0 56304 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1456__CLK
timestamp 1607721120
transform 1 0 56856 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__A2
timestamp 1607721120
transform 1 0 56488 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1455_
timestamp 1607721120
transform 1 0 57040 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_22_639
timestamp 1607721120
transform 1 0 59892 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_631
timestamp 1607721120
transform 1 0 59156 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_627
timestamp 1607721120
transform 1 0 58788 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__A2
timestamp 1607721120
transform 1 0 58972 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_654
timestamp 1607721120
transform 1 0 61272 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_642
timestamp 1607721120
transform 1 0 60168 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1607721120
transform 1 0 60076 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_674
timestamp 1607721120
transform 1 0 63112 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_666
timestamp 1607721120
transform 1 0 62376 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1607721120
transform -1 0 63480 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1607721120
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1607721120
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1607721120
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_42
timestamp 1607721120
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_38
timestamp 1607721120
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_35
timestamp 1607721120
transform 1 0 4324 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_27
timestamp 1607721120
transform 1 0 3588 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1429__CLK
timestamp 1607721120
transform 1 0 4416 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1344__B
timestamp 1607721120
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1344__A
timestamp 1607721120
transform 1 0 5152 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_62
timestamp 1607721120
transform 1 0 6808 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1607721120
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_53
timestamp 1607721120
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1430__CLK
timestamp 1607721120
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0892__A
timestamp 1607721120
transform 1 0 7084 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1429__D
timestamp 1607721120
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1607721120
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1430_
timestamp 1607721120
transform 1 0 7268 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1344_
timestamp 1607721120
transform 1 0 5336 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_23_90
timestamp 1607721120
transform 1 0 9384 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_86
timestamp 1607721120
transform 1 0 9016 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0892__C
timestamp 1607721120
transform 1 0 9200 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_114
timestamp 1607721120
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1607721120
transform 1 0 11224 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_106
timestamp 1607721120
transform 1 0 10856 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1428__D
timestamp 1607721120
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__B1
timestamp 1607721120
transform 1 0 11040 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _0893_
timestamp 1607721120
transform 1 0 9752 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_135
timestamp 1607721120
transform 1 0 13524 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_118
timestamp 1607721120
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1380__CLK
timestamp 1607721120
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1358__CLK
timestamp 1607721120
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__B1
timestamp 1607721120
transform 1 0 13708 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1607721120
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _0878_
timestamp 1607721120
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_159
timestamp 1607721120
transform 1 0 15732 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_151
timestamp 1607721120
transform 1 0 14996 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_147
timestamp 1607721120
transform 1 0 14628 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_139
timestamp 1607721120
transform 1 0 13892 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__A
timestamp 1607721120
transform 1 0 14076 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__A
timestamp 1607721120
transform 1 0 15180 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__A
timestamp 1607721120
transform 1 0 14812 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0871_
timestamp 1607721120
transform 1 0 15364 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0870_
timestamp 1607721120
transform 1 0 14260 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_163
timestamp 1607721120
transform 1 0 16100 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__A
timestamp 1607721120
transform 1 0 15916 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_167
timestamp 1607721120
transform 1 0 16468 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1377__CLK
timestamp 1607721120
transform 1 0 16284 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1378__CLK
timestamp 1607721120
transform 1 0 16652 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0836_
timestamp 1607721120
transform 1 0 16836 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_179
timestamp 1607721120
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_175
timestamp 1607721120
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__A
timestamp 1607721120
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__A
timestamp 1607721120
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_197
timestamp 1607721120
transform 1 0 19228 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_193
timestamp 1607721120
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__A
timestamp 1607721120
transform 1 0 19044 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__A
timestamp 1607721120
transform 1 0 19412 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1607721120
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0858_
timestamp 1607721120
transform 1 0 18032 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_4  _0851_
timestamp 1607721120
transform 1 0 19596 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_217
timestamp 1607721120
transform 1 0 21068 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_213
timestamp 1607721120
transform 1 0 20700 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1381__D
timestamp 1607721120
transform 1 0 21252 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__B1
timestamp 1607721120
transform 1 0 20884 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _0844_
timestamp 1607721120
transform 1 0 21436 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_241
timestamp 1607721120
transform 1 0 23276 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_237
timestamp 1607721120
transform 1 0 22908 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_233
timestamp 1607721120
transform 1 0 22540 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0844__A1
timestamp 1607721120
transform 1 0 23092 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0844__B1
timestamp 1607721120
transform 1 0 22724 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1607721120
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0850_
timestamp 1607721120
transform 1 0 23644 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_23_266
timestamp 1607721120
transform 1 0 25576 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_262
timestamp 1607721120
transform 1 0 25208 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_258
timestamp 1607721120
transform 1 0 24840 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_254
timestamp 1607721120
transform 1 0 24472 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1379__CLK
timestamp 1607721120
transform 1 0 25024 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__A
timestamp 1607721120
transform 1 0 25668 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__A
timestamp 1607721120
transform 1 0 24656 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0822_
timestamp 1607721120
transform 1 0 25852 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_23_283
timestamp 1607721120
transform 1 0 27140 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_280
timestamp 1607721120
transform 1 0 26864 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_276
timestamp 1607721120
transform 1 0 26496 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__C
timestamp 1607721120
transform 1 0 27416 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__A
timestamp 1607721120
transform 1 0 26956 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0829_
timestamp 1607721120
transform 1 0 27600 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_319
timestamp 1607721120
transform 1 0 30452 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_315
timestamp 1607721120
transform 1 0 30084 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_301
timestamp 1607721120
transform 1 0 28796 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_297
timestamp 1607721120
transform 1 0 28428 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__B
timestamp 1607721120
transform 1 0 30268 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__A2
timestamp 1607721120
transform 1 0 28612 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__B1
timestamp 1607721120
transform 1 0 28980 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1607721120
transform 1 0 29164 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0824_
timestamp 1607721120
transform 1 0 29256 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1288__A
timestamp 1607721120
transform 1 0 30636 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1288_
timestamp 1607721120
transform 1 0 30820 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_326
timestamp 1607721120
transform 1 0 31096 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__A
timestamp 1607721120
transform 1 0 31280 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_330
timestamp 1607721120
transform 1 0 31464 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__C
timestamp 1607721120
transform 1 0 31648 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0801_
timestamp 1607721120
transform 1 0 31832 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_338
timestamp 1607721120
transform 1 0 32200 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_342
timestamp 1607721120
transform 1 0 32568 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0801__A
timestamp 1607721120
transform 1 0 32384 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_362
timestamp 1607721120
transform 1 0 34408 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_358
timestamp 1607721120
transform 1 0 34040 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__A
timestamp 1607721120
transform 1 0 32752 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__A1
timestamp 1607721120
transform 1 0 34592 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__B1
timestamp 1607721120
transform 1 0 34224 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _0909_
timestamp 1607721120
transform 1 0 32936 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_382
timestamp 1607721120
transform 1 0 36248 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_378
timestamp 1607721120
transform 1 0 35880 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_374
timestamp 1607721120
transform 1 0 35512 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1311__A
timestamp 1607721120
transform 1 0 36340 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__A
timestamp 1607721120
transform 1 0 35696 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1607721120
transform 1 0 34776 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1311_
timestamp 1607721120
transform 1 0 36524 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _1310_
timestamp 1607721120
transform 1 0 34868 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_23_406
timestamp 1607721120
transform 1 0 38456 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_400
timestamp 1607721120
transform 1 0 37904 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_396
timestamp 1607721120
transform 1 0 37536 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_392
timestamp 1607721120
transform 1 0 37168 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1316__B2
timestamp 1607721120
transform 1 0 37720 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1231__A
timestamp 1607721120
transform 1 0 37352 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__B
timestamp 1607721120
transform 1 0 38272 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1444__D
timestamp 1607721120
transform 1 0 38640 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0789_
timestamp 1607721120
transform 1 0 38824 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_432
timestamp 1607721120
transform 1 0 40848 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_428
timestamp 1607721120
transform 1 0 40480 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_423
timestamp 1607721120
transform 1 0 40020 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_419
timestamp 1607721120
transform 1 0 39652 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__C
timestamp 1607721120
transform 1 0 40204 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0787__B
timestamp 1607721120
transform 1 0 40664 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__A2
timestamp 1607721120
transform 1 0 39836 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1607721120
transform 1 0 40388 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_450
timestamp 1607721120
transform 1 0 42504 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_446
timestamp 1607721120
transform 1 0 42136 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__B1
timestamp 1607721120
transform 1 0 42688 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__B1
timestamp 1607721120
transform 1 0 42320 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0782_
timestamp 1607721120
transform 1 0 42872 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_4  _0776_
timestamp 1607721120
transform 1 0 41032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_479
timestamp 1607721120
transform 1 0 45172 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_467
timestamp 1607721120
transform 1 0 44068 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_463
timestamp 1607721120
transform 1 0 43700 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__A2
timestamp 1607721120
transform 1 0 43884 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_502
timestamp 1607721120
transform 1 0 47288 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_498
timestamp 1607721120
transform 1 0 46920 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_493
timestamp 1607721120
transform 1 0 46460 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_489
timestamp 1607721120
transform 1 0 46092 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_487
timestamp 1607721120
transform 1 0 45908 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__A
timestamp 1607721120
transform 1 0 46276 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__A
timestamp 1607721120
transform 1 0 47104 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1607721120
transform 1 0 46000 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0730_
timestamp 1607721120
transform 1 0 46552 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_522
timestamp 1607721120
transform 1 0 49128 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_518
timestamp 1607721120
transform 1 0 48760 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__A
timestamp 1607721120
transform 1 0 47472 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__A
timestamp 1607721120
transform 1 0 49312 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__B1
timestamp 1607721120
transform 1 0 48944 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _0762_
timestamp 1607721120
transform 1 0 47656 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_547
timestamp 1607721120
transform 1 0 51428 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_543
timestamp 1607721120
transform 1 0 51060 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_539
timestamp 1607721120
transform 1 0 50692 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_535
timestamp 1607721120
transform 1 0 50324 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__B
timestamp 1607721120
transform 1 0 50508 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__A2
timestamp 1607721120
transform 1 0 50876 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__B1
timestamp 1607721120
transform 1 0 51244 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0766_
timestamp 1607721120
transform 1 0 49496 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_558
timestamp 1607721120
transform 1 0 52440 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_554
timestamp 1607721120
transform 1 0 52072 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__A
timestamp 1607721120
transform 1 0 52624 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__A1
timestamp 1607721120
transform 1 0 52256 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1607721120
transform 1 0 51612 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0739_
timestamp 1607721120
transform 1 0 52808 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0693_
timestamp 1607721120
transform 1 0 51704 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_579
timestamp 1607721120
transform 1 0 54372 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_575
timestamp 1607721120
transform 1 0 54004 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_571
timestamp 1607721120
transform 1 0 53636 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__A1
timestamp 1607721120
transform 1 0 54188 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__C
timestamp 1607721120
transform 1 0 55476 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__B1
timestamp 1607721120
transform 1 0 53820 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0724_
timestamp 1607721120
transform 1 0 55660 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_608
timestamp 1607721120
transform 1 0 57040 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_602
timestamp 1607721120
transform 1 0 56488 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__B1
timestamp 1607721120
transform 1 0 56856 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1607721120
transform 1 0 57224 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1456_
timestamp 1607721120
transform 1 0 57316 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_23_630
timestamp 1607721120
transform 1 0 59064 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_654
timestamp 1607721120
transform 1 0 61272 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_642
timestamp 1607721120
transform 1 0 60168 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_672
timestamp 1607721120
transform 1 0 62928 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_670
timestamp 1607721120
transform 1 0 62744 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_666
timestamp 1607721120
transform 1 0 62376 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1607721120
transform 1 0 62836 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1607721120
transform -1 0 63480 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1607721120
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1607721120
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1607721120
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_44
timestamp 1607721120
transform 1 0 5152 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1607721120
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1607721120
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1607721120
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_65
timestamp 1607721120
transform 1 0 7084 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1429_
timestamp 1607721120
transform 1 0 5336 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_24_88
timestamp 1607721120
transform 1 0 9200 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_84
timestamp 1607721120
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_72
timestamp 1607721120
transform 1 0 7728 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_69
timestamp 1607721120
transform 1 0 7452 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0892__B
timestamp 1607721120
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1430__D
timestamp 1607721120
transform 1 0 7544 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0892_
timestamp 1607721120
transform 1 0 8004 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_105
timestamp 1607721120
transform 1 0 10764 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_101
timestamp 1607721120
transform 1 0 10396 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_93
timestamp 1607721120
transform 1 0 9660 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1428__CLK
timestamp 1607721120
transform 1 0 10212 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__A1
timestamp 1607721120
transform 1 0 10580 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1607721120
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1428_
timestamp 1607721120
transform 1 0 10948 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_24_130
timestamp 1607721120
transform 1 0 13064 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_126
timestamp 1607721120
transform 1 0 12696 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1331__C
timestamp 1607721120
transform 1 0 12880 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__A1
timestamp 1607721120
transform 1 0 13248 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0877_
timestamp 1607721120
transform 1 0 13432 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_24_158
timestamp 1607721120
transform 1 0 15640 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_147
timestamp 1607721120
transform 1 0 14628 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_143
timestamp 1607721120
transform 1 0 14260 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__B
timestamp 1607721120
transform 1 0 14444 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1607721120
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0872_
timestamp 1607721120
transform 1 0 15272 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_176
timestamp 1607721120
transform 1 0 17296 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_171
timestamp 1607721120
transform 1 0 16836 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_167
timestamp 1607721120
transform 1 0 16468 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_164
timestamp 1607721120
transform 1 0 16192 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__C
timestamp 1607721120
transform 1 0 16652 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__C
timestamp 1607721120
transform 1 0 17112 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__B
timestamp 1607721120
transform 1 0 17480 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__A
timestamp 1607721120
transform 1 0 16284 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0864_
timestamp 1607721120
transform 1 0 17664 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_193
timestamp 1607721120
transform 1 0 18860 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_189
timestamp 1607721120
transform 1 0 18492 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__A2
timestamp 1607721120
transform 1 0 19044 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1435__D
timestamp 1607721120
transform 1 0 18676 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _0671_
timestamp 1607721120
transform 1 0 19228 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_215
timestamp 1607721120
transform 1 0 20884 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_210
timestamp 1607721120
transform 1 0 20424 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_206
timestamp 1607721120
transform 1 0 20056 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__A1
timestamp 1607721120
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__B
timestamp 1607721120
transform 1 0 20240 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1607721120
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_223
timestamp 1607721120
transform 1 0 21620 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_219
timestamp 1607721120
transform 1 0 21252 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1375__CLK
timestamp 1607721120
transform 1 0 21436 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1382__CLK
timestamp 1607721120
transform 1 0 21068 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1381_
timestamp 1607721120
transform 1 0 21712 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_24_247
timestamp 1607721120
transform 1 0 23828 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_243
timestamp 1607721120
transform 1 0 23460 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__B
timestamp 1607721120
transform 1 0 24012 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__A
timestamp 1607721120
transform 1 0 23644 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0837_
timestamp 1607721120
transform 1 0 24196 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_272
timestamp 1607721120
transform 1 0 26128 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_268
timestamp 1607721120
transform 1 0 25760 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_263
timestamp 1607721120
transform 1 0 25300 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_255
timestamp 1607721120
transform 1 0 24564 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1419__CLK
timestamp 1607721120
transform 1 0 25576 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__B
timestamp 1607721120
transform 1 0 25944 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_294
timestamp 1607721120
transform 1 0 28152 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_290
timestamp 1607721120
transform 1 0 27784 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_276
timestamp 1607721120
transform 1 0 26496 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__C
timestamp 1607721120
transform 1 0 26772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__B
timestamp 1607721120
transform 1 0 28336 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__A
timestamp 1607721120
transform 1 0 27968 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1607721120
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0835_
timestamp 1607721120
transform 1 0 26956 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_319
timestamp 1607721120
transform 1 0 30452 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_314
timestamp 1607721120
transform 1 0 29992 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_310
timestamp 1607721120
transform 1 0 29624 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__A
timestamp 1607721120
transform 1 0 29808 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__B1
timestamp 1607721120
transform 1 0 30268 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _0825_
timestamp 1607721120
transform 1 0 28520 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_332
timestamp 1607721120
transform 1 0 31648 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_328
timestamp 1607721120
transform 1 0 31280 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_323
timestamp 1607721120
transform 1 0 30820 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1427__CLK
timestamp 1607721120
transform 1 0 31464 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1368__CLK
timestamp 1607721120
transform 1 0 31832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__A2
timestamp 1607721120
transform 1 0 30636 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1607721120
transform 1 0 32016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0816_
timestamp 1607721120
transform 1 0 32108 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0803_
timestamp 1607721120
transform 1 0 30912 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_364
timestamp 1607721120
transform 1 0 34592 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_351
timestamp 1607721120
transform 1 0 33396 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_346
timestamp 1607721120
transform 1 0 32936 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__A
timestamp 1607721120
transform 1 0 33212 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__A2
timestamp 1607721120
transform 1 0 33580 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0809_
timestamp 1607721120
transform 1 0 33764 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_383
timestamp 1607721120
transform 1 0 36340 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_380
timestamp 1607721120
transform 1 0 36064 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_376
timestamp 1607721120
transform 1 0 35696 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_368
timestamp 1607721120
transform 1 0 34960 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1349__C
timestamp 1607721120
transform 1 0 36156 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1310__A
timestamp 1607721120
transform 1 0 35144 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__B
timestamp 1607721120
transform 1 0 34776 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1231_
timestamp 1607721120
transform 1 0 36524 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0802_
timestamp 1607721120
transform 1 0 35328 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_404
timestamp 1607721120
transform 1 0 38272 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_398
timestamp 1607721120
transform 1 0 37720 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_393
timestamp 1607721120
transform 1 0 37260 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_389
timestamp 1607721120
transform 1 0 36892 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1444__CLK
timestamp 1607721120
transform 1 0 38364 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1311__B
timestamp 1607721120
transform 1 0 37076 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__A
timestamp 1607721120
transform 1 0 37444 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1607721120
transform 1 0 37628 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1444_
timestamp 1607721120
transform 1 0 38548 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_24_430
timestamp 1607721120
transform 1 0 40664 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_426
timestamp 1607721120
transform 1 0 40296 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1374__CLK
timestamp 1607721120
transform 1 0 40848 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0787__A
timestamp 1607721120
transform 1 0 40480 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_456
timestamp 1607721120
transform 1 0 43056 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_450
timestamp 1607721120
transform 1 0 42504 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_434
timestamp 1607721120
transform 1 0 41032 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__A2
timestamp 1607721120
transform 1 0 41216 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__A
timestamp 1607721120
transform 1 0 42872 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _0770_
timestamp 1607721120
transform 1 0 41400 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_479
timestamp 1607721120
transform 1 0 45172 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_467
timestamp 1607721120
transform 1 0 44068 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_463
timestamp 1607721120
transform 1 0 43700 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_459
timestamp 1607721120
transform 1 0 43332 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__C
timestamp 1607721120
transform 1 0 43884 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__B
timestamp 1607721120
transform 1 0 43516 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1607721120
transform 1 0 43240 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_498
timestamp 1607721120
transform 1 0 46920 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_494
timestamp 1607721120
transform 1 0 46552 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_487
timestamp 1607721120
transform 1 0 45908 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__C
timestamp 1607721120
transform 1 0 46736 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__B
timestamp 1607721120
transform 1 0 47104 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0761_
timestamp 1607721120
transform 1 0 47288 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0732_
timestamp 1607721120
transform 1 0 46184 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_517
timestamp 1607721120
transform 1 0 48668 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_511
timestamp 1607721120
transform 1 0 48116 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__A1
timestamp 1607721120
transform 1 0 48484 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1607721120
transform 1 0 48852 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0756_
timestamp 1607721120
transform 1 0 48944 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_24_537
timestamp 1607721120
transform 1 0 50508 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_533
timestamp 1607721120
transform 1 0 50140 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_529
timestamp 1607721120
transform 1 0 49772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__C
timestamp 1607721120
transform 1 0 50324 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__B
timestamp 1607721120
transform 1 0 49956 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _0694_
timestamp 1607721120
transform 1 0 50784 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_556
timestamp 1607721120
transform 1 0 52256 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_552
timestamp 1607721120
transform 1 0 51888 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__C
timestamp 1607721120
transform 1 0 52440 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__A
timestamp 1607721120
transform 1 0 52072 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _0740_
timestamp 1607721120
transform 1 0 52624 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_581
timestamp 1607721120
transform 1 0 54556 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_576
timestamp 1607721120
transform 1 0 54096 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_572
timestamp 1607721120
transform 1 0 53728 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__A2
timestamp 1607721120
transform 1 0 53912 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__A
timestamp 1607721120
transform 1 0 55660 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1607721120
transform 1 0 54464 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_613
timestamp 1607721120
transform 1 0 57500 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_599
timestamp 1607721120
transform 1 0 56212 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_595
timestamp 1607721120
transform 1 0 55844 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__B
timestamp 1607721120
transform 1 0 56028 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1456__D
timestamp 1607721120
transform 1 0 57684 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _0720_
timestamp 1607721120
transform 1 0 56396 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_633
timestamp 1607721120
transform 1 0 59340 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_621
timestamp 1607721120
transform 1 0 58236 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_617
timestamp 1607721120
transform 1 0 57868 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__A1
timestamp 1607721120
transform 1 0 58052 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_654
timestamp 1607721120
transform 1 0 61272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_642
timestamp 1607721120
transform 1 0 60168 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1607721120
transform 1 0 60076 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_674
timestamp 1607721120
transform 1 0 63112 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_666
timestamp 1607721120
transform 1 0 62376 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1607721120
transform -1 0 63480 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1607721120
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1607721120
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1607721120
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1607721120
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1607721120
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_62
timestamp 1607721120
transform 1 0 6808 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1607721120
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1607721120
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1431__CLK
timestamp 1607721120
transform 1 0 7360 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1607721120
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_74
timestamp 1607721120
transform 1 0 7912 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_70
timestamp 1607721120
transform 1 0 7544 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__A2
timestamp 1607721120
transform 1 0 7728 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__B1
timestamp 1607721120
transform 1 0 8096 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1431_
timestamp 1607721120
transform 1 0 8280 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_25_114
timestamp 1607721120
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_101
timestamp 1607721120
transform 1 0 10396 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_97
timestamp 1607721120
transform 1 0 10028 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0885__C
timestamp 1607721120
transform 1 0 10212 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0885__B
timestamp 1607721120
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0885_
timestamp 1607721120
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_131
timestamp 1607721120
transform 1 0 13156 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_123
timestamp 1607721120
transform 1 0 12420 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_118
timestamp 1607721120
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1432__CLK
timestamp 1607721120
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1432__D
timestamp 1607721120
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1607721120
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _0873_
timestamp 1607721120
transform 1 0 13340 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_157
timestamp 1607721120
transform 1 0 15548 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_153
timestamp 1607721120
transform 1 0 15180 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_149
timestamp 1607721120
transform 1 0 14812 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_145
timestamp 1607721120
transform 1 0 14444 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1434__CLK
timestamp 1607721120
transform 1 0 15640 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__A1
timestamp 1607721120
transform 1 0 14996 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__B1
timestamp 1607721120
transform 1 0 14628 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_178
timestamp 1607721120
transform 1 0 17480 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_174
timestamp 1607721120
transform 1 0 17112 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_164
timestamp 1607721120
transform 1 0 16192 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_160
timestamp 1607721120
transform 1 0 15824 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1376__CLK
timestamp 1607721120
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__B
timestamp 1607721120
transform 1 0 17296 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1434__D
timestamp 1607721120
transform 1 0 16008 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0869_
timestamp 1607721120
transform 1 0 16284 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_204
timestamp 1607721120
transform 1 0 19872 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_200
timestamp 1607721120
transform 1 0 19504 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_196
timestamp 1607721120
transform 1 0 19136 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__A1
timestamp 1607721120
transform 1 0 19688 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__B1
timestamp 1607721120
transform 1 0 19320 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1607721120
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _0865_
timestamp 1607721120
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1607721120
transform 1 0 21804 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1437__D
timestamp 1607721120
transform 1 0 21988 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1436_
timestamp 1607721120
transform 1 0 20056 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_25_240
timestamp 1607721120
transform 1 0 23184 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_237
timestamp 1607721120
transform 1 0 22908 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_233
timestamp 1607721120
transform 1 0 22540 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_229
timestamp 1607721120
transform 1 0 22172 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__C
timestamp 1607721120
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0844__A2
timestamp 1607721120
transform 1 0 22356 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__A
timestamp 1607721120
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1607721120
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0843_
timestamp 1607721120
transform 1 0 23644 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_25_270
timestamp 1607721120
transform 1 0 25944 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_266
timestamp 1607721120
transform 1 0 25576 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_258
timestamp 1607721120
transform 1 0 24840 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_254
timestamp 1607721120
transform 1 0 24472 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1438__CLK
timestamp 1607721120
transform 1 0 25024 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__A
timestamp 1607721120
transform 1 0 25760 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1438__D
timestamp 1607721120
transform 1 0 24656 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0838_
timestamp 1607721120
transform 1 0 25208 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_284
timestamp 1607721120
transform 1 0 27232 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_280
timestamp 1607721120
transform 1 0 26864 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1439__CLK
timestamp 1607721120
transform 1 0 26680 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__A
timestamp 1607721120
transform 1 0 27048 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1439__D
timestamp 1607721120
transform 1 0 27416 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0830_
timestamp 1607721120
transform 1 0 27600 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_301
timestamp 1607721120
transform 1 0 28796 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_297
timestamp 1607721120
transform 1 0 28428 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__C
timestamp 1607721120
transform 1 0 28980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__B
timestamp 1607721120
transform 1 0 28612 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1607721120
transform 1 0 29164 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1441_
timestamp 1607721120
transform 1 0 29256 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_25_336
timestamp 1607721120
transform 1 0 32016 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_333
timestamp 1607721120
transform 1 0 31740 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_329
timestamp 1607721120
transform 1 0 31372 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_325
timestamp 1607721120
transform 1 0 31004 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1442__CLK
timestamp 1607721120
transform 1 0 31832 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__A1
timestamp 1607721120
transform 1 0 31188 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1442__D
timestamp 1607721120
transform 1 0 32200 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _0810_
timestamp 1607721120
transform 1 0 32384 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_360
timestamp 1607721120
transform 1 0 34224 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_356
timestamp 1607721120
transform 1 0 33856 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_352
timestamp 1607721120
transform 1 0 33488 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1443__CLK
timestamp 1607721120
transform 1 0 34592 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__A1
timestamp 1607721120
transform 1 0 34040 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__B1
timestamp 1607721120
transform 1 0 33672 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_371
timestamp 1607721120
transform 1 0 35236 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_367
timestamp 1607721120
transform 1 0 34868 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1443__D
timestamp 1607721120
transform 1 0 35052 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1607721120
transform 1 0 34776 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_375
timestamp 1607721120
transform 1 0 35604 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1310__B
timestamp 1607721120
transform 1 0 35420 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1349__D
timestamp 1607721120
transform 1 0 35972 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_381
timestamp 1607721120
transform 1 0 36156 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1369__CLK
timestamp 1607721120
transform 1 0 36432 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_386
timestamp 1607721120
transform 1 0 36616 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_403
timestamp 1607721120
transform 1 0 38180 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_398
timestamp 1607721120
transform 1 0 37720 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1445__CLK
timestamp 1607721120
transform 1 0 37168 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__A1
timestamp 1607721120
transform 1 0 38364 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1445__D
timestamp 1607721120
transform 1 0 37996 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _0783_
timestamp 1607721120
transform 1 0 38548 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0767_
timestamp 1607721120
transform 1 0 37352 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_432
timestamp 1607721120
transform 1 0 40848 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_423
timestamp 1607721120
transform 1 0 40020 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_419
timestamp 1607721120
transform 1 0 39652 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0768__A
timestamp 1607721120
transform 1 0 40204 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__B1
timestamp 1607721120
transform 1 0 39836 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1607721120
transform 1 0 40388 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0768_
timestamp 1607721120
transform 1 0 40480 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_442
timestamp 1607721120
transform 1 0 41768 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_436
timestamp 1607721120
transform 1 0 41216 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1371__CLK
timestamp 1607721120
transform 1 0 41584 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1446__D
timestamp 1607721120
transform 1 0 41032 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1448_
timestamp 1607721120
transform 1 0 41860 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_25_474
timestamp 1607721120
transform 1 0 44712 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_462
timestamp 1607721120
transform 1 0 43608 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_498
timestamp 1607721120
transform 1 0 46920 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_494
timestamp 1607721120
transform 1 0 46552 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_489
timestamp 1607721120
transform 1 0 46092 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_486
timestamp 1607721120
transform 1 0 45816 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__A
timestamp 1607721120
transform 1 0 46736 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__B1
timestamp 1607721120
transform 1 0 47104 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1607721120
transform 1 0 46000 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1450_
timestamp 1607721120
transform 1 0 47288 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _0734_
timestamp 1607721120
transform 1 0 46184 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_525
timestamp 1607721120
transform 1 0 49404 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_521
timestamp 1607721120
transform 1 0 49036 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1451__D
timestamp 1607721120
transform 1 0 49220 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__A2
timestamp 1607721120
transform 1 0 49588 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0684_
timestamp 1607721120
transform 1 0 49772 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_533
timestamp 1607721120
transform 1 0 50140 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_537
timestamp 1607721120
transform 1 0 50508 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1451__CLK
timestamp 1607721120
transform 1 0 50692 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__A
timestamp 1607721120
transform 1 0 50324 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_541
timestamp 1607721120
transform 1 0 50876 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__B
timestamp 1607721120
transform 1 0 51060 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_545
timestamp 1607721120
transform 1 0 51244 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__A
timestamp 1607721120
transform 1 0 51428 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_563
timestamp 1607721120
transform 1 0 52900 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_559
timestamp 1607721120
transform 1 0 52532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1452__CLK
timestamp 1607721120
transform 1 0 53084 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1452__D
timestamp 1607721120
transform 1 0 52716 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1607721120
transform 1 0 51612 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1453_
timestamp 1607721120
transform 1 0 53268 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__and3_4  _0748_
timestamp 1607721120
transform 1 0 51704 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_25_586
timestamp 1607721120
transform 1 0 55016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_615
timestamp 1607721120
transform 1 0 57684 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_611
timestamp 1607721120
transform 1 0 57316 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_598
timestamp 1607721120
transform 1 0 56120 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__A2
timestamp 1607721120
transform 1 0 57500 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1607721120
transform 1 0 57224 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_639
timestamp 1607721120
transform 1 0 59892 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_627
timestamp 1607721120
transform 1 0 58788 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_651
timestamp 1607721120
transform 1 0 60996 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_672
timestamp 1607721120
transform 1 0 62928 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_663
timestamp 1607721120
transform 1 0 62100 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1607721120
transform 1 0 62836 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1607721120
transform -1 0 63480 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1607721120
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1607721120
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1607721120
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1607721120
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1607721120
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1607721120
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_44
timestamp 1607721120
transform 1 0 5152 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_32
timestamp 1607721120
transform 1 0 4048 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_27
timestamp 1607721120
transform 1 0 3588 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1607721120
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1607721120
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1607721120
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1607721120
transform 1 0 3956 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1607721120
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_63
timestamp 1607721120
transform 1 0 6900 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_56
timestamp 1607721120
transform 1 0 6256 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_68
timestamp 1607721120
transform 1 0 7360 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1607721120
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1607721120
transform 1 0 6808 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_87
timestamp 1607721120
transform 1 0 9108 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_75
timestamp 1607721120
transform 1 0 8004 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_88
timestamp 1607721120
transform 1 0 9200 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_84
timestamp 1607721120
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__A1
timestamp 1607721120
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1431__D
timestamp 1607721120
transform 1 0 9016 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _0886_
timestamp 1607721120
transform 1 0 7728 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_106
timestamp 1607721120
transform 1 0 10856 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_94
timestamp 1607721120
transform 1 0 9752 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_107
timestamp 1607721120
transform 1 0 10948 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1607721120
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0885__A
timestamp 1607721120
transform 1 0 10764 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1607721120
transform 1 0 9660 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1607721120
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1432_
timestamp 1607721120
transform 1 0 11040 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_27_125
timestamp 1607721120
transform 1 0 12604 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_118
timestamp 1607721120
transform 1 0 11960 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_132
timestamp 1607721120
transform 1 0 13248 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_127
timestamp 1607721120
transform 1 0 12788 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1433__CLK
timestamp 1607721120
transform 1 0 12328 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1433__D
timestamp 1607721120
transform 1 0 13064 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1607721120
transform 1 0 12512 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1433_
timestamp 1607721120
transform 1 0 12788 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_27_146
timestamp 1607721120
transform 1 0 14536 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_144
timestamp 1607721120
transform 1 0 14352 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_140
timestamp 1607721120
transform 1 0 13984 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__A2
timestamp 1607721120
transform 1 0 14168 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_154
timestamp 1607721120
transform 1 0 15272 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_158
timestamp 1607721120
transform 1 0 15640 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_154
timestamp 1607721120
transform 1 0 15272 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_152
timestamp 1607721120
transform 1 0 15088 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1607721120
transform 1 0 15364 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1607721120
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_156
timestamp 1607721120
transform 1 0 15456 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1434_
timestamp 1607721120
transform 1 0 15732 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_27_180
timestamp 1607721120
transform 1 0 17664 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_168
timestamp 1607721120
transform 1 0 16560 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_178
timestamp 1607721120
transform 1 0 17480 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_203
timestamp 1607721120
transform 1 0 19780 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_199
timestamp 1607721120
transform 1 0 19412 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_205
timestamp 1607721120
transform 1 0 19964 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1435__CLK
timestamp 1607721120
transform 1 0 18032 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0859__A1
timestamp 1607721120
transform 1 0 19964 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0859__B1
timestamp 1607721120
transform 1 0 19596 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1607721120
transform 1 0 18216 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1435_
timestamp 1607721120
transform 1 0 18216 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__a21o_4  _0859_
timestamp 1607721120
transform 1 0 18308 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_215
timestamp 1607721120
transform 1 0 20884 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_211
timestamp 1607721120
transform 1 0 20516 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_207
timestamp 1607721120
transform 1 0 20148 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_215
timestamp 1607721120
transform 1 0 20884 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_211
timestamp 1607721120
transform 1 0 20516 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1436__CLK
timestamp 1607721120
transform 1 0 20700 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0859__A2
timestamp 1607721120
transform 1 0 20332 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1436__D
timestamp 1607721120
transform 1 0 20332 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1607721120
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_226
timestamp 1607721120
transform 1 0 21896 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1607721120
transform 1 0 21528 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_218
timestamp 1607721120
transform 1 0 21160 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1437__CLK
timestamp 1607721120
transform 1 0 21344 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1381__CLK
timestamp 1607721120
transform 1 0 21712 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1607721120
transform 1 0 21068 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1437_
timestamp 1607721120
transform 1 0 21068 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__a21o_4  _0839_
timestamp 1607721120
transform 1 0 22080 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_236
timestamp 1607721120
transform 1 0 22816 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__A2
timestamp 1607721120
transform 1 0 23000 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_244
timestamp 1607721120
transform 1 0 23552 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_240
timestamp 1607721120
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_240
timestamp 1607721120
transform 1 0 23184 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__A1
timestamp 1607721120
transform 1 0 23736 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__B1
timestamp 1607721120
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1607721120
transform 1 0 23920 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_249
timestamp 1607721120
transform 1 0 24012 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1438_
timestamp 1607721120
transform 1 0 23552 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_27_273
timestamp 1607721120
transform 1 0 26220 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_261
timestamp 1607721120
transform 1 0 25116 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_263
timestamp 1607721120
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_280
timestamp 1607721120
transform 1 0 26864 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_282
timestamp 1607721120
transform 1 0 27048 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_276
timestamp 1607721120
transform 1 0 26496 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1440__CLK
timestamp 1607721120
transform 1 0 27140 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1440__D
timestamp 1607721120
transform 1 0 26588 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1607721120
transform 1 0 26772 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1607721120
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1440_
timestamp 1607721120
transform 1 0 27140 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1439_
timestamp 1607721120
transform 1 0 27324 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_27_308
timestamp 1607721120
transform 1 0 29440 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_302
timestamp 1607721120
transform 1 0 28888 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_308
timestamp 1607721120
transform 1 0 29440 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_304
timestamp 1607721120
transform 1 0 29072 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1441__CLK
timestamp 1607721120
transform 1 0 29256 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_311
timestamp 1607721120
transform 1 0 29716 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1441__D
timestamp 1607721120
transform 1 0 29532 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1607721120
transform 1 0 29624 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _0831_
timestamp 1607721120
transform 1 0 29716 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_4  _0817_
timestamp 1607721120
transform 1 0 29808 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_331
timestamp 1607721120
transform 1 0 31556 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_327
timestamp 1607721120
transform 1 0 31188 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_323
timestamp 1607721120
transform 1 0 30820 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_328
timestamp 1607721120
transform 1 0 31280 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_324
timestamp 1607721120
transform 1 0 30912 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__A2
timestamp 1607721120
transform 1 0 31096 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__A1
timestamp 1607721120
transform 1 0 31372 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__B1
timestamp 1607721120
transform 1 0 31004 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_342
timestamp 1607721120
transform 1 0 32568 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_339
timestamp 1607721120
transform 1 0 32292 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1607721120
transform 1 0 32476 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1607721120
transform 1 0 32016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1442_
timestamp 1607721120
transform 1 0 32108 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_27_364
timestamp 1607721120
transform 1 0 34592 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_350
timestamp 1607721120
transform 1 0 33304 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_360
timestamp 1607721120
transform 1 0 34224 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_356
timestamp 1607721120
transform 1 0 33856 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__A2
timestamp 1607721120
transform 1 0 34408 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__A2
timestamp 1607721120
transform 1 0 34040 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1443_
timestamp 1607721120
transform 1 0 34592 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__a21o_4  _0804_
timestamp 1607721120
transform 1 0 33488 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_385
timestamp 1607721120
transform 1 0 36524 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_373
timestamp 1607721120
transform 1 0 35420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_368
timestamp 1607721120
transform 1 0 34960 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_383
timestamp 1607721120
transform 1 0 36340 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__A1
timestamp 1607721120
transform 1 0 35144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__B1
timestamp 1607721120
transform 1 0 34776 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1607721120
transform 1 0 35328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_404
timestamp 1607721120
transform 1 0 38272 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_397
timestamp 1607721120
transform 1 0 37628 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_396
timestamp 1607721120
transform 1 0 37536 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_391
timestamp 1607721120
transform 1 0 37076 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__A2
timestamp 1607721120
transform 1 0 38824 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__A
timestamp 1607721120
transform 1 0 37352 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1607721120
transform 1 0 38180 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1607721120
transform 1 0 37628 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1445_
timestamp 1607721120
transform 1 0 37720 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_27_428
timestamp 1607721120
transform 1 0 40480 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_424
timestamp 1607721120
transform 1 0 40112 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_423
timestamp 1607721120
transform 1 0 40020 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_417
timestamp 1607721120
transform 1 0 39468 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__A1
timestamp 1607721120
transform 1 0 39836 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1447__D
timestamp 1607721120
transform 1 0 40848 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__B1
timestamp 1607721120
transform 1 0 40296 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1446_
timestamp 1607721120
transform 1 0 40204 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__a21o_4  _0790_
timestamp 1607721120
transform 1 0 39008 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_444
timestamp 1607721120
transform 1 0 41952 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1607721120
transform 1 0 41032 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_454
timestamp 1607721120
transform 1 0 42872 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_456
timestamp 1607721120
transform 1 0 43056 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_452
timestamp 1607721120
transform 1 0 42688 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_448
timestamp 1607721120
transform 1 0 42320 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1448__CLK
timestamp 1607721120
transform 1 0 42872 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1447__CLK
timestamp 1607721120
transform 1 0 43056 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1446__CLK
timestamp 1607721120
transform 1 0 42504 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1448__D
timestamp 1607721120
transform 1 0 42136 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1447_
timestamp 1607721120
transform 1 0 41124 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_27_478
timestamp 1607721120
transform 1 0 45080 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_466
timestamp 1607721120
transform 1 0 43976 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_464
timestamp 1607721120
transform 1 0 43792 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_458
timestamp 1607721120
transform 1 0 43240 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_471
timestamp 1607721120
transform 1 0 44436 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_459
timestamp 1607721120
transform 1 0 43332 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1607721120
transform 1 0 43884 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1607721120
transform 1 0 43240 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_490
timestamp 1607721120
transform 1 0 46184 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_483
timestamp 1607721120
transform 1 0 45540 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_495
timestamp 1607721120
transform 1 0 46644 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_491
timestamp 1607721120
transform 1 0 46276 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1450__CLK
timestamp 1607721120
transform 1 0 46460 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1449__CLK
timestamp 1607721120
transform 1 0 46828 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1449__D
timestamp 1607721120
transform 1 0 46552 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1607721120
transform 1 0 46736 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1449_
timestamp 1607721120
transform 1 0 46828 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__a21o_4  _0757_
timestamp 1607721120
transform 1 0 47012 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_524
timestamp 1607721120
transform 1 0 49312 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_516
timestamp 1607721120
transform 1 0 48576 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_515
timestamp 1607721120
transform 1 0 48484 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_511
timestamp 1607721120
transform 1 0 48116 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__A1
timestamp 1607721120
transform 1 0 48668 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1450__D
timestamp 1607721120
transform 1 0 48300 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1607721120
transform 1 0 48852 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1451_
timestamp 1607721120
transform 1 0 48944 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1607721120
transform 1 0 49588 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_548
timestamp 1607721120
transform 1 0 51520 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_544
timestamp 1607721120
transform 1 0 51152 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_540
timestamp 1607721120
transform 1 0 50784 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_543
timestamp 1607721120
transform 1 0 51060 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_539
timestamp 1607721120
transform 1 0 50692 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__A2
timestamp 1607721120
transform 1 0 50876 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__A1
timestamp 1607721120
transform 1 0 51336 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__B1
timestamp 1607721120
transform 1 0 50968 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _0749_
timestamp 1607721120
transform 1 0 49680 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1607721120
transform 1 0 52532 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_556
timestamp 1607721120
transform 1 0 52256 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_570
timestamp 1607721120
transform 1 0 53544 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1607721120
transform 1 0 52440 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1452_
timestamp 1607721120
transform 1 0 51796 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__a21o_4  _0735_
timestamp 1607721120
transform 1 0 52624 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_576
timestamp 1607721120
transform 1 0 54096 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_572
timestamp 1607721120
transform 1 0 53728 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_574
timestamp 1607721120
transform 1 0 53912 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__A2
timestamp 1607721120
transform 1 0 54096 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1453__D
timestamp 1607721120
transform 1 0 53728 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__B1
timestamp 1607721120
transform 1 0 53912 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_581
timestamp 1607721120
transform 1 0 54556 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_578
timestamp 1607721120
transform 1 0 54280 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__A1
timestamp 1607721120
transform 1 0 54280 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1607721120
transform 1 0 54464 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_580
timestamp 1607721120
transform 1 0 54464 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_588
timestamp 1607721120
transform 1 0 55200 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1453__CLK
timestamp 1607721120
transform 1 0 54740 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1607721120
transform 1 0 55292 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_590
timestamp 1607721120
transform 1 0 55384 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_585
timestamp 1607721120
transform 1 0 54924 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_614
timestamp 1607721120
transform 1 0 57592 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_602
timestamp 1607721120
transform 1 0 56488 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_609
timestamp 1607721120
transform 1 0 57132 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_597
timestamp 1607721120
transform 1 0 56028 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_633
timestamp 1607721120
transform 1 0 59340 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_621
timestamp 1607721120
transform 1 0 58236 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_633
timestamp 1607721120
transform 1 0 59340 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_621
timestamp 1607721120
transform 1 0 58236 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382
timestamp 1607721120
transform 1 0 58144 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_652
timestamp 1607721120
transform 1 0 61088 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_645
timestamp 1607721120
transform 1 0 60444 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_654
timestamp 1607721120
transform 1 0 61272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_642
timestamp 1607721120
transform 1 0 60168 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1607721120
transform 1 0 60996 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1607721120
transform 1 0 60076 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_672
timestamp 1607721120
transform 1 0 62928 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_664
timestamp 1607721120
transform 1 0 62192 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_674
timestamp 1607721120
transform 1 0 63112 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_666
timestamp 1607721120
transform 1 0 62376 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1607721120
transform -1 0 63480 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1607721120
transform -1 0 63480 0 -1 16864
box -38 -48 314 592
<< labels >>
rlabel metal3 s 0 1096 800 1216 6 cen
port 0 nsew default tristate
rlabel metal3 s 0 3272 800 3392 6 set_out[0]
port 1 nsew default tristate
rlabel metal3 s 0 5448 800 5568 6 set_out[1]
port 2 nsew default tristate
rlabel metal3 s 0 7760 800 7880 6 set_out[2]
port 3 nsew default tristate
rlabel metal3 s 0 9936 800 10056 6 set_out[3]
port 4 nsew default tristate
rlabel metal3 s 0 12112 800 12232 6 shift_out[0]
port 5 nsew default tristate
rlabel metal3 s 0 14424 800 14544 6 shift_out[1]
port 6 nsew default tristate
rlabel metal3 s 0 16600 800 16720 6 shift_out[2]
port 7 nsew default tristate
rlabel metal3 s 0 18776 800 18896 6 shift_out[3]
port 8 nsew default tristate
rlabel metal2 s 386 0 442 800 6 wb_clk_i
port 9 nsew default input
rlabel metal2 s 1214 0 1270 800 6 wb_rst_i
port 10 nsew default input
rlabel metal2 s 938 19162 994 19962 6 wbs_ack_o
port 11 nsew default tristate
rlabel metal2 s 36634 0 36690 800 6 wbs_addr_i[0]
port 12 nsew default input
rlabel metal2 s 45558 0 45614 800 6 wbs_addr_i[10]
port 13 nsew default input
rlabel metal2 s 46386 0 46442 800 6 wbs_addr_i[11]
port 14 nsew default input
rlabel metal2 s 47306 0 47362 800 6 wbs_addr_i[12]
port 15 nsew default input
rlabel metal2 s 48226 0 48282 800 6 wbs_addr_i[13]
port 16 nsew default input
rlabel metal2 s 49054 0 49110 800 6 wbs_addr_i[14]
port 17 nsew default input
rlabel metal2 s 49974 0 50030 800 6 wbs_addr_i[15]
port 18 nsew default input
rlabel metal2 s 50802 0 50858 800 6 wbs_addr_i[16]
port 19 nsew default input
rlabel metal2 s 51722 0 51778 800 6 wbs_addr_i[17]
port 20 nsew default input
rlabel metal2 s 52642 0 52698 800 6 wbs_addr_i[18]
port 21 nsew default input
rlabel metal2 s 53470 0 53526 800 6 wbs_addr_i[19]
port 22 nsew default input
rlabel metal2 s 37554 0 37610 800 6 wbs_addr_i[1]
port 23 nsew default input
rlabel metal2 s 54390 0 54446 800 6 wbs_addr_i[20]
port 24 nsew default input
rlabel metal2 s 55310 0 55366 800 6 wbs_addr_i[21]
port 25 nsew default input
rlabel metal2 s 56138 0 56194 800 6 wbs_addr_i[22]
port 26 nsew default input
rlabel metal2 s 57058 0 57114 800 6 wbs_addr_i[23]
port 27 nsew default input
rlabel metal2 s 57886 0 57942 800 6 wbs_addr_i[24]
port 28 nsew default input
rlabel metal2 s 58806 0 58862 800 6 wbs_addr_i[25]
port 29 nsew default input
rlabel metal2 s 59726 0 59782 800 6 wbs_addr_i[26]
port 30 nsew default input
rlabel metal2 s 60554 0 60610 800 6 wbs_addr_i[27]
port 31 nsew default input
rlabel metal2 s 61474 0 61530 800 6 wbs_addr_i[28]
port 32 nsew default input
rlabel metal2 s 62394 0 62450 800 6 wbs_addr_i[29]
port 33 nsew default input
rlabel metal2 s 38474 0 38530 800 6 wbs_addr_i[2]
port 34 nsew default input
rlabel metal2 s 63222 0 63278 800 6 wbs_addr_i[30]
port 35 nsew default input
rlabel metal2 s 64142 0 64198 800 6 wbs_addr_i[31]
port 36 nsew default input
rlabel metal2 s 39302 0 39358 800 6 wbs_addr_i[3]
port 37 nsew default input
rlabel metal2 s 40222 0 40278 800 6 wbs_addr_i[4]
port 38 nsew default input
rlabel metal2 s 41050 0 41106 800 6 wbs_addr_i[5]
port 39 nsew default input
rlabel metal2 s 41970 0 42026 800 6 wbs_addr_i[6]
port 40 nsew default input
rlabel metal2 s 42890 0 42946 800 6 wbs_addr_i[7]
port 41 nsew default input
rlabel metal2 s 43718 0 43774 800 6 wbs_addr_i[8]
port 42 nsew default input
rlabel metal2 s 44638 0 44694 800 6 wbs_addr_i[9]
port 43 nsew default input
rlabel metal2 s 2962 0 3018 800 6 wbs_cyc_i
port 44 nsew default input
rlabel metal2 s 8298 0 8354 800 6 wbs_data_i[0]
port 45 nsew default input
rlabel metal2 s 17130 0 17186 800 6 wbs_data_i[10]
port 46 nsew default input
rlabel metal2 s 18050 0 18106 800 6 wbs_data_i[11]
port 47 nsew default input
rlabel metal2 s 18970 0 19026 800 6 wbs_data_i[12]
port 48 nsew default input
rlabel metal2 s 19798 0 19854 800 6 wbs_data_i[13]
port 49 nsew default input
rlabel metal2 s 20718 0 20774 800 6 wbs_data_i[14]
port 50 nsew default input
rlabel metal2 s 21638 0 21694 800 6 wbs_data_i[15]
port 51 nsew default input
rlabel metal2 s 22466 0 22522 800 6 wbs_data_i[16]
port 52 nsew default input
rlabel metal2 s 23386 0 23442 800 6 wbs_data_i[17]
port 53 nsew default input
rlabel metal2 s 24306 0 24362 800 6 wbs_data_i[18]
port 54 nsew default input
rlabel metal2 s 25134 0 25190 800 6 wbs_data_i[19]
port 55 nsew default input
rlabel metal2 s 9218 0 9274 800 6 wbs_data_i[1]
port 56 nsew default input
rlabel metal2 s 26054 0 26110 800 6 wbs_data_i[20]
port 57 nsew default input
rlabel metal2 s 26882 0 26938 800 6 wbs_data_i[21]
port 58 nsew default input
rlabel metal2 s 27802 0 27858 800 6 wbs_data_i[22]
port 59 nsew default input
rlabel metal2 s 28722 0 28778 800 6 wbs_data_i[23]
port 60 nsew default input
rlabel metal2 s 29550 0 29606 800 6 wbs_data_i[24]
port 61 nsew default input
rlabel metal2 s 30470 0 30526 800 6 wbs_data_i[25]
port 62 nsew default input
rlabel metal2 s 31390 0 31446 800 6 wbs_data_i[26]
port 63 nsew default input
rlabel metal2 s 32218 0 32274 800 6 wbs_data_i[27]
port 64 nsew default input
rlabel metal2 s 33138 0 33194 800 6 wbs_data_i[28]
port 65 nsew default input
rlabel metal2 s 33966 0 34022 800 6 wbs_data_i[29]
port 66 nsew default input
rlabel metal2 s 10046 0 10102 800 6 wbs_data_i[2]
port 67 nsew default input
rlabel metal2 s 34886 0 34942 800 6 wbs_data_i[30]
port 68 nsew default input
rlabel metal2 s 35806 0 35862 800 6 wbs_data_i[31]
port 69 nsew default input
rlabel metal2 s 10966 0 11022 800 6 wbs_data_i[3]
port 70 nsew default input
rlabel metal2 s 11886 0 11942 800 6 wbs_data_i[4]
port 71 nsew default input
rlabel metal2 s 12714 0 12770 800 6 wbs_data_i[5]
port 72 nsew default input
rlabel metal2 s 13634 0 13690 800 6 wbs_data_i[6]
port 73 nsew default input
rlabel metal2 s 14554 0 14610 800 6 wbs_data_i[7]
port 74 nsew default input
rlabel metal2 s 15382 0 15438 800 6 wbs_data_i[8]
port 75 nsew default input
rlabel metal2 s 16302 0 16358 800 6 wbs_data_i[9]
port 76 nsew default input
rlabel metal2 s 2870 19162 2926 19962 6 wbs_data_o[0]
port 77 nsew default tristate
rlabel metal2 s 22466 19162 22522 19962 6 wbs_data_o[10]
port 78 nsew default tristate
rlabel metal2 s 24398 19162 24454 19962 6 wbs_data_o[11]
port 79 nsew default tristate
rlabel metal2 s 26330 19162 26386 19962 6 wbs_data_o[12]
port 80 nsew default tristate
rlabel metal2 s 28354 19162 28410 19962 6 wbs_data_o[13]
port 81 nsew default tristate
rlabel metal2 s 30286 19162 30342 19962 6 wbs_data_o[14]
port 82 nsew default tristate
rlabel metal2 s 32218 19162 32274 19962 6 wbs_data_o[15]
port 83 nsew default tristate
rlabel metal2 s 34242 19162 34298 19962 6 wbs_data_o[16]
port 84 nsew default tristate
rlabel metal2 s 36174 19162 36230 19962 6 wbs_data_o[17]
port 85 nsew default tristate
rlabel metal2 s 38106 19162 38162 19962 6 wbs_data_o[18]
port 86 nsew default tristate
rlabel metal2 s 40130 19162 40186 19962 6 wbs_data_o[19]
port 87 nsew default tristate
rlabel metal2 s 4802 19162 4858 19962 6 wbs_data_o[1]
port 88 nsew default tristate
rlabel metal2 s 42062 19162 42118 19962 6 wbs_data_o[20]
port 89 nsew default tristate
rlabel metal2 s 43994 19162 44050 19962 6 wbs_data_o[21]
port 90 nsew default tristate
rlabel metal2 s 45926 19162 45982 19962 6 wbs_data_o[22]
port 91 nsew default tristate
rlabel metal2 s 47950 19162 48006 19962 6 wbs_data_o[23]
port 92 nsew default tristate
rlabel metal2 s 49882 19162 49938 19962 6 wbs_data_o[24]
port 93 nsew default tristate
rlabel metal2 s 51814 19162 51870 19962 6 wbs_data_o[25]
port 94 nsew default tristate
rlabel metal2 s 53838 19162 53894 19962 6 wbs_data_o[26]
port 95 nsew default tristate
rlabel metal2 s 55770 19162 55826 19962 6 wbs_data_o[27]
port 96 nsew default tristate
rlabel metal2 s 57702 19162 57758 19962 6 wbs_data_o[28]
port 97 nsew default tristate
rlabel metal2 s 59726 19162 59782 19962 6 wbs_data_o[29]
port 98 nsew default tristate
rlabel metal2 s 6734 19162 6790 19962 6 wbs_data_o[2]
port 99 nsew default tristate
rlabel metal2 s 61658 19162 61714 19962 6 wbs_data_o[30]
port 100 nsew default tristate
rlabel metal2 s 63590 19162 63646 19962 6 wbs_data_o[31]
port 101 nsew default tristate
rlabel metal2 s 8758 19162 8814 19962 6 wbs_data_o[3]
port 102 nsew default tristate
rlabel metal2 s 10690 19162 10746 19962 6 wbs_data_o[4]
port 103 nsew default tristate
rlabel metal2 s 12622 19162 12678 19962 6 wbs_data_o[5]
port 104 nsew default tristate
rlabel metal2 s 14646 19162 14702 19962 6 wbs_data_o[6]
port 105 nsew default tristate
rlabel metal2 s 16578 19162 16634 19962 6 wbs_data_o[7]
port 106 nsew default tristate
rlabel metal2 s 18510 19162 18566 19962 6 wbs_data_o[8]
port 107 nsew default tristate
rlabel metal2 s 20534 19162 20590 19962 6 wbs_data_o[9]
port 108 nsew default tristate
rlabel metal2 s 4802 0 4858 800 6 wbs_sel_i[0]
port 109 nsew default input
rlabel metal2 s 5630 0 5686 800 6 wbs_sel_i[1]
port 110 nsew default input
rlabel metal2 s 6550 0 6606 800 6 wbs_sel_i[2]
port 111 nsew default input
rlabel metal2 s 7470 0 7526 800 6 wbs_sel_i[3]
port 112 nsew default input
rlabel metal2 s 2134 0 2190 800 6 wbs_stb_i
port 113 nsew default input
rlabel metal2 s 3882 0 3938 800 6 wbs_we_i
port 114 nsew default input
rlabel metal4 s 11340 2128 11660 17456 6 VPWR
port 115 nsew default input
rlabel metal4 s 21736 2128 22056 17456 6 VGND
port 116 nsew default input
<< properties >>
string FIXED_BBOX 0 0 64202 19962
<< end >>

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga
  CLASS BLOCK ;
  FOREIGN fpga ;
  ORIGIN 0.000 0.000 ;
  SIZE 2850.000 BY 3400.000 ;
  PIN gpio_east[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 60.560 2850.000 61.160 ;
    END
  END gpio_east[0]
  PIN gpio_east[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 181.600 2850.000 182.200 ;
    END
  END gpio_east[1]
  PIN gpio_east[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 303.320 2850.000 303.920 ;
    END
  END gpio_east[2]
  PIN gpio_east[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 424.360 2850.000 424.960 ;
    END
  END gpio_east[3]
  PIN gpio_east[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 546.080 2850.000 546.680 ;
    END
  END gpio_east[4]
  PIN gpio_east[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 667.120 2850.000 667.720 ;
    END
  END gpio_east[5]
  PIN gpio_east[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 788.840 2850.000 789.440 ;
    END
  END gpio_east[6]
  PIN gpio_east[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 910.560 2850.000 911.160 ;
    END
  END gpio_east[7]
  PIN gpio_east[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1031.600 2850.000 1032.200 ;
    END
  END gpio_east[8]
  PIN gpio_east[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1153.320 2850.000 1153.920 ;
    END
  END gpio_east[9]
  PIN gpio_north[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 52.530 3396.000 52.810 3400.000 ;
    END
  END gpio_north[0]
  PIN gpio_north[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 157.870 3396.000 158.150 3400.000 ;
    END
  END gpio_north[1]
  PIN gpio_north[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 263.210 3396.000 263.490 3400.000 ;
    END
  END gpio_north[2]
  PIN gpio_north[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 369.010 3396.000 369.290 3400.000 ;
    END
  END gpio_north[3]
  PIN gpio_north[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 474.350 3396.000 474.630 3400.000 ;
    END
  END gpio_north[4]
  PIN gpio_north[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 580.150 3396.000 580.430 3400.000 ;
    END
  END gpio_north[5]
  PIN gpio_north[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 685.490 3396.000 685.770 3400.000 ;
    END
  END gpio_north[6]
  PIN gpio_north[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 791.290 3396.000 791.570 3400.000 ;
    END
  END gpio_north[7]
  PIN gpio_north[8]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 896.630 3396.000 896.910 3400.000 ;
    END
  END gpio_north[8]
  PIN gpio_north[9]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1002.430 3396.000 1002.710 3400.000 ;
    END
  END gpio_north[9]
  PIN gpio_south[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END gpio_south[0]
  PIN gpio_south[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END gpio_south[1]
  PIN gpio_south[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END gpio_south[2]
  PIN gpio_south[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 177.650 0.000 177.930 4.000 ;
    END
  END gpio_south[3]
  PIN gpio_south[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END gpio_south[4]
  PIN gpio_south[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END gpio_south[5]
  PIN gpio_south[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 330.370 0.000 330.650 4.000 ;
    END
  END gpio_south[6]
  PIN gpio_south[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 381.430 0.000 381.710 4.000 ;
    END
  END gpio_south[7]
  PIN gpio_west[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END gpio_west[0]
  PIN gpio_west[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END gpio_west[1]
  PIN gpio_west[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END gpio_west[2]
  PIN gpio_west[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.760 4.000 360.360 ;
    END
  END gpio_west[3]
  PIN gpio_west[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.120 4.000 463.720 ;
    END
  END gpio_west[4]
  PIN gpio_west[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 565.800 4.000 566.400 ;
    END
  END gpio_west[5]
  PIN gpio_west[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.160 4.000 669.760 ;
    END
  END gpio_west[6]
  PIN gpio_west[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 771.840 4.000 772.440 ;
    END
  END gpio_west[7]
  PIN gpio_west[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 875.200 4.000 875.800 ;
    END
  END gpio_west[8]
  PIN gpio_west[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 977.880 4.000 978.480 ;
    END
  END gpio_west[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2060.890 0.000 2061.170 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1107.770 3396.000 1108.050 3400.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2111.950 0.000 2112.230 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_addr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1081.240 4.000 1081.840 ;
    END
  END wbs_addr_i[0]
  PIN wbs_addr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2213.610 0.000 2213.890 4.000 ;
    END
  END wbs_addr_i[10]
  PIN wbs_addr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1596.000 4.000 1596.600 ;
    END
  END wbs_addr_i[11]
  PIN wbs_addr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1699.360 4.000 1699.960 ;
    END
  END wbs_addr_i[12]
  PIN wbs_addr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1424.710 3396.000 1424.990 3400.000 ;
    END
  END wbs_addr_i[13]
  PIN wbs_addr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1530.050 3396.000 1530.330 3400.000 ;
    END
  END wbs_addr_i[14]
  PIN wbs_addr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2264.670 0.000 2264.950 4.000 ;
    END
  END wbs_addr_i[15]
  PIN wbs_addr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2315.270 0.000 2315.550 4.000 ;
    END
  END wbs_addr_i[16]
  PIN wbs_addr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2366.330 0.000 2366.610 4.000 ;
    END
  END wbs_addr_i[17]
  PIN wbs_addr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1635.850 3396.000 1636.130 3400.000 ;
    END
  END wbs_addr_i[18]
  PIN wbs_addr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1741.190 3396.000 1741.470 3400.000 ;
    END
  END wbs_addr_i[19]
  PIN wbs_addr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2163.010 0.000 2163.290 4.000 ;
    END
  END wbs_addr_i[1]
  PIN wbs_addr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2417.390 0.000 2417.670 4.000 ;
    END
  END wbs_addr_i[20]
  PIN wbs_addr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1802.040 4.000 1802.640 ;
    END
  END wbs_addr_i[21]
  PIN wbs_addr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1905.400 4.000 1906.000 ;
    END
  END wbs_addr_i[22]
  PIN wbs_addr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1517.120 2850.000 1517.720 ;
    END
  END wbs_addr_i[23]
  PIN wbs_addr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2467.990 0.000 2468.270 4.000 ;
    END
  END wbs_addr_i[24]
  PIN wbs_addr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2008.080 4.000 2008.680 ;
    END
  END wbs_addr_i[25]
  PIN wbs_addr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2111.440 4.000 2112.040 ;
    END
  END wbs_addr_i[26]
  PIN wbs_addr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1638.840 2850.000 1639.440 ;
    END
  END wbs_addr_i[27]
  PIN wbs_addr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1760.560 2850.000 1761.160 ;
    END
  END wbs_addr_i[28]
  PIN wbs_addr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2214.120 4.000 2214.720 ;
    END
  END wbs_addr_i[29]
  PIN wbs_addr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1213.570 3396.000 1213.850 3400.000 ;
    END
  END wbs_addr_i[2]
  PIN wbs_addr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1881.600 2850.000 1882.200 ;
    END
  END wbs_addr_i[30]
  PIN wbs_addr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2317.480 4.000 2318.080 ;
    END
  END wbs_addr_i[31]
  PIN wbs_addr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1318.910 3396.000 1319.190 3400.000 ;
    END
  END wbs_addr_i[3]
  PIN wbs_addr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1183.920 4.000 1184.520 ;
    END
  END wbs_addr_i[4]
  PIN wbs_addr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1274.360 2850.000 1274.960 ;
    END
  END wbs_addr_i[5]
  PIN wbs_addr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1396.080 2850.000 1396.680 ;
    END
  END wbs_addr_i[6]
  PIN wbs_addr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1287.280 4.000 1287.880 ;
    END
  END wbs_addr_i[7]
  PIN wbs_addr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1389.960 4.000 1390.560 ;
    END
  END wbs_addr_i[8]
  PIN wbs_addr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1493.320 4.000 1493.920 ;
    END
  END wbs_addr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1846.990 3396.000 1847.270 3400.000 ;
    END
  END wbs_cyc_i
  PIN wbs_data_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2420.160 4.000 2420.760 ;
    END
  END wbs_data_i[0]
  PIN wbs_data_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2626.200 4.000 2626.800 ;
    END
  END wbs_data_i[10]
  PIN wbs_data_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2367.120 2850.000 2367.720 ;
    END
  END wbs_data_i[11]
  PIN wbs_data_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2488.840 2850.000 2489.440 ;
    END
  END wbs_data_i[12]
  PIN wbs_data_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2163.470 3396.000 2163.750 3400.000 ;
    END
  END wbs_data_i[13]
  PIN wbs_data_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2671.770 0.000 2672.050 4.000 ;
    END
  END wbs_data_i[14]
  PIN wbs_data_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2269.270 3396.000 2269.550 3400.000 ;
    END
  END wbs_data_i[15]
  PIN wbs_data_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2729.560 4.000 2730.160 ;
    END
  END wbs_data_i[16]
  PIN wbs_data_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2374.610 3396.000 2374.890 3400.000 ;
    END
  END wbs_data_i[17]
  PIN wbs_data_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2480.410 3396.000 2480.690 3400.000 ;
    END
  END wbs_data_i[18]
  PIN wbs_data_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2610.560 2850.000 2611.160 ;
    END
  END wbs_data_i[19]
  PIN wbs_data_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2519.050 0.000 2519.330 4.000 ;
    END
  END wbs_data_i[1]
  PIN wbs_data_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2731.600 2850.000 2732.200 ;
    END
  END wbs_data_i[20]
  PIN wbs_data_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2832.240 4.000 2832.840 ;
    END
  END wbs_data_i[21]
  PIN wbs_data_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2853.320 2850.000 2853.920 ;
    END
  END wbs_data_i[22]
  PIN wbs_data_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2974.360 2850.000 2974.960 ;
    END
  END wbs_data_i[23]
  PIN wbs_data_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 3096.080 2850.000 3096.680 ;
    END
  END wbs_data_i[24]
  PIN wbs_data_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2722.830 0.000 2723.110 4.000 ;
    END
  END wbs_data_i[25]
  PIN wbs_data_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2585.750 3396.000 2586.030 3400.000 ;
    END
  END wbs_data_i[26]
  PIN wbs_data_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2691.550 3396.000 2691.830 3400.000 ;
    END
  END wbs_data_i[27]
  PIN wbs_data_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2773.430 0.000 2773.710 4.000 ;
    END
  END wbs_data_i[28]
  PIN wbs_data_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2935.600 4.000 2936.200 ;
    END
  END wbs_data_i[29]
  PIN wbs_data_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1952.330 3396.000 1952.610 3400.000 ;
    END
  END wbs_data_i[2]
  PIN wbs_data_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3038.280 4.000 3038.880 ;
    END
  END wbs_data_i[30]
  PIN wbs_data_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3141.640 4.000 3142.240 ;
    END
  END wbs_data_i[31]
  PIN wbs_data_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2058.130 3396.000 2058.410 3400.000 ;
    END
  END wbs_data_i[3]
  PIN wbs_data_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2003.320 2850.000 2003.920 ;
    END
  END wbs_data_i[4]
  PIN wbs_data_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2124.360 2850.000 2124.960 ;
    END
  END wbs_data_i[5]
  PIN wbs_data_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2570.110 0.000 2570.390 4.000 ;
    END
  END wbs_data_i[6]
  PIN wbs_data_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2620.710 0.000 2620.990 4.000 ;
    END
  END wbs_data_i[7]
  PIN wbs_data_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2246.080 2850.000 2246.680 ;
    END
  END wbs_data_i[8]
  PIN wbs_data_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2523.520 4.000 2524.120 ;
    END
  END wbs_data_i[9]
  PIN wbs_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 432.490 0.000 432.770 4.000 ;
    END
  END wbs_data_o[0]
  PIN wbs_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 941.250 0.000 941.530 4.000 ;
    END
  END wbs_data_o[10]
  PIN wbs_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 992.310 0.000 992.590 4.000 ;
    END
  END wbs_data_o[11]
  PIN wbs_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1042.910 0.000 1043.190 4.000 ;
    END
  END wbs_data_o[12]
  PIN wbs_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1093.970 0.000 1094.250 4.000 ;
    END
  END wbs_data_o[13]
  PIN wbs_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1145.030 0.000 1145.310 4.000 ;
    END
  END wbs_data_o[14]
  PIN wbs_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1195.630 0.000 1195.910 4.000 ;
    END
  END wbs_data_o[15]
  PIN wbs_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1246.690 0.000 1246.970 4.000 ;
    END
  END wbs_data_o[16]
  PIN wbs_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1297.750 0.000 1298.030 4.000 ;
    END
  END wbs_data_o[17]
  PIN wbs_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1348.350 0.000 1348.630 4.000 ;
    END
  END wbs_data_o[18]
  PIN wbs_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1399.410 0.000 1399.690 4.000 ;
    END
  END wbs_data_o[19]
  PIN wbs_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END wbs_data_o[1]
  PIN wbs_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1450.470 0.000 1450.750 4.000 ;
    END
  END wbs_data_o[20]
  PIN wbs_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1501.070 0.000 1501.350 4.000 ;
    END
  END wbs_data_o[21]
  PIN wbs_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1552.130 0.000 1552.410 4.000 ;
    END
  END wbs_data_o[22]
  PIN wbs_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1602.730 0.000 1603.010 4.000 ;
    END
  END wbs_data_o[23]
  PIN wbs_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1653.790 0.000 1654.070 4.000 ;
    END
  END wbs_data_o[24]
  PIN wbs_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1704.850 0.000 1705.130 4.000 ;
    END
  END wbs_data_o[25]
  PIN wbs_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1755.450 0.000 1755.730 4.000 ;
    END
  END wbs_data_o[26]
  PIN wbs_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1806.510 0.000 1806.790 4.000 ;
    END
  END wbs_data_o[27]
  PIN wbs_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1857.570 0.000 1857.850 4.000 ;
    END
  END wbs_data_o[28]
  PIN wbs_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1908.170 0.000 1908.450 4.000 ;
    END
  END wbs_data_o[29]
  PIN wbs_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 534.150 0.000 534.430 4.000 ;
    END
  END wbs_data_o[2]
  PIN wbs_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1959.230 0.000 1959.510 4.000 ;
    END
  END wbs_data_o[30]
  PIN wbs_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2010.290 0.000 2010.570 4.000 ;
    END
  END wbs_data_o[31]
  PIN wbs_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 585.210 0.000 585.490 4.000 ;
    END
  END wbs_data_o[3]
  PIN wbs_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 635.810 0.000 636.090 4.000 ;
    END
  END wbs_data_o[4]
  PIN wbs_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 686.870 0.000 687.150 4.000 ;
    END
  END wbs_data_o[5]
  PIN wbs_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 737.930 0.000 738.210 4.000 ;
    END
  END wbs_data_o[6]
  PIN wbs_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 788.530 0.000 788.810 4.000 ;
    END
  END wbs_data_o[7]
  PIN wbs_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 839.590 0.000 839.870 4.000 ;
    END
  END wbs_data_o[8]
  PIN wbs_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 890.190 0.000 890.470 4.000 ;
    END
  END wbs_data_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3244.320 4.000 3244.920 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3347.680 4.000 3348.280 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 3217.120 2850.000 3217.720 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2796.890 3396.000 2797.170 3400.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 3338.840 2850.000 3339.440 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2824.490 0.000 2824.770 4.000 ;
    END
  END wbs_we_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 2844.180 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 64.785 2844.180 66.385 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2844.180 3389.205 ;
      LAYER met1 ;
        RECT 5.520 10.640 2844.180 3389.360 ;
      LAYER met2 ;
        RECT 13.780 3395.720 52.250 3396.000 ;
        RECT 53.090 3395.720 157.590 3396.000 ;
        RECT 158.430 3395.720 262.930 3396.000 ;
        RECT 263.770 3395.720 368.730 3396.000 ;
        RECT 369.570 3395.720 474.070 3396.000 ;
        RECT 474.910 3395.720 579.870 3396.000 ;
        RECT 580.710 3395.720 685.210 3396.000 ;
        RECT 686.050 3395.720 791.010 3396.000 ;
        RECT 791.850 3395.720 896.350 3396.000 ;
        RECT 897.190 3395.720 1002.150 3396.000 ;
        RECT 1002.990 3395.720 1107.490 3396.000 ;
        RECT 1108.330 3395.720 1213.290 3396.000 ;
        RECT 1214.130 3395.720 1318.630 3396.000 ;
        RECT 1319.470 3395.720 1424.430 3396.000 ;
        RECT 1425.270 3395.720 1529.770 3396.000 ;
        RECT 1530.610 3395.720 1635.570 3396.000 ;
        RECT 1636.410 3395.720 1740.910 3396.000 ;
        RECT 1741.750 3395.720 1846.710 3396.000 ;
        RECT 1847.550 3395.720 1952.050 3396.000 ;
        RECT 1952.890 3395.720 2057.850 3396.000 ;
        RECT 2058.690 3395.720 2163.190 3396.000 ;
        RECT 2164.030 3395.720 2268.990 3396.000 ;
        RECT 2269.830 3395.720 2374.330 3396.000 ;
        RECT 2375.170 3395.720 2480.130 3396.000 ;
        RECT 2480.970 3395.720 2585.470 3396.000 ;
        RECT 2586.310 3395.720 2691.270 3396.000 ;
        RECT 2692.110 3395.720 2796.610 3396.000 ;
        RECT 2797.450 3395.720 2835.810 3396.000 ;
        RECT 13.780 4.280 2835.810 3395.720 ;
        RECT 13.780 4.000 25.110 4.280 ;
        RECT 25.950 4.000 75.710 4.280 ;
        RECT 76.550 4.000 126.770 4.280 ;
        RECT 127.610 4.000 177.370 4.280 ;
        RECT 178.210 4.000 228.430 4.280 ;
        RECT 229.270 4.000 279.490 4.280 ;
        RECT 280.330 4.000 330.090 4.280 ;
        RECT 330.930 4.000 381.150 4.280 ;
        RECT 381.990 4.000 432.210 4.280 ;
        RECT 433.050 4.000 482.810 4.280 ;
        RECT 483.650 4.000 533.870 4.280 ;
        RECT 534.710 4.000 584.930 4.280 ;
        RECT 585.770 4.000 635.530 4.280 ;
        RECT 636.370 4.000 686.590 4.280 ;
        RECT 687.430 4.000 737.650 4.280 ;
        RECT 738.490 4.000 788.250 4.280 ;
        RECT 789.090 4.000 839.310 4.280 ;
        RECT 840.150 4.000 889.910 4.280 ;
        RECT 890.750 4.000 940.970 4.280 ;
        RECT 941.810 4.000 992.030 4.280 ;
        RECT 992.870 4.000 1042.630 4.280 ;
        RECT 1043.470 4.000 1093.690 4.280 ;
        RECT 1094.530 4.000 1144.750 4.280 ;
        RECT 1145.590 4.000 1195.350 4.280 ;
        RECT 1196.190 4.000 1246.410 4.280 ;
        RECT 1247.250 4.000 1297.470 4.280 ;
        RECT 1298.310 4.000 1348.070 4.280 ;
        RECT 1348.910 4.000 1399.130 4.280 ;
        RECT 1399.970 4.000 1450.190 4.280 ;
        RECT 1451.030 4.000 1500.790 4.280 ;
        RECT 1501.630 4.000 1551.850 4.280 ;
        RECT 1552.690 4.000 1602.450 4.280 ;
        RECT 1603.290 4.000 1653.510 4.280 ;
        RECT 1654.350 4.000 1704.570 4.280 ;
        RECT 1705.410 4.000 1755.170 4.280 ;
        RECT 1756.010 4.000 1806.230 4.280 ;
        RECT 1807.070 4.000 1857.290 4.280 ;
        RECT 1858.130 4.000 1907.890 4.280 ;
        RECT 1908.730 4.000 1958.950 4.280 ;
        RECT 1959.790 4.000 2010.010 4.280 ;
        RECT 2010.850 4.000 2060.610 4.280 ;
        RECT 2061.450 4.000 2111.670 4.280 ;
        RECT 2112.510 4.000 2162.730 4.280 ;
        RECT 2163.570 4.000 2213.330 4.280 ;
        RECT 2214.170 4.000 2264.390 4.280 ;
        RECT 2265.230 4.000 2314.990 4.280 ;
        RECT 2315.830 4.000 2366.050 4.280 ;
        RECT 2366.890 4.000 2417.110 4.280 ;
        RECT 2417.950 4.000 2467.710 4.280 ;
        RECT 2468.550 4.000 2518.770 4.280 ;
        RECT 2519.610 4.000 2569.830 4.280 ;
        RECT 2570.670 4.000 2620.430 4.280 ;
        RECT 2621.270 4.000 2671.490 4.280 ;
        RECT 2672.330 4.000 2722.550 4.280 ;
        RECT 2723.390 4.000 2773.150 4.280 ;
        RECT 2773.990 4.000 2824.210 4.280 ;
        RECT 2825.050 4.000 2835.810 4.280 ;
      LAYER met3 ;
        RECT 4.000 3348.680 2846.000 3389.285 ;
        RECT 4.400 3347.280 2846.000 3348.680 ;
        RECT 4.000 3339.840 2846.000 3347.280 ;
        RECT 4.000 3338.440 2845.600 3339.840 ;
        RECT 4.000 3245.320 2846.000 3338.440 ;
        RECT 4.400 3243.920 2846.000 3245.320 ;
        RECT 4.000 3218.120 2846.000 3243.920 ;
        RECT 4.000 3216.720 2845.600 3218.120 ;
        RECT 4.000 3142.640 2846.000 3216.720 ;
        RECT 4.400 3141.240 2846.000 3142.640 ;
        RECT 4.000 3097.080 2846.000 3141.240 ;
        RECT 4.000 3095.680 2845.600 3097.080 ;
        RECT 4.000 3039.280 2846.000 3095.680 ;
        RECT 4.400 3037.880 2846.000 3039.280 ;
        RECT 4.000 2975.360 2846.000 3037.880 ;
        RECT 4.000 2973.960 2845.600 2975.360 ;
        RECT 4.000 2936.600 2846.000 2973.960 ;
        RECT 4.400 2935.200 2846.000 2936.600 ;
        RECT 4.000 2854.320 2846.000 2935.200 ;
        RECT 4.000 2852.920 2845.600 2854.320 ;
        RECT 4.000 2833.240 2846.000 2852.920 ;
        RECT 4.400 2831.840 2846.000 2833.240 ;
        RECT 4.000 2732.600 2846.000 2831.840 ;
        RECT 4.000 2731.200 2845.600 2732.600 ;
        RECT 4.000 2730.560 2846.000 2731.200 ;
        RECT 4.400 2729.160 2846.000 2730.560 ;
        RECT 4.000 2627.200 2846.000 2729.160 ;
        RECT 4.400 2625.800 2846.000 2627.200 ;
        RECT 4.000 2611.560 2846.000 2625.800 ;
        RECT 4.000 2610.160 2845.600 2611.560 ;
        RECT 4.000 2524.520 2846.000 2610.160 ;
        RECT 4.400 2523.120 2846.000 2524.520 ;
        RECT 4.000 2489.840 2846.000 2523.120 ;
        RECT 4.000 2488.440 2845.600 2489.840 ;
        RECT 4.000 2421.160 2846.000 2488.440 ;
        RECT 4.400 2419.760 2846.000 2421.160 ;
        RECT 4.000 2368.120 2846.000 2419.760 ;
        RECT 4.000 2366.720 2845.600 2368.120 ;
        RECT 4.000 2318.480 2846.000 2366.720 ;
        RECT 4.400 2317.080 2846.000 2318.480 ;
        RECT 4.000 2247.080 2846.000 2317.080 ;
        RECT 4.000 2245.680 2845.600 2247.080 ;
        RECT 4.000 2215.120 2846.000 2245.680 ;
        RECT 4.400 2213.720 2846.000 2215.120 ;
        RECT 4.000 2125.360 2846.000 2213.720 ;
        RECT 4.000 2123.960 2845.600 2125.360 ;
        RECT 4.000 2112.440 2846.000 2123.960 ;
        RECT 4.400 2111.040 2846.000 2112.440 ;
        RECT 4.000 2009.080 2846.000 2111.040 ;
        RECT 4.400 2007.680 2846.000 2009.080 ;
        RECT 4.000 2004.320 2846.000 2007.680 ;
        RECT 4.000 2002.920 2845.600 2004.320 ;
        RECT 4.000 1906.400 2846.000 2002.920 ;
        RECT 4.400 1905.000 2846.000 1906.400 ;
        RECT 4.000 1882.600 2846.000 1905.000 ;
        RECT 4.000 1881.200 2845.600 1882.600 ;
        RECT 4.000 1803.040 2846.000 1881.200 ;
        RECT 4.400 1801.640 2846.000 1803.040 ;
        RECT 4.000 1761.560 2846.000 1801.640 ;
        RECT 4.000 1760.160 2845.600 1761.560 ;
        RECT 4.000 1700.360 2846.000 1760.160 ;
        RECT 4.400 1698.960 2846.000 1700.360 ;
        RECT 4.000 1639.840 2846.000 1698.960 ;
        RECT 4.000 1638.440 2845.600 1639.840 ;
        RECT 4.000 1597.000 2846.000 1638.440 ;
        RECT 4.400 1595.600 2846.000 1597.000 ;
        RECT 4.000 1518.120 2846.000 1595.600 ;
        RECT 4.000 1516.720 2845.600 1518.120 ;
        RECT 4.000 1494.320 2846.000 1516.720 ;
        RECT 4.400 1492.920 2846.000 1494.320 ;
        RECT 4.000 1397.080 2846.000 1492.920 ;
        RECT 4.000 1395.680 2845.600 1397.080 ;
        RECT 4.000 1390.960 2846.000 1395.680 ;
        RECT 4.400 1389.560 2846.000 1390.960 ;
        RECT 4.000 1288.280 2846.000 1389.560 ;
        RECT 4.400 1286.880 2846.000 1288.280 ;
        RECT 4.000 1275.360 2846.000 1286.880 ;
        RECT 4.000 1273.960 2845.600 1275.360 ;
        RECT 4.000 1184.920 2846.000 1273.960 ;
        RECT 4.400 1183.520 2846.000 1184.920 ;
        RECT 4.000 1154.320 2846.000 1183.520 ;
        RECT 4.000 1152.920 2845.600 1154.320 ;
        RECT 4.000 1082.240 2846.000 1152.920 ;
        RECT 4.400 1080.840 2846.000 1082.240 ;
        RECT 4.000 1032.600 2846.000 1080.840 ;
        RECT 4.000 1031.200 2845.600 1032.600 ;
        RECT 4.000 978.880 2846.000 1031.200 ;
        RECT 4.400 977.480 2846.000 978.880 ;
        RECT 4.000 911.560 2846.000 977.480 ;
        RECT 4.000 910.160 2845.600 911.560 ;
        RECT 4.000 876.200 2846.000 910.160 ;
        RECT 4.400 874.800 2846.000 876.200 ;
        RECT 4.000 789.840 2846.000 874.800 ;
        RECT 4.000 788.440 2845.600 789.840 ;
        RECT 4.000 772.840 2846.000 788.440 ;
        RECT 4.400 771.440 2846.000 772.840 ;
        RECT 4.000 670.160 2846.000 771.440 ;
        RECT 4.400 668.760 2846.000 670.160 ;
        RECT 4.000 668.120 2846.000 668.760 ;
        RECT 4.000 666.720 2845.600 668.120 ;
        RECT 4.000 566.800 2846.000 666.720 ;
        RECT 4.400 565.400 2846.000 566.800 ;
        RECT 4.000 547.080 2846.000 565.400 ;
        RECT 4.000 545.680 2845.600 547.080 ;
        RECT 4.000 464.120 2846.000 545.680 ;
        RECT 4.400 462.720 2846.000 464.120 ;
        RECT 4.000 425.360 2846.000 462.720 ;
        RECT 4.000 423.960 2845.600 425.360 ;
        RECT 4.000 360.760 2846.000 423.960 ;
        RECT 4.400 359.360 2846.000 360.760 ;
        RECT 4.000 304.320 2846.000 359.360 ;
        RECT 4.000 302.920 2845.600 304.320 ;
        RECT 4.000 258.080 2846.000 302.920 ;
        RECT 4.400 256.680 2846.000 258.080 ;
        RECT 4.000 182.600 2846.000 256.680 ;
        RECT 4.000 181.200 2845.600 182.600 ;
        RECT 4.000 154.720 2846.000 181.200 ;
        RECT 4.400 153.320 2846.000 154.720 ;
        RECT 4.000 61.560 2846.000 153.320 ;
        RECT 4.000 60.160 2845.600 61.560 ;
        RECT 4.000 52.040 2846.000 60.160 ;
        RECT 4.400 50.640 2846.000 52.040 ;
        RECT 4.000 10.715 2846.000 50.640 ;
      LAYER met4 ;
        RECT 13.720 10.640 2813.505 3389.360 ;
      LAYER met5 ;
        RECT 5.520 103.080 2844.180 3359.755 ;
  END
END fpga
END LIBRARY


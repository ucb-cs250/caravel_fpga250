VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga
  CLASS BLOCK ;
  FOREIGN fpga ;
  ORIGIN 0.000 0.000 ;
  SIZE 2850.000 BY 3400.000 ;
  PIN gpio_east[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 53.080 2850.000 53.680 ;
    END
  END gpio_east[0]
  PIN gpio_east[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 159.160 2850.000 159.760 ;
    END
  END gpio_east[1]
  PIN gpio_east[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 265.240 2850.000 265.840 ;
    END
  END gpio_east[2]
  PIN gpio_east[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 371.320 2850.000 371.920 ;
    END
  END gpio_east[3]
  PIN gpio_east[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 478.080 2850.000 478.680 ;
    END
  END gpio_east[4]
  PIN gpio_east[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 584.160 2850.000 584.760 ;
    END
  END gpio_east[5]
  PIN gpio_east[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 690.240 2850.000 690.840 ;
    END
  END gpio_east[6]
  PIN gpio_east[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 796.320 2850.000 796.920 ;
    END
  END gpio_east[7]
  PIN gpio_east[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 903.080 2850.000 903.680 ;
    END
  END gpio_east[8]
  PIN gpio_east[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1009.160 2850.000 1009.760 ;
    END
  END gpio_east[9]
  PIN gpio_north[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 70.930 3396.000 71.210 3400.000 ;
    END
  END gpio_north[0]
  PIN gpio_north[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 213.070 3396.000 213.350 3400.000 ;
    END
  END gpio_north[1]
  PIN gpio_north[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 355.670 3396.000 355.950 3400.000 ;
    END
  END gpio_north[2]
  PIN gpio_north[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 498.270 3396.000 498.550 3400.000 ;
    END
  END gpio_north[3]
  PIN gpio_north[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 640.870 3396.000 641.150 3400.000 ;
    END
  END gpio_north[4]
  PIN gpio_north[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 783.470 3396.000 783.750 3400.000 ;
    END
  END gpio_north[5]
  PIN gpio_north[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 925.610 3396.000 925.890 3400.000 ;
    END
  END gpio_north[6]
  PIN gpio_north[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1068.210 3396.000 1068.490 3400.000 ;
    END
  END gpio_north[7]
  PIN gpio_north[8]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1210.810 3396.000 1211.090 3400.000 ;
    END
  END gpio_north[8]
  PIN gpio_north[9]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1353.410 3396.000 1353.690 3400.000 ;
    END
  END gpio_north[9]
  PIN gpio_south[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END gpio_south[0]
  PIN gpio_south[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END gpio_south[1]
  PIN gpio_south[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END gpio_south[2]
  PIN gpio_south[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 168.910 0.000 169.190 4.000 ;
    END
  END gpio_south[3]
  PIN gpio_south[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END gpio_south[4]
  PIN gpio_south[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 265.510 0.000 265.790 4.000 ;
    END
  END gpio_south[5]
  PIN gpio_south[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 313.810 0.000 314.090 4.000 ;
    END
  END gpio_south[6]
  PIN gpio_south[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 362.110 0.000 362.390 4.000 ;
    END
  END gpio_south[7]
  PIN gpio_west[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END gpio_west[0]
  PIN gpio_west[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END gpio_west[1]
  PIN gpio_west[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END gpio_west[2]
  PIN gpio_west[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.760 4.000 360.360 ;
    END
  END gpio_west[3]
  PIN gpio_west[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.120 4.000 463.720 ;
    END
  END gpio_west[4]
  PIN gpio_west[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 565.800 4.000 566.400 ;
    END
  END gpio_west[5]
  PIN gpio_west[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.160 4.000 669.760 ;
    END
  END gpio_west[6]
  PIN gpio_west[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 771.840 4.000 772.440 ;
    END
  END gpio_west[7]
  PIN gpio_west[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 875.200 4.000 875.800 ;
    END
  END gpio_west[8]
  PIN gpio_west[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 977.880 4.000 978.480 ;
    END
  END gpio_west[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1115.240 2850.000 1115.840 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1956.010 0.000 1956.290 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2004.310 0.000 2004.590 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_addr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1221.320 2850.000 1221.920 ;
    END
  END wbs_addr_i[0]
  PIN wbs_addr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1540.240 2850.000 1540.840 ;
    END
  END wbs_addr_i[10]
  PIN wbs_addr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1389.960 4.000 1390.560 ;
    END
  END wbs_addr_i[11]
  PIN wbs_addr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1646.320 2850.000 1646.920 ;
    END
  END wbs_addr_i[12]
  PIN wbs_addr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2149.210 0.000 2149.490 4.000 ;
    END
  END wbs_addr_i[13]
  PIN wbs_addr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1780.750 3396.000 1781.030 3400.000 ;
    END
  END wbs_addr_i[14]
  PIN wbs_addr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1753.080 2850.000 1753.680 ;
    END
  END wbs_addr_i[15]
  PIN wbs_addr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1493.320 4.000 1493.920 ;
    END
  END wbs_addr_i[16]
  PIN wbs_addr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1596.000 4.000 1596.600 ;
    END
  END wbs_addr_i[17]
  PIN wbs_addr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1859.160 2850.000 1859.760 ;
    END
  END wbs_addr_i[18]
  PIN wbs_addr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1699.360 4.000 1699.960 ;
    END
  END wbs_addr_i[19]
  PIN wbs_addr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1496.010 3396.000 1496.290 3400.000 ;
    END
  END wbs_addr_i[1]
  PIN wbs_addr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1923.350 3396.000 1923.630 3400.000 ;
    END
  END wbs_addr_i[20]
  PIN wbs_addr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1965.240 2850.000 1965.840 ;
    END
  END wbs_addr_i[21]
  PIN wbs_addr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2065.950 3396.000 2066.230 3400.000 ;
    END
  END wbs_addr_i[22]
  PIN wbs_addr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1802.040 4.000 1802.640 ;
    END
  END wbs_addr_i[23]
  PIN wbs_addr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1905.400 4.000 1906.000 ;
    END
  END wbs_addr_i[24]
  PIN wbs_addr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2008.080 4.000 2008.680 ;
    END
  END wbs_addr_i[25]
  PIN wbs_addr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2071.320 2850.000 2071.920 ;
    END
  END wbs_addr_i[26]
  PIN wbs_addr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2178.080 2850.000 2178.680 ;
    END
  END wbs_addr_i[27]
  PIN wbs_addr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2111.440 4.000 2112.040 ;
    END
  END wbs_addr_i[28]
  PIN wbs_addr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2284.160 2850.000 2284.760 ;
    END
  END wbs_addr_i[29]
  PIN wbs_addr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1328.080 2850.000 1328.680 ;
    END
  END wbs_addr_i[2]
  PIN wbs_addr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2390.240 2850.000 2390.840 ;
    END
  END wbs_addr_i[30]
  PIN wbs_addr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2496.320 2850.000 2496.920 ;
    END
  END wbs_addr_i[31]
  PIN wbs_addr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1081.240 4.000 1081.840 ;
    END
  END wbs_addr_i[3]
  PIN wbs_addr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1638.150 3396.000 1638.430 3400.000 ;
    END
  END wbs_addr_i[4]
  PIN wbs_addr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1183.920 4.000 1184.520 ;
    END
  END wbs_addr_i[5]
  PIN wbs_addr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1434.160 2850.000 1434.760 ;
    END
  END wbs_addr_i[6]
  PIN wbs_addr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2052.610 0.000 2052.890 4.000 ;
    END
  END wbs_addr_i[7]
  PIN wbs_addr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1287.280 4.000 1287.880 ;
    END
  END wbs_addr_i[8]
  PIN wbs_addr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2100.910 0.000 2101.190 4.000 ;
    END
  END wbs_addr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2197.510 0.000 2197.790 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_data_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2245.810 0.000 2246.090 4.000 ;
    END
  END wbs_data_i[0]
  PIN wbs_data_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2350.690 3396.000 2350.970 3400.000 ;
    END
  END wbs_data_i[10]
  PIN wbs_data_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2493.290 3396.000 2493.570 3400.000 ;
    END
  END wbs_data_i[11]
  PIN wbs_data_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2523.520 4.000 2524.120 ;
    END
  END wbs_data_i[12]
  PIN wbs_data_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2439.010 0.000 2439.290 4.000 ;
    END
  END wbs_data_i[13]
  PIN wbs_data_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2815.240 2850.000 2815.840 ;
    END
  END wbs_data_i[14]
  PIN wbs_data_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2487.310 0.000 2487.590 4.000 ;
    END
  END wbs_data_i[15]
  PIN wbs_data_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2626.200 4.000 2626.800 ;
    END
  END wbs_data_i[16]
  PIN wbs_data_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2921.320 2850.000 2921.920 ;
    END
  END wbs_data_i[17]
  PIN wbs_data_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2635.890 3396.000 2636.170 3400.000 ;
    END
  END wbs_data_i[18]
  PIN wbs_data_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 3028.080 2850.000 3028.680 ;
    END
  END wbs_data_i[19]
  PIN wbs_data_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2214.120 4.000 2214.720 ;
    END
  END wbs_data_i[1]
  PIN wbs_data_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 3134.160 2850.000 3134.760 ;
    END
  END wbs_data_i[20]
  PIN wbs_data_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2729.560 4.000 2730.160 ;
    END
  END wbs_data_i[21]
  PIN wbs_data_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2535.610 0.000 2535.890 4.000 ;
    END
  END wbs_data_i[22]
  PIN wbs_data_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2832.240 4.000 2832.840 ;
    END
  END wbs_data_i[23]
  PIN wbs_data_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2583.910 0.000 2584.190 4.000 ;
    END
  END wbs_data_i[24]
  PIN wbs_data_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 3240.240 2850.000 3240.840 ;
    END
  END wbs_data_i[25]
  PIN wbs_data_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2935.600 4.000 2936.200 ;
    END
  END wbs_data_i[26]
  PIN wbs_data_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3038.280 4.000 3038.880 ;
    END
  END wbs_data_i[27]
  PIN wbs_data_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3141.640 4.000 3142.240 ;
    END
  END wbs_data_i[28]
  PIN wbs_data_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2632.210 0.000 2632.490 4.000 ;
    END
  END wbs_data_i[29]
  PIN wbs_data_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2317.480 4.000 2318.080 ;
    END
  END wbs_data_i[2]
  PIN wbs_data_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2680.510 0.000 2680.790 4.000 ;
    END
  END wbs_data_i[30]
  PIN wbs_data_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2728.810 0.000 2729.090 4.000 ;
    END
  END wbs_data_i[31]
  PIN wbs_data_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2420.160 4.000 2420.760 ;
    END
  END wbs_data_i[3]
  PIN wbs_data_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2603.080 2850.000 2603.680 ;
    END
  END wbs_data_i[4]
  PIN wbs_data_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2294.110 0.000 2294.390 4.000 ;
    END
  END wbs_data_i[5]
  PIN wbs_data_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2709.160 2850.000 2709.760 ;
    END
  END wbs_data_i[6]
  PIN wbs_data_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2342.410 0.000 2342.690 4.000 ;
    END
  END wbs_data_i[7]
  PIN wbs_data_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2390.710 0.000 2390.990 4.000 ;
    END
  END wbs_data_i[8]
  PIN wbs_data_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2208.550 3396.000 2208.830 3400.000 ;
    END
  END wbs_data_i[9]
  PIN wbs_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 410.410 0.000 410.690 4.000 ;
    END
  END wbs_data_o[0]
  PIN wbs_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 893.410 0.000 893.690 4.000 ;
    END
  END wbs_data_o[10]
  PIN wbs_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 941.710 0.000 941.990 4.000 ;
    END
  END wbs_data_o[11]
  PIN wbs_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 990.010 0.000 990.290 4.000 ;
    END
  END wbs_data_o[12]
  PIN wbs_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1038.310 0.000 1038.590 4.000 ;
    END
  END wbs_data_o[13]
  PIN wbs_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1086.610 0.000 1086.890 4.000 ;
    END
  END wbs_data_o[14]
  PIN wbs_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1134.910 0.000 1135.190 4.000 ;
    END
  END wbs_data_o[15]
  PIN wbs_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1183.210 0.000 1183.490 4.000 ;
    END
  END wbs_data_o[16]
  PIN wbs_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1231.510 0.000 1231.790 4.000 ;
    END
  END wbs_data_o[17]
  PIN wbs_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1279.810 0.000 1280.090 4.000 ;
    END
  END wbs_data_o[18]
  PIN wbs_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1328.110 0.000 1328.390 4.000 ;
    END
  END wbs_data_o[19]
  PIN wbs_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 458.710 0.000 458.990 4.000 ;
    END
  END wbs_data_o[1]
  PIN wbs_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1376.410 0.000 1376.690 4.000 ;
    END
  END wbs_data_o[20]
  PIN wbs_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1424.710 0.000 1424.990 4.000 ;
    END
  END wbs_data_o[21]
  PIN wbs_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1473.010 0.000 1473.290 4.000 ;
    END
  END wbs_data_o[22]
  PIN wbs_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1521.310 0.000 1521.590 4.000 ;
    END
  END wbs_data_o[23]
  PIN wbs_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1569.610 0.000 1569.890 4.000 ;
    END
  END wbs_data_o[24]
  PIN wbs_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1617.910 0.000 1618.190 4.000 ;
    END
  END wbs_data_o[25]
  PIN wbs_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1666.210 0.000 1666.490 4.000 ;
    END
  END wbs_data_o[26]
  PIN wbs_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1714.510 0.000 1714.790 4.000 ;
    END
  END wbs_data_o[27]
  PIN wbs_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1762.810 0.000 1763.090 4.000 ;
    END
  END wbs_data_o[28]
  PIN wbs_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1811.110 0.000 1811.390 4.000 ;
    END
  END wbs_data_o[29]
  PIN wbs_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 507.010 0.000 507.290 4.000 ;
    END
  END wbs_data_o[2]
  PIN wbs_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1859.410 0.000 1859.690 4.000 ;
    END
  END wbs_data_o[30]
  PIN wbs_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1907.710 0.000 1907.990 4.000 ;
    END
  END wbs_data_o[31]
  PIN wbs_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 555.310 0.000 555.590 4.000 ;
    END
  END wbs_data_o[3]
  PIN wbs_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 603.610 0.000 603.890 4.000 ;
    END
  END wbs_data_o[4]
  PIN wbs_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 651.910 0.000 652.190 4.000 ;
    END
  END wbs_data_o[5]
  PIN wbs_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 700.210 0.000 700.490 4.000 ;
    END
  END wbs_data_o[6]
  PIN wbs_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 748.510 0.000 748.790 4.000 ;
    END
  END wbs_data_o[7]
  PIN wbs_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 796.810 0.000 797.090 4.000 ;
    END
  END wbs_data_o[8]
  PIN wbs_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 845.110 0.000 845.390 4.000 ;
    END
  END wbs_data_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2778.490 3396.000 2778.770 3400.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 3346.320 2850.000 3346.920 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3244.320 4.000 3244.920 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2777.110 0.000 2777.390 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2825.410 0.000 2825.690 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3347.680 4.000 3348.280 ;
    END
  END wbs_we_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 2844.180 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 64.785 2844.180 66.385 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2844.180 3389.205 ;
      LAYER met1 ;
        RECT 5.520 10.640 2844.180 3389.360 ;
      LAYER met2 ;
        RECT 13.780 3395.720 70.650 3396.000 ;
        RECT 71.490 3395.720 212.790 3396.000 ;
        RECT 213.630 3395.720 355.390 3396.000 ;
        RECT 356.230 3395.720 497.990 3396.000 ;
        RECT 498.830 3395.720 640.590 3396.000 ;
        RECT 641.430 3395.720 783.190 3396.000 ;
        RECT 784.030 3395.720 925.330 3396.000 ;
        RECT 926.170 3395.720 1067.930 3396.000 ;
        RECT 1068.770 3395.720 1210.530 3396.000 ;
        RECT 1211.370 3395.720 1353.130 3396.000 ;
        RECT 1353.970 3395.720 1495.730 3396.000 ;
        RECT 1496.570 3395.720 1637.870 3396.000 ;
        RECT 1638.710 3395.720 1780.470 3396.000 ;
        RECT 1781.310 3395.720 1923.070 3396.000 ;
        RECT 1923.910 3395.720 2065.670 3396.000 ;
        RECT 2066.510 3395.720 2208.270 3396.000 ;
        RECT 2209.110 3395.720 2350.410 3396.000 ;
        RECT 2351.250 3395.720 2493.010 3396.000 ;
        RECT 2493.850 3395.720 2635.610 3396.000 ;
        RECT 2636.450 3395.720 2778.210 3396.000 ;
        RECT 2779.050 3395.720 2835.810 3396.000 ;
        RECT 13.780 4.280 2835.810 3395.720 ;
        RECT 13.780 4.000 23.730 4.280 ;
        RECT 24.570 4.000 72.030 4.280 ;
        RECT 72.870 4.000 120.330 4.280 ;
        RECT 121.170 4.000 168.630 4.280 ;
        RECT 169.470 4.000 216.930 4.280 ;
        RECT 217.770 4.000 265.230 4.280 ;
        RECT 266.070 4.000 313.530 4.280 ;
        RECT 314.370 4.000 361.830 4.280 ;
        RECT 362.670 4.000 410.130 4.280 ;
        RECT 410.970 4.000 458.430 4.280 ;
        RECT 459.270 4.000 506.730 4.280 ;
        RECT 507.570 4.000 555.030 4.280 ;
        RECT 555.870 4.000 603.330 4.280 ;
        RECT 604.170 4.000 651.630 4.280 ;
        RECT 652.470 4.000 699.930 4.280 ;
        RECT 700.770 4.000 748.230 4.280 ;
        RECT 749.070 4.000 796.530 4.280 ;
        RECT 797.370 4.000 844.830 4.280 ;
        RECT 845.670 4.000 893.130 4.280 ;
        RECT 893.970 4.000 941.430 4.280 ;
        RECT 942.270 4.000 989.730 4.280 ;
        RECT 990.570 4.000 1038.030 4.280 ;
        RECT 1038.870 4.000 1086.330 4.280 ;
        RECT 1087.170 4.000 1134.630 4.280 ;
        RECT 1135.470 4.000 1182.930 4.280 ;
        RECT 1183.770 4.000 1231.230 4.280 ;
        RECT 1232.070 4.000 1279.530 4.280 ;
        RECT 1280.370 4.000 1327.830 4.280 ;
        RECT 1328.670 4.000 1376.130 4.280 ;
        RECT 1376.970 4.000 1424.430 4.280 ;
        RECT 1425.270 4.000 1472.730 4.280 ;
        RECT 1473.570 4.000 1521.030 4.280 ;
        RECT 1521.870 4.000 1569.330 4.280 ;
        RECT 1570.170 4.000 1617.630 4.280 ;
        RECT 1618.470 4.000 1665.930 4.280 ;
        RECT 1666.770 4.000 1714.230 4.280 ;
        RECT 1715.070 4.000 1762.530 4.280 ;
        RECT 1763.370 4.000 1810.830 4.280 ;
        RECT 1811.670 4.000 1859.130 4.280 ;
        RECT 1859.970 4.000 1907.430 4.280 ;
        RECT 1908.270 4.000 1955.730 4.280 ;
        RECT 1956.570 4.000 2004.030 4.280 ;
        RECT 2004.870 4.000 2052.330 4.280 ;
        RECT 2053.170 4.000 2100.630 4.280 ;
        RECT 2101.470 4.000 2148.930 4.280 ;
        RECT 2149.770 4.000 2197.230 4.280 ;
        RECT 2198.070 4.000 2245.530 4.280 ;
        RECT 2246.370 4.000 2293.830 4.280 ;
        RECT 2294.670 4.000 2342.130 4.280 ;
        RECT 2342.970 4.000 2390.430 4.280 ;
        RECT 2391.270 4.000 2438.730 4.280 ;
        RECT 2439.570 4.000 2487.030 4.280 ;
        RECT 2487.870 4.000 2535.330 4.280 ;
        RECT 2536.170 4.000 2583.630 4.280 ;
        RECT 2584.470 4.000 2631.930 4.280 ;
        RECT 2632.770 4.000 2680.230 4.280 ;
        RECT 2681.070 4.000 2728.530 4.280 ;
        RECT 2729.370 4.000 2776.830 4.280 ;
        RECT 2777.670 4.000 2825.130 4.280 ;
        RECT 2825.970 4.000 2835.810 4.280 ;
      LAYER met3 ;
        RECT 4.000 3348.680 2846.000 3389.285 ;
        RECT 4.400 3347.320 2846.000 3348.680 ;
        RECT 4.400 3347.280 2845.600 3347.320 ;
        RECT 4.000 3345.920 2845.600 3347.280 ;
        RECT 4.000 3245.320 2846.000 3345.920 ;
        RECT 4.400 3243.920 2846.000 3245.320 ;
        RECT 4.000 3241.240 2846.000 3243.920 ;
        RECT 4.000 3239.840 2845.600 3241.240 ;
        RECT 4.000 3142.640 2846.000 3239.840 ;
        RECT 4.400 3141.240 2846.000 3142.640 ;
        RECT 4.000 3135.160 2846.000 3141.240 ;
        RECT 4.000 3133.760 2845.600 3135.160 ;
        RECT 4.000 3039.280 2846.000 3133.760 ;
        RECT 4.400 3037.880 2846.000 3039.280 ;
        RECT 4.000 3029.080 2846.000 3037.880 ;
        RECT 4.000 3027.680 2845.600 3029.080 ;
        RECT 4.000 2936.600 2846.000 3027.680 ;
        RECT 4.400 2935.200 2846.000 2936.600 ;
        RECT 4.000 2922.320 2846.000 2935.200 ;
        RECT 4.000 2920.920 2845.600 2922.320 ;
        RECT 4.000 2833.240 2846.000 2920.920 ;
        RECT 4.400 2831.840 2846.000 2833.240 ;
        RECT 4.000 2816.240 2846.000 2831.840 ;
        RECT 4.000 2814.840 2845.600 2816.240 ;
        RECT 4.000 2730.560 2846.000 2814.840 ;
        RECT 4.400 2729.160 2846.000 2730.560 ;
        RECT 4.000 2710.160 2846.000 2729.160 ;
        RECT 4.000 2708.760 2845.600 2710.160 ;
        RECT 4.000 2627.200 2846.000 2708.760 ;
        RECT 4.400 2625.800 2846.000 2627.200 ;
        RECT 4.000 2604.080 2846.000 2625.800 ;
        RECT 4.000 2602.680 2845.600 2604.080 ;
        RECT 4.000 2524.520 2846.000 2602.680 ;
        RECT 4.400 2523.120 2846.000 2524.520 ;
        RECT 4.000 2497.320 2846.000 2523.120 ;
        RECT 4.000 2495.920 2845.600 2497.320 ;
        RECT 4.000 2421.160 2846.000 2495.920 ;
        RECT 4.400 2419.760 2846.000 2421.160 ;
        RECT 4.000 2391.240 2846.000 2419.760 ;
        RECT 4.000 2389.840 2845.600 2391.240 ;
        RECT 4.000 2318.480 2846.000 2389.840 ;
        RECT 4.400 2317.080 2846.000 2318.480 ;
        RECT 4.000 2285.160 2846.000 2317.080 ;
        RECT 4.000 2283.760 2845.600 2285.160 ;
        RECT 4.000 2215.120 2846.000 2283.760 ;
        RECT 4.400 2213.720 2846.000 2215.120 ;
        RECT 4.000 2179.080 2846.000 2213.720 ;
        RECT 4.000 2177.680 2845.600 2179.080 ;
        RECT 4.000 2112.440 2846.000 2177.680 ;
        RECT 4.400 2111.040 2846.000 2112.440 ;
        RECT 4.000 2072.320 2846.000 2111.040 ;
        RECT 4.000 2070.920 2845.600 2072.320 ;
        RECT 4.000 2009.080 2846.000 2070.920 ;
        RECT 4.400 2007.680 2846.000 2009.080 ;
        RECT 4.000 1966.240 2846.000 2007.680 ;
        RECT 4.000 1964.840 2845.600 1966.240 ;
        RECT 4.000 1906.400 2846.000 1964.840 ;
        RECT 4.400 1905.000 2846.000 1906.400 ;
        RECT 4.000 1860.160 2846.000 1905.000 ;
        RECT 4.000 1858.760 2845.600 1860.160 ;
        RECT 4.000 1803.040 2846.000 1858.760 ;
        RECT 4.400 1801.640 2846.000 1803.040 ;
        RECT 4.000 1754.080 2846.000 1801.640 ;
        RECT 4.000 1752.680 2845.600 1754.080 ;
        RECT 4.000 1700.360 2846.000 1752.680 ;
        RECT 4.400 1698.960 2846.000 1700.360 ;
        RECT 4.000 1647.320 2846.000 1698.960 ;
        RECT 4.000 1645.920 2845.600 1647.320 ;
        RECT 4.000 1597.000 2846.000 1645.920 ;
        RECT 4.400 1595.600 2846.000 1597.000 ;
        RECT 4.000 1541.240 2846.000 1595.600 ;
        RECT 4.000 1539.840 2845.600 1541.240 ;
        RECT 4.000 1494.320 2846.000 1539.840 ;
        RECT 4.400 1492.920 2846.000 1494.320 ;
        RECT 4.000 1435.160 2846.000 1492.920 ;
        RECT 4.000 1433.760 2845.600 1435.160 ;
        RECT 4.000 1390.960 2846.000 1433.760 ;
        RECT 4.400 1389.560 2846.000 1390.960 ;
        RECT 4.000 1329.080 2846.000 1389.560 ;
        RECT 4.000 1327.680 2845.600 1329.080 ;
        RECT 4.000 1288.280 2846.000 1327.680 ;
        RECT 4.400 1286.880 2846.000 1288.280 ;
        RECT 4.000 1222.320 2846.000 1286.880 ;
        RECT 4.000 1220.920 2845.600 1222.320 ;
        RECT 4.000 1184.920 2846.000 1220.920 ;
        RECT 4.400 1183.520 2846.000 1184.920 ;
        RECT 4.000 1116.240 2846.000 1183.520 ;
        RECT 4.000 1114.840 2845.600 1116.240 ;
        RECT 4.000 1082.240 2846.000 1114.840 ;
        RECT 4.400 1080.840 2846.000 1082.240 ;
        RECT 4.000 1010.160 2846.000 1080.840 ;
        RECT 4.000 1008.760 2845.600 1010.160 ;
        RECT 4.000 978.880 2846.000 1008.760 ;
        RECT 4.400 977.480 2846.000 978.880 ;
        RECT 4.000 904.080 2846.000 977.480 ;
        RECT 4.000 902.680 2845.600 904.080 ;
        RECT 4.000 876.200 2846.000 902.680 ;
        RECT 4.400 874.800 2846.000 876.200 ;
        RECT 4.000 797.320 2846.000 874.800 ;
        RECT 4.000 795.920 2845.600 797.320 ;
        RECT 4.000 772.840 2846.000 795.920 ;
        RECT 4.400 771.440 2846.000 772.840 ;
        RECT 4.000 691.240 2846.000 771.440 ;
        RECT 4.000 689.840 2845.600 691.240 ;
        RECT 4.000 670.160 2846.000 689.840 ;
        RECT 4.400 668.760 2846.000 670.160 ;
        RECT 4.000 585.160 2846.000 668.760 ;
        RECT 4.000 583.760 2845.600 585.160 ;
        RECT 4.000 566.800 2846.000 583.760 ;
        RECT 4.400 565.400 2846.000 566.800 ;
        RECT 4.000 479.080 2846.000 565.400 ;
        RECT 4.000 477.680 2845.600 479.080 ;
        RECT 4.000 464.120 2846.000 477.680 ;
        RECT 4.400 462.720 2846.000 464.120 ;
        RECT 4.000 372.320 2846.000 462.720 ;
        RECT 4.000 370.920 2845.600 372.320 ;
        RECT 4.000 360.760 2846.000 370.920 ;
        RECT 4.400 359.360 2846.000 360.760 ;
        RECT 4.000 266.240 2846.000 359.360 ;
        RECT 4.000 264.840 2845.600 266.240 ;
        RECT 4.000 258.080 2846.000 264.840 ;
        RECT 4.400 256.680 2846.000 258.080 ;
        RECT 4.000 160.160 2846.000 256.680 ;
        RECT 4.000 158.760 2845.600 160.160 ;
        RECT 4.000 154.720 2846.000 158.760 ;
        RECT 4.400 153.320 2846.000 154.720 ;
        RECT 4.000 54.080 2846.000 153.320 ;
        RECT 4.000 52.680 2845.600 54.080 ;
        RECT 4.000 52.040 2846.000 52.680 ;
        RECT 4.400 50.640 2846.000 52.040 ;
        RECT 4.000 10.715 2846.000 50.640 ;
      LAYER met4 ;
        RECT 13.720 10.640 2813.505 3389.360 ;
      LAYER met5 ;
        RECT 5.520 103.080 2844.180 3359.755 ;
  END
END fpga
END LIBRARY


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2881.000 88.210 2885.000 88.680 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2881.000 88.080 2924.800 88.210 ;
        RECT 2884.510 87.910 2924.800 88.080 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1388.350 3445.460 1388.670 3445.520 ;
        RECT 2880.590 3445.460 2880.910 3445.520 ;
        RECT 1388.350 3445.320 2880.910 3445.460 ;
        RECT 1388.350 3445.260 1388.670 3445.320 ;
        RECT 2880.590 3445.260 2880.910 3445.320 ;
        RECT 2880.590 2435.660 2880.910 2435.720 ;
        RECT 2898.530 2435.660 2898.850 2435.720 ;
        RECT 2880.590 2435.520 2898.850 2435.660 ;
        RECT 2880.590 2435.460 2880.910 2435.520 ;
        RECT 2898.530 2435.460 2898.850 2435.520 ;
      LAYER via ;
        RECT 1388.380 3445.260 1388.640 3445.520 ;
        RECT 2880.620 3445.260 2880.880 3445.520 ;
        RECT 2880.620 2435.460 2880.880 2435.720 ;
        RECT 2898.560 2435.460 2898.820 2435.720 ;
      LAYER met2 ;
        RECT 1388.380 3445.230 1388.640 3445.550 ;
        RECT 2880.620 3445.230 2880.880 3445.550 ;
        RECT 1388.440 3435.000 1388.580 3445.230 ;
        RECT 1388.410 3431.000 1388.690 3435.000 ;
        RECT 2880.680 2435.750 2880.820 3445.230 ;
        RECT 2880.620 2435.430 2880.880 2435.750 ;
        RECT 2898.560 2435.430 2898.820 2435.750 ;
        RECT 2898.620 2434.245 2898.760 2435.430 ;
        RECT 2898.550 2433.875 2898.830 2434.245 ;
      LAYER via2 ;
        RECT 2898.550 2433.920 2898.830 2434.200 ;
      LAYER met3 ;
        RECT 2898.525 2434.210 2898.855 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2898.525 2433.910 2924.800 2434.210 ;
        RECT 2898.525 2433.895 2898.855 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 252.150 34.240 252.470 34.300 ;
        RECT 2902.670 34.240 2902.990 34.300 ;
        RECT 252.150 34.100 2902.990 34.240 ;
        RECT 252.150 34.040 252.470 34.100 ;
        RECT 2902.670 34.040 2902.990 34.100 ;
      LAYER via ;
        RECT 252.180 34.040 252.440 34.300 ;
        RECT 2902.700 34.040 2902.960 34.300 ;
      LAYER met2 ;
        RECT 2902.690 2669.155 2902.970 2669.525 ;
        RECT 252.210 35.000 252.490 39.000 ;
        RECT 252.240 34.330 252.380 35.000 ;
        RECT 2902.760 34.330 2902.900 2669.155 ;
        RECT 252.180 34.010 252.440 34.330 ;
        RECT 2902.700 34.010 2902.960 34.330 ;
      LAYER via2 ;
        RECT 2902.690 2669.200 2902.970 2669.480 ;
      LAYER met3 ;
        RECT 2902.665 2669.490 2902.995 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2902.665 2669.190 2924.800 2669.490 ;
        RECT 2902.665 2669.175 2902.995 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 300.450 33.900 300.770 33.960 ;
        RECT 2902.210 33.900 2902.530 33.960 ;
        RECT 300.450 33.760 2902.530 33.900 ;
        RECT 300.450 33.700 300.770 33.760 ;
        RECT 2902.210 33.700 2902.530 33.760 ;
      LAYER via ;
        RECT 300.480 33.700 300.740 33.960 ;
        RECT 2902.240 33.700 2902.500 33.960 ;
      LAYER met2 ;
        RECT 2902.230 2903.755 2902.510 2904.125 ;
        RECT 300.510 35.000 300.790 39.000 ;
        RECT 300.540 33.990 300.680 35.000 ;
        RECT 2902.300 33.990 2902.440 2903.755 ;
        RECT 300.480 33.670 300.740 33.990 ;
        RECT 2902.240 33.670 2902.500 33.990 ;
      LAYER via2 ;
        RECT 2902.230 2903.800 2902.510 2904.080 ;
      LAYER met3 ;
        RECT 2902.205 2904.090 2902.535 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2902.205 2903.790 2924.800 2904.090 ;
        RECT 2902.205 2903.775 2902.535 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 348.750 33.560 349.070 33.620 ;
        RECT 2901.750 33.560 2902.070 33.620 ;
        RECT 348.750 33.420 2902.070 33.560 ;
        RECT 348.750 33.360 349.070 33.420 ;
        RECT 2901.750 33.360 2902.070 33.420 ;
      LAYER via ;
        RECT 348.780 33.360 349.040 33.620 ;
        RECT 2901.780 33.360 2902.040 33.620 ;
      LAYER met2 ;
        RECT 2901.770 3138.355 2902.050 3138.725 ;
        RECT 348.810 35.000 349.090 39.000 ;
        RECT 348.840 33.650 348.980 35.000 ;
        RECT 2901.840 33.650 2901.980 3138.355 ;
        RECT 348.780 33.330 349.040 33.650 ;
        RECT 2901.780 33.330 2902.040 33.650 ;
      LAYER via2 ;
        RECT 2901.770 3138.400 2902.050 3138.680 ;
      LAYER met3 ;
        RECT 2901.745 3138.690 2902.075 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2901.745 3138.390 2924.800 3138.690 ;
        RECT 2901.745 3138.375 2902.075 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 397.050 33.220 397.370 33.280 ;
        RECT 2901.290 33.220 2901.610 33.280 ;
        RECT 397.050 33.080 2901.610 33.220 ;
        RECT 397.050 33.020 397.370 33.080 ;
        RECT 2901.290 33.020 2901.610 33.080 ;
      LAYER via ;
        RECT 397.080 33.020 397.340 33.280 ;
        RECT 2901.320 33.020 2901.580 33.280 ;
      LAYER met2 ;
        RECT 2901.310 3372.955 2901.590 3373.325 ;
        RECT 397.110 35.000 397.390 39.000 ;
        RECT 397.140 33.310 397.280 35.000 ;
        RECT 2901.380 33.310 2901.520 3372.955 ;
        RECT 397.080 32.990 397.340 33.310 ;
        RECT 2901.320 32.990 2901.580 33.310 ;
      LAYER via2 ;
        RECT 2901.310 3373.000 2901.590 3373.280 ;
      LAYER met3 ;
        RECT 2901.285 3373.290 2901.615 3373.305 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2901.285 3372.990 2924.800 3373.290 ;
        RECT 2901.285 3372.975 2901.615 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 110.010 3501.560 110.330 3501.620 ;
        RECT 2798.250 3501.560 2798.570 3501.620 ;
        RECT 110.010 3501.420 2798.570 3501.560 ;
        RECT 110.010 3501.360 110.330 3501.420 ;
        RECT 2798.250 3501.360 2798.570 3501.420 ;
        RECT 105.870 3447.840 106.190 3447.900 ;
        RECT 110.010 3447.840 110.330 3447.900 ;
        RECT 105.870 3447.700 110.330 3447.840 ;
        RECT 105.870 3447.640 106.190 3447.700 ;
        RECT 110.010 3447.640 110.330 3447.700 ;
      LAYER via ;
        RECT 110.040 3501.360 110.300 3501.620 ;
        RECT 2798.280 3501.360 2798.540 3501.620 ;
        RECT 105.900 3447.640 106.160 3447.900 ;
        RECT 110.040 3447.640 110.300 3447.900 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3501.650 2798.480 3517.600 ;
        RECT 110.040 3501.330 110.300 3501.650 ;
        RECT 2798.280 3501.330 2798.540 3501.650 ;
        RECT 110.100 3447.930 110.240 3501.330 ;
        RECT 105.900 3447.610 106.160 3447.930 ;
        RECT 110.040 3447.610 110.300 3447.930 ;
        RECT 105.960 3435.000 106.100 3447.610 ;
        RECT 105.930 3431.000 106.210 3435.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 248.010 3501.900 248.330 3501.960 ;
        RECT 2473.950 3501.900 2474.270 3501.960 ;
        RECT 248.010 3501.760 2474.270 3501.900 ;
        RECT 248.010 3501.700 248.330 3501.760 ;
        RECT 2473.950 3501.700 2474.270 3501.760 ;
      LAYER via ;
        RECT 248.040 3501.700 248.300 3501.960 ;
        RECT 2473.980 3501.700 2474.240 3501.960 ;
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3501.990 2474.180 3517.600 ;
        RECT 248.040 3501.670 248.300 3501.990 ;
        RECT 2473.980 3501.670 2474.240 3501.990 ;
        RECT 248.100 3435.000 248.240 3501.670 ;
        RECT 248.070 3431.000 248.350 3435.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 392.910 3502.240 393.230 3502.300 ;
        RECT 2149.190 3502.240 2149.510 3502.300 ;
        RECT 392.910 3502.100 2149.510 3502.240 ;
        RECT 392.910 3502.040 393.230 3502.100 ;
        RECT 2149.190 3502.040 2149.510 3502.100 ;
      LAYER via ;
        RECT 392.940 3502.040 393.200 3502.300 ;
        RECT 2149.220 3502.040 2149.480 3502.300 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3502.330 2149.420 3517.600 ;
        RECT 392.940 3502.010 393.200 3502.330 ;
        RECT 2149.220 3502.010 2149.480 3502.330 ;
        RECT 390.670 3434.410 390.950 3435.000 ;
        RECT 393.000 3434.410 393.140 3502.010 ;
        RECT 390.670 3434.270 393.140 3434.410 ;
        RECT 390.670 3431.000 390.950 3434.270 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 537.810 3502.580 538.130 3502.640 ;
        RECT 1824.890 3502.580 1825.210 3502.640 ;
        RECT 537.810 3502.440 1825.210 3502.580 ;
        RECT 537.810 3502.380 538.130 3502.440 ;
        RECT 1824.890 3502.380 1825.210 3502.440 ;
        RECT 533.210 3447.840 533.530 3447.900 ;
        RECT 537.810 3447.840 538.130 3447.900 ;
        RECT 533.210 3447.700 538.130 3447.840 ;
        RECT 533.210 3447.640 533.530 3447.700 ;
        RECT 537.810 3447.640 538.130 3447.700 ;
      LAYER via ;
        RECT 537.840 3502.380 538.100 3502.640 ;
        RECT 1824.920 3502.380 1825.180 3502.640 ;
        RECT 533.240 3447.640 533.500 3447.900 ;
        RECT 537.840 3447.640 538.100 3447.900 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3502.670 1825.120 3517.600 ;
        RECT 537.840 3502.350 538.100 3502.670 ;
        RECT 1824.920 3502.350 1825.180 3502.670 ;
        RECT 537.900 3447.930 538.040 3502.350 ;
        RECT 533.240 3447.610 533.500 3447.930 ;
        RECT 537.840 3447.610 538.100 3447.930 ;
        RECT 533.300 3435.000 533.440 3447.610 ;
        RECT 533.270 3431.000 533.550 3435.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 675.810 3502.920 676.130 3502.980 ;
        RECT 1500.590 3502.920 1500.910 3502.980 ;
        RECT 675.810 3502.780 1500.910 3502.920 ;
        RECT 675.810 3502.720 676.130 3502.780 ;
        RECT 1500.590 3502.720 1500.910 3502.780 ;
      LAYER via ;
        RECT 675.840 3502.720 676.100 3502.980 ;
        RECT 1500.620 3502.720 1500.880 3502.980 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3503.010 1500.820 3517.600 ;
        RECT 675.840 3502.690 676.100 3503.010 ;
        RECT 1500.620 3502.690 1500.880 3503.010 ;
        RECT 675.900 3435.000 676.040 3502.690 ;
        RECT 675.870 3431.000 676.150 3435.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2890.710 197.780 2891.030 197.840 ;
        RECT 2903.130 197.780 2903.450 197.840 ;
        RECT 2890.710 197.640 2903.450 197.780 ;
        RECT 2890.710 197.580 2891.030 197.640 ;
        RECT 2903.130 197.580 2903.450 197.640 ;
      LAYER via ;
        RECT 2890.740 197.580 2891.000 197.840 ;
        RECT 2903.160 197.580 2903.420 197.840 ;
      LAYER met2 ;
        RECT 2903.150 322.475 2903.430 322.845 ;
        RECT 2903.220 197.870 2903.360 322.475 ;
        RECT 2890.740 197.725 2891.000 197.870 ;
        RECT 2890.730 197.355 2891.010 197.725 ;
        RECT 2903.160 197.550 2903.420 197.870 ;
      LAYER via2 ;
        RECT 2903.150 322.520 2903.430 322.800 ;
        RECT 2890.730 197.400 2891.010 197.680 ;
      LAYER met3 ;
        RECT 2903.125 322.810 2903.455 322.825 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2903.125 322.510 2924.800 322.810 ;
        RECT 2903.125 322.495 2903.455 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
        RECT 2890.705 197.690 2891.035 197.705 ;
        RECT 2884.510 197.390 2891.035 197.690 ;
        RECT 2884.510 194.760 2884.810 197.390 ;
        RECT 2890.705 197.375 2891.035 197.390 ;
        RECT 2881.000 194.160 2885.000 194.760 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 820.710 3503.260 821.030 3503.320 ;
        RECT 1175.830 3503.260 1176.150 3503.320 ;
        RECT 820.710 3503.120 1176.150 3503.260 ;
        RECT 820.710 3503.060 821.030 3503.120 ;
        RECT 1175.830 3503.060 1176.150 3503.120 ;
      LAYER via ;
        RECT 820.740 3503.060 821.000 3503.320 ;
        RECT 1175.860 3503.060 1176.120 3503.320 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3503.350 1176.060 3517.600 ;
        RECT 820.740 3503.030 821.000 3503.350 ;
        RECT 1175.860 3503.030 1176.120 3503.350 ;
        RECT 818.470 3434.410 818.750 3435.000 ;
        RECT 820.800 3434.410 820.940 3503.030 ;
        RECT 818.470 3434.270 820.940 3434.410 ;
        RECT 818.470 3431.000 818.750 3434.270 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 851.530 3498.500 851.850 3498.560 ;
        RECT 855.210 3498.500 855.530 3498.560 ;
        RECT 851.530 3498.360 855.530 3498.500 ;
        RECT 851.530 3498.300 851.850 3498.360 ;
        RECT 855.210 3498.300 855.530 3498.360 ;
        RECT 855.210 3447.160 855.530 3447.220 ;
        RECT 960.550 3447.160 960.870 3447.220 ;
        RECT 855.210 3447.020 960.870 3447.160 ;
        RECT 855.210 3446.960 855.530 3447.020 ;
        RECT 960.550 3446.960 960.870 3447.020 ;
      LAYER via ;
        RECT 851.560 3498.300 851.820 3498.560 ;
        RECT 855.240 3498.300 855.500 3498.560 ;
        RECT 855.240 3446.960 855.500 3447.220 ;
        RECT 960.580 3446.960 960.840 3447.220 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3498.590 851.760 3517.600 ;
        RECT 851.560 3498.270 851.820 3498.590 ;
        RECT 855.240 3498.270 855.500 3498.590 ;
        RECT 855.300 3447.250 855.440 3498.270 ;
        RECT 855.240 3446.930 855.500 3447.250 ;
        RECT 960.580 3446.930 960.840 3447.250 ;
        RECT 960.640 3435.000 960.780 3446.930 ;
        RECT 960.610 3431.000 960.890 3435.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 527.230 3502.580 527.550 3502.640 ;
        RECT 530.910 3502.580 531.230 3502.640 ;
        RECT 527.230 3502.440 531.230 3502.580 ;
        RECT 527.230 3502.380 527.550 3502.440 ;
        RECT 530.910 3502.380 531.230 3502.440 ;
        RECT 530.910 3446.820 531.230 3446.880 ;
        RECT 1103.150 3446.820 1103.470 3446.880 ;
        RECT 530.910 3446.680 1103.470 3446.820 ;
        RECT 530.910 3446.620 531.230 3446.680 ;
        RECT 1103.150 3446.620 1103.470 3446.680 ;
      LAYER via ;
        RECT 527.260 3502.380 527.520 3502.640 ;
        RECT 530.940 3502.380 531.200 3502.640 ;
        RECT 530.940 3446.620 531.200 3446.880 ;
        RECT 1103.180 3446.620 1103.440 3446.880 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3502.670 527.460 3517.600 ;
        RECT 527.260 3502.350 527.520 3502.670 ;
        RECT 530.940 3502.350 531.200 3502.670 ;
        RECT 531.000 3446.910 531.140 3502.350 ;
        RECT 530.940 3446.590 531.200 3446.910 ;
        RECT 1103.180 3446.590 1103.440 3446.910 ;
        RECT 1103.240 3435.000 1103.380 3446.590 ;
        RECT 1103.210 3431.000 1103.490 3435.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 202.470 3502.240 202.790 3502.300 ;
        RECT 206.610 3502.240 206.930 3502.300 ;
        RECT 202.470 3502.100 206.930 3502.240 ;
        RECT 202.470 3502.040 202.790 3502.100 ;
        RECT 206.610 3502.040 206.930 3502.100 ;
        RECT 206.610 3446.480 206.930 3446.540 ;
        RECT 1245.750 3446.480 1246.070 3446.540 ;
        RECT 206.610 3446.340 1246.070 3446.480 ;
        RECT 206.610 3446.280 206.930 3446.340 ;
        RECT 1245.750 3446.280 1246.070 3446.340 ;
      LAYER via ;
        RECT 202.500 3502.040 202.760 3502.300 ;
        RECT 206.640 3502.040 206.900 3502.300 ;
        RECT 206.640 3446.280 206.900 3446.540 ;
        RECT 1245.780 3446.280 1246.040 3446.540 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3502.330 202.700 3517.600 ;
        RECT 202.500 3502.010 202.760 3502.330 ;
        RECT 206.640 3502.010 206.900 3502.330 ;
        RECT 206.700 3446.570 206.840 3502.010 ;
        RECT 206.640 3446.250 206.900 3446.570 ;
        RECT 1245.780 3446.250 1246.040 3446.570 ;
        RECT 1245.840 3435.000 1245.980 3446.250 ;
        RECT 1245.810 3431.000 1246.090 3435.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 3408.740 17.870 3408.800 ;
        RECT 37.790 3408.740 38.110 3408.800 ;
        RECT 17.550 3408.600 38.110 3408.740 ;
        RECT 17.550 3408.540 17.870 3408.600 ;
        RECT 37.790 3408.540 38.110 3408.600 ;
        RECT 37.790 27.440 38.110 27.500 ;
        RECT 58.950 27.440 59.270 27.500 ;
        RECT 37.790 27.300 59.270 27.440 ;
        RECT 37.790 27.240 38.110 27.300 ;
        RECT 58.950 27.240 59.270 27.300 ;
      LAYER via ;
        RECT 17.580 3408.540 17.840 3408.800 ;
        RECT 37.820 3408.540 38.080 3408.800 ;
        RECT 37.820 27.240 38.080 27.500 ;
        RECT 58.980 27.240 59.240 27.500 ;
      LAYER met2 ;
        RECT 17.570 3411.035 17.850 3411.405 ;
        RECT 17.640 3408.830 17.780 3411.035 ;
        RECT 17.580 3408.510 17.840 3408.830 ;
        RECT 37.820 3408.510 38.080 3408.830 ;
        RECT 37.880 27.530 38.020 3408.510 ;
        RECT 59.010 35.000 59.290 39.000 ;
        RECT 59.040 27.530 59.180 35.000 ;
        RECT 37.820 27.210 38.080 27.530 ;
        RECT 58.980 27.210 59.240 27.530 ;
      LAYER via2 ;
        RECT 17.570 3411.080 17.850 3411.360 ;
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 17.545 3411.370 17.875 3411.385 ;
        RECT -4.800 3411.070 17.875 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 17.545 3411.055 17.875 3411.070 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 30.965 2995.145 31.135 3042.915 ;
        RECT 30.965 2958.765 31.135 2994.635 ;
        RECT 30.965 2898.585 31.135 2946.355 ;
        RECT 30.505 2849.625 30.675 2898.075 ;
        RECT 30.505 2801.345 30.675 2825.655 ;
        RECT 30.505 2753.065 30.675 2767.175 ;
        RECT 30.505 2704.785 30.675 2752.555 ;
        RECT 30.045 2656.505 30.215 2670.615 ;
        RECT 30.505 2415.445 30.675 2439.075 ;
        RECT 29.585 2367.165 29.755 2380.935 ;
        RECT 30.505 2283.525 30.675 2359.855 ;
        RECT 30.505 2222.325 30.675 2260.915 ;
        RECT 30.505 2173.705 30.675 2221.815 ;
        RECT 30.505 2125.425 30.675 2158.235 ;
        RECT 30.965 2077.145 31.135 2125.255 ;
        RECT 30.505 2028.525 30.675 2052.835 ;
        RECT 30.965 1883.685 31.135 1931.795 ;
        RECT 30.965 1739.185 31.135 1786.275 ;
        RECT 31.885 1638.885 32.055 1683.595 ;
        RECT 30.965 1546.065 31.135 1593.835 ;
        RECT 30.965 1509.685 31.135 1545.555 ;
        RECT 30.965 1449.505 31.135 1497.275 ;
        RECT 30.965 1413.805 31.135 1448.995 ;
        RECT 30.965 1352.945 31.135 1400.715 ;
        RECT 30.965 1316.565 31.135 1352.435 ;
        RECT 30.965 1256.385 31.135 1304.155 ;
        RECT 30.505 1207.425 30.675 1255.875 ;
        RECT 30.505 1159.145 30.675 1183.455 ;
        RECT 30.505 1110.865 30.675 1124.975 ;
        RECT 30.505 1062.585 30.675 1110.355 ;
        RECT 30.505 773.245 30.675 796.875 ;
        RECT 30.505 531.505 30.675 579.615 ;
        RECT 30.505 483.225 30.675 507.195 ;
        RECT 30.965 434.945 31.135 483.055 ;
        RECT 30.505 386.325 30.675 410.635 ;
        RECT 30.965 241.485 31.135 289.595 ;
        RECT 30.965 193.205 31.135 237.235 ;
        RECT 31.425 96.645 31.595 144.755 ;
      LAYER mcon ;
        RECT 30.965 3042.745 31.135 3042.915 ;
        RECT 30.965 2994.465 31.135 2994.635 ;
        RECT 30.965 2946.185 31.135 2946.355 ;
        RECT 30.505 2897.905 30.675 2898.075 ;
        RECT 30.505 2825.485 30.675 2825.655 ;
        RECT 30.505 2767.005 30.675 2767.175 ;
        RECT 30.505 2752.385 30.675 2752.555 ;
        RECT 30.045 2670.445 30.215 2670.615 ;
        RECT 30.505 2438.905 30.675 2439.075 ;
        RECT 29.585 2380.765 29.755 2380.935 ;
        RECT 30.505 2359.685 30.675 2359.855 ;
        RECT 30.505 2260.745 30.675 2260.915 ;
        RECT 30.505 2221.645 30.675 2221.815 ;
        RECT 30.505 2158.065 30.675 2158.235 ;
        RECT 30.965 2125.085 31.135 2125.255 ;
        RECT 30.505 2052.665 30.675 2052.835 ;
        RECT 30.965 1931.625 31.135 1931.795 ;
        RECT 30.965 1786.105 31.135 1786.275 ;
        RECT 31.885 1683.425 32.055 1683.595 ;
        RECT 30.965 1593.665 31.135 1593.835 ;
        RECT 30.965 1545.385 31.135 1545.555 ;
        RECT 30.965 1497.105 31.135 1497.275 ;
        RECT 30.965 1448.825 31.135 1448.995 ;
        RECT 30.965 1400.545 31.135 1400.715 ;
        RECT 30.965 1352.265 31.135 1352.435 ;
        RECT 30.965 1303.985 31.135 1304.155 ;
        RECT 30.505 1255.705 30.675 1255.875 ;
        RECT 30.505 1183.285 30.675 1183.455 ;
        RECT 30.505 1124.805 30.675 1124.975 ;
        RECT 30.505 1110.185 30.675 1110.355 ;
        RECT 30.505 796.705 30.675 796.875 ;
        RECT 30.505 579.445 30.675 579.615 ;
        RECT 30.505 507.025 30.675 507.195 ;
        RECT 30.965 482.885 31.135 483.055 ;
        RECT 30.505 410.465 30.675 410.635 ;
        RECT 30.965 289.425 31.135 289.595 ;
        RECT 30.965 237.065 31.135 237.235 ;
        RECT 31.425 144.585 31.595 144.755 ;
      LAYER met1 ;
        RECT 15.710 3084.380 16.030 3084.440 ;
        RECT 31.810 3084.380 32.130 3084.440 ;
        RECT 15.710 3084.240 32.130 3084.380 ;
        RECT 15.710 3084.180 16.030 3084.240 ;
        RECT 31.810 3084.180 32.130 3084.240 ;
        RECT 30.890 3042.900 31.210 3042.960 ;
        RECT 30.695 3042.760 31.210 3042.900 ;
        RECT 30.890 3042.700 31.210 3042.760 ;
        RECT 30.890 2995.300 31.210 2995.360 ;
        RECT 30.695 2995.160 31.210 2995.300 ;
        RECT 30.890 2995.100 31.210 2995.160 ;
        RECT 30.890 2994.620 31.210 2994.680 ;
        RECT 30.695 2994.480 31.210 2994.620 ;
        RECT 30.890 2994.420 31.210 2994.480 ;
        RECT 30.890 2958.920 31.210 2958.980 ;
        RECT 30.695 2958.780 31.210 2958.920 ;
        RECT 30.890 2958.720 31.210 2958.780 ;
        RECT 30.890 2946.340 31.210 2946.400 ;
        RECT 30.695 2946.200 31.210 2946.340 ;
        RECT 30.890 2946.140 31.210 2946.200 ;
        RECT 30.890 2898.740 31.210 2898.800 ;
        RECT 30.695 2898.600 31.210 2898.740 ;
        RECT 30.890 2898.540 31.210 2898.600 ;
        RECT 30.445 2898.060 30.735 2898.105 ;
        RECT 30.890 2898.060 31.210 2898.120 ;
        RECT 30.445 2897.920 31.210 2898.060 ;
        RECT 30.445 2897.875 30.735 2897.920 ;
        RECT 30.890 2897.860 31.210 2897.920 ;
        RECT 30.430 2849.780 30.750 2849.840 ;
        RECT 30.235 2849.640 30.750 2849.780 ;
        RECT 30.430 2849.580 30.750 2849.640 ;
        RECT 30.430 2825.640 30.750 2825.700 ;
        RECT 30.235 2825.500 30.750 2825.640 ;
        RECT 30.430 2825.440 30.750 2825.500 ;
        RECT 30.430 2801.500 30.750 2801.560 ;
        RECT 30.235 2801.360 30.750 2801.500 ;
        RECT 30.430 2801.300 30.750 2801.360 ;
        RECT 30.430 2767.160 30.750 2767.220 ;
        RECT 30.235 2767.020 30.750 2767.160 ;
        RECT 30.430 2766.960 30.750 2767.020 ;
        RECT 30.430 2753.220 30.750 2753.280 ;
        RECT 30.235 2753.080 30.750 2753.220 ;
        RECT 30.430 2753.020 30.750 2753.080 ;
        RECT 30.430 2752.540 30.750 2752.600 ;
        RECT 30.235 2752.400 30.750 2752.540 ;
        RECT 30.430 2752.340 30.750 2752.400 ;
        RECT 30.430 2704.940 30.750 2705.000 ;
        RECT 30.235 2704.800 30.750 2704.940 ;
        RECT 30.430 2704.740 30.750 2704.800 ;
        RECT 29.985 2670.600 30.275 2670.645 ;
        RECT 30.430 2670.600 30.750 2670.660 ;
        RECT 29.985 2670.460 30.750 2670.600 ;
        RECT 29.985 2670.415 30.275 2670.460 ;
        RECT 30.430 2670.400 30.750 2670.460 ;
        RECT 29.970 2656.660 30.290 2656.720 ;
        RECT 29.775 2656.520 30.290 2656.660 ;
        RECT 29.970 2656.460 30.290 2656.520 ;
        RECT 29.050 2608.380 29.370 2608.440 ;
        RECT 30.430 2608.380 30.750 2608.440 ;
        RECT 29.050 2608.240 30.750 2608.380 ;
        RECT 29.050 2608.180 29.370 2608.240 ;
        RECT 30.430 2608.180 30.750 2608.240 ;
        RECT 30.430 2573.840 30.750 2574.100 ;
        RECT 30.520 2573.700 30.660 2573.840 ;
        RECT 30.890 2573.700 31.210 2573.760 ;
        RECT 30.520 2573.560 31.210 2573.700 ;
        RECT 30.890 2573.500 31.210 2573.560 ;
        RECT 31.350 2511.820 31.670 2511.880 ;
        RECT 32.270 2511.820 32.590 2511.880 ;
        RECT 31.350 2511.680 32.590 2511.820 ;
        RECT 31.350 2511.620 31.670 2511.680 ;
        RECT 32.270 2511.620 32.590 2511.680 ;
        RECT 30.430 2439.060 30.750 2439.120 ;
        RECT 30.235 2438.920 30.750 2439.060 ;
        RECT 30.430 2438.860 30.750 2438.920 ;
        RECT 30.445 2415.600 30.735 2415.645 ;
        RECT 30.890 2415.600 31.210 2415.660 ;
        RECT 30.445 2415.460 31.210 2415.600 ;
        RECT 30.445 2415.415 30.735 2415.460 ;
        RECT 30.890 2415.400 31.210 2415.460 ;
        RECT 29.525 2380.920 29.815 2380.965 ;
        RECT 30.890 2380.920 31.210 2380.980 ;
        RECT 29.525 2380.780 31.210 2380.920 ;
        RECT 29.525 2380.735 29.815 2380.780 ;
        RECT 30.890 2380.720 31.210 2380.780 ;
        RECT 29.510 2367.320 29.830 2367.380 ;
        RECT 29.315 2367.180 29.830 2367.320 ;
        RECT 29.510 2367.120 29.830 2367.180 ;
        RECT 29.510 2359.840 29.830 2359.900 ;
        RECT 30.445 2359.840 30.735 2359.885 ;
        RECT 29.510 2359.700 30.735 2359.840 ;
        RECT 29.510 2359.640 29.830 2359.700 ;
        RECT 30.445 2359.655 30.735 2359.700 ;
        RECT 30.430 2283.680 30.750 2283.740 ;
        RECT 30.235 2283.540 30.750 2283.680 ;
        RECT 30.430 2283.480 30.750 2283.540 ;
        RECT 30.430 2260.900 30.750 2260.960 ;
        RECT 30.235 2260.760 30.750 2260.900 ;
        RECT 30.430 2260.700 30.750 2260.760 ;
        RECT 30.445 2222.480 30.735 2222.525 ;
        RECT 30.890 2222.480 31.210 2222.540 ;
        RECT 30.445 2222.340 31.210 2222.480 ;
        RECT 30.445 2222.295 30.735 2222.340 ;
        RECT 30.890 2222.280 31.210 2222.340 ;
        RECT 30.445 2221.800 30.735 2221.845 ;
        RECT 30.890 2221.800 31.210 2221.860 ;
        RECT 30.445 2221.660 31.210 2221.800 ;
        RECT 30.445 2221.615 30.735 2221.660 ;
        RECT 30.890 2221.600 31.210 2221.660 ;
        RECT 30.430 2173.860 30.750 2173.920 ;
        RECT 30.235 2173.720 30.750 2173.860 ;
        RECT 30.430 2173.660 30.750 2173.720 ;
        RECT 30.430 2158.220 30.750 2158.280 ;
        RECT 30.235 2158.080 30.750 2158.220 ;
        RECT 30.430 2158.020 30.750 2158.080 ;
        RECT 30.430 2125.580 30.750 2125.640 ;
        RECT 30.235 2125.440 30.750 2125.580 ;
        RECT 30.430 2125.380 30.750 2125.440 ;
        RECT 30.890 2125.240 31.210 2125.300 ;
        RECT 30.695 2125.100 31.210 2125.240 ;
        RECT 30.890 2125.040 31.210 2125.100 ;
        RECT 30.430 2077.300 30.750 2077.360 ;
        RECT 30.905 2077.300 31.195 2077.345 ;
        RECT 30.430 2077.160 31.195 2077.300 ;
        RECT 30.430 2077.100 30.750 2077.160 ;
        RECT 30.905 2077.115 31.195 2077.160 ;
        RECT 30.430 2052.820 30.750 2052.880 ;
        RECT 30.235 2052.680 30.750 2052.820 ;
        RECT 30.430 2052.620 30.750 2052.680 ;
        RECT 30.430 2028.680 30.750 2028.740 ;
        RECT 30.235 2028.540 30.750 2028.680 ;
        RECT 30.430 2028.480 30.750 2028.540 ;
        RECT 30.430 1994.140 30.750 1994.400 ;
        RECT 30.520 1994.000 30.660 1994.140 ;
        RECT 30.890 1994.000 31.210 1994.060 ;
        RECT 30.520 1993.860 31.210 1994.000 ;
        RECT 30.890 1993.800 31.210 1993.860 ;
        RECT 30.890 1945.860 31.210 1946.120 ;
        RECT 30.430 1945.720 30.750 1945.780 ;
        RECT 30.980 1945.720 31.120 1945.860 ;
        RECT 30.430 1945.580 31.120 1945.720 ;
        RECT 30.430 1945.520 30.750 1945.580 ;
        RECT 30.890 1931.780 31.210 1931.840 ;
        RECT 30.695 1931.640 31.210 1931.780 ;
        RECT 30.890 1931.580 31.210 1931.640 ;
        RECT 30.890 1883.840 31.210 1883.900 ;
        RECT 30.695 1883.700 31.210 1883.840 ;
        RECT 30.890 1883.640 31.210 1883.700 ;
        RECT 30.890 1849.500 31.210 1849.560 ;
        RECT 30.520 1849.360 31.210 1849.500 ;
        RECT 30.520 1849.220 30.660 1849.360 ;
        RECT 30.890 1849.300 31.210 1849.360 ;
        RECT 30.430 1848.960 30.750 1849.220 ;
        RECT 30.430 1801.020 30.750 1801.280 ;
        RECT 30.520 1800.880 30.660 1801.020 ;
        RECT 30.890 1800.880 31.210 1800.940 ;
        RECT 30.520 1800.740 31.210 1800.880 ;
        RECT 30.890 1800.680 31.210 1800.740 ;
        RECT 30.890 1786.260 31.210 1786.320 ;
        RECT 30.695 1786.120 31.210 1786.260 ;
        RECT 30.890 1786.060 31.210 1786.120 ;
        RECT 30.890 1739.340 31.210 1739.400 ;
        RECT 30.695 1739.200 31.210 1739.340 ;
        RECT 30.890 1739.140 31.210 1739.200 ;
        RECT 30.890 1704.460 31.210 1704.720 ;
        RECT 30.980 1703.700 31.120 1704.460 ;
        RECT 30.890 1703.440 31.210 1703.700 ;
        RECT 30.890 1690.380 31.210 1690.440 ;
        RECT 31.810 1690.380 32.130 1690.440 ;
        RECT 30.890 1690.240 32.130 1690.380 ;
        RECT 30.890 1690.180 31.210 1690.240 ;
        RECT 31.810 1690.180 32.130 1690.240 ;
        RECT 31.810 1683.580 32.130 1683.640 ;
        RECT 31.615 1683.440 32.130 1683.580 ;
        RECT 31.810 1683.380 32.130 1683.440 ;
        RECT 31.810 1639.040 32.130 1639.100 ;
        RECT 31.615 1638.900 32.130 1639.040 ;
        RECT 31.810 1638.840 32.130 1638.900 ;
        RECT 30.890 1593.820 31.210 1593.880 ;
        RECT 30.695 1593.680 31.210 1593.820 ;
        RECT 30.890 1593.620 31.210 1593.680 ;
        RECT 30.890 1546.220 31.210 1546.280 ;
        RECT 30.695 1546.080 31.210 1546.220 ;
        RECT 30.890 1546.020 31.210 1546.080 ;
        RECT 30.890 1545.540 31.210 1545.600 ;
        RECT 30.695 1545.400 31.210 1545.540 ;
        RECT 30.890 1545.340 31.210 1545.400 ;
        RECT 30.890 1509.840 31.210 1509.900 ;
        RECT 30.695 1509.700 31.210 1509.840 ;
        RECT 30.890 1509.640 31.210 1509.700 ;
        RECT 30.890 1497.260 31.210 1497.320 ;
        RECT 30.695 1497.120 31.210 1497.260 ;
        RECT 30.890 1497.060 31.210 1497.120 ;
        RECT 30.890 1449.660 31.210 1449.720 ;
        RECT 30.695 1449.520 31.210 1449.660 ;
        RECT 30.890 1449.460 31.210 1449.520 ;
        RECT 30.890 1448.980 31.210 1449.040 ;
        RECT 30.695 1448.840 31.210 1448.980 ;
        RECT 30.890 1448.780 31.210 1448.840 ;
        RECT 30.890 1413.960 31.210 1414.020 ;
        RECT 30.695 1413.820 31.210 1413.960 ;
        RECT 30.890 1413.760 31.210 1413.820 ;
        RECT 30.890 1400.700 31.210 1400.760 ;
        RECT 30.695 1400.560 31.210 1400.700 ;
        RECT 30.890 1400.500 31.210 1400.560 ;
        RECT 30.890 1353.100 31.210 1353.160 ;
        RECT 30.695 1352.960 31.210 1353.100 ;
        RECT 30.890 1352.900 31.210 1352.960 ;
        RECT 30.890 1352.420 31.210 1352.480 ;
        RECT 30.695 1352.280 31.210 1352.420 ;
        RECT 30.890 1352.220 31.210 1352.280 ;
        RECT 30.890 1316.720 31.210 1316.780 ;
        RECT 30.695 1316.580 31.210 1316.720 ;
        RECT 30.890 1316.520 31.210 1316.580 ;
        RECT 30.890 1304.140 31.210 1304.200 ;
        RECT 30.695 1304.000 31.210 1304.140 ;
        RECT 30.890 1303.940 31.210 1304.000 ;
        RECT 30.890 1256.540 31.210 1256.600 ;
        RECT 30.695 1256.400 31.210 1256.540 ;
        RECT 30.890 1256.340 31.210 1256.400 ;
        RECT 30.445 1255.860 30.735 1255.905 ;
        RECT 30.890 1255.860 31.210 1255.920 ;
        RECT 30.445 1255.720 31.210 1255.860 ;
        RECT 30.445 1255.675 30.735 1255.720 ;
        RECT 30.890 1255.660 31.210 1255.720 ;
        RECT 30.430 1207.580 30.750 1207.640 ;
        RECT 30.235 1207.440 30.750 1207.580 ;
        RECT 30.430 1207.380 30.750 1207.440 ;
        RECT 30.430 1183.440 30.750 1183.500 ;
        RECT 30.235 1183.300 30.750 1183.440 ;
        RECT 30.430 1183.240 30.750 1183.300 ;
        RECT 30.430 1159.300 30.750 1159.360 ;
        RECT 30.235 1159.160 30.750 1159.300 ;
        RECT 30.430 1159.100 30.750 1159.160 ;
        RECT 30.430 1124.960 30.750 1125.020 ;
        RECT 30.235 1124.820 30.750 1124.960 ;
        RECT 30.430 1124.760 30.750 1124.820 ;
        RECT 30.430 1111.020 30.750 1111.080 ;
        RECT 30.235 1110.880 30.750 1111.020 ;
        RECT 30.430 1110.820 30.750 1110.880 ;
        RECT 30.430 1110.340 30.750 1110.400 ;
        RECT 30.235 1110.200 30.750 1110.340 ;
        RECT 30.430 1110.140 30.750 1110.200 ;
        RECT 30.430 1062.740 30.750 1062.800 ;
        RECT 30.235 1062.600 30.750 1062.740 ;
        RECT 30.430 1062.540 30.750 1062.600 ;
        RECT 30.430 1028.200 30.750 1028.460 ;
        RECT 30.520 1028.060 30.660 1028.200 ;
        RECT 30.890 1028.060 31.210 1028.120 ;
        RECT 30.520 1027.920 31.210 1028.060 ;
        RECT 30.890 1027.860 31.210 1027.920 ;
        RECT 31.350 966.180 31.670 966.240 ;
        RECT 32.270 966.180 32.590 966.240 ;
        RECT 31.350 966.040 32.590 966.180 ;
        RECT 31.350 965.980 31.670 966.040 ;
        RECT 32.270 965.980 32.590 966.040 ;
        RECT 30.430 917.900 30.750 917.960 ;
        RECT 31.350 917.900 31.670 917.960 ;
        RECT 30.430 917.760 31.670 917.900 ;
        RECT 30.430 917.700 30.750 917.760 ;
        RECT 31.350 917.700 31.670 917.760 ;
        RECT 31.350 869.620 31.670 869.680 ;
        RECT 32.270 869.620 32.590 869.680 ;
        RECT 31.350 869.480 32.590 869.620 ;
        RECT 31.350 869.420 31.670 869.480 ;
        RECT 32.270 869.420 32.590 869.480 ;
        RECT 30.430 796.860 30.750 796.920 ;
        RECT 30.235 796.720 30.750 796.860 ;
        RECT 30.430 796.660 30.750 796.720 ;
        RECT 30.445 773.400 30.735 773.445 ;
        RECT 30.890 773.400 31.210 773.460 ;
        RECT 30.445 773.260 31.210 773.400 ;
        RECT 30.445 773.215 30.735 773.260 ;
        RECT 30.890 773.200 31.210 773.260 ;
        RECT 29.510 772.720 29.830 772.780 ;
        RECT 30.890 772.720 31.210 772.780 ;
        RECT 29.510 772.580 31.210 772.720 ;
        RECT 29.510 772.520 29.830 772.580 ;
        RECT 30.890 772.520 31.210 772.580 ;
        RECT 30.430 690.240 30.750 690.500 ;
        RECT 30.520 689.820 30.660 690.240 ;
        RECT 30.430 689.560 30.750 689.820 ;
        RECT 29.510 676.160 29.830 676.220 ;
        RECT 30.890 676.160 31.210 676.220 ;
        RECT 29.510 676.020 31.210 676.160 ;
        RECT 29.510 675.960 29.830 676.020 ;
        RECT 30.890 675.960 31.210 676.020 ;
        RECT 30.430 593.340 30.750 593.600 ;
        RECT 30.520 593.200 30.660 593.340 ;
        RECT 30.890 593.200 31.210 593.260 ;
        RECT 30.520 593.060 31.210 593.200 ;
        RECT 30.890 593.000 31.210 593.060 ;
        RECT 30.445 579.600 30.735 579.645 ;
        RECT 30.890 579.600 31.210 579.660 ;
        RECT 30.445 579.460 31.210 579.600 ;
        RECT 30.445 579.415 30.735 579.460 ;
        RECT 30.890 579.400 31.210 579.460 ;
        RECT 30.430 531.660 30.750 531.720 ;
        RECT 30.235 531.520 30.750 531.660 ;
        RECT 30.430 531.460 30.750 531.520 ;
        RECT 30.430 507.180 30.750 507.240 ;
        RECT 30.235 507.040 30.750 507.180 ;
        RECT 30.430 506.980 30.750 507.040 ;
        RECT 30.430 483.380 30.750 483.440 ;
        RECT 30.235 483.240 30.750 483.380 ;
        RECT 30.430 483.180 30.750 483.240 ;
        RECT 30.890 483.040 31.210 483.100 ;
        RECT 30.695 482.900 31.210 483.040 ;
        RECT 30.890 482.840 31.210 482.900 ;
        RECT 30.430 435.100 30.750 435.160 ;
        RECT 30.905 435.100 31.195 435.145 ;
        RECT 30.430 434.960 31.195 435.100 ;
        RECT 30.430 434.900 30.750 434.960 ;
        RECT 30.905 434.915 31.195 434.960 ;
        RECT 30.430 410.620 30.750 410.680 ;
        RECT 30.235 410.480 30.750 410.620 ;
        RECT 30.430 410.420 30.750 410.480 ;
        RECT 30.430 386.480 30.750 386.540 ;
        RECT 30.235 386.340 30.750 386.480 ;
        RECT 30.430 386.280 30.750 386.340 ;
        RECT 30.430 351.940 30.750 352.200 ;
        RECT 30.520 351.800 30.660 351.940 ;
        RECT 30.890 351.800 31.210 351.860 ;
        RECT 30.520 351.660 31.210 351.800 ;
        RECT 30.890 351.600 31.210 351.660 ;
        RECT 30.890 303.660 31.210 303.920 ;
        RECT 30.430 303.520 30.750 303.580 ;
        RECT 30.980 303.520 31.120 303.660 ;
        RECT 30.430 303.380 31.120 303.520 ;
        RECT 30.430 303.320 30.750 303.380 ;
        RECT 30.890 289.580 31.210 289.640 ;
        RECT 30.695 289.440 31.210 289.580 ;
        RECT 30.890 289.380 31.210 289.440 ;
        RECT 30.890 241.640 31.210 241.700 ;
        RECT 30.695 241.500 31.210 241.640 ;
        RECT 30.890 241.440 31.210 241.500 ;
        RECT 30.890 237.220 31.210 237.280 ;
        RECT 30.695 237.080 31.210 237.220 ;
        RECT 30.890 237.020 31.210 237.080 ;
        RECT 30.890 193.360 31.210 193.420 ;
        RECT 30.695 193.220 31.210 193.360 ;
        RECT 30.890 193.160 31.210 193.220 ;
        RECT 30.890 158.680 31.210 158.740 ;
        RECT 31.810 158.680 32.130 158.740 ;
        RECT 30.890 158.540 32.130 158.680 ;
        RECT 30.890 158.480 31.210 158.540 ;
        RECT 31.810 158.480 32.130 158.540 ;
        RECT 31.365 144.740 31.655 144.785 ;
        RECT 31.810 144.740 32.130 144.800 ;
        RECT 31.365 144.600 32.130 144.740 ;
        RECT 31.365 144.555 31.655 144.600 ;
        RECT 31.810 144.540 32.130 144.600 ;
        RECT 31.350 96.800 31.670 96.860 ;
        RECT 31.155 96.660 31.670 96.800 ;
        RECT 31.350 96.600 31.670 96.660 ;
        RECT 33.190 24.040 33.510 24.100 ;
        RECT 107.250 24.040 107.570 24.100 ;
        RECT 33.190 23.900 107.570 24.040 ;
        RECT 33.190 23.840 33.510 23.900 ;
        RECT 107.250 23.840 107.570 23.900 ;
      LAYER via ;
        RECT 15.740 3084.180 16.000 3084.440 ;
        RECT 31.840 3084.180 32.100 3084.440 ;
        RECT 30.920 3042.700 31.180 3042.960 ;
        RECT 30.920 2995.100 31.180 2995.360 ;
        RECT 30.920 2994.420 31.180 2994.680 ;
        RECT 30.920 2958.720 31.180 2958.980 ;
        RECT 30.920 2946.140 31.180 2946.400 ;
        RECT 30.920 2898.540 31.180 2898.800 ;
        RECT 30.920 2897.860 31.180 2898.120 ;
        RECT 30.460 2849.580 30.720 2849.840 ;
        RECT 30.460 2825.440 30.720 2825.700 ;
        RECT 30.460 2801.300 30.720 2801.560 ;
        RECT 30.460 2766.960 30.720 2767.220 ;
        RECT 30.460 2753.020 30.720 2753.280 ;
        RECT 30.460 2752.340 30.720 2752.600 ;
        RECT 30.460 2704.740 30.720 2705.000 ;
        RECT 30.460 2670.400 30.720 2670.660 ;
        RECT 30.000 2656.460 30.260 2656.720 ;
        RECT 29.080 2608.180 29.340 2608.440 ;
        RECT 30.460 2608.180 30.720 2608.440 ;
        RECT 30.460 2573.840 30.720 2574.100 ;
        RECT 30.920 2573.500 31.180 2573.760 ;
        RECT 31.380 2511.620 31.640 2511.880 ;
        RECT 32.300 2511.620 32.560 2511.880 ;
        RECT 30.460 2438.860 30.720 2439.120 ;
        RECT 30.920 2415.400 31.180 2415.660 ;
        RECT 30.920 2380.720 31.180 2380.980 ;
        RECT 29.540 2367.120 29.800 2367.380 ;
        RECT 29.540 2359.640 29.800 2359.900 ;
        RECT 30.460 2283.480 30.720 2283.740 ;
        RECT 30.460 2260.700 30.720 2260.960 ;
        RECT 30.920 2222.280 31.180 2222.540 ;
        RECT 30.920 2221.600 31.180 2221.860 ;
        RECT 30.460 2173.660 30.720 2173.920 ;
        RECT 30.460 2158.020 30.720 2158.280 ;
        RECT 30.460 2125.380 30.720 2125.640 ;
        RECT 30.920 2125.040 31.180 2125.300 ;
        RECT 30.460 2077.100 30.720 2077.360 ;
        RECT 30.460 2052.620 30.720 2052.880 ;
        RECT 30.460 2028.480 30.720 2028.740 ;
        RECT 30.460 1994.140 30.720 1994.400 ;
        RECT 30.920 1993.800 31.180 1994.060 ;
        RECT 30.920 1945.860 31.180 1946.120 ;
        RECT 30.460 1945.520 30.720 1945.780 ;
        RECT 30.920 1931.580 31.180 1931.840 ;
        RECT 30.920 1883.640 31.180 1883.900 ;
        RECT 30.920 1849.300 31.180 1849.560 ;
        RECT 30.460 1848.960 30.720 1849.220 ;
        RECT 30.460 1801.020 30.720 1801.280 ;
        RECT 30.920 1800.680 31.180 1800.940 ;
        RECT 30.920 1786.060 31.180 1786.320 ;
        RECT 30.920 1739.140 31.180 1739.400 ;
        RECT 30.920 1704.460 31.180 1704.720 ;
        RECT 30.920 1703.440 31.180 1703.700 ;
        RECT 30.920 1690.180 31.180 1690.440 ;
        RECT 31.840 1690.180 32.100 1690.440 ;
        RECT 31.840 1683.380 32.100 1683.640 ;
        RECT 31.840 1638.840 32.100 1639.100 ;
        RECT 30.920 1593.620 31.180 1593.880 ;
        RECT 30.920 1546.020 31.180 1546.280 ;
        RECT 30.920 1545.340 31.180 1545.600 ;
        RECT 30.920 1509.640 31.180 1509.900 ;
        RECT 30.920 1497.060 31.180 1497.320 ;
        RECT 30.920 1449.460 31.180 1449.720 ;
        RECT 30.920 1448.780 31.180 1449.040 ;
        RECT 30.920 1413.760 31.180 1414.020 ;
        RECT 30.920 1400.500 31.180 1400.760 ;
        RECT 30.920 1352.900 31.180 1353.160 ;
        RECT 30.920 1352.220 31.180 1352.480 ;
        RECT 30.920 1316.520 31.180 1316.780 ;
        RECT 30.920 1303.940 31.180 1304.200 ;
        RECT 30.920 1256.340 31.180 1256.600 ;
        RECT 30.920 1255.660 31.180 1255.920 ;
        RECT 30.460 1207.380 30.720 1207.640 ;
        RECT 30.460 1183.240 30.720 1183.500 ;
        RECT 30.460 1159.100 30.720 1159.360 ;
        RECT 30.460 1124.760 30.720 1125.020 ;
        RECT 30.460 1110.820 30.720 1111.080 ;
        RECT 30.460 1110.140 30.720 1110.400 ;
        RECT 30.460 1062.540 30.720 1062.800 ;
        RECT 30.460 1028.200 30.720 1028.460 ;
        RECT 30.920 1027.860 31.180 1028.120 ;
        RECT 31.380 965.980 31.640 966.240 ;
        RECT 32.300 965.980 32.560 966.240 ;
        RECT 30.460 917.700 30.720 917.960 ;
        RECT 31.380 917.700 31.640 917.960 ;
        RECT 31.380 869.420 31.640 869.680 ;
        RECT 32.300 869.420 32.560 869.680 ;
        RECT 30.460 796.660 30.720 796.920 ;
        RECT 30.920 773.200 31.180 773.460 ;
        RECT 29.540 772.520 29.800 772.780 ;
        RECT 30.920 772.520 31.180 772.780 ;
        RECT 30.460 690.240 30.720 690.500 ;
        RECT 30.460 689.560 30.720 689.820 ;
        RECT 29.540 675.960 29.800 676.220 ;
        RECT 30.920 675.960 31.180 676.220 ;
        RECT 30.460 593.340 30.720 593.600 ;
        RECT 30.920 593.000 31.180 593.260 ;
        RECT 30.920 579.400 31.180 579.660 ;
        RECT 30.460 531.460 30.720 531.720 ;
        RECT 30.460 506.980 30.720 507.240 ;
        RECT 30.460 483.180 30.720 483.440 ;
        RECT 30.920 482.840 31.180 483.100 ;
        RECT 30.460 434.900 30.720 435.160 ;
        RECT 30.460 410.420 30.720 410.680 ;
        RECT 30.460 386.280 30.720 386.540 ;
        RECT 30.460 351.940 30.720 352.200 ;
        RECT 30.920 351.600 31.180 351.860 ;
        RECT 30.920 303.660 31.180 303.920 ;
        RECT 30.460 303.320 30.720 303.580 ;
        RECT 30.920 289.380 31.180 289.640 ;
        RECT 30.920 241.440 31.180 241.700 ;
        RECT 30.920 237.020 31.180 237.280 ;
        RECT 30.920 193.160 31.180 193.420 ;
        RECT 30.920 158.480 31.180 158.740 ;
        RECT 31.840 158.480 32.100 158.740 ;
        RECT 31.840 144.540 32.100 144.800 ;
        RECT 31.380 96.600 31.640 96.860 ;
        RECT 33.220 23.840 33.480 24.100 ;
        RECT 107.280 23.840 107.540 24.100 ;
      LAYER met2 ;
        RECT 15.730 3124.075 16.010 3124.445 ;
        RECT 15.800 3084.470 15.940 3124.075 ;
        RECT 15.740 3084.150 16.000 3084.470 ;
        RECT 31.840 3084.150 32.100 3084.470 ;
        RECT 31.900 3043.410 32.040 3084.150 ;
        RECT 30.980 3043.270 32.040 3043.410 ;
        RECT 30.980 3042.990 31.120 3043.270 ;
        RECT 30.920 3042.670 31.180 3042.990 ;
        RECT 30.920 2995.070 31.180 2995.390 ;
        RECT 30.980 2994.710 31.120 2995.070 ;
        RECT 30.920 2994.390 31.180 2994.710 ;
        RECT 30.920 2958.690 31.180 2959.010 ;
        RECT 30.980 2946.430 31.120 2958.690 ;
        RECT 30.920 2946.110 31.180 2946.430 ;
        RECT 30.920 2898.510 31.180 2898.830 ;
        RECT 30.980 2898.150 31.120 2898.510 ;
        RECT 30.920 2897.830 31.180 2898.150 ;
        RECT 30.460 2849.550 30.720 2849.870 ;
        RECT 30.520 2825.730 30.660 2849.550 ;
        RECT 30.460 2825.410 30.720 2825.730 ;
        RECT 30.460 2801.270 30.720 2801.590 ;
        RECT 30.520 2767.250 30.660 2801.270 ;
        RECT 30.460 2766.930 30.720 2767.250 ;
        RECT 30.460 2752.990 30.720 2753.310 ;
        RECT 30.520 2752.630 30.660 2752.990 ;
        RECT 30.460 2752.310 30.720 2752.630 ;
        RECT 30.460 2704.710 30.720 2705.030 ;
        RECT 30.520 2670.690 30.660 2704.710 ;
        RECT 30.460 2670.370 30.720 2670.690 ;
        RECT 30.000 2656.605 30.260 2656.750 ;
        RECT 29.070 2656.235 29.350 2656.605 ;
        RECT 29.990 2656.235 30.270 2656.605 ;
        RECT 29.140 2608.470 29.280 2656.235 ;
        RECT 29.080 2608.150 29.340 2608.470 ;
        RECT 30.460 2608.150 30.720 2608.470 ;
        RECT 30.520 2574.130 30.660 2608.150 ;
        RECT 30.460 2573.810 30.720 2574.130 ;
        RECT 30.920 2573.470 31.180 2573.790 ;
        RECT 30.980 2560.045 31.120 2573.470 ;
        RECT 30.910 2559.675 31.190 2560.045 ;
        RECT 32.290 2559.675 32.570 2560.045 ;
        RECT 32.360 2511.910 32.500 2559.675 ;
        RECT 31.380 2511.590 31.640 2511.910 ;
        RECT 32.300 2511.590 32.560 2511.910 ;
        RECT 31.440 2463.485 31.580 2511.590 ;
        RECT 30.450 2463.115 30.730 2463.485 ;
        RECT 31.370 2463.115 31.650 2463.485 ;
        RECT 30.520 2439.150 30.660 2463.115 ;
        RECT 30.460 2438.830 30.720 2439.150 ;
        RECT 30.920 2415.370 31.180 2415.690 ;
        RECT 30.980 2381.010 31.120 2415.370 ;
        RECT 30.920 2380.690 31.180 2381.010 ;
        RECT 29.540 2367.090 29.800 2367.410 ;
        RECT 29.600 2359.930 29.740 2367.090 ;
        RECT 29.540 2359.610 29.800 2359.930 ;
        RECT 30.460 2283.450 30.720 2283.770 ;
        RECT 30.520 2260.990 30.660 2283.450 ;
        RECT 30.460 2260.670 30.720 2260.990 ;
        RECT 30.920 2222.250 31.180 2222.570 ;
        RECT 30.980 2221.890 31.120 2222.250 ;
        RECT 30.920 2221.570 31.180 2221.890 ;
        RECT 30.460 2173.630 30.720 2173.950 ;
        RECT 30.520 2158.310 30.660 2173.630 ;
        RECT 30.460 2157.990 30.720 2158.310 ;
        RECT 30.460 2125.410 30.720 2125.670 ;
        RECT 30.460 2125.350 31.120 2125.410 ;
        RECT 30.520 2125.330 31.120 2125.350 ;
        RECT 30.520 2125.270 31.180 2125.330 ;
        RECT 30.920 2125.010 31.180 2125.270 ;
        RECT 30.980 2124.855 31.120 2125.010 ;
        RECT 30.460 2077.070 30.720 2077.390 ;
        RECT 30.520 2052.910 30.660 2077.070 ;
        RECT 30.460 2052.590 30.720 2052.910 ;
        RECT 30.460 2028.450 30.720 2028.770 ;
        RECT 30.520 1994.430 30.660 2028.450 ;
        RECT 30.460 1994.110 30.720 1994.430 ;
        RECT 30.920 1993.770 31.180 1994.090 ;
        RECT 30.980 1946.150 31.120 1993.770 ;
        RECT 30.920 1945.830 31.180 1946.150 ;
        RECT 30.460 1945.490 30.720 1945.810 ;
        RECT 30.520 1932.290 30.660 1945.490 ;
        RECT 30.520 1932.150 31.120 1932.290 ;
        RECT 30.980 1931.870 31.120 1932.150 ;
        RECT 30.920 1931.550 31.180 1931.870 ;
        RECT 30.920 1883.610 31.180 1883.930 ;
        RECT 30.980 1849.590 31.120 1883.610 ;
        RECT 30.920 1849.270 31.180 1849.590 ;
        RECT 30.460 1848.930 30.720 1849.250 ;
        RECT 30.520 1801.310 30.660 1848.930 ;
        RECT 30.460 1800.990 30.720 1801.310 ;
        RECT 30.920 1800.650 31.180 1800.970 ;
        RECT 30.980 1786.350 31.120 1800.650 ;
        RECT 30.920 1786.030 31.180 1786.350 ;
        RECT 30.920 1739.110 31.180 1739.430 ;
        RECT 30.980 1704.750 31.120 1739.110 ;
        RECT 30.920 1704.430 31.180 1704.750 ;
        RECT 30.920 1703.410 31.180 1703.730 ;
        RECT 30.980 1690.470 31.120 1703.410 ;
        RECT 30.920 1690.150 31.180 1690.470 ;
        RECT 31.840 1690.150 32.100 1690.470 ;
        RECT 31.900 1683.670 32.040 1690.150 ;
        RECT 31.840 1683.350 32.100 1683.670 ;
        RECT 31.840 1638.810 32.100 1639.130 ;
        RECT 31.900 1607.250 32.040 1638.810 ;
        RECT 30.980 1607.110 32.040 1607.250 ;
        RECT 30.980 1593.910 31.120 1607.110 ;
        RECT 30.920 1593.590 31.180 1593.910 ;
        RECT 30.920 1545.990 31.180 1546.310 ;
        RECT 30.980 1545.630 31.120 1545.990 ;
        RECT 30.920 1545.310 31.180 1545.630 ;
        RECT 30.920 1509.610 31.180 1509.930 ;
        RECT 30.980 1497.350 31.120 1509.610 ;
        RECT 30.920 1497.030 31.180 1497.350 ;
        RECT 30.920 1449.430 31.180 1449.750 ;
        RECT 30.980 1449.070 31.120 1449.430 ;
        RECT 30.920 1448.750 31.180 1449.070 ;
        RECT 30.920 1413.730 31.180 1414.050 ;
        RECT 30.980 1400.790 31.120 1413.730 ;
        RECT 30.920 1400.470 31.180 1400.790 ;
        RECT 30.920 1352.870 31.180 1353.190 ;
        RECT 30.980 1352.510 31.120 1352.870 ;
        RECT 30.920 1352.190 31.180 1352.510 ;
        RECT 30.920 1316.490 31.180 1316.810 ;
        RECT 30.980 1304.230 31.120 1316.490 ;
        RECT 30.920 1303.910 31.180 1304.230 ;
        RECT 30.920 1256.310 31.180 1256.630 ;
        RECT 30.980 1255.950 31.120 1256.310 ;
        RECT 30.920 1255.630 31.180 1255.950 ;
        RECT 30.460 1207.350 30.720 1207.670 ;
        RECT 30.520 1183.530 30.660 1207.350 ;
        RECT 30.460 1183.210 30.720 1183.530 ;
        RECT 30.460 1159.070 30.720 1159.390 ;
        RECT 30.520 1125.050 30.660 1159.070 ;
        RECT 30.460 1124.730 30.720 1125.050 ;
        RECT 30.460 1110.790 30.720 1111.110 ;
        RECT 30.520 1110.430 30.660 1110.790 ;
        RECT 30.460 1110.110 30.720 1110.430 ;
        RECT 30.460 1062.510 30.720 1062.830 ;
        RECT 30.520 1028.490 30.660 1062.510 ;
        RECT 30.460 1028.170 30.720 1028.490 ;
        RECT 30.920 1027.830 31.180 1028.150 ;
        RECT 30.980 1014.405 31.120 1027.830 ;
        RECT 30.910 1014.035 31.190 1014.405 ;
        RECT 32.290 1014.035 32.570 1014.405 ;
        RECT 32.360 966.270 32.500 1014.035 ;
        RECT 31.380 965.950 31.640 966.270 ;
        RECT 32.300 965.950 32.560 966.270 ;
        RECT 30.520 917.990 30.660 918.145 ;
        RECT 31.440 917.990 31.580 965.950 ;
        RECT 30.460 917.730 30.720 917.990 ;
        RECT 30.910 917.730 31.190 917.845 ;
        RECT 30.460 917.670 31.190 917.730 ;
        RECT 31.380 917.670 31.640 917.990 ;
        RECT 30.520 917.590 31.190 917.670 ;
        RECT 30.910 917.475 31.190 917.590 ;
        RECT 32.290 917.475 32.570 917.845 ;
        RECT 32.360 869.710 32.500 917.475 ;
        RECT 31.380 869.390 31.640 869.710 ;
        RECT 32.300 869.390 32.560 869.710 ;
        RECT 31.440 821.285 31.580 869.390 ;
        RECT 30.450 820.915 30.730 821.285 ;
        RECT 31.370 820.915 31.650 821.285 ;
        RECT 30.520 796.950 30.660 820.915 ;
        RECT 30.460 796.630 30.720 796.950 ;
        RECT 30.920 773.170 31.180 773.490 ;
        RECT 30.980 772.810 31.120 773.170 ;
        RECT 29.540 772.490 29.800 772.810 ;
        RECT 30.920 772.490 31.180 772.810 ;
        RECT 29.600 724.725 29.740 772.490 ;
        RECT 29.530 724.355 29.810 724.725 ;
        RECT 30.450 724.355 30.730 724.725 ;
        RECT 30.520 690.530 30.660 724.355 ;
        RECT 30.460 690.210 30.720 690.530 ;
        RECT 30.460 689.530 30.720 689.850 ;
        RECT 30.520 676.330 30.660 689.530 ;
        RECT 30.520 676.250 31.120 676.330 ;
        RECT 29.540 675.930 29.800 676.250 ;
        RECT 30.520 676.190 31.180 676.250 ;
        RECT 30.920 675.930 31.180 676.190 ;
        RECT 29.600 628.165 29.740 675.930 ;
        RECT 30.980 675.775 31.120 675.930 ;
        RECT 29.530 627.795 29.810 628.165 ;
        RECT 30.450 627.795 30.730 628.165 ;
        RECT 30.520 593.630 30.660 627.795 ;
        RECT 30.460 593.310 30.720 593.630 ;
        RECT 30.920 592.970 31.180 593.290 ;
        RECT 30.980 579.690 31.120 592.970 ;
        RECT 30.920 579.370 31.180 579.690 ;
        RECT 30.460 531.430 30.720 531.750 ;
        RECT 30.520 507.270 30.660 531.430 ;
        RECT 30.460 506.950 30.720 507.270 ;
        RECT 30.460 483.210 30.720 483.470 ;
        RECT 30.460 483.150 31.120 483.210 ;
        RECT 30.520 483.130 31.120 483.150 ;
        RECT 30.520 483.070 31.180 483.130 ;
        RECT 30.920 482.810 31.180 483.070 ;
        RECT 30.980 482.655 31.120 482.810 ;
        RECT 30.460 434.870 30.720 435.190 ;
        RECT 30.520 410.710 30.660 434.870 ;
        RECT 30.460 410.390 30.720 410.710 ;
        RECT 30.460 386.250 30.720 386.570 ;
        RECT 30.520 352.230 30.660 386.250 ;
        RECT 30.460 351.910 30.720 352.230 ;
        RECT 30.920 351.570 31.180 351.890 ;
        RECT 30.980 303.950 31.120 351.570 ;
        RECT 30.920 303.630 31.180 303.950 ;
        RECT 30.460 303.290 30.720 303.610 ;
        RECT 30.520 290.090 30.660 303.290 ;
        RECT 30.520 289.950 31.120 290.090 ;
        RECT 30.980 289.670 31.120 289.950 ;
        RECT 30.920 289.350 31.180 289.670 ;
        RECT 30.920 241.410 31.180 241.730 ;
        RECT 30.980 237.310 31.120 241.410 ;
        RECT 30.920 236.990 31.180 237.310 ;
        RECT 30.920 193.130 31.180 193.450 ;
        RECT 30.980 158.770 31.120 193.130 ;
        RECT 30.920 158.450 31.180 158.770 ;
        RECT 31.840 158.450 32.100 158.770 ;
        RECT 31.900 144.830 32.040 158.450 ;
        RECT 31.840 144.510 32.100 144.830 ;
        RECT 31.380 96.570 31.640 96.890 ;
        RECT 31.440 62.290 31.580 96.570 ;
        RECT 31.440 62.150 33.420 62.290 ;
        RECT 33.280 24.130 33.420 62.150 ;
        RECT 107.310 35.000 107.590 39.000 ;
        RECT 107.340 24.130 107.480 35.000 ;
        RECT 33.220 23.810 33.480 24.130 ;
        RECT 107.280 23.810 107.540 24.130 ;
      LAYER via2 ;
        RECT 15.730 3124.120 16.010 3124.400 ;
        RECT 29.070 2656.280 29.350 2656.560 ;
        RECT 29.990 2656.280 30.270 2656.560 ;
        RECT 30.910 2559.720 31.190 2560.000 ;
        RECT 32.290 2559.720 32.570 2560.000 ;
        RECT 30.450 2463.160 30.730 2463.440 ;
        RECT 31.370 2463.160 31.650 2463.440 ;
        RECT 30.910 1014.080 31.190 1014.360 ;
        RECT 32.290 1014.080 32.570 1014.360 ;
        RECT 30.910 917.520 31.190 917.800 ;
        RECT 32.290 917.520 32.570 917.800 ;
        RECT 30.450 820.960 30.730 821.240 ;
        RECT 31.370 820.960 31.650 821.240 ;
        RECT 29.530 724.400 29.810 724.680 ;
        RECT 30.450 724.400 30.730 724.680 ;
        RECT 29.530 627.840 29.810 628.120 ;
        RECT 30.450 627.840 30.730 628.120 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 15.705 3124.410 16.035 3124.425 ;
        RECT -4.800 3124.110 16.035 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 15.705 3124.095 16.035 3124.110 ;
        RECT 29.045 2656.570 29.375 2656.585 ;
        RECT 29.965 2656.570 30.295 2656.585 ;
        RECT 29.045 2656.270 30.295 2656.570 ;
        RECT 29.045 2656.255 29.375 2656.270 ;
        RECT 29.965 2656.255 30.295 2656.270 ;
        RECT 30.885 2560.010 31.215 2560.025 ;
        RECT 32.265 2560.010 32.595 2560.025 ;
        RECT 30.885 2559.710 32.595 2560.010 ;
        RECT 30.885 2559.695 31.215 2559.710 ;
        RECT 32.265 2559.695 32.595 2559.710 ;
        RECT 30.425 2463.450 30.755 2463.465 ;
        RECT 31.345 2463.450 31.675 2463.465 ;
        RECT 30.425 2463.150 31.675 2463.450 ;
        RECT 30.425 2463.135 30.755 2463.150 ;
        RECT 31.345 2463.135 31.675 2463.150 ;
        RECT 30.885 1014.370 31.215 1014.385 ;
        RECT 32.265 1014.370 32.595 1014.385 ;
        RECT 30.885 1014.070 32.595 1014.370 ;
        RECT 30.885 1014.055 31.215 1014.070 ;
        RECT 32.265 1014.055 32.595 1014.070 ;
        RECT 30.885 917.810 31.215 917.825 ;
        RECT 32.265 917.810 32.595 917.825 ;
        RECT 30.885 917.510 32.595 917.810 ;
        RECT 30.885 917.495 31.215 917.510 ;
        RECT 32.265 917.495 32.595 917.510 ;
        RECT 30.425 821.250 30.755 821.265 ;
        RECT 31.345 821.250 31.675 821.265 ;
        RECT 30.425 820.950 31.675 821.250 ;
        RECT 30.425 820.935 30.755 820.950 ;
        RECT 31.345 820.935 31.675 820.950 ;
        RECT 29.505 724.690 29.835 724.705 ;
        RECT 30.425 724.690 30.755 724.705 ;
        RECT 29.505 724.390 30.755 724.690 ;
        RECT 29.505 724.375 29.835 724.390 ;
        RECT 30.425 724.375 30.755 724.390 ;
        RECT 29.505 628.130 29.835 628.145 ;
        RECT 30.425 628.130 30.755 628.145 ;
        RECT 29.505 627.830 30.755 628.130 ;
        RECT 29.505 627.815 29.835 627.830 ;
        RECT 30.425 627.815 30.755 627.830 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.630 2836.520 16.950 2836.580 ;
        RECT 38.250 2836.520 38.570 2836.580 ;
        RECT 16.630 2836.380 38.570 2836.520 ;
        RECT 16.630 2836.320 16.950 2836.380 ;
        RECT 38.250 2836.320 38.570 2836.380 ;
        RECT 38.250 25.740 38.570 25.800 ;
        RECT 155.550 25.740 155.870 25.800 ;
        RECT 38.250 25.600 155.870 25.740 ;
        RECT 38.250 25.540 38.570 25.600 ;
        RECT 155.550 25.540 155.870 25.600 ;
      LAYER via ;
        RECT 16.660 2836.320 16.920 2836.580 ;
        RECT 38.280 2836.320 38.540 2836.580 ;
        RECT 38.280 25.540 38.540 25.800 ;
        RECT 155.580 25.540 155.840 25.800 ;
      LAYER met2 ;
        RECT 16.650 2836.435 16.930 2836.805 ;
        RECT 16.660 2836.290 16.920 2836.435 ;
        RECT 38.280 2836.290 38.540 2836.610 ;
        RECT 38.340 25.830 38.480 2836.290 ;
        RECT 155.610 35.000 155.890 39.000 ;
        RECT 155.640 25.830 155.780 35.000 ;
        RECT 38.280 25.510 38.540 25.830 ;
        RECT 155.580 25.510 155.840 25.830 ;
      LAYER via2 ;
        RECT 16.650 2836.480 16.930 2836.760 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 16.625 2836.770 16.955 2836.785 ;
        RECT -4.800 2836.470 16.955 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 16.625 2836.455 16.955 2836.470 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 15.710 2546.500 16.030 2546.560 ;
        RECT 38.710 2546.500 39.030 2546.560 ;
        RECT 15.710 2546.360 39.030 2546.500 ;
        RECT 15.710 2546.300 16.030 2546.360 ;
        RECT 38.710 2546.300 39.030 2546.360 ;
        RECT 38.710 25.400 39.030 25.460 ;
        RECT 203.850 25.400 204.170 25.460 ;
        RECT 38.710 25.260 204.170 25.400 ;
        RECT 38.710 25.200 39.030 25.260 ;
        RECT 203.850 25.200 204.170 25.260 ;
      LAYER via ;
        RECT 15.740 2546.300 16.000 2546.560 ;
        RECT 38.740 2546.300 39.000 2546.560 ;
        RECT 38.740 25.200 39.000 25.460 ;
        RECT 203.880 25.200 204.140 25.460 ;
      LAYER met2 ;
        RECT 15.730 2549.475 16.010 2549.845 ;
        RECT 15.800 2546.590 15.940 2549.475 ;
        RECT 15.740 2546.270 16.000 2546.590 ;
        RECT 38.740 2546.270 39.000 2546.590 ;
        RECT 38.800 25.490 38.940 2546.270 ;
        RECT 203.910 35.000 204.190 39.000 ;
        RECT 203.940 25.490 204.080 35.000 ;
        RECT 38.740 25.170 39.000 25.490 ;
        RECT 203.880 25.170 204.140 25.490 ;
      LAYER via2 ;
        RECT 15.730 2549.520 16.010 2549.800 ;
      LAYER met3 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 15.705 2549.810 16.035 2549.825 ;
        RECT -4.800 2549.510 16.035 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 15.705 2549.495 16.035 2549.510 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.110 2261.835 17.390 2262.205 ;
        RECT 17.180 89.605 17.320 2261.835 ;
        RECT 17.110 89.235 17.390 89.605 ;
      LAYER via2 ;
        RECT 17.110 2261.880 17.390 2262.160 ;
        RECT 17.110 89.280 17.390 89.560 ;
      LAYER met3 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 17.085 2262.170 17.415 2262.185 ;
        RECT -4.800 2261.870 17.415 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 17.085 2261.855 17.415 2261.870 ;
        RECT 17.085 89.570 17.415 89.585 ;
        RECT 17.085 89.270 35.570 89.570 ;
        RECT 17.085 89.255 17.415 89.270 ;
        RECT 35.270 86.640 35.570 89.270 ;
        RECT 35.000 86.040 39.000 86.640 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.570 1974.875 17.850 1975.245 ;
        RECT 17.640 191.605 17.780 1974.875 ;
        RECT 17.570 191.235 17.850 191.605 ;
      LAYER via2 ;
        RECT 17.570 1974.920 17.850 1975.200 ;
        RECT 17.570 191.280 17.850 191.560 ;
      LAYER met3 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 17.545 1975.210 17.875 1975.225 ;
        RECT -4.800 1974.910 17.875 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 17.545 1974.895 17.875 1974.910 ;
        RECT 17.545 191.570 17.875 191.585 ;
        RECT 17.545 191.270 35.570 191.570 ;
        RECT 17.545 191.255 17.875 191.270 ;
        RECT 35.270 189.320 35.570 191.270 ;
        RECT 35.000 188.720 39.000 189.320 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2890.710 303.180 2891.030 303.240 ;
        RECT 2904.050 303.180 2904.370 303.240 ;
        RECT 2890.710 303.040 2904.370 303.180 ;
        RECT 2890.710 302.980 2891.030 303.040 ;
        RECT 2904.050 302.980 2904.370 303.040 ;
      LAYER via ;
        RECT 2890.740 302.980 2891.000 303.240 ;
        RECT 2904.080 302.980 2904.340 303.240 ;
      LAYER met2 ;
        RECT 2904.070 557.075 2904.350 557.445 ;
        RECT 2904.140 303.270 2904.280 557.075 ;
        RECT 2890.740 303.125 2891.000 303.270 ;
        RECT 2890.730 302.755 2891.010 303.125 ;
        RECT 2904.080 302.950 2904.340 303.270 ;
      LAYER via2 ;
        RECT 2904.070 557.120 2904.350 557.400 ;
        RECT 2890.730 302.800 2891.010 303.080 ;
      LAYER met3 ;
        RECT 2904.045 557.410 2904.375 557.425 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2904.045 557.110 2924.800 557.410 ;
        RECT 2904.045 557.095 2904.375 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
        RECT 2890.705 303.090 2891.035 303.105 ;
        RECT 2884.510 302.790 2891.035 303.090 ;
        RECT 2884.510 300.840 2884.810 302.790 ;
        RECT 2890.705 302.775 2891.035 302.790 ;
        RECT 2881.000 300.240 2885.000 300.840 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.030 1687.235 18.310 1687.605 ;
        RECT 18.100 295.645 18.240 1687.235 ;
        RECT 18.030 295.275 18.310 295.645 ;
      LAYER via2 ;
        RECT 18.030 1687.280 18.310 1687.560 ;
        RECT 18.030 295.320 18.310 295.600 ;
      LAYER met3 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 18.005 1687.570 18.335 1687.585 ;
        RECT -4.800 1687.270 18.335 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
        RECT 18.005 1687.255 18.335 1687.270 ;
        RECT 18.005 295.610 18.335 295.625 ;
        RECT 18.005 295.310 35.570 295.610 ;
        RECT 18.005 295.295 18.335 295.310 ;
        RECT 35.270 292.680 35.570 295.310 ;
        RECT 35.000 292.080 39.000 292.680 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 1471.675 18.770 1472.045 ;
        RECT 18.560 398.325 18.700 1471.675 ;
        RECT 18.490 397.955 18.770 398.325 ;
      LAYER via2 ;
        RECT 18.490 1471.720 18.770 1472.000 ;
        RECT 18.490 398.000 18.770 398.280 ;
      LAYER met3 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 18.465 1472.010 18.795 1472.025 ;
        RECT -4.800 1471.710 18.795 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 18.465 1471.695 18.795 1471.710 ;
        RECT 18.465 398.290 18.795 398.305 ;
        RECT 18.465 397.990 35.570 398.290 ;
        RECT 18.465 397.975 18.795 397.990 ;
        RECT 35.270 395.360 35.570 397.990 ;
        RECT 35.000 394.760 39.000 395.360 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.410 1256.115 19.690 1256.485 ;
        RECT 19.480 501.685 19.620 1256.115 ;
        RECT 19.410 501.315 19.690 501.685 ;
      LAYER via2 ;
        RECT 19.410 1256.160 19.690 1256.440 ;
        RECT 19.410 501.360 19.690 501.640 ;
      LAYER met3 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 19.385 1256.450 19.715 1256.465 ;
        RECT -4.800 1256.150 19.715 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 19.385 1256.135 19.715 1256.150 ;
        RECT 19.385 501.650 19.715 501.665 ;
        RECT 19.385 501.350 35.570 501.650 ;
        RECT 19.385 501.335 19.715 501.350 ;
        RECT 35.270 498.720 35.570 501.350 ;
        RECT 35.000 498.120 39.000 498.720 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.330 1040.555 20.610 1040.925 ;
        RECT 20.400 604.365 20.540 1040.555 ;
        RECT 20.330 603.995 20.610 604.365 ;
      LAYER via2 ;
        RECT 20.330 1040.600 20.610 1040.880 ;
        RECT 20.330 604.040 20.610 604.320 ;
      LAYER met3 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 20.305 1040.890 20.635 1040.905 ;
        RECT -4.800 1040.590 20.635 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
        RECT 20.305 1040.575 20.635 1040.590 ;
        RECT 20.305 604.330 20.635 604.345 ;
        RECT 20.305 604.030 35.570 604.330 ;
        RECT 20.305 604.015 20.635 604.030 ;
        RECT 35.270 601.400 35.570 604.030 ;
        RECT 35.000 600.800 39.000 601.400 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.190 824.995 16.470 825.365 ;
        RECT 16.260 707.725 16.400 824.995 ;
        RECT 16.190 707.355 16.470 707.725 ;
      LAYER via2 ;
        RECT 16.190 825.040 16.470 825.320 ;
        RECT 16.190 707.400 16.470 707.680 ;
      LAYER met3 ;
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 16.165 825.330 16.495 825.345 ;
        RECT -4.800 825.030 16.495 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
        RECT 16.165 825.015 16.495 825.030 ;
        RECT 16.165 707.690 16.495 707.705 ;
        RECT 16.165 707.390 35.570 707.690 ;
        RECT 16.165 707.375 16.495 707.390 ;
        RECT 35.270 704.760 35.570 707.390 ;
        RECT 35.000 704.160 39.000 704.760 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.650 803.915 16.930 804.285 ;
        RECT 16.720 610.485 16.860 803.915 ;
        RECT 16.650 610.115 16.930 610.485 ;
      LAYER via2 ;
        RECT 16.650 803.960 16.930 804.240 ;
        RECT 16.650 610.160 16.930 610.440 ;
      LAYER met3 ;
        RECT 35.000 806.840 39.000 807.440 ;
        RECT 16.625 804.250 16.955 804.265 ;
        RECT 35.270 804.250 35.570 806.840 ;
        RECT 16.625 803.950 35.570 804.250 ;
        RECT 16.625 803.935 16.955 803.950 ;
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 16.625 610.450 16.955 610.465 ;
        RECT -4.800 610.150 16.955 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 16.625 610.135 16.955 610.150 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.870 907.275 20.150 907.645 ;
        RECT 19.940 394.925 20.080 907.275 ;
        RECT 19.870 394.555 20.150 394.925 ;
      LAYER via2 ;
        RECT 19.870 907.320 20.150 907.600 ;
        RECT 19.870 394.600 20.150 394.880 ;
      LAYER met3 ;
        RECT 35.000 910.200 39.000 910.800 ;
        RECT 19.845 907.610 20.175 907.625 ;
        RECT 35.270 907.610 35.570 910.200 ;
        RECT 19.845 907.310 35.570 907.610 ;
        RECT 19.845 907.295 20.175 907.310 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 19.845 394.890 20.175 394.905 ;
        RECT -4.800 394.590 20.175 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 19.845 394.575 20.175 394.590 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.950 1009.955 19.230 1010.325 ;
        RECT 19.020 179.365 19.160 1009.955 ;
        RECT 18.950 178.995 19.230 179.365 ;
      LAYER via2 ;
        RECT 18.950 1010.000 19.230 1010.280 ;
        RECT 18.950 179.040 19.230 179.320 ;
      LAYER met3 ;
        RECT 35.000 1012.880 39.000 1013.480 ;
        RECT 18.925 1010.290 19.255 1010.305 ;
        RECT 35.270 1010.290 35.570 1012.880 ;
        RECT 18.925 1009.990 35.570 1010.290 ;
        RECT 18.925 1009.975 19.255 1009.990 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 18.925 179.330 19.255 179.345 ;
        RECT -4.800 179.030 19.255 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 18.925 179.015 19.255 179.030 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2890.710 406.880 2891.030 406.940 ;
        RECT 2903.590 406.880 2903.910 406.940 ;
        RECT 2890.710 406.740 2903.910 406.880 ;
        RECT 2890.710 406.680 2891.030 406.740 ;
        RECT 2903.590 406.680 2903.910 406.740 ;
      LAYER via ;
        RECT 2890.740 406.680 2891.000 406.940 ;
        RECT 2903.620 406.680 2903.880 406.940 ;
      LAYER met2 ;
        RECT 2903.610 791.675 2903.890 792.045 ;
        RECT 2890.730 406.795 2891.010 407.165 ;
        RECT 2903.680 406.970 2903.820 791.675 ;
        RECT 2890.740 406.650 2891.000 406.795 ;
        RECT 2903.620 406.650 2903.880 406.970 ;
      LAYER via2 ;
        RECT 2903.610 791.720 2903.890 792.000 ;
        RECT 2890.730 406.840 2891.010 407.120 ;
      LAYER met3 ;
        RECT 2903.585 792.010 2903.915 792.025 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2903.585 791.710 2924.800 792.010 ;
        RECT 2903.585 791.695 2903.915 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
        RECT 2890.705 407.130 2891.035 407.145 ;
        RECT 2884.510 406.920 2891.035 407.130 ;
        RECT 2881.000 406.830 2891.035 406.920 ;
        RECT 2881.000 406.320 2885.000 406.830 ;
        RECT 2890.705 406.815 2891.035 406.830 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2890.710 516.020 2891.030 516.080 ;
        RECT 2903.130 516.020 2903.450 516.080 ;
        RECT 2890.710 515.880 2903.450 516.020 ;
        RECT 2890.710 515.820 2891.030 515.880 ;
        RECT 2903.130 515.820 2903.450 515.880 ;
      LAYER via ;
        RECT 2890.740 515.820 2891.000 516.080 ;
        RECT 2903.160 515.820 2903.420 516.080 ;
      LAYER met2 ;
        RECT 2903.150 1026.275 2903.430 1026.645 ;
        RECT 2903.220 516.110 2903.360 1026.275 ;
        RECT 2890.740 515.965 2891.000 516.110 ;
        RECT 2890.730 515.595 2891.010 515.965 ;
        RECT 2903.160 515.790 2903.420 516.110 ;
      LAYER via2 ;
        RECT 2903.150 1026.320 2903.430 1026.600 ;
        RECT 2890.730 515.640 2891.010 515.920 ;
      LAYER met3 ;
        RECT 2903.125 1026.610 2903.455 1026.625 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2903.125 1026.310 2924.800 1026.610 ;
        RECT 2903.125 1026.295 2903.455 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
        RECT 2890.705 515.930 2891.035 515.945 ;
        RECT 2884.510 515.630 2891.035 515.930 ;
        RECT 2884.510 513.680 2884.810 515.630 ;
        RECT 2890.705 515.615 2891.035 515.630 ;
        RECT 2881.000 513.080 2885.000 513.680 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2900.850 1260.875 2901.130 1261.245 ;
        RECT 2900.920 620.685 2901.060 1260.875 ;
        RECT 2900.850 620.315 2901.130 620.685 ;
      LAYER via2 ;
        RECT 2900.850 1260.920 2901.130 1261.200 ;
        RECT 2900.850 620.360 2901.130 620.640 ;
      LAYER met3 ;
        RECT 2900.825 1261.210 2901.155 1261.225 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2900.825 1260.910 2924.800 1261.210 ;
        RECT 2900.825 1260.895 2901.155 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
        RECT 2900.825 620.650 2901.155 620.665 ;
        RECT 2884.510 620.350 2901.155 620.650 ;
        RECT 2884.510 619.760 2884.810 620.350 ;
        RECT 2900.825 620.335 2901.155 620.350 ;
        RECT 2881.000 619.160 2885.000 619.760 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2890.710 728.860 2891.030 728.920 ;
        RECT 2904.510 728.860 2904.830 728.920 ;
        RECT 2890.710 728.720 2904.830 728.860 ;
        RECT 2890.710 728.660 2891.030 728.720 ;
        RECT 2904.510 728.660 2904.830 728.720 ;
      LAYER via ;
        RECT 2890.740 728.660 2891.000 728.920 ;
        RECT 2904.540 728.660 2904.800 728.920 ;
      LAYER met2 ;
        RECT 2904.530 1495.475 2904.810 1495.845 ;
        RECT 2904.600 728.950 2904.740 1495.475 ;
        RECT 2890.740 728.805 2891.000 728.950 ;
        RECT 2890.730 728.435 2891.010 728.805 ;
        RECT 2904.540 728.630 2904.800 728.950 ;
      LAYER via2 ;
        RECT 2904.530 1495.520 2904.810 1495.800 ;
        RECT 2890.730 728.480 2891.010 728.760 ;
      LAYER met3 ;
        RECT 2904.505 1495.810 2904.835 1495.825 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2904.505 1495.510 2924.800 1495.810 ;
        RECT 2904.505 1495.495 2904.835 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
        RECT 2890.705 728.770 2891.035 728.785 ;
        RECT 2884.510 728.470 2891.035 728.770 ;
        RECT 2884.510 725.840 2884.810 728.470 ;
        RECT 2890.705 728.455 2891.035 728.470 ;
        RECT 2881.000 725.240 2885.000 725.840 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2890.710 834.940 2891.030 835.000 ;
        RECT 2904.050 834.940 2904.370 835.000 ;
        RECT 2890.710 834.800 2904.370 834.940 ;
        RECT 2890.710 834.740 2891.030 834.800 ;
        RECT 2904.050 834.740 2904.370 834.800 ;
      LAYER via ;
        RECT 2890.740 834.740 2891.000 835.000 ;
        RECT 2904.080 834.740 2904.340 835.000 ;
      LAYER met2 ;
        RECT 2904.070 1730.075 2904.350 1730.445 ;
        RECT 2904.140 835.030 2904.280 1730.075 ;
        RECT 2890.740 834.885 2891.000 835.030 ;
        RECT 2890.730 834.515 2891.010 834.885 ;
        RECT 2904.080 834.710 2904.340 835.030 ;
      LAYER via2 ;
        RECT 2904.070 1730.120 2904.350 1730.400 ;
        RECT 2890.730 834.560 2891.010 834.840 ;
      LAYER met3 ;
        RECT 2904.045 1730.410 2904.375 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2904.045 1730.110 2924.800 1730.410 ;
        RECT 2904.045 1730.095 2904.375 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
        RECT 2890.705 834.850 2891.035 834.865 ;
        RECT 2884.510 834.550 2891.035 834.850 ;
        RECT 2884.510 831.920 2884.810 834.550 ;
        RECT 2890.705 834.535 2891.035 834.550 ;
        RECT 2881.000 831.320 2885.000 831.920 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2890.710 938.300 2891.030 938.360 ;
        RECT 2903.590 938.300 2903.910 938.360 ;
        RECT 2890.710 938.160 2903.910 938.300 ;
        RECT 2890.710 938.100 2891.030 938.160 ;
        RECT 2903.590 938.100 2903.910 938.160 ;
      LAYER via ;
        RECT 2890.740 938.100 2891.000 938.360 ;
        RECT 2903.620 938.100 2903.880 938.360 ;
      LAYER met2 ;
        RECT 2903.610 1964.675 2903.890 1965.045 ;
        RECT 2903.680 938.390 2903.820 1964.675 ;
        RECT 2890.740 938.245 2891.000 938.390 ;
        RECT 2890.730 937.875 2891.010 938.245 ;
        RECT 2903.620 938.070 2903.880 938.390 ;
      LAYER via2 ;
        RECT 2903.610 1964.720 2903.890 1965.000 ;
        RECT 2890.730 937.920 2891.010 938.200 ;
      LAYER met3 ;
        RECT 2903.585 1965.010 2903.915 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2903.585 1964.710 2924.800 1965.010 ;
        RECT 2903.585 1964.695 2903.915 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
        RECT 2881.000 938.210 2885.000 938.680 ;
        RECT 2890.705 938.210 2891.035 938.225 ;
        RECT 2881.000 938.080 2891.035 938.210 ;
        RECT 2884.510 937.910 2891.035 938.080 ;
        RECT 2890.705 937.895 2891.035 937.910 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2890.710 1047.100 2891.030 1047.160 ;
        RECT 2903.130 1047.100 2903.450 1047.160 ;
        RECT 2890.710 1046.960 2903.450 1047.100 ;
        RECT 2890.710 1046.900 2891.030 1046.960 ;
        RECT 2903.130 1046.900 2903.450 1046.960 ;
      LAYER via ;
        RECT 2890.740 1046.900 2891.000 1047.160 ;
        RECT 2903.160 1046.900 2903.420 1047.160 ;
      LAYER met2 ;
        RECT 2903.150 2199.275 2903.430 2199.645 ;
        RECT 2903.220 1047.190 2903.360 2199.275 ;
        RECT 2890.740 1047.045 2891.000 1047.190 ;
        RECT 2890.730 1046.675 2891.010 1047.045 ;
        RECT 2903.160 1046.870 2903.420 1047.190 ;
      LAYER via2 ;
        RECT 2903.150 2199.320 2903.430 2199.600 ;
        RECT 2890.730 1046.720 2891.010 1047.000 ;
      LAYER met3 ;
        RECT 2903.125 2199.610 2903.455 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2903.125 2199.310 2924.800 2199.610 ;
        RECT 2903.125 2199.295 2903.455 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
        RECT 2890.705 1047.010 2891.035 1047.025 ;
        RECT 2884.510 1046.710 2891.035 1047.010 ;
        RECT 2884.510 1044.760 2884.810 1046.710 ;
        RECT 2890.705 1046.695 2891.035 1046.710 ;
        RECT 2881.000 1044.160 2885.000 1044.760 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 204.420 2924.800 205.620 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2551.100 2924.800 2552.300 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2785.700 2924.800 2786.900 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3020.300 2924.800 3021.500 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3254.900 2924.800 3256.100 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3489.500 2924.800 3490.700 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 439.020 2924.800 440.220 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 3267.140 2.400 3268.340 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2979.500 2.400 2980.700 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2692.540 2.400 2693.740 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2404.900 2.400 2406.100 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2117.940 2.400 2119.140 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1830.300 2.400 1831.500 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 673.620 2924.800 674.820 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1543.340 2.400 1544.540 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1327.780 2.400 1328.980 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1112.220 2.400 1113.420 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 896.660 2.400 897.860 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 681.100 2.400 682.300 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 465.540 2.400 466.740 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 249.980 2.400 251.180 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 35.100 2.400 36.300 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 908.900 2924.800 910.100 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1143.500 2924.800 1144.700 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1378.100 2924.800 1379.300 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1612.700 2924.800 1613.900 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1847.300 2924.800 1848.500 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2081.900 2924.800 2083.100 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2316.500 2924.800 2317.700 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 145.940 2924.800 147.140 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2492.620 2924.800 2493.820 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2727.220 2924.800 2728.420 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2961.820 2924.800 2963.020 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3196.420 2924.800 3197.620 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3431.020 2924.800 3432.220 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 380.540 2924.800 381.740 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 3339.220 2.400 3340.420 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 3051.580 2.400 3052.780 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2764.620 2.400 2765.820 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2476.980 2.400 2478.180 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2189.340 2.400 2190.540 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1902.380 2.400 1903.580 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 615.140 2924.800 616.340 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1614.740 2.400 1615.940 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1399.860 2.400 1401.060 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1184.300 2.400 1185.500 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 968.740 2.400 969.940 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 753.180 2.400 754.380 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 537.620 2.400 538.820 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 322.060 2.400 323.260 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 106.500 2.400 107.700 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 849.740 2924.800 850.940 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1084.340 2924.800 1085.540 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1318.940 2924.800 1320.140 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1553.540 2924.800 1554.740 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1788.820 2924.800 1790.020 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2023.420 2924.800 2024.620 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2258.020 2924.800 2259.220 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 674.310 -4.800 674.870 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2.830 30.840 3.150 30.900 ;
        RECT 2897.610 30.840 2897.930 30.900 ;
        RECT 2.830 30.700 2897.930 30.840 ;
        RECT 2.830 30.640 3.150 30.700 ;
        RECT 2897.610 30.640 2897.930 30.700 ;
      LAYER via ;
        RECT 2.860 30.640 3.120 30.900 ;
        RECT 2897.640 30.640 2897.900 30.900 ;
      LAYER met2 ;
        RECT 2897.630 1147.995 2897.910 1148.365 ;
        RECT 2897.700 30.930 2897.840 1147.995 ;
        RECT 2.860 30.610 3.120 30.930 ;
        RECT 2897.640 30.610 2897.900 30.930 ;
        RECT 2.920 2.400 3.060 30.610 ;
        RECT 2.710 -4.800 3.270 2.400 ;
      LAYER via2 ;
        RECT 2897.630 1148.040 2897.910 1148.320 ;
      LAYER met3 ;
        RECT 2881.000 1150.240 2885.000 1150.840 ;
        RECT 2884.510 1148.330 2884.810 1150.240 ;
        RECT 2897.605 1148.330 2897.935 1148.345 ;
        RECT 2884.510 1148.030 2897.935 1148.330 ;
        RECT 2897.605 1148.015 2897.935 1148.030 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 8.350 10.440 8.670 10.500 ;
        RECT 1990.950 10.440 1991.270 10.500 ;
        RECT 8.350 10.300 1991.270 10.440 ;
        RECT 8.350 10.240 8.670 10.300 ;
        RECT 1990.950 10.240 1991.270 10.300 ;
      LAYER via ;
        RECT 8.380 10.240 8.640 10.500 ;
        RECT 1990.980 10.240 1991.240 10.500 ;
      LAYER met2 ;
        RECT 1991.010 35.000 1991.290 39.000 ;
        RECT 1991.040 10.530 1991.180 35.000 ;
        RECT 8.380 10.210 8.640 10.530 ;
        RECT 1990.980 10.210 1991.240 10.530 ;
        RECT 8.440 2.400 8.580 10.210 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.330 25.060 14.650 25.120 ;
        RECT 2039.250 25.060 2039.570 25.120 ;
        RECT 14.330 24.920 2039.570 25.060 ;
        RECT 14.330 24.860 14.650 24.920 ;
        RECT 2039.250 24.860 2039.570 24.920 ;
      LAYER via ;
        RECT 14.360 24.860 14.620 25.120 ;
        RECT 2039.280 24.860 2039.540 25.120 ;
      LAYER met2 ;
        RECT 2039.310 35.000 2039.590 39.000 ;
        RECT 2039.340 25.150 2039.480 35.000 ;
        RECT 14.360 24.830 14.620 25.150 ;
        RECT 2039.280 24.830 2039.540 25.150 ;
        RECT 14.420 2.400 14.560 24.830 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 37.330 31.180 37.650 31.240 ;
        RECT 2897.150 31.180 2897.470 31.240 ;
        RECT 37.330 31.040 2897.470 31.180 ;
        RECT 37.330 30.980 37.650 31.040 ;
        RECT 2897.150 30.980 2897.470 31.040 ;
      LAYER via ;
        RECT 37.360 30.980 37.620 31.240 ;
        RECT 2897.180 30.980 2897.440 31.240 ;
      LAYER met2 ;
        RECT 2897.170 1256.115 2897.450 1256.485 ;
        RECT 2897.240 31.270 2897.380 1256.115 ;
        RECT 37.360 30.950 37.620 31.270 ;
        RECT 2897.180 30.950 2897.440 31.270 ;
        RECT 37.420 14.010 37.560 30.950 ;
        RECT 37.420 13.870 38.480 14.010 ;
        RECT 38.340 2.400 38.480 13.870 ;
        RECT 38.130 -4.800 38.690 2.400 ;
      LAYER via2 ;
        RECT 2897.170 1256.160 2897.450 1256.440 ;
      LAYER met3 ;
        RECT 2881.000 1256.450 2885.000 1256.920 ;
        RECT 2897.145 1256.450 2897.475 1256.465 ;
        RECT 2881.000 1256.320 2897.475 1256.450 ;
        RECT 2884.510 1256.150 2897.475 1256.320 ;
        RECT 2897.145 1256.135 2897.475 1256.150 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 240.650 31.520 240.970 31.580 ;
        RECT 2895.770 31.520 2896.090 31.580 ;
        RECT 240.650 31.380 2896.090 31.520 ;
        RECT 240.650 31.320 240.970 31.380 ;
        RECT 2895.770 31.320 2896.090 31.380 ;
      LAYER via ;
        RECT 240.680 31.320 240.940 31.580 ;
        RECT 2895.800 31.320 2896.060 31.580 ;
      LAYER met2 ;
        RECT 2895.790 1573.675 2896.070 1574.045 ;
        RECT 2895.860 31.610 2896.000 1573.675 ;
        RECT 240.680 31.290 240.940 31.610 ;
        RECT 2895.800 31.290 2896.060 31.610 ;
        RECT 240.740 2.400 240.880 31.290 ;
        RECT 240.530 -4.800 241.090 2.400 ;
      LAYER via2 ;
        RECT 2895.790 1573.720 2896.070 1574.000 ;
      LAYER met3 ;
        RECT 2881.000 1575.240 2885.000 1575.840 ;
        RECT 2884.510 1574.010 2884.810 1575.240 ;
        RECT 2895.765 1574.010 2896.095 1574.025 ;
        RECT 2884.510 1573.710 2896.095 1574.010 ;
        RECT 2895.765 1573.695 2896.095 1573.710 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 21.230 15.880 21.550 15.940 ;
        RECT 258.130 15.880 258.450 15.940 ;
        RECT 21.230 15.740 258.450 15.880 ;
        RECT 21.230 15.680 21.550 15.740 ;
        RECT 258.130 15.680 258.450 15.740 ;
      LAYER via ;
        RECT 21.260 15.680 21.520 15.940 ;
        RECT 258.160 15.680 258.420 15.940 ;
      LAYER met2 ;
        RECT 21.250 1422.035 21.530 1422.405 ;
        RECT 21.320 15.970 21.460 1422.035 ;
        RECT 21.260 15.650 21.520 15.970 ;
        RECT 258.160 15.650 258.420 15.970 ;
        RECT 258.220 2.400 258.360 15.650 ;
        RECT 258.010 -4.800 258.570 2.400 ;
      LAYER via2 ;
        RECT 21.250 1422.080 21.530 1422.360 ;
      LAYER met3 ;
        RECT 35.000 1424.960 39.000 1425.560 ;
        RECT 21.225 1422.370 21.555 1422.385 ;
        RECT 35.270 1422.370 35.570 1424.960 ;
        RECT 21.225 1422.070 35.570 1422.370 ;
        RECT 21.225 1422.055 21.555 1422.070 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 276.070 31.860 276.390 31.920 ;
        RECT 2895.310 31.860 2895.630 31.920 ;
        RECT 276.070 31.720 2895.630 31.860 ;
        RECT 276.070 31.660 276.390 31.720 ;
        RECT 2895.310 31.660 2895.630 31.720 ;
      LAYER via ;
        RECT 276.100 31.660 276.360 31.920 ;
        RECT 2895.340 31.660 2895.600 31.920 ;
      LAYER met2 ;
        RECT 2895.330 1679.075 2895.610 1679.445 ;
        RECT 2895.400 31.950 2895.540 1679.075 ;
        RECT 276.100 31.630 276.360 31.950 ;
        RECT 2895.340 31.630 2895.600 31.950 ;
        RECT 276.160 2.400 276.300 31.630 ;
        RECT 275.950 -4.800 276.510 2.400 ;
      LAYER via2 ;
        RECT 2895.330 1679.120 2895.610 1679.400 ;
      LAYER met3 ;
        RECT 2881.000 1681.320 2885.000 1681.920 ;
        RECT 2884.510 1679.410 2884.810 1681.320 ;
        RECT 2895.305 1679.410 2895.635 1679.425 ;
        RECT 2884.510 1679.110 2895.635 1679.410 ;
        RECT 2895.305 1679.095 2895.635 1679.110 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 294.010 25.400 294.330 25.460 ;
        RECT 2184.150 25.400 2184.470 25.460 ;
        RECT 294.010 25.260 2184.470 25.400 ;
        RECT 294.010 25.200 294.330 25.260 ;
        RECT 2184.150 25.200 2184.470 25.260 ;
      LAYER via ;
        RECT 294.040 25.200 294.300 25.460 ;
        RECT 2184.180 25.200 2184.440 25.460 ;
      LAYER met2 ;
        RECT 2184.210 35.000 2184.490 39.000 ;
        RECT 2184.240 25.490 2184.380 35.000 ;
        RECT 294.040 25.170 294.300 25.490 ;
        RECT 2184.180 25.170 2184.440 25.490 ;
        RECT 294.100 2.400 294.240 25.170 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 45.150 3444.780 45.470 3444.840 ;
        RECT 1815.690 3444.780 1816.010 3444.840 ;
        RECT 45.150 3444.640 1816.010 3444.780 ;
        RECT 45.150 3444.580 45.470 3444.640 ;
        RECT 1815.690 3444.580 1816.010 3444.640 ;
        RECT 311.950 37.980 312.270 38.040 ;
        RECT 62.720 37.840 312.270 37.980 ;
        RECT 45.150 36.960 45.470 37.020 ;
        RECT 62.720 36.960 62.860 37.840 ;
        RECT 311.950 37.780 312.270 37.840 ;
        RECT 45.150 36.820 62.860 36.960 ;
        RECT 45.150 36.760 45.470 36.820 ;
      LAYER via ;
        RECT 45.180 3444.580 45.440 3444.840 ;
        RECT 1815.720 3444.580 1815.980 3444.840 ;
        RECT 45.180 36.760 45.440 37.020 ;
        RECT 311.980 37.780 312.240 38.040 ;
      LAYER met2 ;
        RECT 45.180 3444.550 45.440 3444.870 ;
        RECT 1815.720 3444.550 1815.980 3444.870 ;
        RECT 45.240 37.050 45.380 3444.550 ;
        RECT 1815.780 3435.000 1815.920 3444.550 ;
        RECT 1815.750 3431.000 1816.030 3435.000 ;
        RECT 311.980 37.750 312.240 38.070 ;
        RECT 45.180 36.730 45.440 37.050 ;
        RECT 312.040 2.400 312.180 37.750 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 329.890 32.200 330.210 32.260 ;
        RECT 2894.850 32.200 2895.170 32.260 ;
        RECT 329.890 32.060 2895.170 32.200 ;
        RECT 329.890 32.000 330.210 32.060 ;
        RECT 2894.850 32.000 2895.170 32.060 ;
      LAYER via ;
        RECT 329.920 32.000 330.180 32.260 ;
        RECT 2894.880 32.000 2895.140 32.260 ;
      LAYER met2 ;
        RECT 2894.870 1787.195 2895.150 1787.565 ;
        RECT 2894.940 32.290 2895.080 1787.195 ;
        RECT 329.920 31.970 330.180 32.290 ;
        RECT 2894.880 31.970 2895.140 32.290 ;
        RECT 329.980 2.400 330.120 31.970 ;
        RECT 329.770 -4.800 330.330 2.400 ;
      LAYER via2 ;
        RECT 2894.870 1787.240 2895.150 1787.520 ;
      LAYER met3 ;
        RECT 2881.000 1788.080 2885.000 1788.680 ;
        RECT 2884.510 1787.530 2884.810 1788.080 ;
        RECT 2894.845 1787.530 2895.175 1787.545 ;
        RECT 2884.510 1787.230 2895.175 1787.530 ;
        RECT 2894.845 1787.215 2895.175 1787.230 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 21.690 16.220 22.010 16.280 ;
        RECT 347.370 16.220 347.690 16.280 ;
        RECT 21.690 16.080 347.690 16.220 ;
        RECT 21.690 16.020 22.010 16.080 ;
        RECT 347.370 16.020 347.690 16.080 ;
      LAYER via ;
        RECT 21.720 16.020 21.980 16.280 ;
        RECT 347.400 16.020 347.660 16.280 ;
      LAYER met2 ;
        RECT 21.710 1525.395 21.990 1525.765 ;
        RECT 21.780 16.310 21.920 1525.395 ;
        RECT 21.720 15.990 21.980 16.310 ;
        RECT 347.400 15.990 347.660 16.310 ;
        RECT 347.460 2.400 347.600 15.990 ;
        RECT 347.250 -4.800 347.810 2.400 ;
      LAYER via2 ;
        RECT 21.710 1525.440 21.990 1525.720 ;
      LAYER met3 ;
        RECT 35.000 1528.320 39.000 1528.920 ;
        RECT 21.685 1525.730 22.015 1525.745 ;
        RECT 35.270 1525.730 35.570 1528.320 ;
        RECT 21.685 1525.430 35.570 1525.730 ;
        RECT 21.685 1525.415 22.015 1525.430 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 22.150 16.560 22.470 16.620 ;
        RECT 365.310 16.560 365.630 16.620 ;
        RECT 22.150 16.420 365.630 16.560 ;
        RECT 22.150 16.360 22.470 16.420 ;
        RECT 365.310 16.360 365.630 16.420 ;
      LAYER via ;
        RECT 22.180 16.360 22.440 16.620 ;
        RECT 365.340 16.360 365.600 16.620 ;
      LAYER met2 ;
        RECT 22.170 1628.755 22.450 1629.125 ;
        RECT 22.240 16.650 22.380 1628.755 ;
        RECT 22.180 16.330 22.440 16.650 ;
        RECT 365.340 16.330 365.600 16.650 ;
        RECT 365.400 2.400 365.540 16.330 ;
        RECT 365.190 -4.800 365.750 2.400 ;
      LAYER via2 ;
        RECT 22.170 1628.800 22.450 1629.080 ;
      LAYER met3 ;
        RECT 35.000 1631.000 39.000 1631.600 ;
        RECT 22.145 1629.090 22.475 1629.105 ;
        RECT 35.270 1629.090 35.570 1631.000 ;
        RECT 22.145 1628.790 35.570 1629.090 ;
        RECT 22.145 1628.775 22.475 1628.790 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 383.250 32.540 383.570 32.600 ;
        RECT 2894.390 32.540 2894.710 32.600 ;
        RECT 383.250 32.400 2894.710 32.540 ;
        RECT 383.250 32.340 383.570 32.400 ;
        RECT 2894.390 32.340 2894.710 32.400 ;
      LAYER via ;
        RECT 383.280 32.340 383.540 32.600 ;
        RECT 2894.420 32.340 2894.680 32.600 ;
      LAYER met2 ;
        RECT 2894.410 1891.235 2894.690 1891.605 ;
        RECT 2894.480 32.630 2894.620 1891.235 ;
        RECT 383.280 32.310 383.540 32.630 ;
        RECT 2894.420 32.310 2894.680 32.630 ;
        RECT 383.340 2.400 383.480 32.310 ;
        RECT 383.130 -4.800 383.690 2.400 ;
      LAYER via2 ;
        RECT 2894.410 1891.280 2894.690 1891.560 ;
      LAYER met3 ;
        RECT 2881.000 1894.160 2885.000 1894.760 ;
        RECT 2884.510 1891.570 2884.810 1894.160 ;
        RECT 2894.385 1891.570 2894.715 1891.585 ;
        RECT 2884.510 1891.270 2894.715 1891.570 ;
        RECT 2894.385 1891.255 2894.715 1891.270 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 22.610 16.900 22.930 16.960 ;
        RECT 401.190 16.900 401.510 16.960 ;
        RECT 22.610 16.760 401.510 16.900 ;
        RECT 22.610 16.700 22.930 16.760 ;
        RECT 401.190 16.700 401.510 16.760 ;
      LAYER via ;
        RECT 22.640 16.700 22.900 16.960 ;
        RECT 401.220 16.700 401.480 16.960 ;
      LAYER met2 ;
        RECT 22.630 1732.115 22.910 1732.485 ;
        RECT 22.700 16.990 22.840 1732.115 ;
        RECT 22.640 16.670 22.900 16.990 ;
        RECT 401.220 16.670 401.480 16.990 ;
        RECT 401.280 2.400 401.420 16.670 ;
        RECT 401.070 -4.800 401.630 2.400 ;
      LAYER via2 ;
        RECT 22.630 1732.160 22.910 1732.440 ;
      LAYER met3 ;
        RECT 35.000 1734.360 39.000 1734.960 ;
        RECT 22.605 1732.450 22.935 1732.465 ;
        RECT 35.270 1732.450 35.570 1734.360 ;
        RECT 22.605 1732.150 35.570 1732.450 ;
        RECT 22.605 1732.135 22.935 1732.150 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 46.530 3445.800 46.850 3445.860 ;
        RECT 1530.950 3445.800 1531.270 3445.860 ;
        RECT 46.530 3445.660 1531.270 3445.800 ;
        RECT 46.530 3445.600 46.850 3445.660 ;
        RECT 1530.950 3445.600 1531.270 3445.660 ;
        RECT 46.530 38.320 46.850 38.380 ;
        RECT 46.530 38.180 56.880 38.320 ;
        RECT 46.530 38.120 46.850 38.180 ;
        RECT 56.740 37.980 56.880 38.180 ;
        RECT 62.170 37.980 62.490 38.040 ;
        RECT 56.740 37.840 62.490 37.980 ;
        RECT 62.170 37.780 62.490 37.840 ;
      LAYER via ;
        RECT 46.560 3445.600 46.820 3445.860 ;
        RECT 1530.980 3445.600 1531.240 3445.860 ;
        RECT 46.560 38.120 46.820 38.380 ;
        RECT 62.200 37.780 62.460 38.040 ;
      LAYER met2 ;
        RECT 46.560 3445.570 46.820 3445.890 ;
        RECT 1530.980 3445.570 1531.240 3445.890 ;
        RECT 46.620 38.410 46.760 3445.570 ;
        RECT 1531.040 3435.000 1531.180 3445.570 ;
        RECT 1531.010 3431.000 1531.290 3435.000 ;
        RECT 46.560 38.090 46.820 38.410 ;
        RECT 62.200 37.750 62.460 38.070 ;
        RECT 62.260 2.400 62.400 37.750 ;
        RECT 62.050 -4.800 62.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 44.230 34.580 44.550 34.640 ;
        RECT 44.230 34.440 48.600 34.580 ;
        RECT 44.230 34.380 44.550 34.440 ;
        RECT 48.460 34.240 48.600 34.440 ;
        RECT 55.270 34.240 55.590 34.300 ;
        RECT 48.460 34.100 55.590 34.240 ;
        RECT 55.270 34.040 55.590 34.100 ;
        RECT 55.270 26.760 55.590 26.820 ;
        RECT 419.130 26.760 419.450 26.820 ;
        RECT 55.270 26.620 419.450 26.760 ;
        RECT 55.270 26.560 55.590 26.620 ;
        RECT 419.130 26.560 419.450 26.620 ;
      LAYER via ;
        RECT 44.260 34.380 44.520 34.640 ;
        RECT 55.300 34.040 55.560 34.300 ;
        RECT 55.300 26.560 55.560 26.820 ;
        RECT 419.160 26.560 419.420 26.820 ;
      LAYER met2 ;
        RECT 1957.390 3431.690 1957.670 3431.805 ;
        RECT 1958.350 3431.690 1958.630 3435.000 ;
        RECT 1957.390 3431.550 1958.630 3431.690 ;
        RECT 1957.390 3431.435 1957.670 3431.550 ;
        RECT 1958.350 3431.000 1958.630 3431.550 ;
        RECT 44.250 3425.995 44.530 3426.365 ;
        RECT 44.320 34.670 44.460 3425.995 ;
        RECT 44.260 34.350 44.520 34.670 ;
        RECT 55.300 34.010 55.560 34.330 ;
        RECT 55.360 26.850 55.500 34.010 ;
        RECT 55.300 26.530 55.560 26.850 ;
        RECT 419.160 26.530 419.420 26.850 ;
        RECT 419.220 2.400 419.360 26.530 ;
        RECT 419.010 -4.800 419.570 2.400 ;
      LAYER via2 ;
        RECT 1957.390 3431.480 1957.670 3431.760 ;
        RECT 44.250 3426.040 44.530 3426.320 ;
      LAYER met3 ;
        RECT 1957.365 3431.780 1957.695 3431.785 ;
        RECT 1957.110 3431.770 1957.695 3431.780 ;
        RECT 1956.910 3431.470 1957.695 3431.770 ;
        RECT 1957.110 3431.460 1957.695 3431.470 ;
        RECT 1957.365 3431.455 1957.695 3431.460 ;
        RECT 44.225 3426.330 44.555 3426.345 ;
        RECT 1957.110 3426.330 1957.490 3426.340 ;
        RECT 44.225 3426.030 1957.490 3426.330 ;
        RECT 44.225 3426.015 44.555 3426.030 ;
        RECT 1957.110 3426.020 1957.490 3426.030 ;
      LAYER via3 ;
        RECT 1957.140 3431.460 1957.460 3431.780 ;
        RECT 1957.140 3426.020 1957.460 3426.340 ;
      LAYER met4 ;
        RECT 1957.135 3431.455 1957.465 3431.785 ;
        RECT 1957.150 3426.345 1957.450 3431.455 ;
        RECT 1957.135 3426.015 1957.465 3426.345 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 436.610 32.880 436.930 32.940 ;
        RECT 2893.930 32.880 2894.250 32.940 ;
        RECT 436.610 32.740 2894.250 32.880 ;
        RECT 436.610 32.680 436.930 32.740 ;
        RECT 2893.930 32.680 2894.250 32.740 ;
      LAYER via ;
        RECT 436.640 32.680 436.900 32.940 ;
        RECT 2893.960 32.680 2894.220 32.940 ;
      LAYER met2 ;
        RECT 2893.950 1997.315 2894.230 1997.685 ;
        RECT 2894.020 32.970 2894.160 1997.315 ;
        RECT 436.640 32.650 436.900 32.970 ;
        RECT 2893.960 32.650 2894.220 32.970 ;
        RECT 436.700 2.400 436.840 32.650 ;
        RECT 436.490 -4.800 437.050 2.400 ;
      LAYER via2 ;
        RECT 2893.950 1997.360 2894.230 1997.640 ;
      LAYER met3 ;
        RECT 2881.000 2000.240 2885.000 2000.840 ;
        RECT 2884.510 1997.650 2884.810 2000.240 ;
        RECT 2893.925 1997.650 2894.255 1997.665 ;
        RECT 2884.510 1997.350 2894.255 1997.650 ;
        RECT 2893.925 1997.335 2894.255 1997.350 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 44.690 26.420 45.010 26.480 ;
        RECT 454.550 26.420 454.870 26.480 ;
        RECT 44.690 26.280 454.870 26.420 ;
        RECT 44.690 26.220 45.010 26.280 ;
        RECT 454.550 26.220 454.870 26.280 ;
      LAYER via ;
        RECT 44.720 26.220 44.980 26.480 ;
        RECT 454.580 26.220 454.840 26.480 ;
      LAYER met2 ;
        RECT 2099.990 3431.690 2100.270 3431.805 ;
        RECT 2100.950 3431.690 2101.230 3435.000 ;
        RECT 2099.990 3431.550 2101.230 3431.690 ;
        RECT 2099.990 3431.435 2100.270 3431.550 ;
        RECT 2100.950 3431.000 2101.230 3431.550 ;
        RECT 44.710 3425.315 44.990 3425.685 ;
        RECT 44.780 26.510 44.920 3425.315 ;
        RECT 44.720 26.190 44.980 26.510 ;
        RECT 454.580 26.190 454.840 26.510 ;
        RECT 454.640 2.400 454.780 26.190 ;
        RECT 454.430 -4.800 454.990 2.400 ;
      LAYER via2 ;
        RECT 2099.990 3431.480 2100.270 3431.760 ;
        RECT 44.710 3425.360 44.990 3425.640 ;
      LAYER met3 ;
        RECT 2099.965 3431.780 2100.295 3431.785 ;
        RECT 2099.710 3431.770 2100.295 3431.780 ;
        RECT 2099.510 3431.470 2100.295 3431.770 ;
        RECT 2099.710 3431.460 2100.295 3431.470 ;
        RECT 2099.965 3431.455 2100.295 3431.460 ;
        RECT 44.685 3425.650 45.015 3425.665 ;
        RECT 2099.710 3425.650 2100.090 3425.660 ;
        RECT 44.685 3425.350 2100.090 3425.650 ;
        RECT 44.685 3425.335 45.015 3425.350 ;
        RECT 2099.710 3425.340 2100.090 3425.350 ;
      LAYER via3 ;
        RECT 2099.740 3431.460 2100.060 3431.780 ;
        RECT 2099.740 3425.340 2100.060 3425.660 ;
      LAYER met4 ;
        RECT 2099.735 3431.455 2100.065 3431.785 ;
        RECT 2099.750 3425.665 2100.050 3431.455 ;
        RECT 2099.735 3425.335 2100.065 3425.665 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 23.070 24.720 23.390 24.780 ;
        RECT 472.490 24.720 472.810 24.780 ;
        RECT 23.070 24.580 472.810 24.720 ;
        RECT 23.070 24.520 23.390 24.580 ;
        RECT 472.490 24.520 472.810 24.580 ;
      LAYER via ;
        RECT 23.100 24.520 23.360 24.780 ;
        RECT 472.520 24.520 472.780 24.780 ;
      LAYER met2 ;
        RECT 23.090 1836.155 23.370 1836.525 ;
        RECT 23.160 24.810 23.300 1836.155 ;
        RECT 23.100 24.490 23.360 24.810 ;
        RECT 472.520 24.490 472.780 24.810 ;
        RECT 472.580 2.400 472.720 24.490 ;
        RECT 472.370 -4.800 472.930 2.400 ;
      LAYER via2 ;
        RECT 23.090 1836.200 23.370 1836.480 ;
      LAYER met3 ;
        RECT 35.000 1837.040 39.000 1837.640 ;
        RECT 23.065 1836.490 23.395 1836.505 ;
        RECT 35.270 1836.490 35.570 1837.040 ;
        RECT 23.065 1836.190 35.570 1836.490 ;
        RECT 23.065 1836.175 23.395 1836.190 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 23.530 17.920 23.850 17.980 ;
        RECT 490.430 17.920 490.750 17.980 ;
        RECT 23.530 17.780 490.750 17.920 ;
        RECT 23.530 17.720 23.850 17.780 ;
        RECT 490.430 17.720 490.750 17.780 ;
      LAYER via ;
        RECT 23.560 17.720 23.820 17.980 ;
        RECT 490.460 17.720 490.720 17.980 ;
      LAYER met2 ;
        RECT 23.550 1938.835 23.830 1939.205 ;
        RECT 23.620 18.010 23.760 1938.835 ;
        RECT 23.560 17.690 23.820 18.010 ;
        RECT 490.460 17.690 490.720 18.010 ;
        RECT 490.520 2.400 490.660 17.690 ;
        RECT 490.310 -4.800 490.870 2.400 ;
      LAYER via2 ;
        RECT 23.550 1938.880 23.830 1939.160 ;
      LAYER met3 ;
        RECT 35.000 1940.400 39.000 1941.000 ;
        RECT 23.525 1939.170 23.855 1939.185 ;
        RECT 35.270 1939.170 35.570 1940.400 ;
        RECT 23.525 1938.870 35.570 1939.170 ;
        RECT 23.525 1938.855 23.855 1938.870 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 23.990 19.620 24.310 19.680 ;
        RECT 507.910 19.620 508.230 19.680 ;
        RECT 23.990 19.480 508.230 19.620 ;
        RECT 23.990 19.420 24.310 19.480 ;
        RECT 507.910 19.420 508.230 19.480 ;
      LAYER via ;
        RECT 24.020 19.420 24.280 19.680 ;
        RECT 507.940 19.420 508.200 19.680 ;
      LAYER met2 ;
        RECT 24.010 2042.875 24.290 2043.245 ;
        RECT 24.080 19.710 24.220 2042.875 ;
        RECT 24.020 19.390 24.280 19.710 ;
        RECT 507.940 19.390 508.200 19.710 ;
        RECT 508.000 2.400 508.140 19.390 ;
        RECT 507.790 -4.800 508.350 2.400 ;
      LAYER via2 ;
        RECT 24.010 2042.920 24.290 2043.200 ;
      LAYER met3 ;
        RECT 23.985 2043.210 24.315 2043.225 ;
        RECT 35.000 2043.210 39.000 2043.680 ;
        RECT 23.985 2043.080 39.000 2043.210 ;
        RECT 23.985 2042.910 35.570 2043.080 ;
        RECT 23.985 2042.895 24.315 2042.910 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 525.850 30.500 526.170 30.560 ;
        RECT 2893.470 30.500 2893.790 30.560 ;
        RECT 525.850 30.360 2893.790 30.500 ;
        RECT 525.850 30.300 526.170 30.360 ;
        RECT 2893.470 30.300 2893.790 30.360 ;
      LAYER via ;
        RECT 525.880 30.300 526.140 30.560 ;
        RECT 2893.500 30.300 2893.760 30.560 ;
      LAYER met2 ;
        RECT 2893.490 2104.755 2893.770 2105.125 ;
        RECT 2893.560 30.590 2893.700 2104.755 ;
        RECT 525.880 30.270 526.140 30.590 ;
        RECT 2893.500 30.270 2893.760 30.590 ;
        RECT 525.940 2.400 526.080 30.270 ;
        RECT 525.730 -4.800 526.290 2.400 ;
      LAYER via2 ;
        RECT 2893.490 2104.800 2893.770 2105.080 ;
      LAYER met3 ;
        RECT 2881.000 2106.320 2885.000 2106.920 ;
        RECT 2884.510 2105.090 2884.810 2106.320 ;
        RECT 2893.465 2105.090 2893.795 2105.105 ;
        RECT 2884.510 2104.790 2893.795 2105.090 ;
        RECT 2893.465 2104.775 2893.795 2104.790 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 543.790 30.160 544.110 30.220 ;
        RECT 2893.010 30.160 2893.330 30.220 ;
        RECT 543.790 30.020 2893.330 30.160 ;
        RECT 543.790 29.960 544.110 30.020 ;
        RECT 2893.010 29.960 2893.330 30.020 ;
      LAYER via ;
        RECT 543.820 29.960 544.080 30.220 ;
        RECT 2893.040 29.960 2893.300 30.220 ;
      LAYER met2 ;
        RECT 2893.030 2210.835 2893.310 2211.205 ;
        RECT 2893.100 30.250 2893.240 2210.835 ;
        RECT 543.820 29.930 544.080 30.250 ;
        RECT 2893.040 29.930 2893.300 30.250 ;
        RECT 543.880 2.400 544.020 29.930 ;
        RECT 543.670 -4.800 544.230 2.400 ;
      LAYER via2 ;
        RECT 2893.030 2210.880 2893.310 2211.160 ;
      LAYER met3 ;
        RECT 2881.000 2213.080 2885.000 2213.680 ;
        RECT 2884.510 2211.170 2884.810 2213.080 ;
        RECT 2893.005 2211.170 2893.335 2211.185 ;
        RECT 2884.510 2210.870 2893.335 2211.170 ;
        RECT 2893.005 2210.855 2893.335 2210.870 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 24.450 19.280 24.770 19.340 ;
        RECT 561.730 19.280 562.050 19.340 ;
        RECT 24.450 19.140 562.050 19.280 ;
        RECT 24.450 19.080 24.770 19.140 ;
        RECT 561.730 19.080 562.050 19.140 ;
      LAYER via ;
        RECT 24.480 19.080 24.740 19.340 ;
        RECT 561.760 19.080 562.020 19.340 ;
      LAYER met2 ;
        RECT 24.470 2146.235 24.750 2146.605 ;
        RECT 24.540 19.370 24.680 2146.235 ;
        RECT 24.480 19.050 24.740 19.370 ;
        RECT 561.760 19.050 562.020 19.370 ;
        RECT 561.820 2.400 561.960 19.050 ;
        RECT 561.610 -4.800 562.170 2.400 ;
      LAYER via2 ;
        RECT 24.470 2146.280 24.750 2146.560 ;
      LAYER met3 ;
        RECT 24.445 2146.570 24.775 2146.585 ;
        RECT 35.000 2146.570 39.000 2147.040 ;
        RECT 24.445 2146.440 39.000 2146.570 ;
        RECT 24.445 2146.270 35.570 2146.440 ;
        RECT 24.445 2146.255 24.775 2146.270 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 579.670 29.820 579.990 29.880 ;
        RECT 2892.550 29.820 2892.870 29.880 ;
        RECT 579.670 29.680 2892.870 29.820 ;
        RECT 579.670 29.620 579.990 29.680 ;
        RECT 2892.550 29.620 2892.870 29.680 ;
      LAYER via ;
        RECT 579.700 29.620 579.960 29.880 ;
        RECT 2892.580 29.620 2892.840 29.880 ;
      LAYER met2 ;
        RECT 2892.570 2318.275 2892.850 2318.645 ;
        RECT 2892.640 29.910 2892.780 2318.275 ;
        RECT 579.700 29.590 579.960 29.910 ;
        RECT 2892.580 29.590 2892.840 29.910 ;
        RECT 579.760 2.400 579.900 29.590 ;
        RECT 579.550 -4.800 580.110 2.400 ;
      LAYER via2 ;
        RECT 2892.570 2318.320 2892.850 2318.600 ;
      LAYER met3 ;
        RECT 2881.000 2319.160 2885.000 2319.760 ;
        RECT 2884.510 2318.610 2884.810 2319.160 ;
        RECT 2892.545 2318.610 2892.875 2318.625 ;
        RECT 2884.510 2318.310 2892.875 2318.610 ;
        RECT 2892.545 2318.295 2892.875 2318.310 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2896.710 1360.155 2896.990 1360.525 ;
        RECT 2896.780 17.525 2896.920 1360.155 ;
        RECT 86.110 17.155 86.390 17.525 ;
        RECT 2896.710 17.155 2896.990 17.525 ;
        RECT 86.180 2.400 86.320 17.155 ;
        RECT 85.970 -4.800 86.530 2.400 ;
      LAYER via2 ;
        RECT 2896.710 1360.200 2896.990 1360.480 ;
        RECT 86.110 17.200 86.390 17.480 ;
        RECT 2896.710 17.200 2896.990 17.480 ;
      LAYER met3 ;
        RECT 2881.000 1363.080 2885.000 1363.680 ;
        RECT 2884.510 1360.490 2884.810 1363.080 ;
        RECT 2896.685 1360.490 2897.015 1360.505 ;
        RECT 2884.510 1360.190 2897.015 1360.490 ;
        RECT 2896.685 1360.175 2897.015 1360.190 ;
        RECT 86.085 17.490 86.415 17.505 ;
        RECT 2896.685 17.490 2897.015 17.505 ;
        RECT 86.085 17.190 2897.015 17.490 ;
        RECT 86.085 17.175 86.415 17.190 ;
        RECT 2896.685 17.175 2897.015 17.190 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 597.150 29.480 597.470 29.540 ;
        RECT 2892.090 29.480 2892.410 29.540 ;
        RECT 597.150 29.340 2892.410 29.480 ;
        RECT 597.150 29.280 597.470 29.340 ;
        RECT 2892.090 29.280 2892.410 29.340 ;
      LAYER via ;
        RECT 597.180 29.280 597.440 29.540 ;
        RECT 2892.120 29.280 2892.380 29.540 ;
      LAYER met2 ;
        RECT 2892.110 2422.315 2892.390 2422.685 ;
        RECT 2892.180 29.570 2892.320 2422.315 ;
        RECT 597.180 29.250 597.440 29.570 ;
        RECT 2892.120 29.250 2892.380 29.570 ;
        RECT 597.240 2.400 597.380 29.250 ;
        RECT 597.030 -4.800 597.590 2.400 ;
      LAYER via2 ;
        RECT 2892.110 2422.360 2892.390 2422.640 ;
      LAYER met3 ;
        RECT 2881.000 2425.240 2885.000 2425.840 ;
        RECT 2884.510 2422.650 2884.810 2425.240 ;
        RECT 2892.085 2422.650 2892.415 2422.665 ;
        RECT 2884.510 2422.350 2892.415 2422.650 ;
        RECT 2892.085 2422.335 2892.415 2422.350 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2891.650 2528.395 2891.930 2528.765 ;
        RECT 2891.720 20.245 2891.860 2528.395 ;
        RECT 615.110 19.875 615.390 20.245 ;
        RECT 2891.650 19.875 2891.930 20.245 ;
        RECT 615.180 2.400 615.320 19.875 ;
        RECT 614.970 -4.800 615.530 2.400 ;
      LAYER via2 ;
        RECT 2891.650 2528.440 2891.930 2528.720 ;
        RECT 615.110 19.920 615.390 20.200 ;
        RECT 2891.650 19.920 2891.930 20.200 ;
      LAYER met3 ;
        RECT 2881.000 2531.320 2885.000 2531.920 ;
        RECT 2884.510 2528.730 2884.810 2531.320 ;
        RECT 2891.625 2528.730 2891.955 2528.745 ;
        RECT 2884.510 2528.430 2891.955 2528.730 ;
        RECT 2891.625 2528.415 2891.955 2528.430 ;
        RECT 615.085 20.210 615.415 20.225 ;
        RECT 2891.625 20.210 2891.955 20.225 ;
        RECT 615.085 19.910 2891.955 20.210 ;
        RECT 615.085 19.895 615.415 19.910 ;
        RECT 2891.625 19.895 2891.955 19.910 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 35.490 14.180 35.810 14.240 ;
        RECT 109.550 14.180 109.870 14.240 ;
        RECT 35.490 14.040 109.870 14.180 ;
        RECT 35.490 13.980 35.810 14.040 ;
        RECT 109.550 13.980 109.870 14.040 ;
      LAYER via ;
        RECT 35.520 13.980 35.780 14.240 ;
        RECT 109.580 13.980 109.840 14.240 ;
      LAYER met2 ;
        RECT 35.510 1113.315 35.790 1113.685 ;
        RECT 35.580 14.270 35.720 1113.315 ;
        RECT 35.520 13.950 35.780 14.270 ;
        RECT 109.580 13.950 109.840 14.270 ;
        RECT 109.640 2.400 109.780 13.950 ;
        RECT 109.430 -4.800 109.990 2.400 ;
      LAYER via2 ;
        RECT 35.510 1113.360 35.790 1113.640 ;
      LAYER met3 ;
        RECT 35.000 1116.240 39.000 1116.840 ;
        RECT 35.270 1113.665 35.570 1116.240 ;
        RECT 35.270 1113.350 35.815 1113.665 ;
        RECT 35.485 1113.335 35.815 1113.350 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 47.910 3445.120 48.230 3445.180 ;
        RECT 1673.090 3445.120 1673.410 3445.180 ;
        RECT 47.910 3444.980 1673.410 3445.120 ;
        RECT 47.910 3444.920 48.230 3444.980 ;
        RECT 1673.090 3444.920 1673.410 3444.980 ;
        RECT 47.910 15.200 48.230 15.260 ;
        RECT 133.470 15.200 133.790 15.260 ;
        RECT 47.910 15.060 133.790 15.200 ;
        RECT 47.910 15.000 48.230 15.060 ;
        RECT 133.470 15.000 133.790 15.060 ;
      LAYER via ;
        RECT 47.940 3444.920 48.200 3445.180 ;
        RECT 1673.120 3444.920 1673.380 3445.180 ;
        RECT 47.940 15.000 48.200 15.260 ;
        RECT 133.500 15.000 133.760 15.260 ;
      LAYER met2 ;
        RECT 47.940 3444.890 48.200 3445.210 ;
        RECT 1673.120 3444.890 1673.380 3445.210 ;
        RECT 48.000 15.290 48.140 3444.890 ;
        RECT 1673.180 3435.000 1673.320 3444.890 ;
        RECT 1673.150 3431.000 1673.430 3435.000 ;
        RECT 47.940 14.970 48.200 15.290 ;
        RECT 133.500 14.970 133.760 15.290 ;
        RECT 133.560 2.400 133.700 14.970 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 68.685 18.785 68.855 19.975 ;
      LAYER mcon ;
        RECT 68.685 19.805 68.855 19.975 ;
      LAYER met1 ;
        RECT 35.030 19.960 35.350 20.020 ;
        RECT 68.625 19.960 68.915 20.005 ;
        RECT 35.030 19.820 68.915 19.960 ;
        RECT 35.030 19.760 35.350 19.820 ;
        RECT 68.625 19.775 68.915 19.820 ;
        RECT 68.625 18.940 68.915 18.985 ;
        RECT 151.410 18.940 151.730 19.000 ;
        RECT 68.625 18.800 151.730 18.940 ;
        RECT 68.625 18.755 68.915 18.800 ;
        RECT 151.410 18.740 151.730 18.800 ;
      LAYER via ;
        RECT 35.060 19.760 35.320 20.020 ;
        RECT 151.440 18.740 151.700 19.000 ;
      LAYER met2 ;
        RECT 35.050 1215.995 35.330 1216.365 ;
        RECT 35.120 20.050 35.260 1215.995 ;
        RECT 35.060 19.730 35.320 20.050 ;
        RECT 151.440 18.710 151.700 19.030 ;
        RECT 151.500 2.400 151.640 18.710 ;
        RECT 151.290 -4.800 151.850 2.400 ;
      LAYER via2 ;
        RECT 35.050 1216.040 35.330 1216.320 ;
      LAYER met3 ;
        RECT 35.000 1218.920 39.000 1219.520 ;
        RECT 35.270 1216.345 35.570 1218.920 ;
        RECT 35.025 1216.030 35.570 1216.345 ;
        RECT 35.025 1216.015 35.355 1216.030 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2896.250 1466.235 2896.530 1466.605 ;
        RECT 2896.320 18.885 2896.460 1466.235 ;
        RECT 169.370 18.515 169.650 18.885 ;
        RECT 2896.250 18.515 2896.530 18.885 ;
        RECT 169.440 2.400 169.580 18.515 ;
        RECT 169.230 -4.800 169.790 2.400 ;
      LAYER via2 ;
        RECT 2896.250 1466.280 2896.530 1466.560 ;
        RECT 169.370 18.560 169.650 18.840 ;
        RECT 2896.250 18.560 2896.530 18.840 ;
      LAYER met3 ;
        RECT 2881.000 1469.160 2885.000 1469.760 ;
        RECT 2884.510 1466.570 2884.810 1469.160 ;
        RECT 2896.225 1466.570 2896.555 1466.585 ;
        RECT 2884.510 1466.270 2896.555 1466.570 ;
        RECT 2896.225 1466.255 2896.555 1466.270 ;
        RECT 169.345 18.850 169.675 18.865 ;
        RECT 2896.225 18.850 2896.555 18.865 ;
        RECT 169.345 18.550 2896.555 18.850 ;
        RECT 169.345 18.535 169.675 18.550 ;
        RECT 2896.225 18.535 2896.555 18.550 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 186.830 18.940 187.150 19.000 ;
        RECT 2087.550 18.940 2087.870 19.000 ;
        RECT 186.830 18.800 2087.870 18.940 ;
        RECT 186.830 18.740 187.150 18.800 ;
        RECT 2087.550 18.740 2087.870 18.800 ;
      LAYER via ;
        RECT 186.860 18.740 187.120 19.000 ;
        RECT 2087.580 18.740 2087.840 19.000 ;
      LAYER met2 ;
        RECT 2087.610 35.000 2087.890 39.000 ;
        RECT 2087.640 19.030 2087.780 35.000 ;
        RECT 186.860 18.710 187.120 19.030 ;
        RECT 2087.580 18.710 2087.840 19.030 ;
        RECT 186.920 2.400 187.060 18.710 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 20.770 18.600 21.090 18.660 ;
        RECT 204.770 18.600 205.090 18.660 ;
        RECT 20.770 18.460 205.090 18.600 ;
        RECT 20.770 18.400 21.090 18.460 ;
        RECT 204.770 18.400 205.090 18.460 ;
      LAYER via ;
        RECT 20.800 18.400 21.060 18.660 ;
        RECT 204.800 18.400 205.060 18.660 ;
      LAYER met2 ;
        RECT 20.790 1319.355 21.070 1319.725 ;
        RECT 20.860 18.690 21.000 1319.355 ;
        RECT 20.800 18.370 21.060 18.690 ;
        RECT 204.800 18.370 205.060 18.690 ;
        RECT 204.860 2.400 205.000 18.370 ;
        RECT 204.650 -4.800 205.210 2.400 ;
      LAYER via2 ;
        RECT 20.790 1319.400 21.070 1319.680 ;
      LAYER met3 ;
        RECT 35.000 1322.280 39.000 1322.880 ;
        RECT 20.765 1319.690 21.095 1319.705 ;
        RECT 35.270 1319.690 35.570 1322.280 ;
        RECT 20.765 1319.390 35.570 1319.690 ;
        RECT 20.765 1319.375 21.095 1319.390 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 222.710 18.600 223.030 18.660 ;
        RECT 2135.850 18.600 2136.170 18.660 ;
        RECT 222.710 18.460 2136.170 18.600 ;
        RECT 222.710 18.400 223.030 18.460 ;
        RECT 2135.850 18.400 2136.170 18.460 ;
      LAYER via ;
        RECT 222.740 18.400 223.000 18.660 ;
        RECT 2135.880 18.400 2136.140 18.660 ;
      LAYER met2 ;
        RECT 2135.910 35.000 2136.190 39.000 ;
        RECT 2135.940 18.690 2136.080 35.000 ;
        RECT 222.740 18.370 223.000 18.690 ;
        RECT 2135.880 18.370 2136.140 18.690 ;
        RECT 222.800 2.400 222.940 18.370 ;
        RECT 222.590 -4.800 223.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 20.310 17.240 20.630 17.300 ;
        RECT 2232.450 17.240 2232.770 17.300 ;
        RECT 20.310 17.100 2232.770 17.240 ;
        RECT 20.310 17.040 20.630 17.100 ;
        RECT 2232.450 17.040 2232.770 17.100 ;
      LAYER via ;
        RECT 20.340 17.040 20.600 17.300 ;
        RECT 2232.480 17.040 2232.740 17.300 ;
      LAYER met2 ;
        RECT 2232.510 35.000 2232.790 39.000 ;
        RECT 2232.540 17.330 2232.680 35.000 ;
        RECT 20.340 17.010 20.600 17.330 ;
        RECT 2232.480 17.010 2232.740 17.330 ;
        RECT 20.400 2.400 20.540 17.010 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2280.810 35.000 2281.090 39.000 ;
        RECT 2280.840 25.005 2280.980 35.000 ;
        RECT 44.250 24.635 44.530 25.005 ;
        RECT 2280.770 24.635 2281.050 25.005 ;
        RECT 44.320 2.400 44.460 24.635 ;
        RECT 44.110 -4.800 44.670 2.400 ;
      LAYER via2 ;
        RECT 44.250 24.680 44.530 24.960 ;
        RECT 2280.770 24.680 2281.050 24.960 ;
      LAYER met3 ;
        RECT 44.225 24.970 44.555 24.985 ;
        RECT 2280.745 24.970 2281.075 24.985 ;
        RECT 44.225 24.670 2281.075 24.970 ;
        RECT 44.225 24.655 44.555 24.670 ;
        RECT 2280.745 24.655 2281.075 24.670 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 57.645 38.505 57.815 39.355 ;
      LAYER mcon ;
        RECT 57.645 39.185 57.815 39.355 ;
      LAYER met1 ;
        RECT 45.610 3444.100 45.930 3444.160 ;
        RECT 2385.630 3444.100 2385.950 3444.160 ;
        RECT 45.610 3443.960 2385.950 3444.100 ;
        RECT 45.610 3443.900 45.930 3443.960 ;
        RECT 2385.630 3443.900 2385.950 3443.960 ;
        RECT 45.610 39.340 45.930 39.400 ;
        RECT 57.585 39.340 57.875 39.385 ;
        RECT 45.610 39.200 57.875 39.340 ;
        RECT 45.610 39.140 45.930 39.200 ;
        RECT 57.585 39.155 57.875 39.200 ;
        RECT 57.585 38.660 57.875 38.705 ;
        RECT 57.585 38.520 228.460 38.660 ;
        RECT 57.585 38.475 57.875 38.520 ;
        RECT 228.320 38.320 228.460 38.520 ;
        RECT 246.630 38.320 246.950 38.380 ;
        RECT 228.320 38.180 246.950 38.320 ;
        RECT 246.630 38.120 246.950 38.180 ;
      LAYER via ;
        RECT 45.640 3443.900 45.900 3444.160 ;
        RECT 2385.660 3443.900 2385.920 3444.160 ;
        RECT 45.640 39.140 45.900 39.400 ;
        RECT 246.660 38.120 246.920 38.380 ;
      LAYER met2 ;
        RECT 45.640 3443.870 45.900 3444.190 ;
        RECT 2385.660 3443.870 2385.920 3444.190 ;
        RECT 45.700 39.430 45.840 3443.870 ;
        RECT 2385.720 3435.000 2385.860 3443.870 ;
        RECT 2385.690 3431.000 2385.970 3435.000 ;
        RECT 45.640 39.110 45.900 39.430 ;
        RECT 246.660 38.090 246.920 38.410 ;
        RECT 246.720 2.400 246.860 38.090 ;
        RECT 246.510 -4.800 247.070 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 227.845 37.145 228.015 38.335 ;
      LAYER mcon ;
        RECT 227.845 38.165 228.015 38.335 ;
      LAYER met1 ;
        RECT 46.070 3443.760 46.390 3443.820 ;
        RECT 2528.230 3443.760 2528.550 3443.820 ;
        RECT 46.070 3443.620 2528.550 3443.760 ;
        RECT 46.070 3443.560 46.390 3443.620 ;
        RECT 2528.230 3443.560 2528.550 3443.620 ;
        RECT 46.070 38.660 46.390 38.720 ;
        RECT 46.070 38.520 57.340 38.660 ;
        RECT 46.070 38.460 46.390 38.520 ;
        RECT 57.200 38.320 57.340 38.520 ;
        RECT 227.785 38.320 228.075 38.365 ;
        RECT 57.200 38.180 228.075 38.320 ;
        RECT 227.785 38.135 228.075 38.180 ;
        RECT 227.785 37.300 228.075 37.345 ;
        RECT 264.110 37.300 264.430 37.360 ;
        RECT 227.785 37.160 264.430 37.300 ;
        RECT 227.785 37.115 228.075 37.160 ;
        RECT 264.110 37.100 264.430 37.160 ;
      LAYER via ;
        RECT 46.100 3443.560 46.360 3443.820 ;
        RECT 2528.260 3443.560 2528.520 3443.820 ;
        RECT 46.100 38.460 46.360 38.720 ;
        RECT 264.140 37.100 264.400 37.360 ;
      LAYER met2 ;
        RECT 46.100 3443.530 46.360 3443.850 ;
        RECT 2528.260 3443.530 2528.520 3443.850 ;
        RECT 46.160 38.750 46.300 3443.530 ;
        RECT 2528.320 3435.000 2528.460 3443.530 ;
        RECT 2528.290 3431.000 2528.570 3435.000 ;
        RECT 46.100 38.430 46.360 38.750 ;
        RECT 264.140 37.070 264.400 37.390 ;
        RECT 264.200 2.400 264.340 37.070 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 25.830 17.580 26.150 17.640 ;
        RECT 282.050 17.580 282.370 17.640 ;
        RECT 25.830 17.440 282.370 17.580 ;
        RECT 25.830 17.380 26.150 17.440 ;
        RECT 282.050 17.380 282.370 17.440 ;
      LAYER via ;
        RECT 25.860 17.380 26.120 17.640 ;
        RECT 282.080 17.380 282.340 17.640 ;
      LAYER met2 ;
        RECT 25.850 2555.595 26.130 2555.965 ;
        RECT 25.920 17.670 26.060 2555.595 ;
        RECT 25.860 17.350 26.120 17.670 ;
        RECT 282.080 17.350 282.340 17.670 ;
        RECT 282.140 2.400 282.280 17.350 ;
        RECT 281.930 -4.800 282.490 2.400 ;
      LAYER via2 ;
        RECT 25.850 2555.640 26.130 2555.920 ;
      LAYER met3 ;
        RECT 35.000 2558.520 39.000 2559.120 ;
        RECT 25.825 2555.930 26.155 2555.945 ;
        RECT 35.270 2555.930 35.570 2558.520 ;
        RECT 25.825 2555.630 35.570 2555.930 ;
        RECT 25.825 2555.615 26.155 2555.630 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 299.990 17.580 300.310 17.640 ;
        RECT 2473.950 17.580 2474.270 17.640 ;
        RECT 299.990 17.440 2474.270 17.580 ;
        RECT 299.990 17.380 300.310 17.440 ;
        RECT 2473.950 17.380 2474.270 17.440 ;
      LAYER via ;
        RECT 300.020 17.380 300.280 17.640 ;
        RECT 2473.980 17.380 2474.240 17.640 ;
      LAYER met2 ;
        RECT 2474.010 35.000 2474.290 39.000 ;
        RECT 2474.040 17.670 2474.180 35.000 ;
        RECT 300.020 17.350 300.280 17.670 ;
        RECT 2473.980 17.350 2474.240 17.670 ;
        RECT 300.080 2.400 300.220 17.350 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 317.950 30.755 318.230 31.125 ;
        RECT 318.020 2.400 318.160 30.755 ;
        RECT 317.810 -4.800 318.370 2.400 ;
      LAYER via2 ;
        RECT 317.950 30.800 318.230 31.080 ;
      LAYER met3 ;
        RECT 2881.000 2850.370 2885.000 2850.840 ;
        RECT 2895.510 2850.370 2895.890 2850.380 ;
        RECT 2881.000 2850.240 2895.890 2850.370 ;
        RECT 2884.510 2850.070 2895.890 2850.240 ;
        RECT 2895.510 2850.060 2895.890 2850.070 ;
        RECT 317.925 31.090 318.255 31.105 ;
        RECT 2895.510 31.090 2895.890 31.100 ;
        RECT 317.925 30.790 2895.890 31.090 ;
        RECT 317.925 30.775 318.255 30.790 ;
        RECT 2895.510 30.780 2895.890 30.790 ;
      LAYER via3 ;
        RECT 2895.540 2850.060 2895.860 2850.380 ;
        RECT 2895.540 30.780 2895.860 31.100 ;
      LAYER met4 ;
        RECT 2895.535 2850.055 2895.865 2850.385 ;
        RECT 2895.550 31.105 2895.850 2850.055 ;
        RECT 2895.535 30.775 2895.865 31.105 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2522.310 35.000 2522.590 39.000 ;
        RECT 2522.340 26.365 2522.480 35.000 ;
        RECT 335.890 25.995 336.170 26.365 ;
        RECT 2522.270 25.995 2522.550 26.365 ;
        RECT 335.960 2.400 336.100 25.995 ;
        RECT 335.750 -4.800 336.310 2.400 ;
      LAYER via2 ;
        RECT 335.890 26.040 336.170 26.320 ;
        RECT 2522.270 26.040 2522.550 26.320 ;
      LAYER met3 ;
        RECT 335.865 26.330 336.195 26.345 ;
        RECT 2522.245 26.330 2522.575 26.345 ;
        RECT 335.865 26.030 2522.575 26.330 ;
        RECT 335.865 26.015 336.195 26.030 ;
        RECT 2522.245 26.015 2522.575 26.030 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 26.290 27.100 26.610 27.160 ;
        RECT 353.350 27.100 353.670 27.160 ;
        RECT 26.290 26.960 353.670 27.100 ;
        RECT 26.290 26.900 26.610 26.960 ;
        RECT 353.350 26.900 353.670 26.960 ;
      LAYER via ;
        RECT 26.320 26.900 26.580 27.160 ;
        RECT 353.380 26.900 353.640 27.160 ;
      LAYER met2 ;
        RECT 26.310 2658.275 26.590 2658.645 ;
        RECT 26.380 27.190 26.520 2658.275 ;
        RECT 26.320 26.870 26.580 27.190 ;
        RECT 353.380 26.870 353.640 27.190 ;
        RECT 353.440 2.400 353.580 26.870 ;
        RECT 353.230 -4.800 353.790 2.400 ;
      LAYER via2 ;
        RECT 26.310 2658.320 26.590 2658.600 ;
      LAYER met3 ;
        RECT 35.000 2661.200 39.000 2661.800 ;
        RECT 26.285 2658.610 26.615 2658.625 ;
        RECT 35.270 2658.610 35.570 2661.200 ;
        RECT 26.285 2658.310 35.570 2658.610 ;
        RECT 26.285 2658.295 26.615 2658.310 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 371.310 31.435 371.590 31.805 ;
        RECT 371.380 2.400 371.520 31.435 ;
        RECT 371.170 -4.800 371.730 2.400 ;
      LAYER via2 ;
        RECT 371.310 31.480 371.590 31.760 ;
      LAYER met3 ;
        RECT 2881.000 2956.320 2885.000 2956.920 ;
        RECT 2884.510 2953.730 2884.810 2956.320 ;
        RECT 2894.590 2953.730 2894.970 2953.740 ;
        RECT 2884.510 2953.430 2894.970 2953.730 ;
        RECT 2894.590 2953.420 2894.970 2953.430 ;
        RECT 371.285 31.770 371.615 31.785 ;
        RECT 2894.590 31.770 2894.970 31.780 ;
        RECT 371.285 31.470 2894.970 31.770 ;
        RECT 371.285 31.455 371.615 31.470 ;
        RECT 2894.590 31.460 2894.970 31.470 ;
      LAYER via3 ;
        RECT 2894.620 2953.420 2894.940 2953.740 ;
        RECT 2894.620 31.460 2894.940 31.780 ;
      LAYER met4 ;
        RECT 2894.615 2953.415 2894.945 2953.745 ;
        RECT 2894.630 31.785 2894.930 2953.415 ;
        RECT 2894.615 31.455 2894.945 31.785 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2670.850 3442.995 2671.130 3443.365 ;
        RECT 2670.920 3435.000 2671.060 3442.995 ;
        RECT 2670.890 3431.000 2671.170 3435.000 ;
        RECT 389.250 37.555 389.530 37.925 ;
        RECT 389.320 2.400 389.460 37.555 ;
        RECT 389.110 -4.800 389.670 2.400 ;
      LAYER via2 ;
        RECT 2670.850 3443.040 2671.130 3443.320 ;
        RECT 389.250 37.600 389.530 37.880 ;
      LAYER met3 ;
        RECT 2670.825 3443.330 2671.155 3443.345 ;
        RECT 2848.590 3443.330 2848.970 3443.340 ;
        RECT 2670.825 3443.030 2848.970 3443.330 ;
        RECT 2670.825 3443.015 2671.155 3443.030 ;
        RECT 2848.590 3443.020 2848.970 3443.030 ;
        RECT 389.225 37.890 389.555 37.905 ;
        RECT 2848.590 37.890 2848.970 37.900 ;
        RECT 389.225 37.590 2848.970 37.890 ;
        RECT 389.225 37.575 389.555 37.590 ;
        RECT 2848.590 37.580 2848.970 37.590 ;
      LAYER via3 ;
        RECT 2848.620 3443.020 2848.940 3443.340 ;
        RECT 2848.620 37.580 2848.940 37.900 ;
      LAYER met4 ;
        RECT 2848.615 3443.015 2848.945 3443.345 ;
        RECT 2848.630 3429.050 2848.930 3443.015 ;
        RECT 2848.630 3428.750 2850.770 3429.050 ;
        RECT 2850.470 3425.650 2850.770 3428.750 ;
        RECT 2850.470 3425.350 2851.690 3425.650 ;
        RECT 2851.390 3378.050 2851.690 3425.350 ;
        RECT 2851.390 3377.750 2852.610 3378.050 ;
        RECT 2852.310 3371.250 2852.610 3377.750 ;
        RECT 2852.310 3370.950 2853.530 3371.250 ;
        RECT 2853.230 3296.450 2853.530 3370.950 ;
        RECT 2852.310 3296.150 2853.530 3296.450 ;
        RECT 2852.310 3245.450 2852.610 3296.150 ;
        RECT 2850.470 3245.150 2852.610 3245.450 ;
        RECT 2850.470 3211.450 2850.770 3245.150 ;
        RECT 2850.470 3211.150 2851.690 3211.450 ;
        RECT 2851.390 3187.650 2851.690 3211.150 ;
        RECT 2851.390 3187.350 2852.610 3187.650 ;
        RECT 2852.310 3140.050 2852.610 3187.350 ;
        RECT 2852.310 3139.750 2853.530 3140.050 ;
        RECT 2853.230 3106.050 2853.530 3139.750 ;
        RECT 2852.310 3105.750 2853.530 3106.050 ;
        RECT 2852.310 3058.450 2852.610 3105.750 ;
        RECT 2851.390 3058.150 2852.610 3058.450 ;
        RECT 2851.390 3007.450 2851.690 3058.150 ;
        RECT 2851.390 3007.150 2852.610 3007.450 ;
        RECT 2852.310 2959.850 2852.610 3007.150 ;
        RECT 2850.470 2959.550 2852.610 2959.850 ;
        RECT 2850.470 2946.250 2850.770 2959.550 ;
        RECT 2850.470 2945.950 2855.370 2946.250 ;
        RECT 2855.070 2908.850 2855.370 2945.950 ;
        RECT 2849.550 2908.550 2855.370 2908.850 ;
        RECT 2849.550 2895.250 2849.850 2908.550 ;
        RECT 2849.550 2894.950 2851.690 2895.250 ;
        RECT 2851.390 2864.650 2851.690 2894.950 ;
        RECT 2849.550 2864.350 2851.690 2864.650 ;
        RECT 2849.550 2850.370 2849.850 2864.350 ;
        RECT 2849.550 2850.070 2851.690 2850.370 ;
        RECT 2851.390 2813.650 2851.690 2850.070 ;
        RECT 2850.470 2813.350 2851.690 2813.650 ;
        RECT 2850.470 2766.050 2850.770 2813.350 ;
        RECT 2850.470 2765.750 2851.690 2766.050 ;
        RECT 2851.390 2715.050 2851.690 2765.750 ;
        RECT 2849.550 2714.750 2851.690 2715.050 ;
        RECT 2849.550 2704.850 2849.850 2714.750 ;
        RECT 2849.550 2704.550 2855.370 2704.850 ;
        RECT 2855.070 2657.250 2855.370 2704.550 ;
        RECT 2851.390 2656.950 2855.370 2657.250 ;
        RECT 2851.390 2623.250 2851.690 2656.950 ;
        RECT 2850.470 2622.950 2851.690 2623.250 ;
        RECT 2850.470 2606.250 2850.770 2622.950 ;
        RECT 2850.470 2605.950 2851.690 2606.250 ;
        RECT 2851.390 2599.450 2851.690 2605.950 ;
        RECT 2851.390 2599.150 2856.290 2599.450 ;
        RECT 2855.990 2562.050 2856.290 2599.150 ;
        RECT 2851.390 2561.750 2856.290 2562.050 ;
        RECT 2851.390 2521.250 2851.690 2561.750 ;
        RECT 2849.550 2520.950 2851.690 2521.250 ;
        RECT 2849.550 2477.050 2849.850 2520.950 ;
        RECT 2849.550 2476.750 2850.770 2477.050 ;
        RECT 2850.470 2460.050 2850.770 2476.750 ;
        RECT 2850.470 2459.750 2851.690 2460.050 ;
        RECT 2851.390 2426.050 2851.690 2459.750 ;
        RECT 2851.390 2425.750 2853.530 2426.050 ;
        RECT 2853.230 2378.450 2853.530 2425.750 ;
        RECT 2852.310 2378.150 2853.530 2378.450 ;
        RECT 2852.310 2337.650 2852.610 2378.150 ;
        RECT 2852.310 2337.350 2856.290 2337.650 ;
        RECT 2855.990 2330.850 2856.290 2337.350 ;
        RECT 2850.470 2330.550 2856.290 2330.850 ;
        RECT 2850.470 2293.450 2850.770 2330.550 ;
        RECT 2850.470 2293.150 2851.690 2293.450 ;
        RECT 2851.390 2164.250 2851.690 2293.150 ;
        RECT 2851.390 2163.950 2856.290 2164.250 ;
        RECT 2855.990 2157.450 2856.290 2163.950 ;
        RECT 2851.390 2157.150 2856.290 2157.450 ;
        RECT 2851.390 2133.650 2851.690 2157.150 ;
        RECT 2849.550 2133.350 2851.690 2133.650 ;
        RECT 2849.550 2109.850 2849.850 2133.350 ;
        RECT 2849.550 2109.550 2855.370 2109.850 ;
        RECT 2855.070 2065.650 2855.370 2109.550 ;
        RECT 2850.470 2065.350 2855.370 2065.650 ;
        RECT 2850.470 1919.450 2850.770 2065.350 ;
        RECT 2850.470 1919.150 2852.610 1919.450 ;
        RECT 2852.310 1909.250 2852.610 1919.150 ;
        RECT 2852.310 1908.950 2853.530 1909.250 ;
        RECT 2853.230 1848.050 2853.530 1908.950 ;
        RECT 2852.310 1847.750 2853.530 1848.050 ;
        RECT 2852.310 1800.450 2852.610 1847.750 ;
        RECT 2852.310 1800.150 2853.530 1800.450 ;
        RECT 2853.230 1756.250 2853.530 1800.150 ;
        RECT 2852.310 1755.950 2853.530 1756.250 ;
        RECT 2852.310 1739.250 2852.610 1755.950 ;
        RECT 2851.390 1738.950 2852.610 1739.250 ;
        RECT 2851.390 1735.850 2851.690 1738.950 ;
        RECT 2851.390 1735.550 2852.610 1735.850 ;
        RECT 2852.310 1729.050 2852.610 1735.550 ;
        RECT 2852.310 1728.750 2853.530 1729.050 ;
        RECT 2853.230 1654.250 2853.530 1728.750 ;
        RECT 2852.310 1653.950 2853.530 1654.250 ;
        RECT 2852.310 1603.250 2852.610 1653.950 ;
        RECT 2850.470 1602.950 2852.610 1603.250 ;
        RECT 2850.470 1569.250 2850.770 1602.950 ;
        RECT 2850.470 1568.950 2851.690 1569.250 ;
        RECT 2851.390 1545.450 2851.690 1568.950 ;
        RECT 2851.390 1545.150 2852.610 1545.450 ;
        RECT 2852.310 1497.850 2852.610 1545.150 ;
        RECT 2852.310 1497.550 2853.530 1497.850 ;
        RECT 2853.230 1463.850 2853.530 1497.550 ;
        RECT 2852.310 1463.550 2853.530 1463.850 ;
        RECT 2852.310 1416.250 2852.610 1463.550 ;
        RECT 2851.390 1415.950 2852.610 1416.250 ;
        RECT 2851.390 1375.450 2851.690 1415.950 ;
        RECT 2851.390 1375.150 2853.530 1375.450 ;
        RECT 2853.230 1317.650 2853.530 1375.150 ;
        RECT 2850.470 1317.350 2853.530 1317.650 ;
        RECT 2850.470 1304.050 2850.770 1317.350 ;
        RECT 2850.470 1303.750 2855.370 1304.050 ;
        RECT 2855.070 1266.650 2855.370 1303.750 ;
        RECT 2849.550 1266.350 2855.370 1266.650 ;
        RECT 2849.550 1253.050 2849.850 1266.350 ;
        RECT 2849.550 1252.750 2851.690 1253.050 ;
        RECT 2851.390 1249.650 2851.690 1252.750 ;
        RECT 2851.390 1249.350 2856.290 1249.650 ;
        RECT 2855.990 1208.850 2856.290 1249.350 ;
        RECT 2851.390 1208.550 2856.290 1208.850 ;
        RECT 2851.390 1171.450 2851.690 1208.550 ;
        RECT 2850.470 1171.150 2851.690 1171.450 ;
        RECT 2850.470 1123.850 2850.770 1171.150 ;
        RECT 2850.470 1123.550 2851.690 1123.850 ;
        RECT 2851.390 1072.850 2851.690 1123.550 ;
        RECT 2849.550 1072.550 2851.690 1072.850 ;
        RECT 2849.550 1062.650 2849.850 1072.550 ;
        RECT 2849.550 1062.350 2855.370 1062.650 ;
        RECT 2855.070 1015.050 2855.370 1062.350 ;
        RECT 2851.390 1014.750 2855.370 1015.050 ;
        RECT 2851.390 981.050 2851.690 1014.750 ;
        RECT 2850.470 980.750 2851.690 981.050 ;
        RECT 2850.470 964.050 2850.770 980.750 ;
        RECT 2850.470 963.750 2855.370 964.050 ;
        RECT 2855.070 926.650 2855.370 963.750 ;
        RECT 2850.470 926.350 2855.370 926.650 ;
        RECT 2850.470 919.850 2850.770 926.350 ;
        RECT 2849.550 919.550 2850.770 919.850 ;
        RECT 2849.550 882.450 2849.850 919.550 ;
        RECT 2849.550 882.150 2850.770 882.450 ;
        RECT 2850.470 868.850 2850.770 882.150 ;
        RECT 2850.470 868.550 2851.690 868.850 ;
        RECT 2851.390 834.850 2851.690 868.550 ;
        RECT 2850.470 834.550 2851.690 834.850 ;
        RECT 2850.470 821.250 2850.770 834.550 ;
        RECT 2850.470 820.950 2851.690 821.250 ;
        RECT 2851.390 783.850 2851.690 820.950 ;
        RECT 2849.550 783.550 2851.690 783.850 ;
        RECT 2849.550 770.250 2849.850 783.550 ;
        RECT 2849.550 769.950 2851.690 770.250 ;
        RECT 2851.390 766.850 2851.690 769.950 ;
        RECT 2851.390 766.550 2855.370 766.850 ;
        RECT 2855.070 726.050 2855.370 766.550 ;
        RECT 2851.390 725.750 2855.370 726.050 ;
        RECT 2851.390 688.650 2851.690 725.750 ;
        RECT 2850.470 688.350 2851.690 688.650 ;
        RECT 2850.470 651.250 2850.770 688.350 ;
        RECT 2850.470 650.950 2851.690 651.250 ;
        RECT 2851.390 522.050 2851.690 650.950 ;
        RECT 2851.390 521.750 2856.290 522.050 ;
        RECT 2855.990 515.250 2856.290 521.750 ;
        RECT 2851.390 514.950 2856.290 515.250 ;
        RECT 2851.390 491.450 2851.690 514.950 ;
        RECT 2849.550 491.150 2851.690 491.450 ;
        RECT 2849.550 467.650 2849.850 491.150 ;
        RECT 2849.550 467.350 2855.370 467.650 ;
        RECT 2855.070 423.450 2855.370 467.350 ;
        RECT 2850.470 423.150 2855.370 423.450 ;
        RECT 2850.470 324.850 2850.770 423.150 ;
        RECT 2849.550 324.550 2850.770 324.850 ;
        RECT 2849.550 297.650 2849.850 324.550 ;
        RECT 2849.550 297.350 2852.610 297.650 ;
        RECT 2852.310 256.850 2852.610 297.350 ;
        RECT 2851.390 256.550 2852.610 256.850 ;
        RECT 2851.390 188.850 2851.690 256.550 ;
        RECT 2850.470 188.550 2851.690 188.850 ;
        RECT 2850.470 168.450 2850.770 188.550 ;
        RECT 2850.470 168.150 2851.690 168.450 ;
        RECT 2851.390 114.050 2851.690 168.150 ;
        RECT 2850.470 113.750 2851.690 114.050 ;
        RECT 2850.470 97.050 2850.770 113.750 ;
        RECT 2849.550 96.750 2850.770 97.050 ;
        RECT 2849.550 87.290 2849.850 96.750 ;
        RECT 2849.110 86.110 2850.290 87.290 ;
        RECT 2849.110 79.310 2850.290 80.490 ;
        RECT 2849.550 42.650 2849.850 79.310 ;
        RECT 2848.630 42.350 2849.850 42.650 ;
        RECT 2848.630 37.905 2848.930 42.350 ;
        RECT 2848.615 37.575 2848.945 37.905 ;
      LAYER met5 ;
        RECT 2842.460 85.900 2850.500 87.500 ;
        RECT 2842.460 80.700 2844.060 85.900 ;
        RECT 2842.460 79.100 2850.500 80.700 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 407.190 32.115 407.470 32.485 ;
        RECT 407.260 2.400 407.400 32.115 ;
        RECT 407.050 -4.800 407.610 2.400 ;
      LAYER via2 ;
        RECT 407.190 32.160 407.470 32.440 ;
      LAYER met3 ;
        RECT 2881.000 3063.080 2885.000 3063.680 ;
        RECT 2884.510 3060.490 2884.810 3063.080 ;
        RECT 2893.670 3060.490 2894.050 3060.500 ;
        RECT 2884.510 3060.190 2894.050 3060.490 ;
        RECT 2893.670 3060.180 2894.050 3060.190 ;
        RECT 407.165 32.450 407.495 32.465 ;
        RECT 2893.670 32.450 2894.050 32.460 ;
        RECT 407.165 32.150 2894.050 32.450 ;
        RECT 407.165 32.135 407.495 32.150 ;
        RECT 2893.670 32.140 2894.050 32.150 ;
      LAYER via3 ;
        RECT 2893.700 3060.180 2894.020 3060.500 ;
        RECT 2893.700 32.140 2894.020 32.460 ;
      LAYER met4 ;
        RECT 2893.695 3060.175 2894.025 3060.505 ;
        RECT 2893.710 32.465 2894.010 3060.175 ;
        RECT 2893.695 32.135 2894.025 32.465 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 34.570 18.940 34.890 19.000 ;
        RECT 68.150 18.940 68.470 19.000 ;
        RECT 34.570 18.800 68.470 18.940 ;
        RECT 34.570 18.740 34.890 18.800 ;
        RECT 68.150 18.740 68.470 18.800 ;
      LAYER via ;
        RECT 34.600 18.740 34.860 19.000 ;
        RECT 68.180 18.740 68.440 19.000 ;
      LAYER met2 ;
        RECT 34.590 2248.235 34.870 2248.605 ;
        RECT 34.660 19.030 34.800 2248.235 ;
        RECT 34.600 18.710 34.860 19.030 ;
        RECT 68.180 18.710 68.440 19.030 ;
        RECT 68.240 2.400 68.380 18.710 ;
        RECT 68.030 -4.800 68.590 2.400 ;
      LAYER via2 ;
        RECT 34.590 2248.280 34.870 2248.560 ;
      LAYER met3 ;
        RECT 35.000 2249.120 39.000 2249.720 ;
        RECT 34.565 2248.570 34.895 2248.585 ;
        RECT 35.270 2248.570 35.570 2249.120 ;
        RECT 34.565 2248.270 35.570 2248.570 ;
        RECT 34.565 2248.255 34.895 2248.270 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 424.670 32.795 424.950 33.165 ;
        RECT 424.740 2.400 424.880 32.795 ;
        RECT 424.530 -4.800 425.090 2.400 ;
      LAYER via2 ;
        RECT 424.670 32.840 424.950 33.120 ;
      LAYER met3 ;
        RECT 2881.000 3169.160 2885.000 3169.760 ;
        RECT 2884.510 3167.250 2884.810 3169.160 ;
        RECT 2892.750 3167.250 2893.130 3167.260 ;
        RECT 2884.510 3166.950 2893.130 3167.250 ;
        RECT 2892.750 3166.940 2893.130 3166.950 ;
        RECT 424.645 33.130 424.975 33.145 ;
        RECT 2892.750 33.130 2893.130 33.140 ;
        RECT 424.645 32.830 2893.130 33.130 ;
        RECT 424.645 32.815 424.975 32.830 ;
        RECT 2892.750 32.820 2893.130 32.830 ;
      LAYER via3 ;
        RECT 2892.780 3166.940 2893.100 3167.260 ;
        RECT 2892.780 32.820 2893.100 33.140 ;
      LAYER met4 ;
        RECT 2892.775 3166.935 2893.105 3167.265 ;
        RECT 2892.790 33.145 2893.090 3166.935 ;
        RECT 2892.775 32.815 2893.105 33.145 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 26.750 18.260 27.070 18.320 ;
        RECT 442.590 18.260 442.910 18.320 ;
        RECT 26.750 18.120 442.910 18.260 ;
        RECT 26.750 18.060 27.070 18.120 ;
        RECT 442.590 18.060 442.910 18.120 ;
      LAYER via ;
        RECT 26.780 18.060 27.040 18.320 ;
        RECT 442.620 18.060 442.880 18.320 ;
      LAYER met2 ;
        RECT 26.770 2761.635 27.050 2762.005 ;
        RECT 26.840 18.350 26.980 2761.635 ;
        RECT 26.780 18.030 27.040 18.350 ;
        RECT 442.620 18.030 442.880 18.350 ;
        RECT 442.680 2.400 442.820 18.030 ;
        RECT 442.470 -4.800 443.030 2.400 ;
      LAYER via2 ;
        RECT 26.770 2761.680 27.050 2761.960 ;
      LAYER met3 ;
        RECT 35.000 2764.560 39.000 2765.160 ;
        RECT 26.745 2761.970 27.075 2761.985 ;
        RECT 35.270 2761.970 35.570 2764.560 ;
        RECT 26.745 2761.670 35.570 2761.970 ;
        RECT 26.745 2761.655 27.075 2761.670 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 460.530 18.260 460.850 18.320 ;
        RECT 2570.550 18.260 2570.870 18.320 ;
        RECT 460.530 18.120 2570.870 18.260 ;
        RECT 460.530 18.060 460.850 18.120 ;
        RECT 2570.550 18.060 2570.870 18.120 ;
      LAYER via ;
        RECT 460.560 18.060 460.820 18.320 ;
        RECT 2570.580 18.060 2570.840 18.320 ;
      LAYER met2 ;
        RECT 2570.610 35.000 2570.890 39.000 ;
        RECT 2570.640 18.350 2570.780 35.000 ;
        RECT 460.560 18.030 460.820 18.350 ;
        RECT 2570.580 18.030 2570.840 18.350 ;
        RECT 460.620 2.400 460.760 18.030 ;
        RECT 460.410 -4.800 460.970 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 27.210 24.380 27.530 24.440 ;
        RECT 478.470 24.380 478.790 24.440 ;
        RECT 27.210 24.240 478.790 24.380 ;
        RECT 27.210 24.180 27.530 24.240 ;
        RECT 478.470 24.180 478.790 24.240 ;
      LAYER via ;
        RECT 27.240 24.180 27.500 24.440 ;
        RECT 478.500 24.180 478.760 24.440 ;
      LAYER met2 ;
        RECT 27.230 2864.315 27.510 2864.685 ;
        RECT 27.300 24.470 27.440 2864.315 ;
        RECT 27.240 24.150 27.500 24.470 ;
        RECT 478.500 24.150 478.760 24.470 ;
        RECT 478.560 2.400 478.700 24.150 ;
        RECT 478.350 -4.800 478.910 2.400 ;
      LAYER via2 ;
        RECT 27.230 2864.360 27.510 2864.640 ;
      LAYER met3 ;
        RECT 35.000 2867.240 39.000 2867.840 ;
        RECT 27.205 2864.650 27.535 2864.665 ;
        RECT 35.270 2864.650 35.570 2867.240 ;
        RECT 27.205 2864.350 35.570 2864.650 ;
        RECT 27.205 2864.335 27.535 2864.350 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 496.410 17.920 496.730 17.980 ;
        RECT 2618.850 17.920 2619.170 17.980 ;
        RECT 496.410 17.780 2619.170 17.920 ;
        RECT 496.410 17.720 496.730 17.780 ;
        RECT 2618.850 17.720 2619.170 17.780 ;
      LAYER via ;
        RECT 496.440 17.720 496.700 17.980 ;
        RECT 2618.880 17.720 2619.140 17.980 ;
      LAYER met2 ;
        RECT 2618.910 35.000 2619.190 39.000 ;
        RECT 2618.940 18.010 2619.080 35.000 ;
        RECT 496.440 17.690 496.700 18.010 ;
        RECT 2618.880 17.690 2619.140 18.010 ;
        RECT 496.500 2.400 496.640 17.690 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 513.910 33.475 514.190 33.845 ;
        RECT 513.980 2.400 514.120 33.475 ;
        RECT 513.770 -4.800 514.330 2.400 ;
      LAYER via2 ;
        RECT 513.910 33.520 514.190 33.800 ;
      LAYER met3 ;
        RECT 2881.000 3275.240 2885.000 3275.840 ;
        RECT 2884.510 3273.330 2884.810 3275.240 ;
        RECT 2891.830 3273.330 2892.210 3273.340 ;
        RECT 2884.510 3273.030 2892.210 3273.330 ;
        RECT 2891.830 3273.020 2892.210 3273.030 ;
        RECT 513.885 33.810 514.215 33.825 ;
        RECT 2891.830 33.810 2892.210 33.820 ;
        RECT 513.885 33.510 2892.210 33.810 ;
        RECT 513.885 33.495 514.215 33.510 ;
        RECT 2891.830 33.500 2892.210 33.510 ;
      LAYER via3 ;
        RECT 2891.860 3273.020 2892.180 3273.340 ;
        RECT 2891.860 33.500 2892.180 33.820 ;
      LAYER met4 ;
        RECT 2891.855 3273.015 2892.185 3273.345 ;
        RECT 2891.870 33.825 2892.170 3273.015 ;
        RECT 2891.855 33.495 2892.185 33.825 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 531.850 23.275 532.130 23.645 ;
        RECT 531.920 2.400 532.060 23.275 ;
        RECT 531.710 -4.800 532.270 2.400 ;
      LAYER via2 ;
        RECT 531.850 23.320 532.130 23.600 ;
      LAYER met3 ;
        RECT 35.000 2970.600 39.000 2971.200 ;
        RECT 25.110 2968.010 25.490 2968.020 ;
        RECT 35.270 2968.010 35.570 2970.600 ;
        RECT 25.110 2967.710 35.570 2968.010 ;
        RECT 25.110 2967.700 25.490 2967.710 ;
        RECT 25.110 23.610 25.490 23.620 ;
        RECT 531.825 23.610 532.155 23.625 ;
        RECT 25.110 23.310 532.155 23.610 ;
        RECT 25.110 23.300 25.490 23.310 ;
        RECT 531.825 23.295 532.155 23.310 ;
      LAYER via3 ;
        RECT 25.140 2967.700 25.460 2968.020 ;
        RECT 25.140 23.300 25.460 23.620 ;
      LAYER met4 ;
        RECT 25.135 2967.695 25.465 2968.025 ;
        RECT 25.150 23.625 25.450 2967.695 ;
        RECT 25.135 23.295 25.465 23.625 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 549.790 15.795 550.070 16.165 ;
        RECT 549.860 2.400 550.000 15.795 ;
        RECT 549.650 -4.800 550.210 2.400 ;
      LAYER via2 ;
        RECT 549.790 15.840 550.070 16.120 ;
      LAYER met3 ;
        RECT 35.000 3073.280 39.000 3073.880 ;
        RECT 26.030 3070.690 26.410 3070.700 ;
        RECT 35.270 3070.690 35.570 3073.280 ;
        RECT 26.030 3070.390 35.570 3070.690 ;
        RECT 26.030 3070.380 26.410 3070.390 ;
        RECT 26.030 16.130 26.410 16.140 ;
        RECT 549.765 16.130 550.095 16.145 ;
        RECT 26.030 15.830 550.095 16.130 ;
        RECT 26.030 15.820 26.410 15.830 ;
        RECT 549.765 15.815 550.095 15.830 ;
      LAYER via3 ;
        RECT 26.060 3070.380 26.380 3070.700 ;
        RECT 26.060 15.820 26.380 16.140 ;
      LAYER met4 ;
        RECT 26.055 3070.375 26.385 3070.705 ;
        RECT 26.070 16.145 26.370 3070.375 ;
        RECT 26.055 15.815 26.385 16.145 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 567.730 19.875 568.010 20.245 ;
        RECT 567.800 2.400 567.940 19.875 ;
        RECT 567.590 -4.800 568.150 2.400 ;
      LAYER via2 ;
        RECT 567.730 19.920 568.010 20.200 ;
      LAYER met3 ;
        RECT 35.000 3176.640 39.000 3177.240 ;
        RECT 26.950 3174.730 27.330 3174.740 ;
        RECT 35.270 3174.730 35.570 3176.640 ;
        RECT 26.950 3174.430 35.570 3174.730 ;
        RECT 26.950 3174.420 27.330 3174.430 ;
        RECT 26.950 20.210 27.330 20.220 ;
        RECT 567.705 20.210 568.035 20.225 ;
        RECT 26.950 19.910 568.035 20.210 ;
        RECT 26.950 19.900 27.330 19.910 ;
        RECT 567.705 19.895 568.035 19.910 ;
      LAYER via3 ;
        RECT 26.980 3174.420 27.300 3174.740 ;
        RECT 26.980 19.900 27.300 20.220 ;
      LAYER met4 ;
        RECT 26.975 3174.415 27.305 3174.745 ;
        RECT 26.990 20.225 27.290 3174.415 ;
        RECT 26.975 19.895 27.305 20.225 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 585.650 24.720 585.970 24.780 ;
        RECT 2667.150 24.720 2667.470 24.780 ;
        RECT 585.650 24.580 2667.470 24.720 ;
        RECT 585.650 24.520 585.970 24.580 ;
        RECT 2667.150 24.520 2667.470 24.580 ;
      LAYER via ;
        RECT 585.680 24.520 585.940 24.780 ;
        RECT 2667.180 24.520 2667.440 24.780 ;
      LAYER met2 ;
        RECT 2667.210 35.000 2667.490 39.000 ;
        RECT 2667.240 24.810 2667.380 35.000 ;
        RECT 585.680 24.490 585.940 24.810 ;
        RECT 2667.180 24.490 2667.440 24.810 ;
        RECT 585.740 2.400 585.880 24.490 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 24.910 14.520 25.230 14.580 ;
        RECT 91.610 14.520 91.930 14.580 ;
        RECT 24.910 14.380 91.930 14.520 ;
        RECT 24.910 14.320 25.230 14.380 ;
        RECT 91.610 14.320 91.930 14.380 ;
      LAYER via ;
        RECT 24.940 14.320 25.200 14.580 ;
        RECT 91.640 14.320 91.900 14.580 ;
      LAYER met2 ;
        RECT 24.930 2349.555 25.210 2349.925 ;
        RECT 25.000 14.610 25.140 2349.555 ;
        RECT 24.940 14.290 25.200 14.610 ;
        RECT 91.640 14.290 91.900 14.610 ;
        RECT 91.700 2.400 91.840 14.290 ;
        RECT 91.490 -4.800 92.050 2.400 ;
      LAYER via2 ;
        RECT 24.930 2349.600 25.210 2349.880 ;
      LAYER met3 ;
        RECT 35.000 2352.480 39.000 2353.080 ;
        RECT 24.905 2349.890 25.235 2349.905 ;
        RECT 35.270 2349.890 35.570 2352.480 ;
        RECT 24.905 2349.590 35.570 2349.890 ;
        RECT 24.905 2349.575 25.235 2349.590 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 603.130 24.380 603.450 24.440 ;
        RECT 2715.450 24.380 2715.770 24.440 ;
        RECT 603.130 24.240 2715.770 24.380 ;
        RECT 603.130 24.180 603.450 24.240 ;
        RECT 2715.450 24.180 2715.770 24.240 ;
      LAYER via ;
        RECT 603.160 24.180 603.420 24.440 ;
        RECT 2715.480 24.180 2715.740 24.440 ;
      LAYER met2 ;
        RECT 2715.510 35.000 2715.790 39.000 ;
        RECT 2715.540 24.470 2715.680 35.000 ;
        RECT 603.160 24.150 603.420 24.470 ;
        RECT 2715.480 24.150 2715.740 24.470 ;
        RECT 603.220 2.400 603.360 24.150 ;
        RECT 603.010 -4.800 603.570 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 621.070 24.040 621.390 24.100 ;
        RECT 2763.750 24.040 2764.070 24.100 ;
        RECT 621.070 23.900 2764.070 24.040 ;
        RECT 621.070 23.840 621.390 23.900 ;
        RECT 2763.750 23.840 2764.070 23.900 ;
      LAYER via ;
        RECT 621.100 23.840 621.360 24.100 ;
        RECT 2763.780 23.840 2764.040 24.100 ;
      LAYER met2 ;
        RECT 2763.810 35.000 2764.090 39.000 ;
        RECT 2763.840 24.130 2763.980 35.000 ;
        RECT 621.100 23.810 621.360 24.130 ;
        RECT 2763.780 23.810 2764.040 24.130 ;
        RECT 621.160 2.400 621.300 23.810 ;
        RECT 620.950 -4.800 621.510 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 25.370 15.540 25.690 15.600 ;
        RECT 115.530 15.540 115.850 15.600 ;
        RECT 25.370 15.400 115.850 15.540 ;
        RECT 25.370 15.340 25.690 15.400 ;
        RECT 115.530 15.340 115.850 15.400 ;
      LAYER via ;
        RECT 25.400 15.340 25.660 15.600 ;
        RECT 115.560 15.340 115.820 15.600 ;
      LAYER met2 ;
        RECT 25.390 2452.235 25.670 2452.605 ;
        RECT 25.460 15.630 25.600 2452.235 ;
        RECT 25.400 15.310 25.660 15.630 ;
        RECT 115.560 15.310 115.820 15.630 ;
        RECT 115.620 2.400 115.760 15.310 ;
        RECT 115.410 -4.800 115.970 2.400 ;
      LAYER via2 ;
        RECT 25.390 2452.280 25.670 2452.560 ;
      LAYER met3 ;
        RECT 35.000 2455.160 39.000 2455.760 ;
        RECT 25.365 2452.570 25.695 2452.585 ;
        RECT 35.270 2452.570 35.570 2455.160 ;
        RECT 25.365 2452.270 35.570 2452.570 ;
        RECT 25.365 2452.255 25.695 2452.270 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2891.190 2635.835 2891.470 2636.205 ;
        RECT 2891.260 18.205 2891.400 2635.835 ;
        RECT 139.470 17.835 139.750 18.205 ;
        RECT 2891.190 17.835 2891.470 18.205 ;
        RECT 139.540 2.400 139.680 17.835 ;
        RECT 139.330 -4.800 139.890 2.400 ;
      LAYER via2 ;
        RECT 2891.190 2635.880 2891.470 2636.160 ;
        RECT 139.470 17.880 139.750 18.160 ;
        RECT 2891.190 17.880 2891.470 18.160 ;
      LAYER met3 ;
        RECT 2881.000 2638.080 2885.000 2638.680 ;
        RECT 2884.510 2636.170 2884.810 2638.080 ;
        RECT 2891.165 2636.170 2891.495 2636.185 ;
        RECT 2884.510 2635.870 2891.495 2636.170 ;
        RECT 2891.165 2635.855 2891.495 2635.870 ;
        RECT 139.445 18.170 139.775 18.185 ;
        RECT 2891.165 18.170 2891.495 18.185 ;
        RECT 139.445 17.870 2891.495 18.170 ;
        RECT 139.445 17.855 139.775 17.870 ;
        RECT 2891.165 17.855 2891.495 17.870 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2329.110 35.000 2329.390 39.000 ;
        RECT 2329.140 27.725 2329.280 35.000 ;
        RECT 157.410 27.355 157.690 27.725 ;
        RECT 2329.070 27.355 2329.350 27.725 ;
        RECT 157.480 2.400 157.620 27.355 ;
        RECT 157.270 -4.800 157.830 2.400 ;
      LAYER via2 ;
        RECT 157.410 27.400 157.690 27.680 ;
        RECT 2329.070 27.400 2329.350 27.680 ;
      LAYER met3 ;
        RECT 157.385 27.690 157.715 27.705 ;
        RECT 2329.045 27.690 2329.375 27.705 ;
        RECT 157.385 27.390 2329.375 27.690 ;
        RECT 157.385 27.375 157.715 27.390 ;
        RECT 2329.045 27.375 2329.375 27.390 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 174.890 19.195 175.170 19.565 ;
        RECT 174.960 2.400 175.100 19.195 ;
        RECT 174.750 -4.800 175.310 2.400 ;
      LAYER via2 ;
        RECT 174.890 19.240 175.170 19.520 ;
      LAYER met3 ;
        RECT 2881.000 2744.160 2885.000 2744.760 ;
        RECT 2884.510 2742.250 2884.810 2744.160 ;
        RECT 2896.430 2742.250 2896.810 2742.260 ;
        RECT 2884.510 2741.950 2896.810 2742.250 ;
        RECT 2896.430 2741.940 2896.810 2741.950 ;
        RECT 174.865 19.530 175.195 19.545 ;
        RECT 2896.430 19.530 2896.810 19.540 ;
        RECT 174.865 19.230 2896.810 19.530 ;
        RECT 174.865 19.215 175.195 19.230 ;
        RECT 2896.430 19.220 2896.810 19.230 ;
      LAYER via3 ;
        RECT 2896.460 2741.940 2896.780 2742.260 ;
        RECT 2896.460 19.220 2896.780 19.540 ;
      LAYER met4 ;
        RECT 2896.455 2741.935 2896.785 2742.265 ;
        RECT 2896.470 19.545 2896.770 2741.935 ;
        RECT 2896.455 19.215 2896.785 19.545 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2377.410 35.000 2377.690 39.000 ;
        RECT 2377.440 27.045 2377.580 35.000 ;
        RECT 192.830 26.675 193.110 27.045 ;
        RECT 2377.370 26.675 2377.650 27.045 ;
        RECT 192.900 2.400 193.040 26.675 ;
        RECT 192.690 -4.800 193.250 2.400 ;
      LAYER via2 ;
        RECT 192.830 26.720 193.110 27.000 ;
        RECT 2377.370 26.720 2377.650 27.000 ;
      LAYER met3 ;
        RECT 192.805 27.010 193.135 27.025 ;
        RECT 2377.345 27.010 2377.675 27.025 ;
        RECT 192.805 26.710 2377.675 27.010 ;
        RECT 192.805 26.695 193.135 26.710 ;
        RECT 2377.345 26.695 2377.675 26.710 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2425.710 35.000 2425.990 39.000 ;
        RECT 2425.740 25.685 2425.880 35.000 ;
        RECT 210.770 25.315 211.050 25.685 ;
        RECT 2425.670 25.315 2425.950 25.685 ;
        RECT 210.840 2.400 210.980 25.315 ;
        RECT 210.630 -4.800 211.190 2.400 ;
      LAYER via2 ;
        RECT 210.770 25.360 211.050 25.640 ;
        RECT 2425.670 25.360 2425.950 25.640 ;
      LAYER met3 ;
        RECT 210.745 25.650 211.075 25.665 ;
        RECT 2425.645 25.650 2425.975 25.665 ;
        RECT 210.745 25.350 2425.975 25.650 ;
        RECT 210.745 25.335 211.075 25.350 ;
        RECT 2425.645 25.335 2425.975 25.350 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 47.450 3444.440 47.770 3444.500 ;
        RECT 2243.490 3444.440 2243.810 3444.500 ;
        RECT 47.450 3444.300 2243.810 3444.440 ;
        RECT 47.450 3444.240 47.770 3444.300 ;
        RECT 2243.490 3444.240 2243.810 3444.300 ;
        RECT 47.450 39.000 47.770 39.060 ;
        RECT 47.450 38.860 228.920 39.000 ;
        RECT 47.450 38.800 47.770 38.860 ;
        RECT 228.780 38.720 228.920 38.860 ;
        RECT 228.690 38.460 229.010 38.720 ;
      LAYER via ;
        RECT 47.480 3444.240 47.740 3444.500 ;
        RECT 2243.520 3444.240 2243.780 3444.500 ;
        RECT 47.480 38.800 47.740 39.060 ;
        RECT 228.720 38.460 228.980 38.720 ;
      LAYER met2 ;
        RECT 47.480 3444.210 47.740 3444.530 ;
        RECT 2243.520 3444.210 2243.780 3444.530 ;
        RECT 47.540 39.090 47.680 3444.210 ;
        RECT 2243.580 3435.000 2243.720 3444.210 ;
        RECT 2243.550 3431.000 2243.830 3435.000 ;
        RECT 47.480 38.770 47.740 39.090 ;
        RECT 228.720 38.430 228.980 38.750 ;
        RECT 228.780 2.400 228.920 38.430 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 50.210 20.300 50.530 20.360 ;
        RECT 445.350 20.300 445.670 20.360 ;
        RECT 50.210 20.160 445.670 20.300 ;
        RECT 50.210 20.100 50.530 20.160 ;
        RECT 445.350 20.100 445.670 20.160 ;
      LAYER via ;
        RECT 50.240 20.100 50.500 20.360 ;
        RECT 445.380 20.100 445.640 20.360 ;
      LAYER met2 ;
        RECT 445.410 35.000 445.690 39.000 ;
        RECT 445.440 20.390 445.580 35.000 ;
        RECT 50.240 20.070 50.500 20.390 ;
        RECT 445.380 20.070 445.640 20.390 ;
        RECT 50.300 2.400 50.440 20.070 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 252.610 22.000 252.930 22.060 ;
        RECT 928.350 22.000 928.670 22.060 ;
        RECT 252.610 21.860 928.670 22.000 ;
        RECT 252.610 21.800 252.930 21.860 ;
        RECT 928.350 21.800 928.670 21.860 ;
      LAYER via ;
        RECT 252.640 21.800 252.900 22.060 ;
        RECT 928.380 21.800 928.640 22.060 ;
      LAYER met2 ;
        RECT 928.410 35.000 928.690 39.000 ;
        RECT 928.440 22.090 928.580 35.000 ;
        RECT 252.640 21.770 252.900 22.090 ;
        RECT 928.380 21.770 928.640 22.090 ;
        RECT 252.700 2.400 252.840 21.770 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 270.090 22.340 270.410 22.400 ;
        RECT 976.650 22.340 976.970 22.400 ;
        RECT 270.090 22.200 976.970 22.340 ;
        RECT 270.090 22.140 270.410 22.200 ;
        RECT 976.650 22.140 976.970 22.200 ;
      LAYER via ;
        RECT 270.120 22.140 270.380 22.400 ;
        RECT 976.680 22.140 976.940 22.400 ;
      LAYER met2 ;
        RECT 976.710 35.000 976.990 39.000 ;
        RECT 976.740 22.430 976.880 35.000 ;
        RECT 270.120 22.110 270.380 22.430 ;
        RECT 976.680 22.110 976.940 22.430 ;
        RECT 270.180 2.400 270.320 22.110 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 288.030 25.740 288.350 25.800 ;
        RECT 1024.950 25.740 1025.270 25.800 ;
        RECT 288.030 25.600 1025.270 25.740 ;
        RECT 288.030 25.540 288.350 25.600 ;
        RECT 1024.950 25.540 1025.270 25.600 ;
      LAYER via ;
        RECT 288.060 25.540 288.320 25.800 ;
        RECT 1024.980 25.540 1025.240 25.800 ;
      LAYER met2 ;
        RECT 1025.010 35.000 1025.290 39.000 ;
        RECT 1025.040 25.830 1025.180 35.000 ;
        RECT 288.060 25.510 288.320 25.830 ;
        RECT 1024.980 25.510 1025.240 25.830 ;
        RECT 288.120 2.400 288.260 25.510 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 305.970 15.540 306.290 15.600 ;
        RECT 1073.250 15.540 1073.570 15.600 ;
        RECT 305.970 15.400 1073.570 15.540 ;
        RECT 305.970 15.340 306.290 15.400 ;
        RECT 1073.250 15.340 1073.570 15.400 ;
      LAYER via ;
        RECT 306.000 15.340 306.260 15.600 ;
        RECT 1073.280 15.340 1073.540 15.600 ;
      LAYER met2 ;
        RECT 1073.310 35.000 1073.590 39.000 ;
        RECT 1073.340 15.630 1073.480 35.000 ;
        RECT 306.000 15.310 306.260 15.630 ;
        RECT 1073.280 15.310 1073.540 15.630 ;
        RECT 306.060 2.400 306.200 15.310 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 323.910 22.680 324.230 22.740 ;
        RECT 1121.550 22.680 1121.870 22.740 ;
        RECT 323.910 22.540 1121.870 22.680 ;
        RECT 323.910 22.480 324.230 22.540 ;
        RECT 1121.550 22.480 1121.870 22.540 ;
      LAYER via ;
        RECT 323.940 22.480 324.200 22.740 ;
        RECT 1121.580 22.480 1121.840 22.740 ;
      LAYER met2 ;
        RECT 1121.610 35.000 1121.890 39.000 ;
        RECT 1121.640 22.770 1121.780 35.000 ;
        RECT 323.940 22.450 324.200 22.770 ;
        RECT 1121.580 22.450 1121.840 22.770 ;
        RECT 324.000 2.400 324.140 22.450 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 341.390 15.880 341.710 15.940 ;
        RECT 1169.850 15.880 1170.170 15.940 ;
        RECT 341.390 15.740 1170.170 15.880 ;
        RECT 341.390 15.680 341.710 15.740 ;
        RECT 1169.850 15.680 1170.170 15.740 ;
      LAYER via ;
        RECT 341.420 15.680 341.680 15.940 ;
        RECT 1169.880 15.680 1170.140 15.940 ;
      LAYER met2 ;
        RECT 1169.910 35.000 1170.190 39.000 ;
        RECT 1169.940 15.970 1170.080 35.000 ;
        RECT 341.420 15.650 341.680 15.970 ;
        RECT 1169.880 15.650 1170.140 15.970 ;
        RECT 341.480 2.400 341.620 15.650 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 359.330 23.020 359.650 23.080 ;
        RECT 1218.150 23.020 1218.470 23.080 ;
        RECT 359.330 22.880 1218.470 23.020 ;
        RECT 359.330 22.820 359.650 22.880 ;
        RECT 1218.150 22.820 1218.470 22.880 ;
      LAYER via ;
        RECT 359.360 22.820 359.620 23.080 ;
        RECT 1218.180 22.820 1218.440 23.080 ;
      LAYER met2 ;
        RECT 1218.210 35.000 1218.490 39.000 ;
        RECT 1218.240 23.110 1218.380 35.000 ;
        RECT 359.360 22.790 359.620 23.110 ;
        RECT 1218.180 22.790 1218.440 23.110 ;
        RECT 359.420 2.400 359.560 22.790 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 783.910 21.320 784.230 21.380 ;
        RECT 1266.450 21.320 1266.770 21.380 ;
        RECT 783.910 21.180 1266.770 21.320 ;
        RECT 783.910 21.120 784.230 21.180 ;
        RECT 1266.450 21.120 1266.770 21.180 ;
        RECT 377.270 14.180 377.590 14.240 ;
        RECT 783.910 14.180 784.230 14.240 ;
        RECT 377.270 14.040 784.230 14.180 ;
        RECT 377.270 13.980 377.590 14.040 ;
        RECT 783.910 13.980 784.230 14.040 ;
      LAYER via ;
        RECT 783.940 21.120 784.200 21.380 ;
        RECT 1266.480 21.120 1266.740 21.380 ;
        RECT 377.300 13.980 377.560 14.240 ;
        RECT 783.940 13.980 784.200 14.240 ;
      LAYER met2 ;
        RECT 1266.510 35.000 1266.790 39.000 ;
        RECT 1266.540 21.410 1266.680 35.000 ;
        RECT 783.940 21.090 784.200 21.410 ;
        RECT 1266.480 21.090 1266.740 21.410 ;
        RECT 784.000 14.270 784.140 21.090 ;
        RECT 377.300 13.950 377.560 14.270 ;
        RECT 783.940 13.950 784.200 14.270 ;
        RECT 377.360 2.400 377.500 13.950 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 395.210 23.360 395.530 23.420 ;
        RECT 1314.750 23.360 1315.070 23.420 ;
        RECT 395.210 23.220 1315.070 23.360 ;
        RECT 395.210 23.160 395.530 23.220 ;
        RECT 1314.750 23.160 1315.070 23.220 ;
      LAYER via ;
        RECT 395.240 23.160 395.500 23.420 ;
        RECT 1314.780 23.160 1315.040 23.420 ;
      LAYER met2 ;
        RECT 1314.810 35.000 1315.090 39.000 ;
        RECT 1314.840 23.450 1314.980 35.000 ;
        RECT 395.240 23.130 395.500 23.450 ;
        RECT 1314.780 23.130 1315.040 23.450 ;
        RECT 395.300 2.400 395.440 23.130 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 413.150 16.220 413.470 16.280 ;
        RECT 1363.050 16.220 1363.370 16.280 ;
        RECT 413.150 16.080 1363.370 16.220 ;
        RECT 413.150 16.020 413.470 16.080 ;
        RECT 1363.050 16.020 1363.370 16.080 ;
      LAYER via ;
        RECT 413.180 16.020 413.440 16.280 ;
        RECT 1363.080 16.020 1363.340 16.280 ;
      LAYER met2 ;
        RECT 1363.110 35.000 1363.390 39.000 ;
        RECT 1363.140 16.310 1363.280 35.000 ;
        RECT 413.180 15.990 413.440 16.310 ;
        RECT 1363.080 15.990 1363.340 16.310 ;
        RECT 413.240 2.400 413.380 15.990 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 74.130 19.960 74.450 20.020 ;
        RECT 493.650 19.960 493.970 20.020 ;
        RECT 74.130 19.820 493.970 19.960 ;
        RECT 74.130 19.760 74.450 19.820 ;
        RECT 493.650 19.760 493.970 19.820 ;
      LAYER via ;
        RECT 74.160 19.760 74.420 20.020 ;
        RECT 493.680 19.760 493.940 20.020 ;
      LAYER met2 ;
        RECT 493.710 35.000 493.990 39.000 ;
        RECT 493.740 20.050 493.880 35.000 ;
        RECT 74.160 19.730 74.420 20.050 ;
        RECT 493.680 19.730 493.940 20.050 ;
        RECT 74.220 2.400 74.360 19.730 ;
        RECT 74.010 -4.800 74.570 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 430.630 23.700 430.950 23.760 ;
        RECT 1411.350 23.700 1411.670 23.760 ;
        RECT 430.630 23.560 1411.670 23.700 ;
        RECT 430.630 23.500 430.950 23.560 ;
        RECT 1411.350 23.500 1411.670 23.560 ;
      LAYER via ;
        RECT 430.660 23.500 430.920 23.760 ;
        RECT 1411.380 23.500 1411.640 23.760 ;
      LAYER met2 ;
        RECT 1411.410 35.000 1411.690 39.000 ;
        RECT 1411.440 23.790 1411.580 35.000 ;
        RECT 430.660 23.470 430.920 23.790 ;
        RECT 1411.380 23.470 1411.640 23.790 ;
        RECT 430.720 2.400 430.860 23.470 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 448.570 16.560 448.890 16.620 ;
        RECT 1459.650 16.560 1459.970 16.620 ;
        RECT 448.570 16.420 1459.970 16.560 ;
        RECT 448.570 16.360 448.890 16.420 ;
        RECT 1459.650 16.360 1459.970 16.420 ;
      LAYER via ;
        RECT 448.600 16.360 448.860 16.620 ;
        RECT 1459.680 16.360 1459.940 16.620 ;
      LAYER met2 ;
        RECT 1459.710 35.000 1459.990 39.000 ;
        RECT 1459.740 16.650 1459.880 35.000 ;
        RECT 448.600 16.330 448.860 16.650 ;
        RECT 1459.680 16.330 1459.940 16.650 ;
        RECT 448.660 2.400 448.800 16.330 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 466.510 27.440 466.830 27.500 ;
        RECT 1507.950 27.440 1508.270 27.500 ;
        RECT 466.510 27.300 1508.270 27.440 ;
        RECT 466.510 27.240 466.830 27.300 ;
        RECT 1507.950 27.240 1508.270 27.300 ;
      LAYER via ;
        RECT 466.540 27.240 466.800 27.500 ;
        RECT 1507.980 27.240 1508.240 27.500 ;
      LAYER met2 ;
        RECT 1508.010 35.000 1508.290 39.000 ;
        RECT 1508.040 27.530 1508.180 35.000 ;
        RECT 466.540 27.210 466.800 27.530 ;
        RECT 1507.980 27.210 1508.240 27.530 ;
        RECT 466.600 2.400 466.740 27.210 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 484.450 16.900 484.770 16.960 ;
        RECT 1556.250 16.900 1556.570 16.960 ;
        RECT 484.450 16.760 1556.570 16.900 ;
        RECT 484.450 16.700 484.770 16.760 ;
        RECT 1556.250 16.700 1556.570 16.760 ;
      LAYER via ;
        RECT 484.480 16.700 484.740 16.960 ;
        RECT 1556.280 16.700 1556.540 16.960 ;
      LAYER met2 ;
        RECT 1556.310 35.000 1556.590 39.000 ;
        RECT 1556.340 16.990 1556.480 35.000 ;
        RECT 484.480 16.670 484.740 16.990 ;
        RECT 1556.280 16.670 1556.540 16.990 ;
        RECT 484.540 2.400 484.680 16.670 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 502.390 27.100 502.710 27.160 ;
        RECT 1604.550 27.100 1604.870 27.160 ;
        RECT 502.390 26.960 1604.870 27.100 ;
        RECT 502.390 26.900 502.710 26.960 ;
        RECT 1604.550 26.900 1604.870 26.960 ;
      LAYER via ;
        RECT 502.420 26.900 502.680 27.160 ;
        RECT 1604.580 26.900 1604.840 27.160 ;
      LAYER met2 ;
        RECT 1604.610 35.000 1604.890 39.000 ;
        RECT 1604.640 27.190 1604.780 35.000 ;
        RECT 502.420 26.870 502.680 27.190 ;
        RECT 1604.580 26.870 1604.840 27.190 ;
        RECT 502.480 2.400 502.620 26.870 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 519.870 20.300 520.190 20.360 ;
        RECT 1652.850 20.300 1653.170 20.360 ;
        RECT 519.870 20.160 1653.170 20.300 ;
        RECT 519.870 20.100 520.190 20.160 ;
        RECT 1652.850 20.100 1653.170 20.160 ;
      LAYER via ;
        RECT 519.900 20.100 520.160 20.360 ;
        RECT 1652.880 20.100 1653.140 20.360 ;
      LAYER met2 ;
        RECT 1652.910 35.000 1653.190 39.000 ;
        RECT 1652.940 20.390 1653.080 35.000 ;
        RECT 519.900 20.070 520.160 20.390 ;
        RECT 1652.880 20.070 1653.140 20.390 ;
        RECT 519.960 2.400 520.100 20.070 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 537.810 26.760 538.130 26.820 ;
        RECT 1701.150 26.760 1701.470 26.820 ;
        RECT 537.810 26.620 1701.470 26.760 ;
        RECT 537.810 26.560 538.130 26.620 ;
        RECT 1701.150 26.560 1701.470 26.620 ;
      LAYER via ;
        RECT 537.840 26.560 538.100 26.820 ;
        RECT 1701.180 26.560 1701.440 26.820 ;
      LAYER met2 ;
        RECT 1701.210 35.000 1701.490 39.000 ;
        RECT 1701.240 26.850 1701.380 35.000 ;
        RECT 537.840 26.530 538.100 26.850 ;
        RECT 1701.180 26.530 1701.440 26.850 ;
        RECT 537.900 2.400 538.040 26.530 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 555.750 19.960 556.070 20.020 ;
        RECT 1749.450 19.960 1749.770 20.020 ;
        RECT 555.750 19.820 1749.770 19.960 ;
        RECT 555.750 19.760 556.070 19.820 ;
        RECT 1749.450 19.760 1749.770 19.820 ;
      LAYER via ;
        RECT 555.780 19.760 556.040 20.020 ;
        RECT 1749.480 19.760 1749.740 20.020 ;
      LAYER met2 ;
        RECT 1749.510 35.000 1749.790 39.000 ;
        RECT 1749.540 20.050 1749.680 35.000 ;
        RECT 555.780 19.730 556.040 20.050 ;
        RECT 1749.480 19.730 1749.740 20.050 ;
        RECT 555.840 2.400 555.980 19.730 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 573.690 26.420 574.010 26.480 ;
        RECT 1797.750 26.420 1798.070 26.480 ;
        RECT 573.690 26.280 1798.070 26.420 ;
        RECT 573.690 26.220 574.010 26.280 ;
        RECT 1797.750 26.220 1798.070 26.280 ;
      LAYER via ;
        RECT 573.720 26.220 573.980 26.480 ;
        RECT 1797.780 26.220 1798.040 26.480 ;
      LAYER met2 ;
        RECT 1797.810 35.000 1798.090 39.000 ;
        RECT 1797.840 26.510 1797.980 35.000 ;
        RECT 573.720 26.190 573.980 26.510 ;
        RECT 1797.780 26.190 1798.040 26.510 ;
        RECT 573.780 2.400 573.920 26.190 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 591.170 19.620 591.490 19.680 ;
        RECT 1846.050 19.620 1846.370 19.680 ;
        RECT 591.170 19.480 1846.370 19.620 ;
        RECT 591.170 19.420 591.490 19.480 ;
        RECT 1846.050 19.420 1846.370 19.480 ;
      LAYER via ;
        RECT 591.200 19.420 591.460 19.680 ;
        RECT 1846.080 19.420 1846.340 19.680 ;
      LAYER met2 ;
        RECT 1846.110 35.000 1846.390 39.000 ;
        RECT 1846.140 19.710 1846.280 35.000 ;
        RECT 591.200 19.390 591.460 19.710 ;
        RECT 1846.080 19.390 1846.340 19.710 ;
        RECT 591.260 2.400 591.400 19.390 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 97.590 26.080 97.910 26.140 ;
        RECT 541.950 26.080 542.270 26.140 ;
        RECT 97.590 25.940 542.270 26.080 ;
        RECT 97.590 25.880 97.910 25.940 ;
        RECT 541.950 25.880 542.270 25.940 ;
      LAYER via ;
        RECT 97.620 25.880 97.880 26.140 ;
        RECT 541.980 25.880 542.240 26.140 ;
      LAYER met2 ;
        RECT 542.010 35.000 542.290 39.000 ;
        RECT 542.040 26.170 542.180 35.000 ;
        RECT 97.620 25.850 97.880 26.170 ;
        RECT 541.980 25.850 542.240 26.170 ;
        RECT 97.680 2.400 97.820 25.850 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 609.110 26.080 609.430 26.140 ;
        RECT 1894.350 26.080 1894.670 26.140 ;
        RECT 609.110 25.940 1894.670 26.080 ;
        RECT 609.110 25.880 609.430 25.940 ;
        RECT 1894.350 25.880 1894.670 25.940 ;
      LAYER via ;
        RECT 609.140 25.880 609.400 26.140 ;
        RECT 1894.380 25.880 1894.640 26.140 ;
      LAYER met2 ;
        RECT 1894.410 35.000 1894.690 39.000 ;
        RECT 1894.440 26.170 1894.580 35.000 ;
        RECT 609.140 25.850 609.400 26.170 ;
        RECT 1894.380 25.850 1894.640 26.170 ;
        RECT 609.200 2.400 609.340 25.850 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 627.050 19.280 627.370 19.340 ;
        RECT 1942.650 19.280 1942.970 19.340 ;
        RECT 627.050 19.140 1942.970 19.280 ;
        RECT 627.050 19.080 627.370 19.140 ;
        RECT 1942.650 19.080 1942.970 19.140 ;
      LAYER via ;
        RECT 627.080 19.080 627.340 19.340 ;
        RECT 1942.680 19.080 1942.940 19.340 ;
      LAYER met2 ;
        RECT 1942.710 35.000 1942.990 39.000 ;
        RECT 1942.740 19.370 1942.880 35.000 ;
        RECT 627.080 19.050 627.340 19.370 ;
        RECT 1942.680 19.050 1942.940 19.370 ;
        RECT 627.140 2.400 627.280 19.050 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 24.040 121.830 24.100 ;
        RECT 590.250 24.040 590.570 24.100 ;
        RECT 121.510 23.900 590.570 24.040 ;
        RECT 121.510 23.840 121.830 23.900 ;
        RECT 590.250 23.840 590.570 23.900 ;
      LAYER via ;
        RECT 121.540 23.840 121.800 24.100 ;
        RECT 590.280 23.840 590.540 24.100 ;
      LAYER met2 ;
        RECT 590.310 35.000 590.590 39.000 ;
        RECT 590.340 24.130 590.480 35.000 ;
        RECT 121.540 23.810 121.800 24.130 ;
        RECT 590.280 23.810 590.540 24.130 ;
        RECT 121.600 2.400 121.740 23.810 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 145.430 14.520 145.750 14.580 ;
        RECT 638.550 14.520 638.870 14.580 ;
        RECT 145.430 14.380 638.870 14.520 ;
        RECT 145.430 14.320 145.750 14.380 ;
        RECT 638.550 14.320 638.870 14.380 ;
      LAYER via ;
        RECT 145.460 14.320 145.720 14.580 ;
        RECT 638.580 14.320 638.840 14.580 ;
      LAYER met2 ;
        RECT 638.610 35.000 638.890 39.000 ;
        RECT 638.640 14.610 638.780 35.000 ;
        RECT 145.460 14.290 145.720 14.610 ;
        RECT 638.580 14.290 638.840 14.610 ;
        RECT 145.520 2.400 145.660 14.290 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 163.370 20.980 163.690 21.040 ;
        RECT 686.850 20.980 687.170 21.040 ;
        RECT 163.370 20.840 687.170 20.980 ;
        RECT 163.370 20.780 163.690 20.840 ;
        RECT 686.850 20.780 687.170 20.840 ;
      LAYER via ;
        RECT 163.400 20.780 163.660 21.040 ;
        RECT 686.880 20.780 687.140 21.040 ;
      LAYER met2 ;
        RECT 686.910 35.000 687.190 39.000 ;
        RECT 686.940 21.070 687.080 35.000 ;
        RECT 163.400 20.750 163.660 21.070 ;
        RECT 686.880 20.750 687.140 21.070 ;
        RECT 163.460 2.400 163.600 20.750 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 180.850 14.860 181.170 14.920 ;
        RECT 735.150 14.860 735.470 14.920 ;
        RECT 180.850 14.720 735.470 14.860 ;
        RECT 180.850 14.660 181.170 14.720 ;
        RECT 735.150 14.660 735.470 14.720 ;
      LAYER via ;
        RECT 180.880 14.660 181.140 14.920 ;
        RECT 735.180 14.660 735.440 14.920 ;
      LAYER met2 ;
        RECT 735.210 35.000 735.490 39.000 ;
        RECT 735.240 14.950 735.380 35.000 ;
        RECT 180.880 14.630 181.140 14.950 ;
        RECT 735.180 14.630 735.440 14.950 ;
        RECT 180.940 2.400 181.080 14.630 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 198.790 21.320 199.110 21.380 ;
        RECT 783.450 21.320 783.770 21.380 ;
        RECT 198.790 21.180 783.770 21.320 ;
        RECT 198.790 21.120 199.110 21.180 ;
        RECT 783.450 21.120 783.770 21.180 ;
      LAYER via ;
        RECT 198.820 21.120 199.080 21.380 ;
        RECT 783.480 21.120 783.740 21.380 ;
      LAYER met2 ;
        RECT 783.510 35.000 783.790 39.000 ;
        RECT 783.540 21.410 783.680 35.000 ;
        RECT 198.820 21.090 199.080 21.410 ;
        RECT 783.480 21.090 783.740 21.410 ;
        RECT 198.880 2.400 199.020 21.090 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 216.730 15.200 217.050 15.260 ;
        RECT 831.750 15.200 832.070 15.260 ;
        RECT 216.730 15.060 832.070 15.200 ;
        RECT 216.730 15.000 217.050 15.060 ;
        RECT 831.750 15.000 832.070 15.060 ;
      LAYER via ;
        RECT 216.760 15.000 217.020 15.260 ;
        RECT 831.780 15.000 832.040 15.260 ;
      LAYER met2 ;
        RECT 831.810 35.000 832.090 39.000 ;
        RECT 831.840 15.290 831.980 35.000 ;
        RECT 216.760 14.970 217.020 15.290 ;
        RECT 831.780 14.970 832.040 15.290 ;
        RECT 216.820 2.400 216.960 14.970 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 234.670 21.660 234.990 21.720 ;
        RECT 880.050 21.660 880.370 21.720 ;
        RECT 234.670 21.520 880.370 21.660 ;
        RECT 234.670 21.460 234.990 21.520 ;
        RECT 880.050 21.460 880.370 21.520 ;
      LAYER via ;
        RECT 234.700 21.460 234.960 21.720 ;
        RECT 880.080 21.460 880.340 21.720 ;
      LAYER met2 ;
        RECT 880.110 35.000 880.390 39.000 ;
        RECT 880.140 21.750 880.280 35.000 ;
        RECT 234.700 21.430 234.960 21.750 ;
        RECT 880.080 21.430 880.340 21.750 ;
        RECT 234.760 2.400 234.900 21.430 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 46.990 3443.420 47.310 3443.480 ;
        RECT 2813.430 3443.420 2813.750 3443.480 ;
        RECT 46.990 3443.280 2813.750 3443.420 ;
        RECT 46.990 3443.220 47.310 3443.280 ;
        RECT 2813.430 3443.220 2813.750 3443.280 ;
        RECT 46.990 37.980 47.310 38.040 ;
        RECT 56.190 37.980 56.510 38.040 ;
        RECT 46.990 37.840 56.510 37.980 ;
        RECT 46.990 37.780 47.310 37.840 ;
        RECT 56.190 37.780 56.510 37.840 ;
      LAYER via ;
        RECT 47.020 3443.220 47.280 3443.480 ;
        RECT 2813.460 3443.220 2813.720 3443.480 ;
        RECT 47.020 37.780 47.280 38.040 ;
        RECT 56.220 37.780 56.480 38.040 ;
      LAYER met2 ;
        RECT 47.020 3443.190 47.280 3443.510 ;
        RECT 2813.460 3443.190 2813.720 3443.510 ;
        RECT 47.080 38.070 47.220 3443.190 ;
        RECT 2813.520 3435.000 2813.660 3443.190 ;
        RECT 2813.490 3431.000 2813.770 3435.000 ;
        RECT 47.020 37.750 47.280 38.070 ;
        RECT 56.220 37.750 56.480 38.070 ;
        RECT 56.280 2.400 56.420 37.750 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.130 16.475 80.410 16.845 ;
        RECT 80.200 2.400 80.340 16.475 ;
        RECT 79.990 -4.800 80.550 2.400 ;
      LAYER via2 ;
        RECT 80.130 16.520 80.410 16.800 ;
      LAYER met3 ;
        RECT 2881.000 3381.450 2885.000 3381.920 ;
        RECT 2890.910 3381.450 2891.290 3381.460 ;
        RECT 2881.000 3381.320 2891.290 3381.450 ;
        RECT 2884.510 3381.150 2891.290 3381.320 ;
        RECT 2890.910 3381.140 2891.290 3381.150 ;
        RECT 80.105 16.810 80.435 16.825 ;
        RECT 2890.910 16.810 2891.290 16.820 ;
        RECT 80.105 16.510 2891.290 16.810 ;
        RECT 80.105 16.495 80.435 16.510 ;
        RECT 2890.910 16.500 2891.290 16.510 ;
      LAYER via3 ;
        RECT 2890.940 3381.140 2891.260 3381.460 ;
        RECT 2890.940 16.500 2891.260 16.820 ;
      LAYER met4 ;
        RECT 2890.935 3381.135 2891.265 3381.465 ;
        RECT 2890.950 16.825 2891.250 3381.135 ;
        RECT 2890.935 16.495 2891.265 16.825 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 34.110 14.860 34.430 14.920 ;
        RECT 103.570 14.860 103.890 14.920 ;
        RECT 34.110 14.720 103.890 14.860 ;
        RECT 34.110 14.660 34.430 14.720 ;
        RECT 103.570 14.660 103.890 14.720 ;
      LAYER via ;
        RECT 34.140 14.660 34.400 14.920 ;
        RECT 103.600 14.660 103.860 14.920 ;
      LAYER met2 ;
        RECT 34.130 3278.435 34.410 3278.805 ;
        RECT 34.200 14.950 34.340 3278.435 ;
        RECT 34.140 14.630 34.400 14.950 ;
        RECT 103.600 14.630 103.860 14.950 ;
        RECT 103.660 2.400 103.800 14.630 ;
        RECT 103.450 -4.800 104.010 2.400 ;
      LAYER via2 ;
        RECT 34.130 3278.480 34.410 3278.760 ;
      LAYER met3 ;
        RECT 35.000 3279.320 39.000 3279.920 ;
        RECT 34.105 3278.770 34.435 3278.785 ;
        RECT 35.270 3278.770 35.570 3279.320 ;
        RECT 34.105 3278.470 35.570 3278.770 ;
        RECT 34.105 3278.455 34.435 3278.470 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2812.110 35.000 2812.390 39.000 ;
        RECT 2812.140 24.325 2812.280 35.000 ;
        RECT 127.510 23.955 127.790 24.325 ;
        RECT 2812.070 23.955 2812.350 24.325 ;
        RECT 127.580 2.400 127.720 23.955 ;
        RECT 127.370 -4.800 127.930 2.400 ;
      LAYER via2 ;
        RECT 127.510 24.000 127.790 24.280 ;
        RECT 2812.070 24.000 2812.350 24.280 ;
      LAYER met3 ;
        RECT 127.485 24.290 127.815 24.305 ;
        RECT 2812.045 24.290 2812.375 24.305 ;
        RECT 127.485 23.990 2812.375 24.290 ;
        RECT 127.485 23.975 127.815 23.990 ;
        RECT 2812.045 23.975 2812.375 23.990 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1103.610 25.740 1103.930 25.800 ;
        RECT 2860.350 25.740 2860.670 25.800 ;
        RECT 1103.610 25.600 2860.670 25.740 ;
        RECT 1103.610 25.540 1103.930 25.600 ;
        RECT 2860.350 25.540 2860.670 25.600 ;
        RECT 26.290 20.640 26.610 20.700 ;
        RECT 1103.610 20.640 1103.930 20.700 ;
        RECT 26.290 20.500 1103.930 20.640 ;
        RECT 26.290 20.440 26.610 20.500 ;
        RECT 1103.610 20.440 1103.930 20.500 ;
      LAYER via ;
        RECT 1103.640 25.540 1103.900 25.800 ;
        RECT 2860.380 25.540 2860.640 25.800 ;
        RECT 26.320 20.440 26.580 20.700 ;
        RECT 1103.640 20.440 1103.900 20.700 ;
      LAYER met2 ;
        RECT 2860.410 35.000 2860.690 39.000 ;
        RECT 2860.440 25.830 2860.580 35.000 ;
        RECT 1103.640 25.510 1103.900 25.830 ;
        RECT 2860.380 25.510 2860.640 25.830 ;
        RECT 1103.700 20.730 1103.840 25.510 ;
        RECT 26.320 20.410 26.580 20.730 ;
        RECT 1103.640 20.410 1103.900 20.730 ;
        RECT 26.380 2.400 26.520 20.410 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 27.670 2.960 27.990 3.020 ;
        RECT 32.270 2.960 32.590 3.020 ;
        RECT 27.670 2.820 32.590 2.960 ;
        RECT 27.670 2.760 27.990 2.820 ;
        RECT 32.270 2.760 32.590 2.820 ;
      LAYER via ;
        RECT 27.700 2.760 27.960 3.020 ;
        RECT 32.300 2.760 32.560 3.020 ;
      LAYER met2 ;
        RECT 27.690 3381.795 27.970 3382.165 ;
        RECT 27.760 3.050 27.900 3381.795 ;
        RECT 27.700 2.730 27.960 3.050 ;
        RECT 32.300 2.730 32.560 3.050 ;
        RECT 32.360 2.400 32.500 2.730 ;
        RECT 32.150 -4.800 32.710 2.400 ;
      LAYER via2 ;
        RECT 27.690 3381.840 27.970 3382.120 ;
      LAYER met3 ;
        RECT 35.000 3382.680 39.000 3383.280 ;
        RECT 27.665 3382.130 27.995 3382.145 ;
        RECT 35.270 3382.130 35.570 3382.680 ;
        RECT 27.665 3381.830 35.570 3382.130 ;
        RECT 27.665 3381.815 27.995 3381.830 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.380 -14.020 -16.380 3533.700 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 497.120 -18.720 500.120 3538.400 ;
        RECT 1257.120 -18.720 1260.120 3538.400 ;
        RECT 2017.120 -18.720 2020.120 3538.400 ;
        RECT 2777.120 -18.720 2780.120 3538.400 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
        RECT 2936.000 -14.020 2939.000 3533.700 ;
      LAYER via4 ;
        RECT -18.470 3532.410 -17.290 3533.590 ;
        RECT -18.470 3530.810 -17.290 3531.990 ;
        RECT 498.030 3532.410 499.210 3533.590 ;
        RECT 498.030 3530.810 499.210 3531.990 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 498.030 3523.010 499.210 3524.190 ;
        RECT 498.030 3521.410 499.210 3522.590 ;
        RECT 498.030 -2.910 499.210 -1.730 ;
        RECT 498.030 -4.510 499.210 -3.330 ;
        RECT -18.470 -12.310 -17.290 -11.130 ;
        RECT -18.470 -13.910 -17.290 -12.730 ;
        RECT 498.030 -12.310 499.210 -11.130 ;
        RECT 498.030 -13.910 499.210 -12.730 ;
        RECT 1258.030 3532.410 1259.210 3533.590 ;
        RECT 1258.030 3530.810 1259.210 3531.990 ;
        RECT 1258.030 3523.010 1259.210 3524.190 ;
        RECT 1258.030 3521.410 1259.210 3522.590 ;
        RECT 1258.030 -2.910 1259.210 -1.730 ;
        RECT 1258.030 -4.510 1259.210 -3.330 ;
        RECT 1258.030 -12.310 1259.210 -11.130 ;
        RECT 1258.030 -13.910 1259.210 -12.730 ;
        RECT 2018.030 3532.410 2019.210 3533.590 ;
        RECT 2018.030 3530.810 2019.210 3531.990 ;
        RECT 2018.030 3523.010 2019.210 3524.190 ;
        RECT 2018.030 3521.410 2019.210 3522.590 ;
        RECT 2018.030 -2.910 2019.210 -1.730 ;
        RECT 2018.030 -4.510 2019.210 -3.330 ;
        RECT 2018.030 -12.310 2019.210 -11.130 ;
        RECT 2018.030 -13.910 2019.210 -12.730 ;
        RECT 2778.030 3532.410 2779.210 3533.590 ;
        RECT 2778.030 3530.810 2779.210 3531.990 ;
        RECT 2936.910 3532.410 2938.090 3533.590 ;
        RECT 2936.910 3530.810 2938.090 3531.990 ;
        RECT 2778.030 3523.010 2779.210 3524.190 ;
        RECT 2778.030 3521.410 2779.210 3522.590 ;
        RECT 2778.030 -2.910 2779.210 -1.730 ;
        RECT 2778.030 -4.510 2779.210 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
        RECT 2778.030 -12.310 2779.210 -11.130 ;
        RECT 2778.030 -13.910 2779.210 -12.730 ;
        RECT 2936.910 -12.310 2938.090 -11.130 ;
        RECT 2936.910 -13.910 2938.090 -12.730 ;
      LAYER met5 ;
        RECT -19.380 3533.700 -16.380 3533.710 ;
        RECT 497.120 3533.700 500.120 3533.710 ;
        RECT 1257.120 3533.700 1260.120 3533.710 ;
        RECT 2017.120 3533.700 2020.120 3533.710 ;
        RECT 2777.120 3533.700 2780.120 3533.710 ;
        RECT 2936.000 3533.700 2939.000 3533.710 ;
        RECT -19.380 3530.700 2939.000 3533.700 ;
        RECT -19.380 3530.690 -16.380 3530.700 ;
        RECT 497.120 3530.690 500.120 3530.700 ;
        RECT 1257.120 3530.690 1260.120 3530.700 ;
        RECT 2017.120 3530.690 2020.120 3530.700 ;
        RECT 2777.120 3530.690 2780.120 3530.700 ;
        RECT 2936.000 3530.690 2939.000 3530.700 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 497.120 3524.300 500.120 3524.310 ;
        RECT 1257.120 3524.300 1260.120 3524.310 ;
        RECT 2017.120 3524.300 2020.120 3524.310 ;
        RECT 2777.120 3524.300 2780.120 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 497.120 3521.290 500.120 3521.300 ;
        RECT 1257.120 3521.290 1260.120 3521.300 ;
        RECT 2017.120 3521.290 2020.120 3521.300 ;
        RECT 2777.120 3521.290 2780.120 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 497.120 -1.620 500.120 -1.610 ;
        RECT 1257.120 -1.620 1260.120 -1.610 ;
        RECT 2017.120 -1.620 2020.120 -1.610 ;
        RECT 2777.120 -1.620 2780.120 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 497.120 -4.630 500.120 -4.620 ;
        RECT 1257.120 -4.630 1260.120 -4.620 ;
        RECT 2017.120 -4.630 2020.120 -4.620 ;
        RECT 2777.120 -4.630 2780.120 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
        RECT -19.380 -11.020 -16.380 -11.010 ;
        RECT 497.120 -11.020 500.120 -11.010 ;
        RECT 1257.120 -11.020 1260.120 -11.010 ;
        RECT 2017.120 -11.020 2020.120 -11.010 ;
        RECT 2777.120 -11.020 2780.120 -11.010 ;
        RECT 2936.000 -11.020 2939.000 -11.010 ;
        RECT -19.380 -14.020 2939.000 -11.020 ;
        RECT -19.380 -14.030 -16.380 -14.020 ;
        RECT 497.120 -14.030 500.120 -14.020 ;
        RECT 1257.120 -14.030 1260.120 -14.020 ;
        RECT 2017.120 -14.030 2020.120 -14.020 ;
        RECT 2777.120 -14.030 2780.120 -14.020 ;
        RECT 2936.000 -14.030 2939.000 -14.020 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -24.080 -18.720 -21.080 3538.400 ;
        RECT -14.680 -9.320 -11.680 3529.000 ;
        RECT 117.120 -18.720 120.120 3538.400 ;
        RECT 877.120 -18.720 880.120 3538.400 ;
        RECT 1637.120 -18.720 1640.120 3538.400 ;
        RECT 2397.120 -18.720 2400.120 3538.400 ;
        RECT 2931.300 -9.320 2934.300 3529.000 ;
        RECT 2940.700 -18.720 2943.700 3538.400 ;
      LAYER via4 ;
        RECT -23.170 3537.110 -21.990 3538.290 ;
        RECT -23.170 3535.510 -21.990 3536.690 ;
        RECT 118.030 3537.110 119.210 3538.290 ;
        RECT 118.030 3535.510 119.210 3536.690 ;
        RECT -13.770 3527.710 -12.590 3528.890 ;
        RECT -13.770 3526.110 -12.590 3527.290 ;
        RECT -13.770 -7.610 -12.590 -6.430 ;
        RECT -13.770 -9.210 -12.590 -8.030 ;
        RECT 118.030 3527.710 119.210 3528.890 ;
        RECT 118.030 3526.110 119.210 3527.290 ;
        RECT 118.030 -7.610 119.210 -6.430 ;
        RECT 118.030 -9.210 119.210 -8.030 ;
        RECT -23.170 -17.010 -21.990 -15.830 ;
        RECT -23.170 -18.610 -21.990 -17.430 ;
        RECT 118.030 -17.010 119.210 -15.830 ;
        RECT 118.030 -18.610 119.210 -17.430 ;
        RECT 878.030 3537.110 879.210 3538.290 ;
        RECT 878.030 3535.510 879.210 3536.690 ;
        RECT 878.030 3527.710 879.210 3528.890 ;
        RECT 878.030 3526.110 879.210 3527.290 ;
        RECT 878.030 -7.610 879.210 -6.430 ;
        RECT 878.030 -9.210 879.210 -8.030 ;
        RECT 878.030 -17.010 879.210 -15.830 ;
        RECT 878.030 -18.610 879.210 -17.430 ;
        RECT 1638.030 3537.110 1639.210 3538.290 ;
        RECT 1638.030 3535.510 1639.210 3536.690 ;
        RECT 1638.030 3527.710 1639.210 3528.890 ;
        RECT 1638.030 3526.110 1639.210 3527.290 ;
        RECT 1638.030 -7.610 1639.210 -6.430 ;
        RECT 1638.030 -9.210 1639.210 -8.030 ;
        RECT 1638.030 -17.010 1639.210 -15.830 ;
        RECT 1638.030 -18.610 1639.210 -17.430 ;
        RECT 2398.030 3537.110 2399.210 3538.290 ;
        RECT 2398.030 3535.510 2399.210 3536.690 ;
        RECT 2941.610 3537.110 2942.790 3538.290 ;
        RECT 2941.610 3535.510 2942.790 3536.690 ;
        RECT 2398.030 3527.710 2399.210 3528.890 ;
        RECT 2398.030 3526.110 2399.210 3527.290 ;
        RECT 2398.030 -7.610 2399.210 -6.430 ;
        RECT 2398.030 -9.210 2399.210 -8.030 ;
        RECT 2932.210 3527.710 2933.390 3528.890 ;
        RECT 2932.210 3526.110 2933.390 3527.290 ;
        RECT 2932.210 -7.610 2933.390 -6.430 ;
        RECT 2932.210 -9.210 2933.390 -8.030 ;
        RECT 2398.030 -17.010 2399.210 -15.830 ;
        RECT 2398.030 -18.610 2399.210 -17.430 ;
        RECT 2941.610 -17.010 2942.790 -15.830 ;
        RECT 2941.610 -18.610 2942.790 -17.430 ;
      LAYER met5 ;
        RECT -24.080 3538.400 -21.080 3538.410 ;
        RECT 117.120 3538.400 120.120 3538.410 ;
        RECT 877.120 3538.400 880.120 3538.410 ;
        RECT 1637.120 3538.400 1640.120 3538.410 ;
        RECT 2397.120 3538.400 2400.120 3538.410 ;
        RECT 2940.700 3538.400 2943.700 3538.410 ;
        RECT -24.080 3535.400 2943.700 3538.400 ;
        RECT -24.080 3535.390 -21.080 3535.400 ;
        RECT 117.120 3535.390 120.120 3535.400 ;
        RECT 877.120 3535.390 880.120 3535.400 ;
        RECT 1637.120 3535.390 1640.120 3535.400 ;
        RECT 2397.120 3535.390 2400.120 3535.400 ;
        RECT 2940.700 3535.390 2943.700 3535.400 ;
        RECT -14.680 3529.000 -11.680 3529.010 ;
        RECT 117.120 3529.000 120.120 3529.010 ;
        RECT 877.120 3529.000 880.120 3529.010 ;
        RECT 1637.120 3529.000 1640.120 3529.010 ;
        RECT 2397.120 3529.000 2400.120 3529.010 ;
        RECT 2931.300 3529.000 2934.300 3529.010 ;
        RECT -14.680 3526.000 2934.300 3529.000 ;
        RECT -14.680 3525.990 -11.680 3526.000 ;
        RECT 117.120 3525.990 120.120 3526.000 ;
        RECT 877.120 3525.990 880.120 3526.000 ;
        RECT 1637.120 3525.990 1640.120 3526.000 ;
        RECT 2397.120 3525.990 2400.120 3526.000 ;
        RECT 2931.300 3525.990 2934.300 3526.000 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 117.120 -6.320 120.120 -6.310 ;
        RECT 877.120 -6.320 880.120 -6.310 ;
        RECT 1637.120 -6.320 1640.120 -6.310 ;
        RECT 2397.120 -6.320 2400.120 -6.310 ;
        RECT 2931.300 -6.320 2934.300 -6.310 ;
        RECT -14.680 -9.320 2934.300 -6.320 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 117.120 -9.330 120.120 -9.320 ;
        RECT 877.120 -9.330 880.120 -9.320 ;
        RECT 1637.120 -9.330 1640.120 -9.320 ;
        RECT 2397.120 -9.330 2400.120 -9.320 ;
        RECT 2931.300 -9.330 2934.300 -9.320 ;
        RECT -24.080 -15.720 -21.080 -15.710 ;
        RECT 117.120 -15.720 120.120 -15.710 ;
        RECT 877.120 -15.720 880.120 -15.710 ;
        RECT 1637.120 -15.720 1640.120 -15.710 ;
        RECT 2397.120 -15.720 2400.120 -15.710 ;
        RECT 2940.700 -15.720 2943.700 -15.710 ;
        RECT -24.080 -18.720 2943.700 -15.720 ;
        RECT -24.080 -18.730 -21.080 -18.720 ;
        RECT 117.120 -18.730 120.120 -18.720 ;
        RECT 877.120 -18.730 880.120 -18.720 ;
        RECT 1637.120 -18.730 1640.120 -18.720 ;
        RECT 2397.120 -18.730 2400.120 -18.720 ;
        RECT 2940.700 -18.730 2943.700 -18.720 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 40.520 45.795 2879.180 3424.205 ;
      LAYER met1 ;
        RECT 40.520 45.640 2879.180 3424.360 ;
      LAYER met2 ;
        RECT 48.780 3430.720 105.650 3431.000 ;
        RECT 106.490 3430.720 247.790 3431.000 ;
        RECT 248.630 3430.720 390.390 3431.000 ;
        RECT 391.230 3430.720 532.990 3431.000 ;
        RECT 533.830 3430.720 675.590 3431.000 ;
        RECT 676.430 3430.720 818.190 3431.000 ;
        RECT 819.030 3430.720 960.330 3431.000 ;
        RECT 961.170 3430.720 1102.930 3431.000 ;
        RECT 1103.770 3430.720 1245.530 3431.000 ;
        RECT 1246.370 3430.720 1388.130 3431.000 ;
        RECT 1388.970 3430.720 1530.730 3431.000 ;
        RECT 1531.570 3430.720 1672.870 3431.000 ;
        RECT 1673.710 3430.720 1815.470 3431.000 ;
        RECT 1816.310 3430.720 1958.070 3431.000 ;
        RECT 1958.910 3430.720 2100.670 3431.000 ;
        RECT 2101.510 3430.720 2243.270 3431.000 ;
        RECT 2244.110 3430.720 2385.410 3431.000 ;
        RECT 2386.250 3430.720 2528.010 3431.000 ;
        RECT 2528.850 3430.720 2670.610 3431.000 ;
        RECT 2671.450 3430.720 2813.210 3431.000 ;
        RECT 2814.050 3430.720 2870.810 3431.000 ;
        RECT 48.780 39.280 2870.810 3430.720 ;
        RECT 48.780 39.000 58.730 39.280 ;
        RECT 59.570 39.000 107.030 39.280 ;
        RECT 107.870 39.000 155.330 39.280 ;
        RECT 156.170 39.000 203.630 39.280 ;
        RECT 204.470 39.000 251.930 39.280 ;
        RECT 252.770 39.000 300.230 39.280 ;
        RECT 301.070 39.000 348.530 39.280 ;
        RECT 349.370 39.000 396.830 39.280 ;
        RECT 397.670 39.000 445.130 39.280 ;
        RECT 445.970 39.000 493.430 39.280 ;
        RECT 494.270 39.000 541.730 39.280 ;
        RECT 542.570 39.000 590.030 39.280 ;
        RECT 590.870 39.000 638.330 39.280 ;
        RECT 639.170 39.000 686.630 39.280 ;
        RECT 687.470 39.000 734.930 39.280 ;
        RECT 735.770 39.000 783.230 39.280 ;
        RECT 784.070 39.000 831.530 39.280 ;
        RECT 832.370 39.000 879.830 39.280 ;
        RECT 880.670 39.000 928.130 39.280 ;
        RECT 928.970 39.000 976.430 39.280 ;
        RECT 977.270 39.000 1024.730 39.280 ;
        RECT 1025.570 39.000 1073.030 39.280 ;
        RECT 1073.870 39.000 1121.330 39.280 ;
        RECT 1122.170 39.000 1169.630 39.280 ;
        RECT 1170.470 39.000 1217.930 39.280 ;
        RECT 1218.770 39.000 1266.230 39.280 ;
        RECT 1267.070 39.000 1314.530 39.280 ;
        RECT 1315.370 39.000 1362.830 39.280 ;
        RECT 1363.670 39.000 1411.130 39.280 ;
        RECT 1411.970 39.000 1459.430 39.280 ;
        RECT 1460.270 39.000 1507.730 39.280 ;
        RECT 1508.570 39.000 1556.030 39.280 ;
        RECT 1556.870 39.000 1604.330 39.280 ;
        RECT 1605.170 39.000 1652.630 39.280 ;
        RECT 1653.470 39.000 1700.930 39.280 ;
        RECT 1701.770 39.000 1749.230 39.280 ;
        RECT 1750.070 39.000 1797.530 39.280 ;
        RECT 1798.370 39.000 1845.830 39.280 ;
        RECT 1846.670 39.000 1894.130 39.280 ;
        RECT 1894.970 39.000 1942.430 39.280 ;
        RECT 1943.270 39.000 1990.730 39.280 ;
        RECT 1991.570 39.000 2039.030 39.280 ;
        RECT 2039.870 39.000 2087.330 39.280 ;
        RECT 2088.170 39.000 2135.630 39.280 ;
        RECT 2136.470 39.000 2183.930 39.280 ;
        RECT 2184.770 39.000 2232.230 39.280 ;
        RECT 2233.070 39.000 2280.530 39.280 ;
        RECT 2281.370 39.000 2328.830 39.280 ;
        RECT 2329.670 39.000 2377.130 39.280 ;
        RECT 2377.970 39.000 2425.430 39.280 ;
        RECT 2426.270 39.000 2473.730 39.280 ;
        RECT 2474.570 39.000 2522.030 39.280 ;
        RECT 2522.870 39.000 2570.330 39.280 ;
        RECT 2571.170 39.000 2618.630 39.280 ;
        RECT 2619.470 39.000 2666.930 39.280 ;
        RECT 2667.770 39.000 2715.230 39.280 ;
        RECT 2716.070 39.000 2763.530 39.280 ;
        RECT 2764.370 39.000 2811.830 39.280 ;
        RECT 2812.670 39.000 2860.130 39.280 ;
        RECT 2860.970 39.000 2870.810 39.280 ;
      LAYER met3 ;
        RECT 39.000 3383.680 2881.000 3424.285 ;
        RECT 39.400 3382.320 2881.000 3383.680 ;
        RECT 39.400 3382.280 2880.600 3382.320 ;
        RECT 39.000 3380.920 2880.600 3382.280 ;
        RECT 39.000 3280.320 2881.000 3380.920 ;
        RECT 39.400 3278.920 2881.000 3280.320 ;
        RECT 39.000 3276.240 2881.000 3278.920 ;
        RECT 39.000 3274.840 2880.600 3276.240 ;
        RECT 39.000 3177.640 2881.000 3274.840 ;
        RECT 39.400 3176.240 2881.000 3177.640 ;
        RECT 39.000 3170.160 2881.000 3176.240 ;
        RECT 39.000 3168.760 2880.600 3170.160 ;
        RECT 39.000 3074.280 2881.000 3168.760 ;
        RECT 39.400 3072.880 2881.000 3074.280 ;
        RECT 39.000 3064.080 2881.000 3072.880 ;
        RECT 39.000 3062.680 2880.600 3064.080 ;
        RECT 39.000 2971.600 2881.000 3062.680 ;
        RECT 39.400 2970.200 2881.000 2971.600 ;
        RECT 39.000 2957.320 2881.000 2970.200 ;
        RECT 39.000 2955.920 2880.600 2957.320 ;
        RECT 39.000 2868.240 2881.000 2955.920 ;
        RECT 39.400 2866.840 2881.000 2868.240 ;
        RECT 39.000 2851.240 2881.000 2866.840 ;
        RECT 39.000 2849.840 2880.600 2851.240 ;
        RECT 39.000 2765.560 2881.000 2849.840 ;
        RECT 39.400 2764.160 2881.000 2765.560 ;
        RECT 39.000 2745.160 2881.000 2764.160 ;
        RECT 39.000 2743.760 2880.600 2745.160 ;
        RECT 39.000 2662.200 2881.000 2743.760 ;
        RECT 39.400 2660.800 2881.000 2662.200 ;
        RECT 39.000 2639.080 2881.000 2660.800 ;
        RECT 39.000 2637.680 2880.600 2639.080 ;
        RECT 39.000 2559.520 2881.000 2637.680 ;
        RECT 39.400 2558.120 2881.000 2559.520 ;
        RECT 39.000 2532.320 2881.000 2558.120 ;
        RECT 39.000 2530.920 2880.600 2532.320 ;
        RECT 39.000 2456.160 2881.000 2530.920 ;
        RECT 39.400 2454.760 2881.000 2456.160 ;
        RECT 39.000 2426.240 2881.000 2454.760 ;
        RECT 39.000 2424.840 2880.600 2426.240 ;
        RECT 39.000 2353.480 2881.000 2424.840 ;
        RECT 39.400 2352.080 2881.000 2353.480 ;
        RECT 39.000 2320.160 2881.000 2352.080 ;
        RECT 39.000 2318.760 2880.600 2320.160 ;
        RECT 39.000 2250.120 2881.000 2318.760 ;
        RECT 39.400 2248.720 2881.000 2250.120 ;
        RECT 39.000 2214.080 2881.000 2248.720 ;
        RECT 39.000 2212.680 2880.600 2214.080 ;
        RECT 39.000 2147.440 2881.000 2212.680 ;
        RECT 39.400 2146.040 2881.000 2147.440 ;
        RECT 39.000 2107.320 2881.000 2146.040 ;
        RECT 39.000 2105.920 2880.600 2107.320 ;
        RECT 39.000 2044.080 2881.000 2105.920 ;
        RECT 39.400 2042.680 2881.000 2044.080 ;
        RECT 39.000 2001.240 2881.000 2042.680 ;
        RECT 39.000 1999.840 2880.600 2001.240 ;
        RECT 39.000 1941.400 2881.000 1999.840 ;
        RECT 39.400 1940.000 2881.000 1941.400 ;
        RECT 39.000 1895.160 2881.000 1940.000 ;
        RECT 39.000 1893.760 2880.600 1895.160 ;
        RECT 39.000 1838.040 2881.000 1893.760 ;
        RECT 39.400 1836.640 2881.000 1838.040 ;
        RECT 39.000 1789.080 2881.000 1836.640 ;
        RECT 39.000 1787.680 2880.600 1789.080 ;
        RECT 39.000 1735.360 2881.000 1787.680 ;
        RECT 39.400 1733.960 2881.000 1735.360 ;
        RECT 39.000 1682.320 2881.000 1733.960 ;
        RECT 39.000 1680.920 2880.600 1682.320 ;
        RECT 39.000 1632.000 2881.000 1680.920 ;
        RECT 39.400 1630.600 2881.000 1632.000 ;
        RECT 39.000 1576.240 2881.000 1630.600 ;
        RECT 39.000 1574.840 2880.600 1576.240 ;
        RECT 39.000 1529.320 2881.000 1574.840 ;
        RECT 39.400 1527.920 2881.000 1529.320 ;
        RECT 39.000 1470.160 2881.000 1527.920 ;
        RECT 39.000 1468.760 2880.600 1470.160 ;
        RECT 39.000 1425.960 2881.000 1468.760 ;
        RECT 39.400 1424.560 2881.000 1425.960 ;
        RECT 39.000 1364.080 2881.000 1424.560 ;
        RECT 39.000 1362.680 2880.600 1364.080 ;
        RECT 39.000 1323.280 2881.000 1362.680 ;
        RECT 39.400 1321.880 2881.000 1323.280 ;
        RECT 39.000 1257.320 2881.000 1321.880 ;
        RECT 39.000 1255.920 2880.600 1257.320 ;
        RECT 39.000 1219.920 2881.000 1255.920 ;
        RECT 39.400 1218.520 2881.000 1219.920 ;
        RECT 39.000 1151.240 2881.000 1218.520 ;
        RECT 39.000 1149.840 2880.600 1151.240 ;
        RECT 39.000 1117.240 2881.000 1149.840 ;
        RECT 39.400 1115.840 2881.000 1117.240 ;
        RECT 39.000 1045.160 2881.000 1115.840 ;
        RECT 39.000 1043.760 2880.600 1045.160 ;
        RECT 39.000 1013.880 2881.000 1043.760 ;
        RECT 39.400 1012.480 2881.000 1013.880 ;
        RECT 39.000 939.080 2881.000 1012.480 ;
        RECT 39.000 937.680 2880.600 939.080 ;
        RECT 39.000 911.200 2881.000 937.680 ;
        RECT 39.400 909.800 2881.000 911.200 ;
        RECT 39.000 832.320 2881.000 909.800 ;
        RECT 39.000 830.920 2880.600 832.320 ;
        RECT 39.000 807.840 2881.000 830.920 ;
        RECT 39.400 806.440 2881.000 807.840 ;
        RECT 39.000 726.240 2881.000 806.440 ;
        RECT 39.000 724.840 2880.600 726.240 ;
        RECT 39.000 705.160 2881.000 724.840 ;
        RECT 39.400 703.760 2881.000 705.160 ;
        RECT 39.000 620.160 2881.000 703.760 ;
        RECT 39.000 618.760 2880.600 620.160 ;
        RECT 39.000 601.800 2881.000 618.760 ;
        RECT 39.400 600.400 2881.000 601.800 ;
        RECT 39.000 514.080 2881.000 600.400 ;
        RECT 39.000 512.680 2880.600 514.080 ;
        RECT 39.000 499.120 2881.000 512.680 ;
        RECT 39.400 497.720 2881.000 499.120 ;
        RECT 39.000 407.320 2881.000 497.720 ;
        RECT 39.000 405.920 2880.600 407.320 ;
        RECT 39.000 395.760 2881.000 405.920 ;
        RECT 39.400 394.360 2881.000 395.760 ;
        RECT 39.000 301.240 2881.000 394.360 ;
        RECT 39.000 299.840 2880.600 301.240 ;
        RECT 39.000 293.080 2881.000 299.840 ;
        RECT 39.400 291.680 2881.000 293.080 ;
        RECT 39.000 195.160 2881.000 291.680 ;
        RECT 39.000 193.760 2880.600 195.160 ;
        RECT 39.000 189.720 2881.000 193.760 ;
        RECT 39.400 188.320 2881.000 189.720 ;
        RECT 39.000 89.080 2881.000 188.320 ;
        RECT 39.000 87.680 2880.600 89.080 ;
        RECT 39.000 87.040 2881.000 87.680 ;
        RECT 39.400 85.640 2881.000 87.040 ;
        RECT 39.000 45.715 2881.000 85.640 ;
      LAYER met4 ;
        RECT 48.720 45.640 117.120 3424.360 ;
        RECT 120.120 45.640 497.120 3424.360 ;
        RECT 500.120 45.640 877.120 3424.360 ;
        RECT 880.120 45.640 1257.120 3424.360 ;
        RECT 1260.120 45.640 1637.120 3424.360 ;
        RECT 1640.120 45.640 2017.120 3424.360 ;
        RECT 2020.120 45.640 2397.120 3424.360 ;
        RECT 2400.120 45.640 2777.120 3424.360 ;
        RECT 2780.120 45.640 2848.505 3424.360 ;
      LAYER met5 ;
        RECT 40.520 138.080 2879.180 3394.755 ;
      LAYER met5 ;
        RECT 40.520 99.785 2879.180 101.385 ;
        RECT 40.520 61.490 2879.180 63.090 ;
  END
END user_project_wrapper
END LIBRARY


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga
  CLASS BLOCK ;
  FOREIGN fpga ;
  ORIGIN 0.000 0.000 ;
  SIZE 2850.000 BY 3400.000 ;
  PIN gpio_east[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 53.080 2850.000 53.680 ;
    END
  END gpio_east[0]
  PIN gpio_east[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 159.160 2850.000 159.760 ;
    END
  END gpio_east[1]
  PIN gpio_east[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 265.240 2850.000 265.840 ;
    END
  END gpio_east[2]
  PIN gpio_east[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 371.320 2850.000 371.920 ;
    END
  END gpio_east[3]
  PIN gpio_east[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 478.080 2850.000 478.680 ;
    END
  END gpio_east[4]
  PIN gpio_east[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 584.160 2850.000 584.760 ;
    END
  END gpio_east[5]
  PIN gpio_east[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 690.240 2850.000 690.840 ;
    END
  END gpio_east[6]
  PIN gpio_east[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 796.320 2850.000 796.920 ;
    END
  END gpio_east[7]
  PIN gpio_east[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 903.080 2850.000 903.680 ;
    END
  END gpio_east[8]
  PIN gpio_east[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1009.160 2850.000 1009.760 ;
    END
  END gpio_east[9]
  PIN gpio_north[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 59.430 3396.000 59.710 3400.000 ;
    END
  END gpio_north[0]
  PIN gpio_north[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 178.110 3396.000 178.390 3400.000 ;
    END
  END gpio_north[1]
  PIN gpio_north[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 296.790 3396.000 297.070 3400.000 ;
    END
  END gpio_north[2]
  PIN gpio_north[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 415.470 3396.000 415.750 3400.000 ;
    END
  END gpio_north[3]
  PIN gpio_north[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 534.150 3396.000 534.430 3400.000 ;
    END
  END gpio_north[4]
  PIN gpio_north[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 652.830 3396.000 653.110 3400.000 ;
    END
  END gpio_north[5]
  PIN gpio_north[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 771.970 3396.000 772.250 3400.000 ;
    END
  END gpio_north[6]
  PIN gpio_north[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 890.650 3396.000 890.930 3400.000 ;
    END
  END gpio_north[7]
  PIN gpio_north[8]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1009.330 3396.000 1009.610 3400.000 ;
    END
  END gpio_north[8]
  PIN gpio_north[9]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1128.010 3396.000 1128.290 3400.000 ;
    END
  END gpio_north[9]
  PIN gpio_south[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END gpio_south[0]
  PIN gpio_south[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END gpio_south[1]
  PIN gpio_south[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 4.000 ;
    END
  END gpio_south[2]
  PIN gpio_south[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 4.000 ;
    END
  END gpio_south[3]
  PIN gpio_south[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END gpio_south[4]
  PIN gpio_south[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 256.310 0.000 256.590 4.000 ;
    END
  END gpio_south[5]
  PIN gpio_south[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 303.230 0.000 303.510 4.000 ;
    END
  END gpio_south[6]
  PIN gpio_south[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 350.150 0.000 350.430 4.000 ;
    END
  END gpio_south[7]
  PIN gpio_west[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END gpio_west[0]
  PIN gpio_west[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 188.400 4.000 189.000 ;
    END
  END gpio_west[1]
  PIN gpio_west[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.200 4.000 314.800 ;
    END
  END gpio_west[2]
  PIN gpio_west[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.000 4.000 440.600 ;
    END
  END gpio_west[3]
  PIN gpio_west[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 565.800 4.000 566.400 ;
    END
  END gpio_west[4]
  PIN gpio_west[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 691.600 4.000 692.200 ;
    END
  END gpio_west[5]
  PIN gpio_west[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 818.080 4.000 818.680 ;
    END
  END gpio_west[6]
  PIN gpio_west[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 943.880 4.000 944.480 ;
    END
  END gpio_west[7]
  PIN gpio_west[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1069.680 4.000 1070.280 ;
    END
  END gpio_west[8]
  PIN gpio_west[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1195.480 4.000 1196.080 ;
    END
  END gpio_west[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1891.610 0.000 1891.890 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1321.280 4.000 1321.880 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1115.240 2850.000 1115.840 ;
    END
  END wbs_ack_o
  PIN wbs_addr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1246.690 3396.000 1246.970 3400.000 ;
    END
  END wbs_addr_i[0]
  PIN wbs_addr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1985.450 0.000 1985.730 4.000 ;
    END
  END wbs_addr_i[10]
  PIN wbs_addr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2031.910 0.000 2032.190 4.000 ;
    END
  END wbs_addr_i[11]
  PIN wbs_addr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1699.360 4.000 1699.960 ;
    END
  END wbs_addr_i[12]
  PIN wbs_addr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1825.160 4.000 1825.760 ;
    END
  END wbs_addr_i[13]
  PIN wbs_addr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2078.830 0.000 2079.110 4.000 ;
    END
  END wbs_addr_i[14]
  PIN wbs_addr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2125.290 0.000 2125.570 4.000 ;
    END
  END wbs_addr_i[15]
  PIN wbs_addr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1950.960 4.000 1951.560 ;
    END
  END wbs_addr_i[16]
  PIN wbs_addr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2076.760 4.000 2077.360 ;
    END
  END wbs_addr_i[17]
  PIN wbs_addr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2203.240 4.000 2203.840 ;
    END
  END wbs_addr_i[18]
  PIN wbs_addr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1646.320 2850.000 1646.920 ;
    END
  END wbs_addr_i[19]
  PIN wbs_addr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1447.760 4.000 1448.360 ;
    END
  END wbs_addr_i[1]
  PIN wbs_addr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1753.080 2850.000 1753.680 ;
    END
  END wbs_addr_i[20]
  PIN wbs_addr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2172.210 0.000 2172.490 4.000 ;
    END
  END wbs_addr_i[21]
  PIN wbs_addr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2218.670 0.000 2218.950 4.000 ;
    END
  END wbs_addr_i[22]
  PIN wbs_addr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1859.160 2850.000 1859.760 ;
    END
  END wbs_addr_i[23]
  PIN wbs_addr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1603.190 3396.000 1603.470 3400.000 ;
    END
  END wbs_addr_i[24]
  PIN wbs_addr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1965.240 2850.000 1965.840 ;
    END
  END wbs_addr_i[25]
  PIN wbs_addr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2265.590 0.000 2265.870 4.000 ;
    END
  END wbs_addr_i[26]
  PIN wbs_addr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1721.870 3396.000 1722.150 3400.000 ;
    END
  END wbs_addr_i[27]
  PIN wbs_addr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2071.320 2850.000 2071.920 ;
    END
  END wbs_addr_i[28]
  PIN wbs_addr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2178.080 2850.000 2178.680 ;
    END
  END wbs_addr_i[29]
  PIN wbs_addr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1221.320 2850.000 1221.920 ;
    END
  END wbs_addr_i[2]
  PIN wbs_addr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2284.160 2850.000 2284.760 ;
    END
  END wbs_addr_i[30]
  PIN wbs_addr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1840.550 3396.000 1840.830 3400.000 ;
    END
  END wbs_addr_i[31]
  PIN wbs_addr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1573.560 4.000 1574.160 ;
    END
  END wbs_addr_i[3]
  PIN wbs_addr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1328.080 2850.000 1328.680 ;
    END
  END wbs_addr_i[4]
  PIN wbs_addr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1938.530 0.000 1938.810 4.000 ;
    END
  END wbs_addr_i[5]
  PIN wbs_addr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1434.160 2850.000 1434.760 ;
    END
  END wbs_addr_i[6]
  PIN wbs_addr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 1540.240 2850.000 1540.840 ;
    END
  END wbs_addr_i[7]
  PIN wbs_addr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1365.370 3396.000 1365.650 3400.000 ;
    END
  END wbs_addr_i[8]
  PIN wbs_addr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1484.510 3396.000 1484.790 3400.000 ;
    END
  END wbs_addr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2329.040 4.000 2329.640 ;
    END
  END wbs_cyc_i
  PIN wbs_data_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1959.230 3396.000 1959.510 3400.000 ;
    END
  END wbs_data_i[0]
  PIN wbs_data_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2921.320 2850.000 2921.920 ;
    END
  END wbs_data_i[10]
  PIN wbs_data_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2454.840 4.000 2455.440 ;
    END
  END wbs_data_i[11]
  PIN wbs_data_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2315.730 3396.000 2316.010 3400.000 ;
    END
  END wbs_data_i[12]
  PIN wbs_data_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2405.890 0.000 2406.170 4.000 ;
    END
  END wbs_data_i[13]
  PIN wbs_data_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 3028.080 2850.000 3028.680 ;
    END
  END wbs_data_i[14]
  PIN wbs_data_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2434.410 3396.000 2434.690 3400.000 ;
    END
  END wbs_data_i[15]
  PIN wbs_data_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2452.350 0.000 2452.630 4.000 ;
    END
  END wbs_data_i[16]
  PIN wbs_data_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 3134.160 2850.000 3134.760 ;
    END
  END wbs_data_i[17]
  PIN wbs_data_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2499.270 0.000 2499.550 4.000 ;
    END
  END wbs_data_i[18]
  PIN wbs_data_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2545.730 0.000 2546.010 4.000 ;
    END
  END wbs_data_i[19]
  PIN wbs_data_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2312.510 0.000 2312.790 4.000 ;
    END
  END wbs_data_i[1]
  PIN wbs_data_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2553.090 3396.000 2553.370 3400.000 ;
    END
  END wbs_data_i[20]
  PIN wbs_data_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2580.640 4.000 2581.240 ;
    END
  END wbs_data_i[21]
  PIN wbs_data_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2592.650 0.000 2592.930 4.000 ;
    END
  END wbs_data_i[22]
  PIN wbs_data_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 3240.240 2850.000 3240.840 ;
    END
  END wbs_data_i[23]
  PIN wbs_data_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2706.440 4.000 2707.040 ;
    END
  END wbs_data_i[24]
  PIN wbs_data_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2671.770 3396.000 2672.050 3400.000 ;
    END
  END wbs_data_i[25]
  PIN wbs_data_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2639.570 0.000 2639.850 4.000 ;
    END
  END wbs_data_i[26]
  PIN wbs_data_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2686.030 0.000 2686.310 4.000 ;
    END
  END wbs_data_i[27]
  PIN wbs_data_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2732.950 0.000 2733.230 4.000 ;
    END
  END wbs_data_i[28]
  PIN wbs_data_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2832.920 4.000 2833.520 ;
    END
  END wbs_data_i[29]
  PIN wbs_data_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2390.240 2850.000 2390.840 ;
    END
  END wbs_data_i[2]
  PIN wbs_data_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2958.720 4.000 2959.320 ;
    END
  END wbs_data_i[30]
  PIN wbs_data_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2779.410 0.000 2779.690 4.000 ;
    END
  END wbs_data_i[31]
  PIN wbs_data_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2496.320 2850.000 2496.920 ;
    END
  END wbs_data_i[3]
  PIN wbs_data_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2077.910 3396.000 2078.190 3400.000 ;
    END
  END wbs_data_i[4]
  PIN wbs_data_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2197.050 3396.000 2197.330 3400.000 ;
    END
  END wbs_data_i[5]
  PIN wbs_data_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2358.970 0.000 2359.250 4.000 ;
    END
  END wbs_data_i[6]
  PIN wbs_data_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2603.080 2850.000 2603.680 ;
    END
  END wbs_data_i[7]
  PIN wbs_data_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2709.160 2850.000 2709.760 ;
    END
  END wbs_data_i[8]
  PIN wbs_data_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 2815.240 2850.000 2815.840 ;
    END
  END wbs_data_i[9]
  PIN wbs_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 396.610 0.000 396.890 4.000 ;
    END
  END wbs_data_o[0]
  PIN wbs_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 863.970 0.000 864.250 4.000 ;
    END
  END wbs_data_o[10]
  PIN wbs_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 910.430 0.000 910.710 4.000 ;
    END
  END wbs_data_o[11]
  PIN wbs_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 957.350 0.000 957.630 4.000 ;
    END
  END wbs_data_o[12]
  PIN wbs_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1004.270 0.000 1004.550 4.000 ;
    END
  END wbs_data_o[13]
  PIN wbs_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1050.730 0.000 1051.010 4.000 ;
    END
  END wbs_data_o[14]
  PIN wbs_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1097.650 0.000 1097.930 4.000 ;
    END
  END wbs_data_o[15]
  PIN wbs_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1144.110 0.000 1144.390 4.000 ;
    END
  END wbs_data_o[16]
  PIN wbs_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1191.030 0.000 1191.310 4.000 ;
    END
  END wbs_data_o[17]
  PIN wbs_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1237.490 0.000 1237.770 4.000 ;
    END
  END wbs_data_o[18]
  PIN wbs_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1284.410 0.000 1284.690 4.000 ;
    END
  END wbs_data_o[19]
  PIN wbs_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 443.530 0.000 443.810 4.000 ;
    END
  END wbs_data_o[1]
  PIN wbs_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1331.330 0.000 1331.610 4.000 ;
    END
  END wbs_data_o[20]
  PIN wbs_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1377.790 0.000 1378.070 4.000 ;
    END
  END wbs_data_o[21]
  PIN wbs_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1424.710 0.000 1424.990 4.000 ;
    END
  END wbs_data_o[22]
  PIN wbs_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1471.170 0.000 1471.450 4.000 ;
    END
  END wbs_data_o[23]
  PIN wbs_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1518.090 0.000 1518.370 4.000 ;
    END
  END wbs_data_o[24]
  PIN wbs_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1564.550 0.000 1564.830 4.000 ;
    END
  END wbs_data_o[25]
  PIN wbs_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1611.470 0.000 1611.750 4.000 ;
    END
  END wbs_data_o[26]
  PIN wbs_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1658.390 0.000 1658.670 4.000 ;
    END
  END wbs_data_o[27]
  PIN wbs_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1704.850 0.000 1705.130 4.000 ;
    END
  END wbs_data_o[28]
  PIN wbs_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1751.770 0.000 1752.050 4.000 ;
    END
  END wbs_data_o[29]
  PIN wbs_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 489.990 0.000 490.270 4.000 ;
    END
  END wbs_data_o[2]
  PIN wbs_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1798.230 0.000 1798.510 4.000 ;
    END
  END wbs_data_o[30]
  PIN wbs_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1845.150 0.000 1845.430 4.000 ;
    END
  END wbs_data_o[31]
  PIN wbs_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 536.910 0.000 537.190 4.000 ;
    END
  END wbs_data_o[3]
  PIN wbs_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 583.370 0.000 583.650 4.000 ;
    END
  END wbs_data_o[4]
  PIN wbs_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 630.290 0.000 630.570 4.000 ;
    END
  END wbs_data_o[5]
  PIN wbs_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 677.210 0.000 677.490 4.000 ;
    END
  END wbs_data_o[6]
  PIN wbs_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 723.670 0.000 723.950 4.000 ;
    END
  END wbs_data_o[7]
  PIN wbs_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 770.590 0.000 770.870 4.000 ;
    END
  END wbs_data_o[8]
  PIN wbs_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 817.050 0.000 817.330 4.000 ;
    END
  END wbs_data_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3084.520 4.000 3085.120 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3210.320 4.000 3210.920 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3336.120 4.000 3336.720 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2826.330 0.000 2826.610 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2790.450 3396.000 2790.730 3400.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2846.000 3346.320 2850.000 3346.920 ;
    END
  END wbs_we_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 2844.180 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 2844.180 104.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2844.180 3389.205 ;
      LAYER met1 ;
        RECT 5.520 4.460 2844.180 3389.360 ;
      LAYER met2 ;
        RECT 14.350 3395.720 59.150 3396.000 ;
        RECT 59.990 3395.720 177.830 3396.000 ;
        RECT 178.670 3395.720 296.510 3396.000 ;
        RECT 297.350 3395.720 415.190 3396.000 ;
        RECT 416.030 3395.720 533.870 3396.000 ;
        RECT 534.710 3395.720 652.550 3396.000 ;
        RECT 653.390 3395.720 771.690 3396.000 ;
        RECT 772.530 3395.720 890.370 3396.000 ;
        RECT 891.210 3395.720 1009.050 3396.000 ;
        RECT 1009.890 3395.720 1127.730 3396.000 ;
        RECT 1128.570 3395.720 1246.410 3396.000 ;
        RECT 1247.250 3395.720 1365.090 3396.000 ;
        RECT 1365.930 3395.720 1484.230 3396.000 ;
        RECT 1485.070 3395.720 1602.910 3396.000 ;
        RECT 1603.750 3395.720 1721.590 3396.000 ;
        RECT 1722.430 3395.720 1840.270 3396.000 ;
        RECT 1841.110 3395.720 1958.950 3396.000 ;
        RECT 1959.790 3395.720 2077.630 3396.000 ;
        RECT 2078.470 3395.720 2196.770 3396.000 ;
        RECT 2197.610 3395.720 2315.450 3396.000 ;
        RECT 2316.290 3395.720 2434.130 3396.000 ;
        RECT 2434.970 3395.720 2552.810 3396.000 ;
        RECT 2553.650 3395.720 2671.490 3396.000 ;
        RECT 2672.330 3395.720 2790.170 3396.000 ;
        RECT 2791.010 3395.720 2835.810 3396.000 ;
        RECT 14.350 4.280 2835.810 3395.720 ;
        RECT 14.350 4.000 22.810 4.280 ;
        RECT 23.650 4.000 69.270 4.280 ;
        RECT 70.110 4.000 116.190 4.280 ;
        RECT 117.030 4.000 162.650 4.280 ;
        RECT 163.490 4.000 209.570 4.280 ;
        RECT 210.410 4.000 256.030 4.280 ;
        RECT 256.870 4.000 302.950 4.280 ;
        RECT 303.790 4.000 349.870 4.280 ;
        RECT 350.710 4.000 396.330 4.280 ;
        RECT 397.170 4.000 443.250 4.280 ;
        RECT 444.090 4.000 489.710 4.280 ;
        RECT 490.550 4.000 536.630 4.280 ;
        RECT 537.470 4.000 583.090 4.280 ;
        RECT 583.930 4.000 630.010 4.280 ;
        RECT 630.850 4.000 676.930 4.280 ;
        RECT 677.770 4.000 723.390 4.280 ;
        RECT 724.230 4.000 770.310 4.280 ;
        RECT 771.150 4.000 816.770 4.280 ;
        RECT 817.610 4.000 863.690 4.280 ;
        RECT 864.530 4.000 910.150 4.280 ;
        RECT 910.990 4.000 957.070 4.280 ;
        RECT 957.910 4.000 1003.990 4.280 ;
        RECT 1004.830 4.000 1050.450 4.280 ;
        RECT 1051.290 4.000 1097.370 4.280 ;
        RECT 1098.210 4.000 1143.830 4.280 ;
        RECT 1144.670 4.000 1190.750 4.280 ;
        RECT 1191.590 4.000 1237.210 4.280 ;
        RECT 1238.050 4.000 1284.130 4.280 ;
        RECT 1284.970 4.000 1331.050 4.280 ;
        RECT 1331.890 4.000 1377.510 4.280 ;
        RECT 1378.350 4.000 1424.430 4.280 ;
        RECT 1425.270 4.000 1470.890 4.280 ;
        RECT 1471.730 4.000 1517.810 4.280 ;
        RECT 1518.650 4.000 1564.270 4.280 ;
        RECT 1565.110 4.000 1611.190 4.280 ;
        RECT 1612.030 4.000 1658.110 4.280 ;
        RECT 1658.950 4.000 1704.570 4.280 ;
        RECT 1705.410 4.000 1751.490 4.280 ;
        RECT 1752.330 4.000 1797.950 4.280 ;
        RECT 1798.790 4.000 1844.870 4.280 ;
        RECT 1845.710 4.000 1891.330 4.280 ;
        RECT 1892.170 4.000 1938.250 4.280 ;
        RECT 1939.090 4.000 1985.170 4.280 ;
        RECT 1986.010 4.000 2031.630 4.280 ;
        RECT 2032.470 4.000 2078.550 4.280 ;
        RECT 2079.390 4.000 2125.010 4.280 ;
        RECT 2125.850 4.000 2171.930 4.280 ;
        RECT 2172.770 4.000 2218.390 4.280 ;
        RECT 2219.230 4.000 2265.310 4.280 ;
        RECT 2266.150 4.000 2312.230 4.280 ;
        RECT 2313.070 4.000 2358.690 4.280 ;
        RECT 2359.530 4.000 2405.610 4.280 ;
        RECT 2406.450 4.000 2452.070 4.280 ;
        RECT 2452.910 4.000 2498.990 4.280 ;
        RECT 2499.830 4.000 2545.450 4.280 ;
        RECT 2546.290 4.000 2592.370 4.280 ;
        RECT 2593.210 4.000 2639.290 4.280 ;
        RECT 2640.130 4.000 2685.750 4.280 ;
        RECT 2686.590 4.000 2732.670 4.280 ;
        RECT 2733.510 4.000 2779.130 4.280 ;
        RECT 2779.970 4.000 2826.050 4.280 ;
        RECT 2826.890 4.000 2835.810 4.280 ;
      LAYER met3 ;
        RECT 4.000 3347.320 2846.000 3389.285 ;
        RECT 4.000 3345.920 2845.600 3347.320 ;
        RECT 4.000 3337.120 2846.000 3345.920 ;
        RECT 4.400 3335.720 2846.000 3337.120 ;
        RECT 4.000 3241.240 2846.000 3335.720 ;
        RECT 4.000 3239.840 2845.600 3241.240 ;
        RECT 4.000 3211.320 2846.000 3239.840 ;
        RECT 4.400 3209.920 2846.000 3211.320 ;
        RECT 4.000 3135.160 2846.000 3209.920 ;
        RECT 4.000 3133.760 2845.600 3135.160 ;
        RECT 4.000 3085.520 2846.000 3133.760 ;
        RECT 4.400 3084.120 2846.000 3085.520 ;
        RECT 4.000 3029.080 2846.000 3084.120 ;
        RECT 4.000 3027.680 2845.600 3029.080 ;
        RECT 4.000 2959.720 2846.000 3027.680 ;
        RECT 4.400 2958.320 2846.000 2959.720 ;
        RECT 4.000 2922.320 2846.000 2958.320 ;
        RECT 4.000 2920.920 2845.600 2922.320 ;
        RECT 4.000 2833.920 2846.000 2920.920 ;
        RECT 4.400 2832.520 2846.000 2833.920 ;
        RECT 4.000 2816.240 2846.000 2832.520 ;
        RECT 4.000 2814.840 2845.600 2816.240 ;
        RECT 4.000 2710.160 2846.000 2814.840 ;
        RECT 4.000 2708.760 2845.600 2710.160 ;
        RECT 4.000 2707.440 2846.000 2708.760 ;
        RECT 4.400 2706.040 2846.000 2707.440 ;
        RECT 4.000 2604.080 2846.000 2706.040 ;
        RECT 4.000 2602.680 2845.600 2604.080 ;
        RECT 4.000 2581.640 2846.000 2602.680 ;
        RECT 4.400 2580.240 2846.000 2581.640 ;
        RECT 4.000 2497.320 2846.000 2580.240 ;
        RECT 4.000 2495.920 2845.600 2497.320 ;
        RECT 4.000 2455.840 2846.000 2495.920 ;
        RECT 4.400 2454.440 2846.000 2455.840 ;
        RECT 4.000 2391.240 2846.000 2454.440 ;
        RECT 4.000 2389.840 2845.600 2391.240 ;
        RECT 4.000 2330.040 2846.000 2389.840 ;
        RECT 4.400 2328.640 2846.000 2330.040 ;
        RECT 4.000 2285.160 2846.000 2328.640 ;
        RECT 4.000 2283.760 2845.600 2285.160 ;
        RECT 4.000 2204.240 2846.000 2283.760 ;
        RECT 4.400 2202.840 2846.000 2204.240 ;
        RECT 4.000 2179.080 2846.000 2202.840 ;
        RECT 4.000 2177.680 2845.600 2179.080 ;
        RECT 4.000 2077.760 2846.000 2177.680 ;
        RECT 4.400 2076.360 2846.000 2077.760 ;
        RECT 4.000 2072.320 2846.000 2076.360 ;
        RECT 4.000 2070.920 2845.600 2072.320 ;
        RECT 4.000 1966.240 2846.000 2070.920 ;
        RECT 4.000 1964.840 2845.600 1966.240 ;
        RECT 4.000 1951.960 2846.000 1964.840 ;
        RECT 4.400 1950.560 2846.000 1951.960 ;
        RECT 4.000 1860.160 2846.000 1950.560 ;
        RECT 4.000 1858.760 2845.600 1860.160 ;
        RECT 4.000 1826.160 2846.000 1858.760 ;
        RECT 4.400 1824.760 2846.000 1826.160 ;
        RECT 4.000 1754.080 2846.000 1824.760 ;
        RECT 4.000 1752.680 2845.600 1754.080 ;
        RECT 4.000 1700.360 2846.000 1752.680 ;
        RECT 4.400 1698.960 2846.000 1700.360 ;
        RECT 4.000 1647.320 2846.000 1698.960 ;
        RECT 4.000 1645.920 2845.600 1647.320 ;
        RECT 4.000 1574.560 2846.000 1645.920 ;
        RECT 4.400 1573.160 2846.000 1574.560 ;
        RECT 4.000 1541.240 2846.000 1573.160 ;
        RECT 4.000 1539.840 2845.600 1541.240 ;
        RECT 4.000 1448.760 2846.000 1539.840 ;
        RECT 4.400 1447.360 2846.000 1448.760 ;
        RECT 4.000 1435.160 2846.000 1447.360 ;
        RECT 4.000 1433.760 2845.600 1435.160 ;
        RECT 4.000 1329.080 2846.000 1433.760 ;
        RECT 4.000 1327.680 2845.600 1329.080 ;
        RECT 4.000 1322.280 2846.000 1327.680 ;
        RECT 4.400 1320.880 2846.000 1322.280 ;
        RECT 4.000 1222.320 2846.000 1320.880 ;
        RECT 4.000 1220.920 2845.600 1222.320 ;
        RECT 4.000 1196.480 2846.000 1220.920 ;
        RECT 4.400 1195.080 2846.000 1196.480 ;
        RECT 4.000 1116.240 2846.000 1195.080 ;
        RECT 4.000 1114.840 2845.600 1116.240 ;
        RECT 4.000 1070.680 2846.000 1114.840 ;
        RECT 4.400 1069.280 2846.000 1070.680 ;
        RECT 4.000 1010.160 2846.000 1069.280 ;
        RECT 4.000 1008.760 2845.600 1010.160 ;
        RECT 4.000 944.880 2846.000 1008.760 ;
        RECT 4.400 943.480 2846.000 944.880 ;
        RECT 4.000 904.080 2846.000 943.480 ;
        RECT 4.000 902.680 2845.600 904.080 ;
        RECT 4.000 819.080 2846.000 902.680 ;
        RECT 4.400 817.680 2846.000 819.080 ;
        RECT 4.000 797.320 2846.000 817.680 ;
        RECT 4.000 795.920 2845.600 797.320 ;
        RECT 4.000 692.600 2846.000 795.920 ;
        RECT 4.400 691.240 2846.000 692.600 ;
        RECT 4.400 691.200 2845.600 691.240 ;
        RECT 4.000 689.840 2845.600 691.200 ;
        RECT 4.000 585.160 2846.000 689.840 ;
        RECT 4.000 583.760 2845.600 585.160 ;
        RECT 4.000 566.800 2846.000 583.760 ;
        RECT 4.400 565.400 2846.000 566.800 ;
        RECT 4.000 479.080 2846.000 565.400 ;
        RECT 4.000 477.680 2845.600 479.080 ;
        RECT 4.000 441.000 2846.000 477.680 ;
        RECT 4.400 439.600 2846.000 441.000 ;
        RECT 4.000 372.320 2846.000 439.600 ;
        RECT 4.000 370.920 2845.600 372.320 ;
        RECT 4.000 315.200 2846.000 370.920 ;
        RECT 4.400 313.800 2846.000 315.200 ;
        RECT 4.000 266.240 2846.000 313.800 ;
        RECT 4.000 264.840 2845.600 266.240 ;
        RECT 4.000 189.400 2846.000 264.840 ;
        RECT 4.400 188.000 2846.000 189.400 ;
        RECT 4.000 160.160 2846.000 188.000 ;
        RECT 4.000 158.760 2845.600 160.160 ;
        RECT 4.000 63.600 2846.000 158.760 ;
        RECT 4.400 62.200 2846.000 63.600 ;
        RECT 4.000 54.080 2846.000 62.200 ;
        RECT 4.000 52.680 2845.600 54.080 ;
        RECT 4.000 4.255 2846.000 52.680 ;
      LAYER met4 ;
        RECT 21.040 10.640 2788.225 3389.360 ;
      LAYER met5 ;
        RECT 5.520 179.670 2844.180 3321.460 ;
  END
END fpga
END LIBRARY

